magic
tech sky130A
magscale 1 2
timestamp 1725547224
<< viali >>
rect 15209 23613 15243 23647
rect 15301 23613 15335 23647
rect 18061 23613 18095 23647
rect 18245 23613 18279 23647
rect 47593 23613 47627 23647
rect 53297 23613 53331 23647
rect 54033 23613 54067 23647
rect 14565 23477 14599 23511
rect 15945 23477 15979 23511
rect 17417 23477 17451 23511
rect 18889 23477 18923 23511
rect 46857 23477 46891 23511
rect 47409 23477 47443 23511
rect 48237 23477 48271 23511
rect 52469 23477 52503 23511
rect 52745 23477 52779 23511
rect 53481 23477 53515 23511
rect 17785 23273 17819 23307
rect 53297 23273 53331 23307
rect 15485 23205 15519 23239
rect 19625 23205 19659 23239
rect 46949 23205 46983 23239
rect 47777 23205 47811 23239
rect 49985 23205 50019 23239
rect 55045 23205 55079 23239
rect 15577 23137 15611 23171
rect 46857 23137 46891 23171
rect 47593 23137 47627 23171
rect 48329 23137 48363 23171
rect 50721 23137 50755 23171
rect 55873 23137 55907 23171
rect 6653 23069 6687 23103
rect 12081 23069 12115 23103
rect 14105 23069 14139 23103
rect 16405 23069 16439 23103
rect 16672 23069 16706 23103
rect 18613 23069 18647 23103
rect 20361 23069 20395 23103
rect 22753 23069 22787 23103
rect 23581 23069 23615 23103
rect 34069 23069 34103 23103
rect 36461 23069 36495 23103
rect 40417 23069 40451 23103
rect 45569 23069 45603 23103
rect 48237 23069 48271 23103
rect 48605 23069 48639 23103
rect 51549 23069 51583 23103
rect 51917 23069 51951 23103
rect 53665 23069 53699 23103
rect 56609 23069 56643 23103
rect 14372 23001 14406 23035
rect 36829 23001 36863 23035
rect 47317 23001 47351 23035
rect 48872 23001 48906 23035
rect 52184 23001 52218 23035
rect 53932 23001 53966 23035
rect 6101 22933 6135 22967
rect 11529 22933 11563 22967
rect 16221 22933 16255 22967
rect 18061 22933 18095 22967
rect 19809 22933 19843 22967
rect 22201 22933 22235 22967
rect 23029 22933 23063 22967
rect 33425 22933 33459 22967
rect 34345 22933 34379 22967
rect 35909 22933 35943 22967
rect 39865 22933 39899 22967
rect 45017 22933 45051 22967
rect 46213 22933 46247 22967
rect 47409 22933 47443 22967
rect 48145 22933 48179 22967
rect 50169 22933 50203 22967
rect 50905 22933 50939 22967
rect 55321 22933 55355 22967
rect 56057 22933 56091 22967
rect 13001 22729 13035 22763
rect 15117 22729 15151 22763
rect 15577 22729 15611 22763
rect 18061 22729 18095 22763
rect 18153 22729 18187 22763
rect 18613 22729 18647 22763
rect 19901 22729 19935 22763
rect 23213 22729 23247 22763
rect 36093 22729 36127 22763
rect 36553 22729 36587 22763
rect 37933 22729 37967 22763
rect 47409 22729 47443 22763
rect 51549 22729 51583 22763
rect 52561 22729 52595 22763
rect 56609 22729 56643 22763
rect 21373 22661 21407 22695
rect 22100 22661 22134 22695
rect 36001 22661 36035 22695
rect 38844 22661 38878 22695
rect 52101 22661 52135 22695
rect 13645 22593 13679 22627
rect 13912 22593 13946 22627
rect 15485 22593 15519 22627
rect 16681 22593 16715 22627
rect 16948 22593 16982 22627
rect 18521 22593 18555 22627
rect 20269 22593 20303 22627
rect 33425 22593 33459 22627
rect 33885 22593 33919 22627
rect 35173 22593 35207 22627
rect 36461 22593 36495 22627
rect 44088 22593 44122 22627
rect 46285 22593 46319 22627
rect 48881 22593 48915 22627
rect 49157 22593 49191 22627
rect 50077 22593 50111 22627
rect 50169 22593 50203 22627
rect 50436 22593 50470 22627
rect 52193 22593 52227 22627
rect 54953 22593 54987 22627
rect 55229 22593 55263 22627
rect 55496 22593 55530 22627
rect 56701 22593 56735 22627
rect 3709 22525 3743 22559
rect 4445 22525 4479 22559
rect 7113 22525 7147 22559
rect 9781 22525 9815 22559
rect 10057 22525 10091 22559
rect 10701 22525 10735 22559
rect 11989 22525 12023 22559
rect 15761 22525 15795 22559
rect 16129 22525 16163 22559
rect 18705 22525 18739 22559
rect 19533 22525 19567 22559
rect 20361 22525 20395 22559
rect 20453 22525 20487 22559
rect 20729 22525 20763 22559
rect 21833 22525 21867 22559
rect 23857 22525 23891 22559
rect 26341 22525 26375 22559
rect 28457 22525 28491 22559
rect 29193 22525 29227 22559
rect 31585 22525 31619 22559
rect 32137 22525 32171 22559
rect 33241 22525 33275 22559
rect 33333 22525 33367 22559
rect 34437 22525 34471 22559
rect 36737 22525 36771 22559
rect 37381 22525 37415 22559
rect 38577 22525 38611 22559
rect 40601 22525 40635 22559
rect 41429 22525 41463 22559
rect 42073 22525 42107 22559
rect 42441 22525 42475 22559
rect 43821 22525 43855 22559
rect 45845 22525 45879 22559
rect 46029 22525 46063 22559
rect 49019 22525 49053 22559
rect 49893 22525 49927 22559
rect 52009 22525 52043 22559
rect 52929 22525 52963 22559
rect 53941 22525 53975 22559
rect 54079 22525 54113 22559
rect 54217 22525 54251 22559
rect 54493 22525 54527 22559
rect 55137 22525 55171 22559
rect 57253 22525 57287 22559
rect 4905 22457 4939 22491
rect 15025 22457 15059 22491
rect 18981 22457 19015 22491
rect 26801 22457 26835 22491
rect 33793 22457 33827 22491
rect 39957 22457 39991 22491
rect 45201 22457 45235 22491
rect 49433 22457 49467 22491
rect 3065 22389 3099 22423
rect 3893 22389 3927 22423
rect 6469 22389 6503 22423
rect 9229 22389 9263 22423
rect 10609 22389 10643 22423
rect 11345 22389 11379 22423
rect 12633 22389 12667 22423
rect 23305 22389 23339 22423
rect 25789 22389 25823 22423
rect 27261 22389 27295 22423
rect 27905 22389 27939 22423
rect 28641 22389 28675 22423
rect 30573 22389 30607 22423
rect 31033 22389 31067 22423
rect 32781 22389 32815 22423
rect 34621 22389 34655 22423
rect 38301 22389 38335 22423
rect 40049 22389 40083 22423
rect 40785 22389 40819 22423
rect 41521 22389 41555 22423
rect 43085 22389 43119 22423
rect 45293 22389 45327 22423
rect 47961 22389 47995 22423
rect 48237 22389 48271 22423
rect 53297 22389 53331 22423
rect 3801 22185 3835 22219
rect 7113 22185 7147 22219
rect 9597 22185 9631 22219
rect 10517 22185 10551 22219
rect 13829 22185 13863 22219
rect 20729 22185 20763 22219
rect 23397 22185 23431 22219
rect 25973 22185 26007 22219
rect 28917 22185 28951 22219
rect 31493 22185 31527 22219
rect 33885 22185 33919 22219
rect 39865 22185 39899 22219
rect 41797 22185 41831 22219
rect 42625 22185 42659 22219
rect 48973 22185 49007 22219
rect 4445 22049 4479 22083
rect 10149 22049 10183 22083
rect 12173 22049 12207 22083
rect 15025 22049 15059 22083
rect 15209 22049 15243 22083
rect 16359 22049 16393 22083
rect 16497 22049 16531 22083
rect 16773 22049 16807 22083
rect 17417 22049 17451 22083
rect 17693 22049 17727 22083
rect 17785 22049 17819 22083
rect 21373 22049 21407 22083
rect 22109 22049 22143 22083
rect 22385 22049 22419 22083
rect 22661 22049 22695 22083
rect 24041 22049 24075 22083
rect 25789 22049 25823 22083
rect 26525 22049 26559 22083
rect 31309 22049 31343 22083
rect 32045 22049 32079 22083
rect 35449 22049 35483 22083
rect 37473 22049 37507 22083
rect 38531 22049 38565 22083
rect 38669 22049 38703 22083
rect 38945 22049 38979 22083
rect 39405 22049 39439 22083
rect 40509 22049 40543 22083
rect 41705 22049 41739 22083
rect 42441 22049 42475 22083
rect 43177 22049 43211 22083
rect 45109 22049 45143 22083
rect 48605 22049 48639 22083
rect 49709 22049 49743 22083
rect 49893 22049 49927 22083
rect 50261 22049 50295 22083
rect 51549 22049 51583 22083
rect 53573 22049 53607 22083
rect 54585 22049 54619 22083
rect 54677 22049 54711 22083
rect 55413 22049 55447 22083
rect 2973 21981 3007 22015
rect 4721 21981 4755 22015
rect 5733 21981 5767 22015
rect 7757 21981 7791 22015
rect 11897 21981 11931 22015
rect 13369 21981 13403 22015
rect 16221 21981 16255 22015
rect 17233 21981 17267 22015
rect 19349 21981 19383 22015
rect 22247 21981 22281 22015
rect 23121 21981 23155 22015
rect 23305 21981 23339 22015
rect 24961 21981 24995 22015
rect 26341 21981 26375 22015
rect 26801 21981 26835 22015
rect 27537 21981 27571 22015
rect 30113 21981 30147 22015
rect 30573 21981 30607 22015
rect 32505 21981 32539 22015
rect 35265 21981 35299 22015
rect 37289 21981 37323 22015
rect 38393 21981 38427 22015
rect 39589 21981 39623 22015
rect 40325 21981 40359 22015
rect 40693 21981 40727 22015
rect 41245 21981 41279 22015
rect 43453 21981 43487 22015
rect 43720 21981 43754 22015
rect 45845 21981 45879 22015
rect 46397 21981 46431 22015
rect 46581 21981 46615 22015
rect 53389 21981 53423 22015
rect 55689 21981 55723 22015
rect 3617 21913 3651 21947
rect 4169 21913 4203 21947
rect 6000 21913 6034 21947
rect 9413 21913 9447 21947
rect 11630 21913 11664 21947
rect 17877 21913 17911 21947
rect 19616 21913 19650 21947
rect 23765 21913 23799 21947
rect 24409 21913 24443 21947
rect 27804 21913 27838 21947
rect 31033 21913 31067 21947
rect 32772 21913 32806 21947
rect 35716 21913 35750 21947
rect 42165 21913 42199 21947
rect 46848 21913 46882 21947
rect 48053 21913 48087 21947
rect 50537 21913 50571 21947
rect 51816 21913 51850 21947
rect 53481 21913 53515 21947
rect 4261 21845 4295 21879
rect 5273 21845 5307 21879
rect 7205 21845 7239 21879
rect 9965 21845 9999 21879
rect 10057 21845 10091 21879
rect 12265 21845 12299 21879
rect 12357 21845 12391 21879
rect 12725 21845 12759 21879
rect 12817 21845 12851 21879
rect 14381 21845 14415 21879
rect 14565 21845 14599 21879
rect 14933 21845 14967 21879
rect 15577 21845 15611 21879
rect 18245 21845 18279 21879
rect 18613 21845 18647 21879
rect 21465 21845 21499 21879
rect 23857 21845 23891 21879
rect 26433 21845 26467 21879
rect 27445 21845 27479 21879
rect 29285 21845 29319 21879
rect 29561 21845 29595 21879
rect 30665 21845 30699 21879
rect 31125 21845 31159 21879
rect 31861 21845 31895 21879
rect 31953 21845 31987 21879
rect 34161 21845 34195 21879
rect 34713 21845 34747 21879
rect 36829 21845 36863 21879
rect 36921 21845 36955 21879
rect 37381 21845 37415 21879
rect 37749 21845 37783 21879
rect 40233 21845 40267 21879
rect 42257 21845 42291 21879
rect 42993 21845 43027 21879
rect 43085 21845 43119 21879
rect 44833 21845 44867 21879
rect 45293 21845 45327 21879
rect 45385 21845 45419 21879
rect 45753 21845 45787 21879
rect 47961 21845 47995 21879
rect 49249 21845 49283 21879
rect 49617 21845 49651 21879
rect 50445 21845 50479 21879
rect 50905 21845 50939 21879
rect 52929 21845 52963 21879
rect 53021 21845 53055 21879
rect 54125 21845 54159 21879
rect 54493 21845 54527 21879
rect 55597 21845 55631 21879
rect 56057 21845 56091 21879
rect 1961 21641 1995 21675
rect 4813 21641 4847 21675
rect 5733 21641 5767 21675
rect 6193 21641 6227 21675
rect 10241 21641 10275 21675
rect 10609 21641 10643 21675
rect 11069 21641 11103 21675
rect 11529 21641 11563 21675
rect 14473 21641 14507 21675
rect 21373 21641 21407 21675
rect 23857 21641 23891 21675
rect 29285 21641 29319 21675
rect 31585 21641 31619 21675
rect 34069 21641 34103 21675
rect 34529 21641 34563 21675
rect 36829 21641 36863 21675
rect 37933 21641 37967 21675
rect 39589 21641 39623 21675
rect 39681 21641 39715 21675
rect 45201 21641 45235 21675
rect 45569 21641 45603 21675
rect 49065 21641 49099 21675
rect 51181 21641 51215 21675
rect 52561 21641 52595 21675
rect 52745 21641 52779 21675
rect 54125 21641 54159 21675
rect 54217 21641 54251 21675
rect 3074 21573 3108 21607
rect 6736 21573 6770 21607
rect 9128 21573 9162 21607
rect 12664 21573 12698 21607
rect 25596 21573 25630 21607
rect 30472 21573 30506 21607
rect 42717 21573 42751 21607
rect 45661 21573 45695 21607
rect 48789 21573 48823 21607
rect 3341 21505 3375 21539
rect 3433 21505 3467 21539
rect 3700 21505 3734 21539
rect 5825 21505 5859 21539
rect 10977 21505 11011 21539
rect 12909 21505 12943 21539
rect 15025 21505 15059 21539
rect 19165 21505 19199 21539
rect 21005 21505 21039 21539
rect 22477 21505 22511 21539
rect 22744 21505 22778 21539
rect 25329 21505 25363 21539
rect 27905 21505 27939 21539
rect 28825 21505 28859 21539
rect 32781 21505 32815 21539
rect 32940 21505 32974 21539
rect 33057 21505 33091 21539
rect 33793 21505 33827 21539
rect 33977 21505 34011 21539
rect 34437 21505 34471 21539
rect 35449 21505 35483 21539
rect 35716 21505 35750 21539
rect 37289 21505 37323 21539
rect 38476 21505 38510 21539
rect 40049 21505 40083 21539
rect 40877 21505 40911 21539
rect 41144 21505 41178 21539
rect 43683 21505 43717 21539
rect 43821 21505 43855 21539
rect 44557 21505 44591 21539
rect 44741 21505 44775 21539
rect 46213 21505 46247 21539
rect 48145 21505 48179 21539
rect 49617 21505 49651 21539
rect 51733 21505 51767 21539
rect 53297 21505 53331 21539
rect 53481 21505 53515 21539
rect 54769 21505 54803 21539
rect 5365 21437 5399 21471
rect 5641 21437 5675 21471
rect 6469 21437 6503 21471
rect 8493 21437 8527 21471
rect 8861 21437 8895 21471
rect 11253 21437 11287 21471
rect 27619 21437 27653 21471
rect 27767 21437 27801 21471
rect 28641 21437 28675 21471
rect 29377 21437 29411 21471
rect 29469 21437 29503 21471
rect 30205 21437 30239 21471
rect 34621 21437 34655 21471
rect 38209 21437 38243 21471
rect 40141 21437 40175 21471
rect 40325 21437 40359 21471
rect 43545 21437 43579 21471
rect 44925 21437 44959 21471
rect 45109 21437 45143 21471
rect 7849 21369 7883 21403
rect 26709 21369 26743 21403
rect 28181 21369 28215 21403
rect 33333 21369 33367 21403
rect 42257 21369 42291 21403
rect 44097 21369 44131 21403
rect 55229 21369 55263 21403
rect 7941 21301 7975 21335
rect 13277 21301 13311 21335
rect 15393 21301 15427 21335
rect 17417 21301 17451 21335
rect 19533 21301 19567 21335
rect 26985 21301 27019 21335
rect 28917 21301 28951 21335
rect 31861 21301 31895 21335
rect 32137 21301 32171 21335
rect 40785 21301 40819 21335
rect 42901 21301 42935 21335
rect 46673 21301 46707 21335
rect 50077 21301 50111 21335
rect 3985 21097 4019 21131
rect 7205 21097 7239 21131
rect 22201 21097 22235 21131
rect 22293 21097 22327 21131
rect 23397 21097 23431 21131
rect 29377 21097 29411 21131
rect 32229 21097 32263 21131
rect 33977 21097 34011 21131
rect 36369 21097 36403 21131
rect 39221 21097 39255 21131
rect 40417 21097 40451 21131
rect 44189 21097 44223 21131
rect 45201 21097 45235 21131
rect 45569 21097 45603 21131
rect 53941 21097 53975 21131
rect 20637 21029 20671 21063
rect 37657 21029 37691 21063
rect 42717 21029 42751 21063
rect 44741 21029 44775 21063
rect 54953 21029 54987 21063
rect 4445 20961 4479 20995
rect 4537 20961 4571 20995
rect 6055 20961 6089 20995
rect 6193 20961 6227 20995
rect 6469 20961 6503 20995
rect 7113 20961 7147 20995
rect 7849 20961 7883 20995
rect 10793 20961 10827 20995
rect 11253 20961 11287 20995
rect 11529 20961 11563 20995
rect 11805 20961 11839 20995
rect 16405 20961 16439 20995
rect 17049 20961 17083 20995
rect 21189 20961 21223 20995
rect 21281 20961 21315 20995
rect 21557 20961 21591 20995
rect 22937 20961 22971 20995
rect 25053 20961 25087 20995
rect 27077 20961 27111 20995
rect 27997 20961 28031 20995
rect 32597 20961 32631 20995
rect 36921 20961 36955 20995
rect 41337 20961 41371 20995
rect 43361 20961 43395 20995
rect 43545 20961 43579 20995
rect 48145 20961 48179 20995
rect 54585 20961 54619 20995
rect 4997 20893 5031 20927
rect 5917 20893 5951 20927
rect 6929 20893 6963 20927
rect 7573 20893 7607 20927
rect 8953 20893 8987 20927
rect 10609 20893 10643 20927
rect 11646 20893 11680 20927
rect 15025 20893 15059 20927
rect 15301 20893 15335 20927
rect 16865 20893 16899 20927
rect 17969 20893 18003 20927
rect 19257 20893 19291 20927
rect 21097 20893 21131 20927
rect 22753 20893 22787 20927
rect 27537 20893 27571 20927
rect 30113 20893 30147 20927
rect 31585 20893 31619 20927
rect 32864 20893 32898 20927
rect 55873 20893 55907 20927
rect 56057 20893 56091 20927
rect 57345 20893 57379 20927
rect 8309 20825 8343 20859
rect 9220 20825 9254 20859
rect 19524 20825 19558 20859
rect 25320 20825 25354 20859
rect 26893 20825 26927 20859
rect 28264 20825 28298 20859
rect 30380 20825 30414 20859
rect 37933 20825 37967 20859
rect 40049 20825 40083 20859
rect 41604 20825 41638 20859
rect 42809 20825 42843 20859
rect 4353 20757 4387 20791
rect 5273 20757 5307 20791
rect 7665 20757 7699 20791
rect 8677 20757 8711 20791
rect 10333 20757 10367 20791
rect 12449 20757 12483 20791
rect 14473 20757 14507 20791
rect 15853 20757 15887 20791
rect 16497 20757 16531 20791
rect 16957 20757 16991 20791
rect 17417 20757 17451 20791
rect 20729 20757 20763 20791
rect 22661 20757 22695 20791
rect 26433 20757 26467 20791
rect 26525 20757 26559 20791
rect 26985 20757 27019 20791
rect 31493 20757 31527 20791
rect 34253 20757 34287 20791
rect 49065 20757 49099 20791
rect 53113 20757 53147 20791
rect 55321 20757 55355 20791
rect 56701 20757 56735 20791
rect 56793 20757 56827 20791
rect 6929 20553 6963 20587
rect 7941 20553 7975 20587
rect 9781 20553 9815 20587
rect 10885 20553 10919 20587
rect 14473 20553 14507 20587
rect 17325 20553 17359 20587
rect 20177 20553 20211 20587
rect 21097 20553 21131 20587
rect 25973 20553 26007 20587
rect 27629 20553 27663 20587
rect 27905 20553 27939 20587
rect 28365 20553 28399 20587
rect 28733 20553 28767 20587
rect 30573 20553 30607 20587
rect 37657 20553 37691 20587
rect 55321 20553 55355 20587
rect 55689 20553 55723 20587
rect 11253 20485 11287 20519
rect 22201 20485 22235 20519
rect 28273 20485 28307 20519
rect 56600 20485 56634 20519
rect 9873 20417 9907 20451
rect 10333 20417 10367 20451
rect 14841 20417 14875 20451
rect 20729 20417 20763 20451
rect 26525 20417 26559 20451
rect 29285 20417 29319 20451
rect 31125 20417 31159 20451
rect 54585 20417 54619 20451
rect 55965 20417 55999 20451
rect 4537 20349 4571 20383
rect 7021 20349 7055 20383
rect 7205 20349 7239 20383
rect 10057 20349 10091 20383
rect 14933 20349 14967 20383
rect 15025 20349 15059 20383
rect 15485 20349 15519 20383
rect 16497 20349 16531 20383
rect 17049 20349 17083 20383
rect 17233 20349 17267 20383
rect 18245 20349 18279 20383
rect 23489 20349 23523 20383
rect 26985 20349 27019 20383
rect 28457 20349 28491 20383
rect 45569 20349 45603 20383
rect 48237 20349 48271 20383
rect 48421 20349 48455 20383
rect 54217 20349 54251 20383
rect 55045 20349 55079 20383
rect 55229 20349 55263 20383
rect 56333 20349 56367 20383
rect 58449 20349 58483 20383
rect 16129 20281 16163 20315
rect 17693 20281 17727 20315
rect 49341 20281 49375 20315
rect 50077 20281 50111 20315
rect 57713 20281 57747 20315
rect 5089 20213 5123 20247
rect 6561 20213 6595 20247
rect 7573 20213 7607 20247
rect 9413 20213 9447 20247
rect 14289 20213 14323 20247
rect 18889 20213 18923 20247
rect 22845 20213 22879 20247
rect 38393 20213 38427 20247
rect 39773 20213 39807 20247
rect 44833 20213 44867 20247
rect 44925 20213 44959 20247
rect 47685 20213 47719 20247
rect 49065 20213 49099 20247
rect 53665 20213 53699 20247
rect 57897 20213 57931 20247
rect 4537 20009 4571 20043
rect 8677 20009 8711 20043
rect 21741 20009 21775 20043
rect 23581 20009 23615 20043
rect 27813 20009 27847 20043
rect 48237 20009 48271 20043
rect 9321 19941 9355 19975
rect 10701 19941 10735 19975
rect 15485 19941 15519 19975
rect 16773 19941 16807 19975
rect 38577 19941 38611 19975
rect 44005 19941 44039 19975
rect 45753 19941 45787 19975
rect 48145 19941 48179 19975
rect 56517 19941 56551 19975
rect 3985 19873 4019 19907
rect 5733 19873 5767 19907
rect 9873 19873 9907 19907
rect 14105 19873 14139 19907
rect 16359 19873 16393 19907
rect 17233 19873 17267 19907
rect 22753 19873 22787 19907
rect 23029 19873 23063 19907
rect 23121 19873 23155 19907
rect 37473 19873 37507 19907
rect 39129 19873 39163 19907
rect 40049 19873 40083 19907
rect 44649 19873 44683 19907
rect 45109 19873 45143 19907
rect 46397 19873 46431 19907
rect 46765 19873 46799 19907
rect 48697 19873 48731 19907
rect 48789 19873 48823 19907
rect 49801 19873 49835 19907
rect 50261 19873 50295 19907
rect 50445 19873 50479 19907
rect 50997 19873 51031 19907
rect 52929 19873 52963 19907
rect 54953 19873 54987 19907
rect 55965 19873 55999 19907
rect 56241 19873 56275 19907
rect 57437 19873 57471 19907
rect 58265 19873 58299 19907
rect 4813 19805 4847 19839
rect 6561 19805 6595 19839
rect 14372 19805 14406 19839
rect 16221 19805 16255 19839
rect 16497 19805 16531 19839
rect 17417 19805 17451 19839
rect 18889 19805 18923 19839
rect 20269 19805 20303 19839
rect 20545 19805 20579 19839
rect 24961 19805 24995 19839
rect 26249 19805 26283 19839
rect 26525 19805 26559 19839
rect 30665 19805 30699 19839
rect 31401 19805 31435 19839
rect 35449 19805 35483 19839
rect 37657 19805 37691 19839
rect 40233 19805 40267 19839
rect 41981 19805 42015 19839
rect 44465 19805 44499 19839
rect 45293 19805 45327 19839
rect 47032 19805 47066 19839
rect 48605 19805 48639 19839
rect 49617 19805 49651 19839
rect 51549 19805 51583 19839
rect 52285 19805 52319 19839
rect 53196 19805 53230 19839
rect 54769 19805 54803 19839
rect 56124 19805 56158 19839
rect 56977 19805 57011 19839
rect 57161 19805 57195 19839
rect 4077 19737 4111 19771
rect 5457 19737 5491 19771
rect 10333 19737 10367 19771
rect 18622 19737 18656 19771
rect 21097 19737 21131 19771
rect 23213 19737 23247 19771
rect 24409 19737 24443 19771
rect 33793 19737 33827 19771
rect 35716 19737 35750 19771
rect 36921 19737 36955 19771
rect 39589 19737 39623 19771
rect 49709 19737 49743 19771
rect 4169 19669 4203 19703
rect 8033 19669 8067 19703
rect 13829 19669 13863 19703
rect 15577 19669 15611 19703
rect 17509 19669 17543 19703
rect 19717 19669 19751 19703
rect 22109 19669 22143 19703
rect 23857 19669 23891 19703
rect 25605 19669 25639 19703
rect 27077 19669 27111 19703
rect 27445 19669 27479 19703
rect 30113 19669 30147 19703
rect 30849 19669 30883 19703
rect 31769 19669 31803 19703
rect 33517 19669 33551 19703
rect 35357 19669 35391 19703
rect 36829 19669 36863 19703
rect 38301 19669 38335 19703
rect 38945 19669 38979 19703
rect 39037 19669 39071 19703
rect 40141 19669 40175 19703
rect 40601 19669 40635 19703
rect 41429 19669 41463 19703
rect 44097 19669 44131 19703
rect 44557 19669 44591 19703
rect 45385 19669 45419 19703
rect 45845 19669 45879 19703
rect 49249 19669 49283 19703
rect 50537 19669 50571 19703
rect 50905 19669 50939 19703
rect 51733 19669 51767 19703
rect 54309 19669 54343 19703
rect 54401 19669 54435 19703
rect 54861 19669 54895 19703
rect 55321 19669 55355 19703
rect 57529 19669 57563 19703
rect 57621 19669 57655 19703
rect 57989 19669 58023 19703
rect 3985 19465 4019 19499
rect 7757 19465 7791 19499
rect 11713 19465 11747 19499
rect 15209 19465 15243 19499
rect 15761 19465 15795 19499
rect 16681 19465 16715 19499
rect 19809 19465 19843 19499
rect 24133 19465 24167 19499
rect 26525 19465 26559 19499
rect 30297 19465 30331 19499
rect 30757 19465 30791 19499
rect 34069 19465 34103 19499
rect 36921 19465 36955 19499
rect 37749 19465 37783 19499
rect 45661 19465 45695 19499
rect 47409 19465 47443 19499
rect 47961 19465 47995 19499
rect 50353 19465 50387 19499
rect 54033 19465 54067 19499
rect 55965 19465 55999 19499
rect 57713 19465 57747 19499
rect 15669 19397 15703 19431
rect 20177 19397 20211 19431
rect 25412 19397 25446 19431
rect 35808 19397 35842 19431
rect 44548 19397 44582 19431
rect 47869 19397 47903 19431
rect 48421 19397 48455 19431
rect 51488 19397 51522 19431
rect 2513 19329 2547 19363
rect 2780 19329 2814 19363
rect 5098 19329 5132 19363
rect 5365 19329 5399 19363
rect 6377 19329 6411 19363
rect 6644 19329 6678 19363
rect 7849 19329 7883 19363
rect 11161 19329 11195 19363
rect 13829 19329 13863 19363
rect 14096 19329 14130 19363
rect 17805 19329 17839 19363
rect 18061 19329 18095 19363
rect 18705 19329 18739 19363
rect 20269 19329 20303 19363
rect 21833 19329 21867 19363
rect 22017 19329 22051 19363
rect 23673 19329 23707 19363
rect 24041 19329 24075 19363
rect 25145 19329 25179 19363
rect 27813 19329 27847 19363
rect 30665 19329 30699 19363
rect 32956 19329 32990 19363
rect 34161 19329 34195 19363
rect 35541 19329 35575 19363
rect 38531 19329 38565 19363
rect 39405 19329 39439 19363
rect 39681 19329 39715 19363
rect 39948 19329 39982 19363
rect 41153 19329 41187 19363
rect 44281 19329 44315 19363
rect 49203 19329 49237 19363
rect 49341 19329 49375 19363
rect 50261 19329 50295 19363
rect 51733 19329 51767 19363
rect 52745 19329 52779 19363
rect 54585 19329 54619 19363
rect 54852 19329 54886 19363
rect 56333 19329 56367 19363
rect 56600 19329 56634 19363
rect 57897 19329 57931 19363
rect 58449 19329 58483 19363
rect 5457 19261 5491 19295
rect 8401 19261 8435 19295
rect 9137 19261 9171 19295
rect 10241 19261 10275 19295
rect 10609 19261 10643 19295
rect 12633 19261 12667 19295
rect 15853 19261 15887 19295
rect 20361 19261 20395 19295
rect 20821 19261 20855 19295
rect 22753 19261 22787 19295
rect 22870 19261 22904 19295
rect 23029 19261 23063 19295
rect 23857 19261 23891 19295
rect 27169 19261 27203 19295
rect 30205 19261 30239 19295
rect 30941 19261 30975 19295
rect 31309 19261 31343 19295
rect 32689 19261 32723 19295
rect 34713 19261 34747 19295
rect 38393 19261 38427 19295
rect 38669 19261 38703 19295
rect 38945 19261 38979 19295
rect 39589 19261 39623 19295
rect 41705 19261 41739 19295
rect 42441 19261 42475 19295
rect 44189 19261 44223 19295
rect 46305 19261 46339 19295
rect 46765 19261 46799 19295
rect 47777 19261 47811 19295
rect 49065 19261 49099 19295
rect 50077 19261 50111 19295
rect 3893 19193 3927 19227
rect 22477 19193 22511 19227
rect 49617 19193 49651 19227
rect 6101 19125 6135 19159
rect 8585 19125 8619 19159
rect 9689 19125 9723 19159
rect 12081 19125 12115 19159
rect 13093 19125 13127 19159
rect 15301 19125 15335 19159
rect 16405 19125 16439 19159
rect 18153 19125 18187 19159
rect 19625 19125 19659 19159
rect 21465 19125 21499 19159
rect 24501 19125 24535 19159
rect 28089 19125 28123 19159
rect 29561 19125 29595 19159
rect 31953 19125 31987 19159
rect 32413 19125 32447 19159
rect 37565 19125 37599 19159
rect 41061 19125 41095 19159
rect 42073 19125 42107 19159
rect 43085 19125 43119 19159
rect 43361 19125 43395 19159
rect 43545 19125 43579 19159
rect 45753 19125 45787 19159
rect 48329 19125 48363 19159
rect 52469 19125 52503 19159
rect 2973 18921 3007 18955
rect 5181 18921 5215 18955
rect 7941 18921 7975 18955
rect 9689 18921 9723 18955
rect 9873 18921 9907 18955
rect 12357 18921 12391 18955
rect 14749 18921 14783 18955
rect 18153 18921 18187 18955
rect 20637 18921 20671 18955
rect 23949 18921 23983 18955
rect 25789 18921 25823 18955
rect 26985 18921 27019 18955
rect 31033 18921 31067 18955
rect 34345 18921 34379 18955
rect 36921 18921 36955 18955
rect 40601 18921 40635 18955
rect 41705 18921 41739 18955
rect 42809 18921 42843 18955
rect 46673 18921 46707 18955
rect 49985 18921 50019 18955
rect 54125 18921 54159 18955
rect 55965 18921 55999 18955
rect 56793 18921 56827 18955
rect 57713 18921 57747 18955
rect 3801 18853 3835 18887
rect 6377 18853 6411 18887
rect 9137 18853 9171 18887
rect 17417 18853 17451 18887
rect 32873 18853 32907 18887
rect 46305 18853 46339 18887
rect 3617 18785 3651 18819
rect 4445 18785 4479 18819
rect 4813 18785 4847 18819
rect 5963 18785 5997 18819
rect 6101 18785 6135 18819
rect 7297 18785 7331 18819
rect 8493 18785 8527 18819
rect 10425 18785 10459 18819
rect 13093 18785 13127 18819
rect 15301 18785 15335 18819
rect 16589 18785 16623 18819
rect 16773 18785 16807 18819
rect 17509 18785 17543 18819
rect 26341 18785 26375 18819
rect 27537 18785 27571 18819
rect 28365 18785 28399 18819
rect 29653 18785 29687 18819
rect 33701 18785 33735 18819
rect 35265 18785 35299 18819
rect 36001 18785 36035 18819
rect 36645 18785 36679 18819
rect 37473 18785 37507 18819
rect 40049 18785 40083 18819
rect 41245 18785 41279 18819
rect 42257 18785 42291 18819
rect 44097 18785 44131 18819
rect 44741 18785 44775 18819
rect 48053 18785 48087 18819
rect 53849 18785 53883 18819
rect 54677 18785 54711 18819
rect 55321 18785 55355 18819
rect 57345 18785 57379 18819
rect 58265 18785 58299 18819
rect 4169 18717 4203 18751
rect 5825 18717 5859 18751
rect 6837 18717 6871 18751
rect 7021 18717 7055 18751
rect 8401 18717 8435 18751
rect 10977 18717 11011 18751
rect 12909 18717 12943 18751
rect 13829 18717 13863 18751
rect 16957 18717 16991 18751
rect 19073 18717 19107 18751
rect 19257 18717 19291 18751
rect 21005 18717 21039 18751
rect 22477 18717 22511 18751
rect 22569 18717 22603 18751
rect 25605 18717 25639 18751
rect 27445 18717 27479 18751
rect 28181 18717 28215 18751
rect 29909 18717 29943 18751
rect 32321 18717 32355 18751
rect 32480 18717 32514 18751
rect 32597 18717 32631 18751
rect 33333 18717 33367 18751
rect 33517 18717 33551 18751
rect 33885 18717 33919 18751
rect 37381 18717 37415 18751
rect 38117 18717 38151 18751
rect 40233 18717 40267 18751
rect 40693 18717 40727 18751
rect 42073 18717 42107 18751
rect 43545 18717 43579 18751
rect 43704 18717 43738 18751
rect 43821 18717 43855 18751
rect 44557 18717 44591 18751
rect 48697 18717 48731 18751
rect 49341 18717 49375 18751
rect 51549 18717 51583 18751
rect 51825 18717 51859 18751
rect 53665 18717 53699 18751
rect 54493 18717 54527 18751
rect 57161 18717 57195 18751
rect 4261 18649 4295 18683
rect 7481 18649 7515 18683
rect 8309 18649 8343 18683
rect 10333 18649 10367 18683
rect 11222 18649 11256 18683
rect 12817 18649 12851 18683
rect 13277 18649 13311 18683
rect 19524 18649 19558 18683
rect 22210 18649 22244 18683
rect 22836 18649 22870 18683
rect 26157 18649 26191 18683
rect 27353 18649 27387 18683
rect 33977 18649 34011 18683
rect 34713 18649 34747 18683
rect 36461 18649 36495 18683
rect 38384 18649 38418 18683
rect 45017 18649 45051 18683
rect 45753 18649 45787 18683
rect 47808 18649 47842 18683
rect 48145 18649 48179 18683
rect 49065 18649 49099 18683
rect 51304 18649 51338 18683
rect 52092 18649 52126 18683
rect 56609 18649 56643 18683
rect 7389 18581 7423 18615
rect 7849 18581 7883 18615
rect 10241 18581 10275 18615
rect 12449 18581 12483 18615
rect 15669 18581 15703 18615
rect 17049 18581 17083 18615
rect 21097 18581 21131 18615
rect 24869 18581 24903 18615
rect 25053 18581 25087 18615
rect 26249 18581 26283 18615
rect 26801 18581 26835 18615
rect 27813 18581 27847 18615
rect 28273 18581 28307 18615
rect 31401 18581 31435 18615
rect 31677 18581 31711 18615
rect 36093 18581 36127 18615
rect 36553 18581 36587 18615
rect 37289 18581 37323 18615
rect 37933 18581 37967 18615
rect 39497 18581 39531 18615
rect 40141 18581 40175 18615
rect 42165 18581 42199 18615
rect 42901 18581 42935 18615
rect 50169 18581 50203 18615
rect 53205 18581 53239 18615
rect 53297 18581 53331 18615
rect 53757 18581 53791 18615
rect 54585 18581 54619 18615
rect 57253 18581 57287 18615
rect 7849 18377 7883 18411
rect 10609 18377 10643 18411
rect 10701 18377 10735 18411
rect 13829 18377 13863 18411
rect 20545 18377 20579 18411
rect 21097 18377 21131 18411
rect 31033 18377 31067 18411
rect 31401 18377 31435 18411
rect 34069 18377 34103 18411
rect 36001 18377 36035 18411
rect 37933 18377 37967 18411
rect 38485 18377 38519 18411
rect 39313 18377 39347 18411
rect 40693 18377 40727 18411
rect 42257 18377 42291 18411
rect 45109 18377 45143 18411
rect 47777 18377 47811 18411
rect 50169 18377 50203 18411
rect 51641 18377 51675 18411
rect 52745 18377 52779 18411
rect 54125 18377 54159 18411
rect 6193 18309 6227 18343
rect 21005 18309 21039 18343
rect 22201 18309 22235 18343
rect 25044 18309 25078 18343
rect 26709 18309 26743 18343
rect 28825 18309 28859 18343
rect 29828 18309 29862 18343
rect 34437 18309 34471 18343
rect 41144 18309 41178 18343
rect 42809 18309 42843 18343
rect 43974 18309 44008 18343
rect 45385 18309 45419 18343
rect 6377 18241 6411 18275
rect 6644 18241 6678 18275
rect 9229 18241 9263 18275
rect 9496 18241 9530 18275
rect 11713 18241 11747 18275
rect 13369 18241 13403 18275
rect 13737 18241 13771 18275
rect 19165 18241 19199 18275
rect 19432 18241 19466 18275
rect 22293 18241 22327 18275
rect 22661 18241 22695 18275
rect 24777 18241 24811 18275
rect 28181 18241 28215 18275
rect 29561 18241 29595 18275
rect 32137 18241 32171 18275
rect 32404 18241 32438 18275
rect 33977 18241 34011 18275
rect 36553 18241 36587 18275
rect 36921 18241 36955 18275
rect 37381 18241 37415 18275
rect 39037 18241 39071 18275
rect 39865 18241 39899 18275
rect 40877 18241 40911 18275
rect 43729 18241 43763 18275
rect 53297 18241 53331 18275
rect 8401 18173 8435 18207
rect 11253 18173 11287 18207
rect 11529 18173 11563 18207
rect 12449 18173 12483 18207
rect 12566 18173 12600 18207
rect 12725 18173 12759 18207
rect 13645 18173 13679 18207
rect 21189 18173 21223 18207
rect 22385 18173 22419 18207
rect 23213 18173 23247 18207
rect 26985 18173 27019 18207
rect 27169 18173 27203 18207
rect 27905 18173 27939 18207
rect 28022 18173 28056 18207
rect 29101 18173 29135 18207
rect 31493 18173 31527 18207
rect 31585 18173 31619 18207
rect 34253 18173 34287 18207
rect 34989 18173 35023 18207
rect 42533 18173 42567 18207
rect 42717 18173 42751 18207
rect 49893 18173 49927 18207
rect 50077 18173 50111 18207
rect 50997 18173 51031 18207
rect 53481 18173 53515 18207
rect 58449 18173 58483 18207
rect 7757 18105 7791 18139
rect 12173 18105 12207 18139
rect 27629 18105 27663 18139
rect 30941 18105 30975 18139
rect 33517 18105 33551 18139
rect 50537 18105 50571 18139
rect 8769 18037 8803 18071
rect 14197 18037 14231 18071
rect 20637 18037 20671 18071
rect 21833 18037 21867 18071
rect 24041 18037 24075 18071
rect 26157 18037 26191 18071
rect 33609 18037 33643 18071
rect 40233 18037 40267 18071
rect 43177 18037 43211 18071
rect 48145 18037 48179 18071
rect 49709 18037 49743 18071
rect 52561 18037 52595 18071
rect 54493 18037 54527 18071
rect 57897 18037 57931 18071
rect 6929 17833 6963 17867
rect 7941 17833 7975 17867
rect 11253 17833 11287 17867
rect 13461 17833 13495 17867
rect 20085 17833 20119 17867
rect 22293 17833 22327 17867
rect 22569 17833 22603 17867
rect 25329 17833 25363 17867
rect 25513 17833 25547 17867
rect 28457 17833 28491 17867
rect 33333 17833 33367 17867
rect 34529 17833 34563 17867
rect 41153 17833 41187 17867
rect 28365 17765 28399 17799
rect 33241 17765 33275 17799
rect 42717 17765 42751 17799
rect 53849 17765 53883 17799
rect 7573 17697 7607 17731
rect 9137 17697 9171 17731
rect 11161 17697 11195 17731
rect 11805 17697 11839 17731
rect 12081 17697 12115 17731
rect 13737 17697 13771 17731
rect 20729 17697 20763 17731
rect 21741 17697 21775 17731
rect 26157 17697 26191 17731
rect 26985 17697 27019 17731
rect 29009 17697 29043 17731
rect 32689 17697 32723 17731
rect 32781 17697 32815 17731
rect 33885 17697 33919 17731
rect 41337 17697 41371 17731
rect 43361 17697 43395 17731
rect 44465 17697 44499 17731
rect 44557 17697 44591 17731
rect 56885 17697 56919 17731
rect 3525 17629 3559 17663
rect 3801 17629 3835 17663
rect 11713 17629 11747 17663
rect 15669 17629 15703 17663
rect 15945 17629 15979 17663
rect 16957 17629 16991 17663
rect 24961 17629 24995 17663
rect 27252 17629 27286 17663
rect 36369 17629 36403 17663
rect 43821 17629 43855 17663
rect 53021 17629 53055 17663
rect 53113 17629 53147 17663
rect 54401 17629 54435 17663
rect 55873 17629 55907 17663
rect 56057 17629 56091 17663
rect 9404 17561 9438 17595
rect 12348 17561 12382 17595
rect 26801 17561 26835 17595
rect 30021 17561 30055 17595
rect 31769 17561 31803 17595
rect 32045 17561 32079 17595
rect 41604 17561 41638 17595
rect 42809 17561 42843 17595
rect 44373 17561 44407 17595
rect 57152 17561 57186 17595
rect 2973 17493 3007 17527
rect 4445 17493 4479 17527
rect 10517 17493 10551 17527
rect 11621 17493 11655 17527
rect 15117 17493 15151 17527
rect 16497 17493 16531 17527
rect 17601 17493 17635 17527
rect 18153 17493 18187 17527
rect 21005 17493 21039 17527
rect 21557 17493 21591 17527
rect 24409 17493 24443 17527
rect 25881 17493 25915 17527
rect 25973 17493 26007 17527
rect 32873 17493 32907 17527
rect 35817 17493 35851 17527
rect 37473 17493 37507 17527
rect 44005 17493 44039 17527
rect 52193 17493 52227 17527
rect 52377 17493 52411 17527
rect 53757 17493 53791 17527
rect 55321 17493 55355 17527
rect 56701 17493 56735 17527
rect 58265 17493 58299 17527
rect 3801 17289 3835 17323
rect 9689 17289 9723 17323
rect 11805 17289 11839 17323
rect 12449 17289 12483 17323
rect 15301 17289 15335 17323
rect 16681 17289 16715 17323
rect 19809 17289 19843 17323
rect 22753 17289 22787 17323
rect 26709 17289 26743 17323
rect 30941 17289 30975 17323
rect 31861 17289 31895 17323
rect 33425 17289 33459 17323
rect 35265 17289 35299 17323
rect 42809 17289 42843 17323
rect 52561 17289 52595 17323
rect 55965 17289 55999 17323
rect 57529 17289 57563 17323
rect 2688 17221 2722 17255
rect 8401 17221 8435 17255
rect 11253 17221 11287 17255
rect 15669 17221 15703 17255
rect 23664 17221 23698 17255
rect 29009 17221 29043 17255
rect 39497 17221 39531 17255
rect 51448 17221 51482 17255
rect 54852 17221 54886 17255
rect 56793 17221 56827 17255
rect 6653 17153 6687 17187
rect 6920 17153 6954 17187
rect 8125 17153 8159 17187
rect 10149 17153 10183 17187
rect 10609 17153 10643 17187
rect 13001 17153 13035 17187
rect 15761 17153 15795 17187
rect 17805 17153 17839 17187
rect 23397 17153 23431 17187
rect 25789 17153 25823 17187
rect 26157 17153 26191 17187
rect 34069 17153 34103 17187
rect 35357 17153 35391 17187
rect 39773 17153 39807 17187
rect 43453 17153 43487 17187
rect 48145 17153 48179 17187
rect 48412 17153 48446 17187
rect 50353 17153 50387 17187
rect 51181 17153 51215 17187
rect 53113 17153 53147 17187
rect 54585 17153 54619 17187
rect 56885 17153 56919 17187
rect 2421 17085 2455 17119
rect 3893 17085 3927 17119
rect 10241 17085 10275 17119
rect 10333 17085 10367 17119
rect 15853 17085 15887 17119
rect 18061 17085 18095 17119
rect 18889 17085 18923 17119
rect 20913 17085 20947 17119
rect 22385 17085 22419 17119
rect 25421 17085 25455 17119
rect 27813 17085 27847 17119
rect 28641 17085 28675 17119
rect 32321 17085 32355 17119
rect 34897 17085 34931 17119
rect 35173 17085 35207 17119
rect 36369 17085 36403 17119
rect 37933 17085 37967 17119
rect 38669 17085 38703 17119
rect 40049 17085 40083 17119
rect 41245 17085 41279 17119
rect 44189 17085 44223 17119
rect 49617 17085 49651 17119
rect 50905 17085 50939 17119
rect 52837 17085 52871 17119
rect 53021 17085 53055 17119
rect 54125 17085 54159 17119
rect 56701 17085 56735 17119
rect 58449 17085 58483 17119
rect 8033 17017 8067 17051
rect 16313 17017 16347 17051
rect 21649 17017 21683 17051
rect 24777 17017 24811 17051
rect 35725 17017 35759 17051
rect 49525 17017 49559 17051
rect 53481 17017 53515 17051
rect 57253 17017 57287 17051
rect 57897 17017 57931 17051
rect 4537 16949 4571 16983
rect 9781 16949 9815 16983
rect 14841 16949 14875 16983
rect 15209 16949 15243 16983
rect 18337 16949 18371 16983
rect 20361 16949 20395 16983
rect 21833 16949 21867 16983
rect 24869 16949 24903 16983
rect 27261 16949 27295 16983
rect 28089 16949 28123 16983
rect 32965 16949 32999 16983
rect 33793 16949 33827 16983
rect 34529 16949 34563 16983
rect 35817 16949 35851 16983
rect 36737 16949 36771 16983
rect 37289 16949 37323 16983
rect 38025 16949 38059 16983
rect 40693 16949 40727 16983
rect 43545 16949 43579 16983
rect 50261 16949 50295 16983
rect 53573 16949 53607 16983
rect 56333 16949 56367 16983
rect 6837 16745 6871 16779
rect 8585 16745 8619 16779
rect 9597 16745 9631 16779
rect 15945 16745 15979 16779
rect 16313 16745 16347 16779
rect 18245 16745 18279 16779
rect 19257 16745 19291 16779
rect 21833 16745 21867 16779
rect 27261 16745 27295 16779
rect 28457 16745 28491 16779
rect 30481 16745 30515 16779
rect 44557 16745 44591 16779
rect 45477 16745 45511 16779
rect 50169 16745 50203 16779
rect 53205 16745 53239 16779
rect 55137 16745 55171 16779
rect 3893 16677 3927 16711
rect 9229 16677 9263 16711
rect 23489 16677 23523 16711
rect 36093 16677 36127 16711
rect 40601 16677 40635 16711
rect 54309 16677 54343 16711
rect 1593 16609 1627 16643
rect 5273 16609 5307 16643
rect 6745 16609 6779 16643
rect 10149 16609 10183 16643
rect 16957 16609 16991 16643
rect 17233 16609 17267 16643
rect 17509 16609 17543 16643
rect 18153 16609 18187 16643
rect 18705 16609 18739 16643
rect 18797 16609 18831 16643
rect 19809 16609 19843 16643
rect 20545 16609 20579 16643
rect 22477 16609 22511 16643
rect 22845 16609 22879 16643
rect 23029 16609 23063 16643
rect 24133 16609 24167 16643
rect 24869 16609 24903 16643
rect 24961 16609 24995 16643
rect 25513 16609 25547 16643
rect 27721 16609 27755 16643
rect 27905 16609 27939 16643
rect 33333 16609 33367 16643
rect 34713 16609 34747 16643
rect 36185 16609 36219 16643
rect 39037 16609 39071 16643
rect 40049 16609 40083 16643
rect 40141 16609 40175 16643
rect 41245 16609 41279 16643
rect 41429 16609 41463 16643
rect 42901 16609 42935 16643
rect 45661 16609 45695 16643
rect 47869 16609 47903 16643
rect 49893 16609 49927 16643
rect 50721 16609 50755 16643
rect 51733 16609 51767 16643
rect 53665 16609 53699 16643
rect 53757 16609 53791 16643
rect 54493 16609 54527 16643
rect 54677 16609 54711 16643
rect 55505 16609 55539 16643
rect 55689 16609 55723 16643
rect 56885 16609 56919 16643
rect 57529 16609 57563 16643
rect 58081 16609 58115 16643
rect 58173 16609 58207 16643
rect 3249 16541 3283 16575
rect 3525 16541 3559 16575
rect 7021 16541 7055 16575
rect 7205 16541 7239 16575
rect 7297 16541 7331 16575
rect 8309 16541 8343 16575
rect 14565 16541 14599 16575
rect 14832 16541 14866 16575
rect 17095 16541 17129 16575
rect 17969 16541 18003 16575
rect 21097 16541 21131 16575
rect 22293 16541 22327 16575
rect 24777 16541 24811 16575
rect 28733 16541 28767 16575
rect 30205 16541 30239 16575
rect 32137 16541 32171 16575
rect 32505 16541 32539 16575
rect 34161 16541 34195 16575
rect 34980 16541 35014 16575
rect 36452 16541 36486 16575
rect 40233 16541 40267 16575
rect 43168 16541 43202 16575
rect 47685 16541 47719 16575
rect 50997 16541 51031 16575
rect 52000 16541 52034 16575
rect 56333 16541 56367 16575
rect 56471 16541 56505 16575
rect 56609 16541 56643 16575
rect 57345 16541 57379 16575
rect 1860 16473 1894 16507
rect 5006 16473 5040 16507
rect 7573 16473 7607 16507
rect 18613 16473 18647 16507
rect 20361 16473 20395 16507
rect 21741 16473 21775 16507
rect 25780 16473 25814 16507
rect 27629 16473 27663 16507
rect 29561 16473 29595 16507
rect 38792 16473 38826 16507
rect 42073 16473 42107 16507
rect 45928 16473 45962 16507
rect 47133 16473 47167 16507
rect 48136 16473 48170 16507
rect 49341 16473 49375 16507
rect 2973 16405 3007 16439
rect 3065 16405 3099 16439
rect 3433 16405 3467 16439
rect 19993 16405 20027 16439
rect 20453 16405 20487 16439
rect 22201 16405 22235 16439
rect 23121 16405 23155 16439
rect 23581 16405 23615 16439
rect 24409 16405 24443 16439
rect 26893 16405 26927 16439
rect 29377 16405 29411 16439
rect 31309 16405 31343 16439
rect 31493 16405 31527 16439
rect 33609 16405 33643 16439
rect 37565 16405 37599 16439
rect 37657 16405 37691 16439
rect 39589 16405 39623 16439
rect 40693 16405 40727 16439
rect 42349 16405 42383 16439
rect 42717 16405 42751 16439
rect 44281 16405 44315 16439
rect 47041 16405 47075 16439
rect 49249 16405 49283 16439
rect 50537 16405 50571 16439
rect 50629 16405 50663 16439
rect 51641 16405 51675 16439
rect 53113 16405 53147 16439
rect 53573 16405 53607 16439
rect 54769 16405 54803 16439
rect 57621 16405 57655 16439
rect 57989 16405 58023 16439
rect 2513 16201 2547 16235
rect 3893 16201 3927 16235
rect 4905 16201 4939 16235
rect 16129 16201 16163 16235
rect 18613 16201 18647 16235
rect 20821 16201 20855 16235
rect 20913 16201 20947 16235
rect 21281 16201 21315 16235
rect 21373 16201 21407 16235
rect 24961 16201 24995 16235
rect 25881 16201 25915 16235
rect 26433 16201 26467 16235
rect 29929 16201 29963 16235
rect 30389 16201 30423 16235
rect 31953 16201 31987 16235
rect 32137 16201 32171 16235
rect 32597 16201 32631 16235
rect 33701 16201 33735 16235
rect 38025 16201 38059 16235
rect 43821 16201 43855 16235
rect 45201 16201 45235 16235
rect 50445 16201 50479 16235
rect 53205 16201 53239 16235
rect 55873 16201 55907 16235
rect 5273 16133 5307 16167
rect 8401 16133 8435 16167
rect 17408 16133 17442 16167
rect 19708 16133 19742 16167
rect 27252 16133 27286 16167
rect 28816 16133 28850 16167
rect 30840 16133 30874 16167
rect 39120 16133 39154 16167
rect 47317 16133 47351 16167
rect 51580 16133 51614 16167
rect 51917 16133 51951 16167
rect 53113 16133 53147 16167
rect 56324 16133 56358 16167
rect 57897 16133 57931 16167
rect 3065 16065 3099 16099
rect 3249 16065 3283 16099
rect 5181 16065 5215 16099
rect 5365 16065 5399 16099
rect 5549 16065 5583 16099
rect 7113 16065 7147 16099
rect 8217 16065 8251 16099
rect 14556 16065 14590 16099
rect 22477 16065 22511 16099
rect 22753 16065 22787 16099
rect 23489 16065 23523 16099
rect 23765 16065 23799 16099
rect 26985 16065 27019 16099
rect 30573 16065 30607 16099
rect 32505 16065 32539 16099
rect 33241 16065 33275 16099
rect 33333 16065 33367 16099
rect 34060 16065 34094 16099
rect 36185 16065 36219 16099
rect 37105 16065 37139 16099
rect 37657 16065 37691 16099
rect 38669 16065 38703 16099
rect 40785 16065 40819 16099
rect 43913 16065 43947 16099
rect 44281 16065 44315 16099
rect 45661 16065 45695 16099
rect 45928 16065 45962 16099
rect 48237 16065 48271 16099
rect 50077 16065 50111 16099
rect 51825 16065 51859 16099
rect 54125 16065 54159 16099
rect 54392 16065 54426 16099
rect 56057 16065 56091 16099
rect 58449 16065 58483 16099
rect 4353 15997 4387 16031
rect 6745 15997 6779 16031
rect 7481 15997 7515 16031
rect 9045 15997 9079 16031
rect 10885 15997 10919 16031
rect 13001 15997 13035 16031
rect 13737 15997 13771 16031
rect 14289 15997 14323 16031
rect 16221 15997 16255 16031
rect 16313 15997 16347 16031
rect 17141 15997 17175 16031
rect 19165 15997 19199 16031
rect 19441 15997 19475 16031
rect 21465 15997 21499 16031
rect 22615 15997 22649 16031
rect 23673 15997 23707 16031
rect 24317 15997 24351 16031
rect 26157 15997 26191 16031
rect 26341 15997 26375 16031
rect 28549 15997 28583 16031
rect 32689 15997 32723 16031
rect 33149 15997 33183 16031
rect 33793 15997 33827 16031
rect 35909 15997 35943 16031
rect 36047 15997 36081 16031
rect 36921 15997 36955 16031
rect 37381 15997 37415 16031
rect 37565 15997 37599 16031
rect 38853 15997 38887 16031
rect 40509 15997 40543 16031
rect 40693 15997 40727 16031
rect 41797 15997 41831 16031
rect 42441 15997 42475 16031
rect 42993 15997 43027 16031
rect 44005 15997 44039 16031
rect 44925 15997 44959 16031
rect 48396 15997 48430 16031
rect 48513 15997 48547 16031
rect 49249 15997 49283 16031
rect 49433 15997 49467 16031
rect 52561 15997 52595 16031
rect 53297 15997 53331 16031
rect 53757 15997 53791 16031
rect 4997 15929 5031 15963
rect 9781 15929 9815 15963
rect 15669 15929 15703 15963
rect 18521 15929 18555 15963
rect 23029 15929 23063 15963
rect 36461 15929 36495 15963
rect 38117 15929 38151 15963
rect 41153 15929 41187 15963
rect 43453 15929 43487 15963
rect 48789 15929 48823 15963
rect 49525 15929 49559 15963
rect 52745 15929 52779 15963
rect 57437 15929 57471 15963
rect 6193 15861 6227 15895
rect 9413 15861 9447 15895
rect 10333 15861 10367 15895
rect 11805 15861 11839 15895
rect 12449 15861 12483 15895
rect 13185 15861 13219 15895
rect 15761 15861 15795 15895
rect 16865 15861 16899 15895
rect 21833 15861 21867 15895
rect 25513 15861 25547 15895
rect 26801 15861 26835 15895
rect 28365 15861 28399 15895
rect 35173 15861 35207 15895
rect 35265 15861 35299 15895
rect 40233 15861 40267 15895
rect 41245 15861 41279 15895
rect 42165 15861 42199 15895
rect 47041 15861 47075 15895
rect 47593 15861 47627 15895
rect 55505 15861 55539 15895
rect 3249 15657 3283 15691
rect 3985 15657 4019 15691
rect 4813 15657 4847 15691
rect 5549 15657 5583 15691
rect 6561 15657 6595 15691
rect 10425 15657 10459 15691
rect 13461 15657 13495 15691
rect 15209 15657 15243 15691
rect 16589 15657 16623 15691
rect 17509 15657 17543 15691
rect 21097 15657 21131 15691
rect 24133 15657 24167 15691
rect 25973 15657 26007 15691
rect 26709 15657 26743 15691
rect 28549 15657 28583 15691
rect 39037 15657 39071 15691
rect 42533 15657 42567 15691
rect 45937 15657 45971 15691
rect 47041 15657 47075 15691
rect 48145 15657 48179 15691
rect 49065 15657 49099 15691
rect 51457 15657 51491 15691
rect 55965 15657 55999 15691
rect 57897 15657 57931 15691
rect 4261 15589 4295 15623
rect 4353 15589 4387 15623
rect 9229 15589 9263 15623
rect 37013 15589 37047 15623
rect 37933 15589 37967 15623
rect 44005 15589 44039 15623
rect 52929 15589 52963 15623
rect 5457 15521 5491 15555
rect 6285 15521 6319 15555
rect 10333 15521 10367 15555
rect 10977 15521 11011 15555
rect 15761 15521 15795 15555
rect 15945 15521 15979 15555
rect 16865 15521 16899 15555
rect 17049 15521 17083 15555
rect 26617 15521 26651 15555
rect 27261 15521 27295 15555
rect 27997 15521 28031 15555
rect 29193 15521 29227 15555
rect 31861 15521 31895 15555
rect 32505 15521 32539 15555
rect 35265 15521 35299 15555
rect 35541 15521 35575 15555
rect 37289 15521 37323 15555
rect 38393 15521 38427 15555
rect 41521 15521 41555 15555
rect 41705 15521 41739 15555
rect 42625 15521 42659 15555
rect 44741 15521 44775 15555
rect 45569 15521 45603 15555
rect 46857 15521 46891 15555
rect 47501 15521 47535 15555
rect 47593 15521 47627 15555
rect 48513 15521 48547 15555
rect 49249 15521 49283 15555
rect 52377 15521 52411 15555
rect 52653 15521 52687 15555
rect 53389 15521 53423 15555
rect 53573 15521 53607 15555
rect 54953 15521 54987 15555
rect 55413 15521 55447 15555
rect 56885 15521 56919 15555
rect 57069 15521 57103 15555
rect 58449 15521 58483 15555
rect 2697 15453 2731 15487
rect 3065 15453 3099 15487
rect 4169 15453 4203 15487
rect 4445 15453 4479 15487
rect 4629 15453 4663 15487
rect 4721 15453 4755 15487
rect 4905 15453 4939 15487
rect 5825 15453 5859 15487
rect 6101 15453 6135 15487
rect 6929 15453 6963 15487
rect 7665 15453 7699 15487
rect 8953 15453 8987 15487
rect 9045 15453 9079 15487
rect 11805 15453 11839 15487
rect 12081 15453 12115 15487
rect 12348 15453 12382 15487
rect 18613 15453 18647 15487
rect 18981 15453 19015 15487
rect 19257 15453 19291 15487
rect 21281 15453 21315 15487
rect 22753 15453 22787 15487
rect 27721 15453 27755 15487
rect 28181 15453 28215 15487
rect 29561 15453 29595 15487
rect 30389 15453 30423 15487
rect 31309 15453 31343 15487
rect 31447 15453 31481 15487
rect 31585 15453 31619 15487
rect 32321 15453 32355 15487
rect 32597 15453 32631 15487
rect 32864 15453 32898 15487
rect 35081 15453 35115 15487
rect 36185 15453 36219 15487
rect 37565 15453 37599 15487
rect 39957 15453 39991 15487
rect 41797 15453 41831 15487
rect 44465 15453 44499 15487
rect 46673 15453 46707 15487
rect 47409 15453 47443 15487
rect 48605 15453 48639 15487
rect 49801 15453 49835 15487
rect 52536 15453 52570 15487
rect 54217 15453 54251 15487
rect 54769 15453 54803 15487
rect 2881 15385 2915 15419
rect 2973 15385 3007 15419
rect 5549 15385 5583 15419
rect 6377 15385 6411 15419
rect 6593 15385 6627 15419
rect 7389 15385 7423 15419
rect 8493 15385 8527 15419
rect 9229 15385 9263 15419
rect 13737 15385 13771 15419
rect 19524 15385 19558 15419
rect 21548 15385 21582 15419
rect 23020 15385 23054 15419
rect 28089 15385 28123 15419
rect 29009 15385 29043 15419
rect 35173 15385 35207 15419
rect 37473 15385 37507 15419
rect 40224 15385 40258 15419
rect 42892 15385 42926 15419
rect 46581 15385 46615 15419
rect 48697 15385 48731 15419
rect 57161 15385 57195 15419
rect 5733 15317 5767 15351
rect 5917 15317 5951 15351
rect 6745 15317 6779 15351
rect 9873 15317 9907 15351
rect 10793 15317 10827 15351
rect 10885 15317 10919 15351
rect 11253 15317 11287 15351
rect 15025 15317 15059 15351
rect 17141 15317 17175 15351
rect 18153 15317 18187 15351
rect 20637 15317 20671 15351
rect 22661 15317 22695 15351
rect 24593 15317 24627 15351
rect 28641 15317 28675 15351
rect 29101 15317 29135 15351
rect 30665 15317 30699 15351
rect 33977 15317 34011 15351
rect 34345 15317 34379 15351
rect 34713 15317 34747 15351
rect 36645 15317 36679 15351
rect 39589 15317 39623 15351
rect 41337 15317 41371 15351
rect 42165 15317 42199 15351
rect 44097 15317 44131 15351
rect 44557 15317 44591 15351
rect 45017 15317 45051 15351
rect 46213 15317 46247 15351
rect 50353 15317 50387 15351
rect 51733 15317 51767 15351
rect 54401 15317 54435 15351
rect 54861 15317 54895 15351
rect 56701 15317 56735 15351
rect 57529 15317 57563 15351
rect 2605 15113 2639 15147
rect 2697 15113 2731 15147
rect 2973 15113 3007 15147
rect 3893 15113 3927 15147
rect 4629 15113 4663 15147
rect 5825 15113 5859 15147
rect 9597 15113 9631 15147
rect 11529 15113 11563 15147
rect 15761 15113 15795 15147
rect 17969 15113 18003 15147
rect 19073 15113 19107 15147
rect 19809 15113 19843 15147
rect 21189 15113 21223 15147
rect 23121 15113 23155 15147
rect 30205 15113 30239 15147
rect 31953 15113 31987 15147
rect 33701 15113 33735 15147
rect 34437 15113 34471 15147
rect 41337 15113 41371 15147
rect 44373 15113 44407 15147
rect 46121 15113 46155 15147
rect 47133 15113 47167 15147
rect 48237 15113 48271 15147
rect 51641 15113 51675 15147
rect 54401 15113 54435 15147
rect 10140 15045 10174 15079
rect 16681 15045 16715 15079
rect 18797 15045 18831 15079
rect 28641 15045 28675 15079
rect 28978 15045 29012 15079
rect 31125 15045 31159 15079
rect 32137 15045 32171 15079
rect 40132 15045 40166 15079
rect 2789 14977 2823 15011
rect 2881 14977 2915 15011
rect 3157 14977 3191 15011
rect 3249 14977 3283 15011
rect 3801 14977 3835 15011
rect 4077 14977 4111 15011
rect 4721 14977 4755 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 7573 14977 7607 15011
rect 7665 14977 7699 15011
rect 7849 14977 7883 15011
rect 7941 14977 7975 15011
rect 8033 14977 8067 15011
rect 13369 14977 13403 15011
rect 13829 14977 13863 15011
rect 14289 14977 14323 15011
rect 20361 14977 20395 15011
rect 20637 14977 20671 15011
rect 22569 14977 22603 15011
rect 28089 14977 28123 15011
rect 28733 14977 28767 15011
rect 30849 14977 30883 15011
rect 34253 14977 34287 15011
rect 34989 14977 35023 15011
rect 41981 14977 42015 15011
rect 43223 14977 43257 15011
rect 43361 14977 43395 15011
rect 44281 14977 44315 15011
rect 46673 14977 46707 15011
rect 47593 14977 47627 15011
rect 48605 14977 48639 15011
rect 54953 14977 54987 15011
rect 2513 14909 2547 14943
rect 3341 14909 3375 14943
rect 3433 14909 3467 14943
rect 4353 14909 4387 14943
rect 7297 14909 7331 14943
rect 8309 14909 8343 14943
rect 9873 14909 9907 14943
rect 12173 14909 12207 14943
rect 12311 14909 12345 14943
rect 12449 14909 12483 14943
rect 13185 14909 13219 14943
rect 13921 14909 13955 14943
rect 14105 14909 14139 14943
rect 14841 14909 14875 14943
rect 32873 14909 32907 14943
rect 33333 14909 33367 14943
rect 35725 14909 35759 14943
rect 39865 14909 39899 14943
rect 43085 14909 43119 14943
rect 44097 14909 44131 14943
rect 44925 14909 44959 14943
rect 49617 14909 49651 14943
rect 50261 14909 50295 14943
rect 4261 14841 4295 14875
rect 6193 14841 6227 14875
rect 7941 14841 7975 14875
rect 12725 14841 12759 14875
rect 30113 14841 30147 14875
rect 41245 14841 41279 14875
rect 43637 14841 43671 14875
rect 51917 14841 51951 14875
rect 4445 14773 4479 14807
rect 4537 14773 4571 14807
rect 6561 14773 6595 14807
rect 11253 14773 11287 14807
rect 13461 14773 13495 14807
rect 16405 14773 16439 14807
rect 21465 14773 21499 14807
rect 23489 14773 23523 14807
rect 35357 14773 35391 14807
rect 42441 14773 42475 14807
rect 46029 14773 46063 14807
rect 48973 14773 49007 14807
rect 49709 14773 49743 14807
rect 57437 14773 57471 14807
rect 3249 14569 3283 14603
rect 4537 14569 4571 14603
rect 6469 14569 6503 14603
rect 6929 14569 6963 14603
rect 14289 14569 14323 14603
rect 18889 14569 18923 14603
rect 21189 14569 21223 14603
rect 27813 14569 27847 14603
rect 28733 14569 28767 14603
rect 30665 14569 30699 14603
rect 32413 14569 32447 14603
rect 34989 14569 35023 14603
rect 35357 14569 35391 14603
rect 37749 14569 37783 14603
rect 41429 14569 41463 14603
rect 48513 14569 48547 14603
rect 49709 14569 49743 14603
rect 54125 14569 54159 14603
rect 56793 14569 56827 14603
rect 11069 14501 11103 14535
rect 13553 14501 13587 14535
rect 30941 14501 30975 14535
rect 52009 14501 52043 14535
rect 9689 14433 9723 14467
rect 11161 14433 11195 14467
rect 12173 14433 12207 14467
rect 13921 14433 13955 14467
rect 21649 14433 21683 14467
rect 26065 14433 26099 14467
rect 42165 14433 42199 14467
rect 42809 14433 42843 14467
rect 42901 14433 42935 14467
rect 43637 14433 43671 14467
rect 43729 14433 43763 14467
rect 45201 14433 45235 14467
rect 48789 14433 48823 14467
rect 49065 14433 49099 14467
rect 52653 14433 52687 14467
rect 53481 14433 53515 14467
rect 3433 14365 3467 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 4077 14365 4111 14399
rect 4169 14365 4203 14399
rect 4353 14365 4387 14399
rect 6837 14365 6871 14399
rect 7113 14365 7147 14399
rect 8493 14365 8527 14399
rect 15761 14365 15795 14399
rect 16589 14365 16623 14399
rect 17509 14365 17543 14399
rect 17969 14365 18003 14399
rect 22385 14365 22419 14399
rect 24961 14365 24995 14399
rect 25329 14365 25363 14399
rect 29745 14365 29779 14399
rect 32781 14365 32815 14399
rect 36093 14365 36127 14399
rect 37105 14365 37139 14399
rect 38577 14365 38611 14399
rect 46673 14365 46707 14399
rect 49249 14365 49283 14399
rect 49341 14365 49375 14399
rect 50629 14365 50663 14399
rect 54861 14365 54895 14399
rect 58449 14365 58483 14399
rect 3617 14297 3651 14331
rect 7665 14297 7699 14331
rect 9956 14297 9990 14331
rect 12440 14297 12474 14331
rect 20729 14297 20763 14331
rect 26310 14297 26344 14331
rect 30297 14297 30331 14331
rect 33701 14297 33735 14331
rect 36001 14297 36035 14331
rect 41705 14297 41739 14331
rect 44557 14297 44591 14331
rect 50896 14297 50930 14331
rect 52469 14297 52503 14331
rect 52929 14297 52963 14331
rect 7297 14229 7331 14263
rect 9137 14229 9171 14263
rect 11805 14229 11839 14263
rect 15117 14229 15151 14263
rect 15945 14229 15979 14263
rect 16957 14229 16991 14263
rect 18613 14229 18647 14263
rect 21833 14229 21867 14263
rect 24041 14229 24075 14263
rect 24409 14229 24443 14263
rect 25881 14229 25915 14263
rect 27445 14229 27479 14263
rect 29377 14229 29411 14263
rect 36737 14229 36771 14263
rect 37933 14229 37967 14263
rect 42349 14229 42383 14263
rect 42717 14229 42751 14263
rect 43821 14229 43855 14263
rect 44189 14229 44223 14263
rect 46121 14229 46155 14263
rect 50537 14229 50571 14263
rect 52101 14229 52135 14263
rect 52561 14229 52595 14263
rect 54309 14229 54343 14263
rect 57161 14229 57195 14263
rect 57897 14229 57931 14263
rect 3341 14025 3375 14059
rect 3801 14025 3835 14059
rect 6837 14025 6871 14059
rect 8677 14025 8711 14059
rect 9045 14025 9079 14059
rect 10241 14025 10275 14059
rect 10609 14025 10643 14059
rect 10701 14025 10735 14059
rect 11253 14025 11287 14059
rect 12265 14025 12299 14059
rect 12449 14025 12483 14059
rect 12909 14025 12943 14059
rect 13277 14025 13311 14059
rect 15577 14025 15611 14059
rect 16037 14025 16071 14059
rect 16405 14025 16439 14059
rect 18061 14025 18095 14059
rect 18521 14025 18555 14059
rect 18889 14025 18923 14059
rect 22569 14025 22603 14059
rect 25513 14025 25547 14059
rect 26157 14025 26191 14059
rect 27261 14025 27295 14059
rect 28825 14025 28859 14059
rect 29285 14025 29319 14059
rect 35817 14025 35851 14059
rect 37289 14025 37323 14059
rect 38853 14025 38887 14059
rect 40785 14025 40819 14059
rect 42257 14025 42291 14059
rect 45017 14025 45051 14059
rect 46029 14025 46063 14059
rect 46305 14025 46339 14059
rect 46765 14025 46799 14059
rect 49985 14025 50019 14059
rect 51549 14025 51583 14059
rect 54493 14025 54527 14059
rect 57253 14025 57287 14059
rect 57345 14025 57379 14059
rect 57713 14025 57747 14059
rect 5273 13957 5307 13991
rect 7950 13957 7984 13991
rect 9505 13957 9539 13991
rect 15209 13957 15243 13991
rect 16937 13957 16971 13991
rect 30481 13957 30515 13991
rect 33241 13957 33275 13991
rect 37657 13957 37691 13991
rect 42441 13957 42475 13991
rect 3249 13889 3283 13923
rect 3617 13889 3651 13923
rect 3801 13889 3835 13923
rect 5181 13889 5215 13923
rect 5365 13889 5399 13923
rect 8217 13889 8251 13923
rect 9413 13889 9447 13923
rect 10149 13889 10183 13923
rect 12817 13889 12851 13923
rect 13829 13889 13863 13923
rect 15669 13889 15703 13923
rect 18429 13889 18463 13923
rect 19533 13889 19567 13923
rect 22109 13889 22143 13923
rect 22201 13889 22235 13923
rect 23213 13889 23247 13923
rect 24400 13889 24434 13923
rect 27445 13889 27479 13923
rect 28181 13889 28215 13923
rect 29193 13889 29227 13923
rect 29653 13889 29687 13923
rect 31125 13889 31159 13923
rect 32413 13889 32447 13923
rect 34437 13889 34471 13923
rect 34704 13889 34738 13923
rect 35909 13889 35943 13923
rect 38485 13889 38519 13923
rect 39497 13889 39531 13923
rect 44097 13889 44131 13923
rect 44833 13889 44867 13923
rect 46673 13889 46707 13923
rect 48237 13889 48271 13923
rect 48605 13889 48639 13923
rect 48872 13889 48906 13923
rect 52101 13889 52135 13923
rect 54861 13889 54895 13923
rect 54953 13889 54987 13923
rect 55965 13889 55999 13923
rect 58449 13889 58483 13923
rect 10793 13821 10827 13855
rect 13093 13821 13127 13855
rect 14749 13821 14783 13855
rect 15393 13821 15427 13855
rect 16681 13821 16715 13855
rect 18245 13821 18279 13855
rect 20177 13821 20211 13855
rect 20729 13821 20763 13855
rect 21005 13821 21039 13855
rect 22017 13821 22051 13855
rect 23489 13821 23523 13855
rect 24133 13821 24167 13855
rect 25881 13821 25915 13855
rect 26801 13821 26835 13855
rect 27997 13821 28031 13855
rect 29469 13821 29503 13855
rect 31677 13821 31711 13855
rect 33517 13821 33551 13855
rect 34161 13821 34195 13855
rect 36461 13821 36495 13855
rect 37749 13821 37783 13855
rect 37841 13821 37875 13855
rect 38209 13821 38243 13855
rect 38393 13821 38427 13855
rect 41061 13821 41095 13855
rect 41613 13821 41647 13855
rect 45569 13821 45603 13855
rect 46857 13821 46891 13855
rect 47409 13821 47443 13855
rect 47593 13821 47627 13855
rect 50077 13821 50111 13855
rect 52745 13821 52779 13855
rect 53297 13821 53331 13855
rect 53481 13821 53515 13855
rect 55045 13821 55079 13855
rect 55321 13821 55355 13855
rect 56609 13821 56643 13855
rect 57069 13821 57103 13855
rect 22661 13753 22695 13787
rect 36829 13753 36863 13787
rect 52469 13753 52503 13787
rect 11713 13685 11747 13719
rect 18981 13685 19015 13719
rect 20085 13685 20119 13719
rect 21649 13685 21683 13719
rect 24041 13685 24075 13719
rect 28733 13685 28767 13719
rect 38945 13685 38979 13719
rect 44281 13685 44315 13719
rect 50721 13685 50755 13719
rect 54125 13685 54159 13719
rect 56057 13685 56091 13719
rect 57897 13685 57931 13719
rect 2881 13481 2915 13515
rect 3433 13481 3467 13515
rect 4077 13481 4111 13515
rect 4629 13481 4663 13515
rect 6561 13481 6595 13515
rect 7021 13481 7055 13515
rect 7389 13481 7423 13515
rect 11529 13481 11563 13515
rect 12173 13481 12207 13515
rect 13369 13481 13403 13515
rect 18337 13481 18371 13515
rect 20269 13481 20303 13515
rect 21373 13481 21407 13515
rect 23305 13481 23339 13515
rect 23489 13481 23523 13515
rect 24409 13481 24443 13515
rect 27169 13481 27203 13515
rect 29377 13481 29411 13515
rect 34345 13481 34379 13515
rect 35817 13481 35851 13515
rect 41153 13481 41187 13515
rect 44649 13481 44683 13515
rect 47041 13481 47075 13515
rect 53573 13481 53607 13515
rect 55137 13481 55171 13515
rect 58265 13481 58299 13515
rect 5917 13413 5951 13447
rect 9781 13413 9815 13447
rect 16037 13413 16071 13447
rect 17601 13413 17635 13447
rect 20361 13413 20395 13447
rect 26433 13413 26467 13447
rect 37013 13413 37047 13447
rect 47409 13413 47443 13447
rect 48789 13413 48823 13447
rect 49709 13413 49743 13447
rect 52561 13413 52595 13447
rect 2605 13345 2639 13379
rect 5825 13345 5859 13379
rect 9689 13345 9723 13379
rect 10241 13345 10275 13379
rect 10425 13345 10459 13379
rect 12633 13345 12667 13379
rect 14657 13345 14691 13379
rect 17325 13345 17359 13379
rect 18061 13345 18095 13379
rect 18889 13345 18923 13379
rect 19809 13345 19843 13379
rect 20821 13345 20855 13379
rect 21005 13345 21039 13379
rect 22753 13345 22787 13379
rect 24041 13345 24075 13379
rect 24869 13345 24903 13379
rect 24961 13345 24995 13379
rect 26019 13345 26053 13379
rect 26157 13345 26191 13379
rect 27721 13345 27755 13379
rect 32597 13345 32631 13379
rect 33425 13345 33459 13379
rect 35265 13345 35299 13379
rect 35449 13345 35483 13379
rect 36461 13345 36495 13379
rect 36737 13345 36771 13379
rect 37473 13345 37507 13379
rect 42349 13345 42383 13379
rect 48237 13345 48271 13379
rect 48375 13345 48409 13379
rect 49249 13345 49283 13379
rect 50353 13345 50387 13379
rect 50445 13345 50479 13379
rect 53113 13345 53147 13379
rect 53757 13345 53791 13379
rect 2513 13277 2547 13311
rect 3249 13277 3283 13311
rect 3525 13277 3559 13311
rect 3801 13277 3835 13311
rect 4721 13277 4755 13311
rect 6192 13277 6226 13311
rect 6285 13277 6319 13311
rect 6652 13277 6686 13311
rect 6745 13277 6779 13311
rect 10149 13277 10183 13311
rect 10609 13277 10643 13311
rect 14924 13277 14958 13311
rect 17049 13277 17083 13311
rect 17187 13277 17221 13311
rect 18245 13277 18279 13311
rect 19257 13277 19291 13311
rect 22486 13277 22520 13311
rect 23857 13277 23891 13311
rect 25881 13277 25915 13311
rect 26893 13277 26927 13311
rect 27077 13277 27111 13311
rect 27997 13277 28031 13311
rect 28549 13277 28583 13311
rect 31861 13277 31895 13311
rect 32137 13277 32171 13311
rect 33241 13277 33275 13311
rect 36620 13277 36654 13311
rect 37657 13277 37691 13311
rect 39129 13277 39163 13311
rect 39405 13277 39439 13311
rect 43085 13277 43119 13311
rect 43269 13277 43303 13311
rect 45293 13277 45327 13311
rect 45661 13277 45695 13311
rect 45928 13277 45962 13311
rect 48513 13277 48547 13311
rect 49433 13277 49467 13311
rect 51549 13277 51583 13311
rect 52469 13277 52503 13311
rect 55321 13277 55355 13311
rect 56885 13277 56919 13311
rect 57152 13277 57186 13311
rect 3893 13209 3927 13243
rect 4077 13209 4111 13243
rect 8769 13209 8803 13243
rect 12081 13209 12115 13243
rect 13001 13209 13035 13243
rect 18797 13209 18831 13243
rect 27537 13209 27571 13243
rect 29561 13209 29595 13243
rect 38862 13209 38896 13243
rect 39865 13209 39899 13243
rect 42073 13209 42107 13243
rect 43536 13209 43570 13243
rect 50537 13209 50571 13243
rect 52929 13209 52963 13243
rect 54024 13209 54058 13243
rect 55588 13209 55622 13243
rect 9045 13141 9079 13175
rect 11253 13141 11287 13175
rect 16405 13141 16439 13175
rect 18705 13141 18739 13175
rect 20729 13141 20763 13175
rect 23949 13141 23983 13175
rect 24777 13141 24811 13175
rect 25237 13141 25271 13175
rect 27629 13141 27663 13175
rect 30849 13141 30883 13175
rect 34805 13141 34839 13175
rect 35173 13141 35207 13175
rect 37749 13141 37783 13175
rect 41705 13141 41739 13175
rect 42165 13141 42199 13175
rect 42533 13141 42567 13175
rect 47593 13141 47627 13175
rect 50905 13141 50939 13175
rect 50997 13141 51031 13175
rect 51825 13141 51859 13175
rect 53021 13141 53055 13175
rect 56701 13141 56735 13175
rect 3525 12937 3559 12971
rect 7297 12937 7331 12971
rect 7481 12937 7515 12971
rect 16313 12937 16347 12971
rect 16865 12937 16899 12971
rect 17325 12937 17359 12971
rect 21097 12937 21131 12971
rect 22569 12937 22603 12971
rect 23673 12937 23707 12971
rect 26801 12937 26835 12971
rect 29929 12937 29963 12971
rect 33517 12937 33551 12971
rect 35817 12937 35851 12971
rect 36277 12937 36311 12971
rect 36921 12937 36955 12971
rect 38669 12937 38703 12971
rect 38761 12937 38795 12971
rect 39681 12937 39715 12971
rect 41245 12937 41279 12971
rect 42717 12937 42751 12971
rect 45569 12937 45603 12971
rect 49617 12937 49651 12971
rect 52745 12937 52779 12971
rect 53113 12937 53147 12971
rect 55965 12937 55999 12971
rect 6754 12869 6788 12903
rect 7113 12869 7147 12903
rect 11069 12869 11103 12903
rect 18460 12869 18494 12903
rect 28816 12869 28850 12903
rect 36185 12869 36219 12903
rect 40132 12869 40166 12903
rect 41337 12869 41371 12903
rect 47777 12869 47811 12903
rect 50169 12869 50203 12903
rect 51448 12869 51482 12903
rect 6377 12801 6411 12835
rect 7021 12801 7055 12835
rect 9790 12801 9824 12835
rect 10425 12801 10459 12835
rect 11529 12801 11563 12835
rect 12909 12801 12943 12835
rect 14740 12801 14774 12835
rect 18705 12801 18739 12835
rect 19717 12801 19751 12835
rect 19984 12801 20018 12835
rect 22477 12801 22511 12835
rect 23765 12801 23799 12835
rect 24032 12801 24066 12835
rect 25421 12801 25455 12835
rect 25688 12801 25722 12835
rect 27353 12801 27387 12835
rect 27445 12801 27479 12835
rect 28457 12801 28491 12835
rect 28549 12801 28583 12835
rect 30481 12801 30515 12835
rect 30573 12801 30607 12835
rect 30840 12801 30874 12835
rect 32137 12801 32171 12835
rect 32404 12801 32438 12835
rect 34345 12801 34379 12835
rect 34612 12801 34646 12835
rect 37556 12801 37590 12835
rect 39865 12801 39899 12835
rect 43085 12801 43119 12835
rect 43352 12801 43386 12835
rect 44557 12801 44591 12835
rect 46020 12801 46054 12835
rect 48237 12801 48271 12835
rect 48504 12801 48538 12835
rect 50077 12801 50111 12835
rect 53205 12801 53239 12835
rect 54815 12801 54849 12835
rect 55689 12801 55723 12835
rect 56333 12801 56367 12835
rect 57345 12801 57379 12835
rect 3065 12733 3099 12767
rect 3801 12733 3835 12767
rect 8033 12733 8067 12767
rect 10057 12733 10091 12767
rect 12357 12733 12391 12767
rect 13553 12733 13587 12767
rect 14473 12733 14507 12767
rect 18981 12733 19015 12767
rect 22661 12733 22695 12767
rect 27537 12733 27571 12767
rect 34161 12733 34195 12767
rect 36461 12733 36495 12767
rect 37289 12733 37323 12767
rect 39313 12733 39347 12767
rect 41889 12733 41923 12767
rect 45109 12733 45143 12767
rect 45753 12733 45787 12767
rect 50353 12733 50387 12767
rect 51181 12733 51215 12767
rect 53297 12733 53331 12767
rect 53757 12733 53791 12767
rect 54677 12733 54711 12767
rect 54953 12733 54987 12767
rect 55873 12733 55907 12767
rect 56425 12733 56459 12767
rect 56517 12733 56551 12767
rect 56793 12733 56827 12767
rect 3433 12665 3467 12699
rect 8677 12665 8711 12699
rect 21649 12665 21683 12699
rect 47133 12665 47167 12699
rect 55229 12665 55263 12699
rect 6745 12597 6779 12631
rect 7297 12597 7331 12631
rect 8585 12597 8619 12631
rect 15853 12597 15887 12631
rect 22109 12597 22143 12631
rect 23305 12597 23339 12631
rect 25145 12597 25179 12631
rect 26985 12597 27019 12631
rect 31953 12597 31987 12631
rect 33609 12597 33643 12631
rect 35725 12597 35759 12631
rect 44465 12597 44499 12631
rect 49709 12597 49743 12631
rect 50813 12597 50847 12631
rect 52561 12597 52595 12631
rect 54033 12597 54067 12631
rect 8769 12393 8803 12427
rect 10425 12393 10459 12427
rect 16957 12393 16991 12427
rect 22753 12393 22787 12427
rect 24501 12393 24535 12427
rect 26341 12393 26375 12427
rect 27353 12393 27387 12427
rect 44097 12393 44131 12427
rect 47041 12393 47075 12427
rect 48053 12393 48087 12427
rect 49617 12393 49651 12427
rect 53941 12393 53975 12427
rect 55505 12393 55539 12427
rect 3801 12325 3835 12359
rect 5089 12325 5123 12359
rect 16681 12325 16715 12359
rect 28641 12325 28675 12359
rect 34713 12325 34747 12359
rect 36185 12325 36219 12359
rect 37933 12325 37967 12359
rect 41337 12325 41371 12359
rect 41429 12325 41463 12359
rect 42625 12325 42659 12359
rect 53205 12325 53239 12359
rect 2605 12257 2639 12291
rect 5549 12257 5583 12291
rect 7573 12257 7607 12291
rect 11345 12257 11379 12291
rect 11621 12257 11655 12291
rect 11897 12257 11931 12291
rect 12541 12257 12575 12291
rect 13093 12257 13127 12291
rect 13185 12257 13219 12291
rect 14565 12257 14599 12291
rect 14657 12257 14691 12291
rect 15807 12257 15841 12291
rect 16129 12257 16163 12291
rect 17509 12257 17543 12291
rect 19441 12257 19475 12291
rect 20913 12257 20947 12291
rect 21557 12257 21591 12291
rect 21833 12257 21867 12291
rect 25145 12257 25179 12291
rect 26985 12257 27019 12291
rect 27997 12257 28031 12291
rect 29285 12257 29319 12291
rect 31447 12257 31481 12291
rect 31585 12257 31619 12291
rect 31861 12257 31895 12291
rect 32781 12257 32815 12291
rect 32873 12257 32907 12291
rect 34069 12257 34103 12291
rect 35265 12257 35299 12291
rect 35633 12257 35667 12291
rect 37105 12257 37139 12291
rect 37381 12257 37415 12291
rect 38669 12257 38703 12291
rect 42211 12257 42245 12291
rect 42349 12257 42383 12291
rect 43453 12257 43487 12291
rect 44741 12257 44775 12291
rect 46397 12257 46431 12291
rect 47685 12257 47719 12291
rect 48605 12257 48639 12291
rect 53297 12257 53331 12291
rect 3341 12189 3375 12223
rect 3525 12189 3559 12223
rect 4076 12189 4110 12223
rect 4169 12189 4203 12223
rect 5825 12189 5859 12223
rect 6285 12189 6319 12223
rect 6653 12189 6687 12223
rect 6929 12189 6963 12223
rect 8217 12189 8251 12223
rect 9045 12189 9079 12223
rect 11483 12189 11517 12223
rect 12357 12189 12391 12223
rect 14473 12189 14507 12223
rect 15577 12189 15611 12223
rect 17417 12189 17451 12223
rect 21097 12189 21131 12223
rect 21950 12189 21984 12223
rect 22109 12189 22143 12223
rect 27813 12189 27847 12223
rect 29745 12189 29779 12223
rect 30389 12189 30423 12223
rect 31309 12189 31343 12223
rect 32321 12189 32355 12223
rect 32505 12189 32539 12223
rect 32965 12189 32999 12223
rect 33885 12189 33919 12223
rect 37473 12189 37507 12223
rect 38025 12189 38059 12223
rect 39957 12189 39991 12223
rect 42073 12189 42107 12223
rect 43085 12189 43119 12223
rect 43269 12189 43303 12223
rect 48237 12189 48271 12223
rect 51825 12189 51859 12223
rect 52092 12189 52126 12223
rect 56057 12189 56091 12223
rect 56701 12189 56735 12223
rect 5089 12121 5123 12155
rect 9290 12121 9324 12155
rect 10701 12121 10735 12155
rect 13001 12121 13035 12155
rect 19708 12121 19742 12155
rect 33793 12121 33827 12155
rect 37565 12121 37599 12155
rect 40224 12121 40258 12155
rect 43729 12121 43763 12155
rect 44189 12121 44223 12155
rect 46581 12121 46615 12155
rect 47133 12121 47167 12155
rect 56609 12121 56643 12155
rect 56946 12121 56980 12155
rect 4445 12053 4479 12087
rect 5641 12053 5675 12087
rect 12633 12053 12667 12087
rect 13829 12053 13863 12087
rect 14105 12053 14139 12087
rect 15209 12053 15243 12087
rect 15669 12053 15703 12087
rect 17325 12053 17359 12087
rect 20821 12053 20855 12087
rect 28549 12053 28583 12087
rect 29009 12053 29043 12087
rect 29101 12053 29135 12087
rect 30665 12053 30699 12087
rect 33333 12053 33367 12087
rect 33425 12053 33459 12087
rect 34529 12053 34563 12087
rect 36461 12053 36495 12087
rect 38945 12053 38979 12087
rect 39681 12053 39715 12087
rect 43637 12053 43671 12087
rect 46121 12053 46155 12087
rect 46673 12053 46707 12087
rect 49893 12053 49927 12087
rect 50997 12053 51031 12087
rect 51641 12053 51675 12087
rect 54309 12053 54343 12087
rect 54677 12053 54711 12087
rect 58081 12053 58115 12087
rect 2973 11849 3007 11883
rect 3801 11849 3835 11883
rect 5733 11849 5767 11883
rect 8861 11849 8895 11883
rect 9229 11849 9263 11883
rect 11805 11849 11839 11883
rect 15025 11849 15059 11883
rect 20453 11849 20487 11883
rect 21557 11849 21591 11883
rect 32505 11849 32539 11883
rect 35909 11849 35943 11883
rect 41981 11849 42015 11883
rect 46213 11849 46247 11883
rect 49525 11849 49559 11883
rect 50905 11849 50939 11883
rect 52929 11849 52963 11883
rect 56609 11849 56643 11883
rect 56793 11849 56827 11883
rect 6561 11781 6595 11815
rect 7113 11781 7147 11815
rect 9321 11781 9355 11815
rect 28794 11781 28828 11815
rect 32597 11781 32631 11815
rect 40969 11781 41003 11815
rect 42625 11781 42659 11815
rect 55781 11781 55815 11815
rect 3248 11713 3282 11747
rect 3341 11713 3375 11747
rect 5641 11713 5675 11747
rect 6655 11735 6689 11769
rect 7021 11713 7055 11747
rect 9956 11713 9990 11747
rect 11989 11713 12023 11747
rect 12256 11713 12290 11747
rect 13645 11713 13679 11747
rect 14197 11713 14231 11747
rect 15577 11713 15611 11747
rect 20913 11713 20947 11747
rect 30665 11713 30699 11747
rect 32965 11713 32999 11747
rect 33517 11713 33551 11747
rect 34253 11713 34287 11747
rect 35081 11713 35115 11747
rect 40509 11713 40543 11747
rect 41613 11713 41647 11747
rect 46857 11713 46891 11747
rect 49433 11713 49467 11747
rect 52837 11713 52871 11747
rect 57161 11713 57195 11747
rect 57253 11713 57287 11747
rect 57897 11713 57931 11747
rect 9505 11645 9539 11679
rect 9689 11645 9723 11679
rect 19533 11645 19567 11679
rect 20545 11645 20579 11679
rect 20637 11645 20671 11679
rect 23581 11645 23615 11679
rect 25421 11645 25455 11679
rect 28549 11645 28583 11679
rect 30021 11645 30055 11679
rect 32689 11645 32723 11679
rect 33701 11645 33735 11679
rect 40233 11645 40267 11679
rect 40417 11645 40451 11679
rect 43269 11645 43303 11679
rect 51457 11645 51491 11679
rect 56241 11645 56275 11679
rect 57437 11645 57471 11679
rect 58449 11645 58483 11679
rect 25237 11577 25271 11611
rect 29929 11577 29963 11611
rect 34713 11577 34747 11611
rect 38945 11577 38979 11611
rect 40877 11577 40911 11611
rect 50537 11577 50571 11611
rect 4169 11509 4203 11543
rect 11069 11509 11103 11543
rect 13369 11509 13403 11543
rect 14841 11509 14875 11543
rect 16865 11509 16899 11543
rect 19901 11509 19935 11543
rect 20085 11509 20119 11543
rect 23029 11509 23063 11543
rect 25973 11509 26007 11543
rect 28365 11509 28399 11543
rect 31953 11509 31987 11543
rect 32137 11509 32171 11543
rect 35357 11509 35391 11543
rect 40049 11509 40083 11543
rect 45661 11509 45695 11543
rect 3985 11305 4019 11339
rect 5089 11305 5123 11339
rect 9873 11305 9907 11339
rect 13921 11305 13955 11339
rect 15301 11305 15335 11339
rect 19901 11305 19935 11339
rect 23305 11305 23339 11339
rect 25421 11305 25455 11339
rect 29837 11305 29871 11339
rect 32597 11305 32631 11339
rect 32781 11305 32815 11339
rect 40325 11305 40359 11339
rect 42257 11305 42291 11339
rect 42625 11305 42659 11339
rect 57621 11305 57655 11339
rect 57989 11305 58023 11339
rect 4169 11237 4203 11271
rect 6561 11237 6595 11271
rect 6653 11237 6687 11271
rect 47501 11237 47535 11271
rect 6745 11169 6779 11203
rect 7205 11169 7239 11203
rect 10333 11169 10367 11203
rect 11713 11169 11747 11203
rect 13369 11169 13403 11203
rect 20453 11169 20487 11203
rect 26065 11169 26099 11203
rect 36185 11169 36219 11203
rect 50905 11169 50939 11203
rect 56517 11169 56551 11203
rect 56793 11169 56827 11203
rect 4261 11101 4295 11135
rect 4445 11101 4479 11135
rect 5365 11101 5399 11135
rect 6101 11101 6135 11135
rect 6193 11101 6227 11135
rect 10149 11101 10183 11135
rect 11529 11101 11563 11135
rect 12633 11101 12667 11135
rect 14381 11101 14415 11135
rect 15393 11101 15427 11135
rect 17417 11101 17451 11135
rect 21741 11101 21775 11135
rect 22569 11101 22603 11135
rect 24409 11101 24443 11135
rect 25789 11101 25823 11135
rect 25881 11101 25915 11135
rect 26249 11101 26283 11135
rect 26801 11101 26835 11135
rect 29101 11101 29135 11135
rect 33609 11101 33643 11135
rect 34345 11101 34379 11135
rect 35357 11101 35391 11135
rect 37013 11101 37047 11135
rect 37749 11101 37783 11135
rect 38761 11101 38795 11135
rect 39589 11101 39623 11135
rect 40601 11101 40635 11135
rect 41889 11101 41923 11135
rect 43821 11101 43855 11135
rect 44465 11101 44499 11135
rect 45569 11101 45603 11135
rect 45845 11101 45879 11135
rect 47041 11101 47075 11135
rect 50721 11101 50755 11135
rect 52193 11101 52227 11135
rect 56977 11101 57011 11135
rect 3801 11033 3835 11067
rect 4353 11033 4387 11067
rect 5089 11033 5123 11067
rect 5273 11033 5307 11067
rect 7113 11033 7147 11067
rect 9505 11033 9539 11067
rect 11437 11033 11471 11067
rect 12173 11033 12207 11067
rect 13185 11033 13219 11067
rect 20821 11033 20855 11067
rect 23213 11033 23247 11067
rect 24041 11033 24075 11067
rect 28549 11033 28583 11067
rect 32873 11033 32907 11067
rect 40417 11033 40451 11067
rect 42533 11033 42567 11067
rect 46397 11033 46431 11067
rect 49893 11033 49927 11067
rect 51641 11033 51675 11067
rect 55505 11033 55539 11067
rect 4011 10965 4045 10999
rect 5457 10965 5491 10999
rect 7849 10965 7883 10999
rect 11069 10965 11103 10999
rect 14933 10965 14967 10999
rect 16865 10965 16899 10999
rect 22017 10965 22051 10999
rect 25053 10965 25087 10999
rect 33057 10965 33091 10999
rect 33793 10965 33827 10999
rect 34897 10965 34931 10999
rect 36461 10965 36495 10999
rect 37197 10965 37231 10999
rect 38209 10965 38243 10999
rect 38945 10965 38979 10999
rect 41245 10965 41279 10999
rect 41337 10965 41371 10999
rect 43177 10965 43211 10999
rect 43913 10965 43947 10999
rect 45017 10965 45051 10999
rect 46489 10965 46523 10999
rect 50169 10965 50203 10999
rect 51549 10965 51583 10999
rect 55965 10965 55999 10999
rect 56885 10965 56919 10999
rect 57345 10965 57379 10999
rect 5365 10761 5399 10795
rect 6469 10761 6503 10795
rect 9873 10761 9907 10795
rect 10517 10761 10551 10795
rect 13645 10761 13679 10795
rect 14105 10761 14139 10795
rect 16865 10761 16899 10795
rect 18521 10761 18555 10795
rect 39221 10761 39255 10795
rect 41245 10761 41279 10795
rect 42257 10761 42291 10795
rect 43821 10761 43855 10795
rect 45477 10761 45511 10795
rect 50629 10761 50663 10795
rect 50721 10761 50755 10795
rect 51181 10761 51215 10795
rect 51549 10761 51583 10795
rect 55689 10761 55723 10795
rect 2605 10693 2639 10727
rect 7604 10693 7638 10727
rect 19993 10693 20027 10727
rect 33057 10693 33091 10727
rect 34345 10693 34379 10727
rect 35072 10693 35106 10727
rect 36553 10693 36587 10727
rect 37740 10693 37774 10727
rect 45753 10693 45787 10727
rect 46296 10693 46330 10727
rect 49065 10693 49099 10727
rect 51089 10693 51123 10727
rect 3801 10625 3835 10659
rect 5457 10625 5491 10659
rect 7849 10625 7883 10659
rect 11069 10625 11103 10659
rect 12725 10625 12759 10659
rect 13185 10625 13219 10659
rect 13277 10625 13311 10659
rect 14013 10625 14047 10659
rect 15853 10625 15887 10659
rect 16773 10625 16807 10659
rect 21097 10625 21131 10659
rect 21649 10625 21683 10659
rect 22201 10625 22235 10659
rect 23581 10625 23615 10659
rect 23673 10625 23707 10659
rect 24685 10625 24719 10659
rect 26074 10625 26108 10659
rect 29101 10625 29135 10659
rect 30205 10625 30239 10659
rect 30849 10625 30883 10659
rect 33517 10625 33551 10659
rect 34805 10625 34839 10659
rect 36369 10625 36403 10659
rect 39313 10625 39347 10659
rect 39773 10625 39807 10659
rect 40040 10625 40074 10659
rect 42441 10625 42475 10659
rect 42708 10625 42742 10659
rect 44097 10625 44131 10659
rect 44364 10625 44398 10659
rect 46029 10625 46063 10659
rect 49516 10625 49550 10659
rect 51917 10625 51951 10659
rect 52009 10625 52043 10659
rect 52745 10625 52779 10659
rect 57529 10625 57563 10659
rect 3709 10557 3743 10591
rect 4813 10557 4847 10591
rect 5825 10557 5859 10591
rect 10425 10557 10459 10591
rect 12173 10557 12207 10591
rect 13461 10557 13495 10591
rect 14197 10557 14231 10591
rect 15393 10557 15427 10591
rect 15945 10557 15979 10591
rect 16037 10557 16071 10591
rect 20729 10557 20763 10591
rect 21925 10557 21959 10591
rect 22109 10557 22143 10591
rect 23765 10557 23799 10591
rect 24041 10557 24075 10591
rect 26341 10557 26375 10591
rect 29193 10557 29227 10591
rect 29285 10557 29319 10591
rect 29561 10557 29595 10591
rect 32597 10557 32631 10591
rect 32781 10557 32815 10591
rect 32965 10557 32999 10591
rect 37473 10557 37507 10591
rect 39129 10557 39163 10591
rect 41797 10557 41831 10591
rect 47593 10557 47627 10591
rect 49249 10557 49283 10591
rect 51365 10557 51399 10591
rect 52193 10557 52227 10591
rect 53297 10557 53331 10591
rect 54125 10557 54159 10591
rect 54769 10557 54803 10591
rect 55505 10557 55539 10591
rect 56333 10557 56367 10591
rect 56471 10557 56505 10591
rect 56609 10557 56643 10591
rect 56885 10557 56919 10591
rect 57345 10557 57379 10591
rect 58449 10557 58483 10591
rect 2973 10489 3007 10523
rect 5733 10489 5767 10523
rect 12817 10489 12851 10523
rect 15485 10489 15519 10523
rect 23121 10489 23155 10523
rect 28641 10489 28675 10523
rect 33425 10489 33459 10523
rect 36185 10489 36219 10523
rect 41153 10489 41187 10523
rect 47409 10489 47443 10523
rect 2421 10421 2455 10455
rect 2605 10421 2639 10455
rect 3065 10421 3099 10455
rect 4445 10421 4479 10455
rect 5595 10421 5629 10455
rect 6101 10421 6135 10455
rect 11897 10421 11931 10455
rect 14749 10421 14783 10455
rect 20085 10421 20119 10455
rect 22569 10421 22603 10455
rect 23213 10421 23247 10455
rect 24961 10421 24995 10455
rect 26709 10421 26743 10455
rect 28733 10421 28767 10455
rect 30757 10421 30791 10455
rect 31861 10421 31895 10455
rect 38853 10421 38887 10455
rect 39681 10421 39715 10455
rect 48237 10421 48271 10455
rect 48513 10421 48547 10455
rect 53481 10421 53515 10455
rect 54217 10421 54251 10455
rect 54953 10421 54987 10455
rect 57897 10421 57931 10455
rect 3525 10217 3559 10251
rect 4721 10217 4755 10251
rect 4905 10217 4939 10251
rect 5825 10217 5859 10251
rect 9229 10217 9263 10251
rect 11989 10217 12023 10251
rect 12541 10217 12575 10251
rect 16497 10217 16531 10251
rect 20545 10217 20579 10251
rect 20913 10217 20947 10251
rect 23857 10217 23891 10251
rect 24133 10217 24167 10251
rect 32045 10217 32079 10251
rect 38577 10217 38611 10251
rect 39865 10217 39899 10251
rect 42809 10217 42843 10251
rect 50813 10217 50847 10251
rect 54125 10217 54159 10251
rect 54953 10217 54987 10251
rect 6469 10149 6503 10183
rect 6653 10149 6687 10183
rect 12357 10149 12391 10183
rect 19073 10149 19107 10183
rect 33517 10149 33551 10183
rect 44833 10149 44867 10183
rect 47133 10149 47167 10183
rect 52009 10149 52043 10183
rect 1961 10081 1995 10115
rect 2237 10081 2271 10115
rect 5273 10081 5307 10115
rect 6009 10081 6043 10115
rect 6561 10081 6595 10115
rect 11345 10081 11379 10115
rect 13921 10081 13955 10115
rect 15485 10081 15519 10115
rect 15761 10081 15795 10115
rect 16405 10081 16439 10115
rect 24501 10081 24535 10115
rect 25145 10081 25179 10115
rect 25421 10081 25455 10115
rect 25697 10081 25731 10115
rect 26985 10081 27019 10115
rect 27445 10081 27479 10115
rect 31125 10081 31159 10115
rect 32137 10081 32171 10115
rect 34253 10081 34287 10115
rect 35495 10081 35529 10115
rect 35909 10081 35943 10115
rect 36369 10081 36403 10115
rect 37105 10081 37139 10115
rect 39037 10081 39071 10115
rect 39221 10081 39255 10115
rect 41337 10081 41371 10115
rect 41889 10081 41923 10115
rect 42165 10081 42199 10115
rect 42349 10081 42383 10115
rect 45569 10081 45603 10115
rect 46583 10081 46617 10115
rect 46740 10081 46774 10115
rect 47777 10081 47811 10115
rect 51733 10081 51767 10115
rect 52653 10081 52687 10115
rect 54309 10081 54343 10115
rect 56793 10081 56827 10115
rect 4077 10013 4111 10047
rect 5641 10013 5675 10047
rect 6101 10013 6135 10047
rect 10885 10013 10919 10047
rect 14381 10013 14415 10047
rect 15209 10013 15243 10047
rect 15368 10013 15402 10047
rect 16221 10013 16255 10047
rect 17049 10013 17083 10047
rect 17693 10013 17727 10047
rect 20085 10013 20119 10047
rect 22026 10013 22060 10047
rect 22293 10013 22327 10047
rect 22477 10013 22511 10047
rect 24685 10013 24719 10047
rect 25538 10013 25572 10047
rect 26801 10013 26835 10047
rect 27997 10013 28031 10047
rect 32404 10013 32438 10047
rect 33977 10013 34011 10047
rect 35357 10013 35391 10047
rect 35633 10013 35667 10047
rect 36553 10013 36587 10047
rect 36921 10013 36955 10047
rect 40989 10013 41023 10047
rect 41245 10013 41279 10047
rect 42441 10013 42475 10047
rect 43453 10013 43487 10047
rect 46857 10013 46891 10047
rect 47593 10013 47627 10047
rect 49249 10013 49283 10047
rect 49985 10013 50019 10047
rect 51457 10013 51491 10047
rect 51616 10013 51650 10047
rect 52469 10013 52503 10047
rect 52745 10013 52779 10047
rect 53012 10013 53046 10047
rect 55321 10013 55355 10047
rect 58449 10013 58483 10047
rect 4629 9945 4663 9979
rect 4905 9945 4939 9979
rect 5457 9945 5491 9979
rect 13654 9945 13688 9979
rect 17960 9945 17994 9979
rect 22744 9945 22778 9979
rect 26341 9945 26375 9979
rect 26893 9945 26927 9979
rect 28264 9945 28298 9979
rect 30858 9945 30892 9979
rect 34069 9945 34103 9979
rect 37372 9945 37406 9979
rect 43720 9945 43754 9979
rect 45385 9945 45419 9979
rect 49004 9945 49038 9979
rect 50353 9945 50387 9979
rect 54493 9945 54527 9979
rect 55588 9945 55622 9979
rect 57060 9945 57094 9979
rect 10333 9877 10367 9911
rect 14565 9877 14599 9911
rect 19533 9877 19567 9911
rect 26433 9877 26467 9911
rect 27905 9877 27939 9911
rect 29377 9877 29411 9911
rect 29745 9877 29779 9911
rect 33609 9877 33643 9911
rect 34713 9877 34747 9911
rect 38485 9877 38519 9911
rect 38945 9877 38979 9911
rect 39681 9877 39715 9911
rect 45017 9877 45051 9911
rect 45477 9877 45511 9911
rect 45937 9877 45971 9911
rect 47869 9877 47903 9911
rect 49341 9877 49375 9911
rect 54585 9877 54619 9911
rect 56701 9877 56735 9911
rect 58173 9877 58207 9911
rect 4261 9673 4295 9707
rect 5365 9673 5399 9707
rect 13001 9673 13035 9707
rect 29469 9673 29503 9707
rect 36369 9673 36403 9707
rect 40969 9673 41003 9707
rect 41613 9673 41647 9707
rect 43913 9673 43947 9707
rect 44097 9673 44131 9707
rect 45201 9673 45235 9707
rect 46305 9673 46339 9707
rect 47041 9673 47075 9707
rect 53113 9673 53147 9707
rect 56057 9673 56091 9707
rect 57253 9673 57287 9707
rect 57897 9673 57931 9707
rect 2228 9605 2262 9639
rect 4997 9605 5031 9639
rect 5181 9605 5215 9639
rect 6377 9605 6411 9639
rect 6929 9605 6963 9639
rect 10232 9605 10266 9639
rect 15200 9605 15234 9639
rect 19432 9605 19466 9639
rect 22293 9605 22327 9639
rect 24225 9605 24259 9639
rect 27353 9605 27387 9639
rect 28356 9605 28390 9639
rect 37105 9605 37139 9639
rect 38117 9605 38151 9639
rect 40877 9605 40911 9639
rect 41981 9605 42015 9639
rect 45293 9605 45327 9639
rect 48596 9605 48630 9639
rect 54024 9605 54058 9639
rect 55505 9605 55539 9639
rect 1961 9537 1995 9571
rect 3525 9537 3559 9571
rect 4445 9537 4479 9571
rect 4629 9537 4663 9571
rect 4721 9537 4755 9571
rect 4813 9537 4847 9571
rect 5273 9537 5307 9571
rect 5457 9537 5491 9571
rect 6561 9537 6595 9571
rect 9413 9537 9447 9571
rect 12357 9537 12391 9571
rect 13093 9537 13127 9571
rect 13349 9537 13383 9571
rect 14933 9537 14967 9571
rect 17805 9537 17839 9571
rect 18061 9537 18095 9571
rect 18521 9537 18555 9571
rect 19165 9537 19199 9571
rect 22385 9537 22419 9571
rect 22652 9537 22686 9571
rect 24317 9537 24351 9571
rect 26361 9537 26395 9571
rect 27169 9537 27203 9571
rect 29561 9537 29595 9571
rect 30598 9537 30632 9571
rect 32680 9537 32714 9571
rect 34529 9537 34563 9571
rect 34796 9537 34830 9571
rect 36277 9537 36311 9571
rect 37473 9537 37507 9571
rect 38025 9537 38059 9571
rect 39313 9537 39347 9571
rect 39589 9537 39623 9571
rect 40325 9537 40359 9571
rect 44741 9537 44775 9571
rect 45661 9537 45695 9571
rect 46949 9537 46983 9571
rect 48145 9537 48179 9571
rect 48329 9537 48363 9571
rect 49801 9537 49835 9571
rect 53021 9537 53055 9571
rect 55597 9537 55631 9571
rect 58449 9537 58483 9571
rect 8217 9469 8251 9503
rect 8953 9469 8987 9503
rect 9965 9469 9999 9503
rect 12081 9469 12115 9503
rect 18613 9469 18647 9503
rect 18797 9469 18831 9503
rect 20637 9469 20671 9503
rect 24409 9469 24443 9503
rect 26617 9469 26651 9503
rect 27905 9469 27939 9503
rect 28089 9469 28123 9503
rect 29745 9469 29779 9503
rect 30481 9469 30515 9503
rect 30757 9469 30791 9503
rect 31401 9469 31435 9503
rect 32413 9469 32447 9503
rect 36185 9469 36219 9503
rect 38209 9469 38243 9503
rect 39451 9469 39485 9503
rect 40509 9469 40543 9503
rect 40693 9469 40727 9503
rect 45477 9469 45511 9503
rect 47133 9469 47167 9503
rect 52193 9469 52227 9503
rect 52929 9469 52963 9503
rect 53757 9469 53791 9503
rect 55321 9469 55355 9503
rect 56609 9469 56643 9503
rect 57345 9469 57379 9503
rect 57437 9469 57471 9503
rect 3341 9401 3375 9435
rect 3709 9401 3743 9435
rect 11345 9401 11379 9435
rect 20545 9401 20579 9435
rect 23765 9401 23799 9435
rect 24869 9401 24903 9435
rect 30205 9401 30239 9435
rect 34345 9401 34379 9435
rect 39865 9401 39899 9435
rect 44833 9401 44867 9435
rect 49709 9401 49743 9435
rect 55965 9401 55999 9435
rect 7205 9333 7239 9367
rect 7665 9333 7699 9367
rect 8401 9333 8435 9367
rect 9781 9333 9815 9367
rect 11529 9333 11563 9367
rect 14473 9333 14507 9367
rect 14841 9333 14875 9367
rect 16313 9333 16347 9367
rect 16681 9333 16715 9367
rect 18153 9333 18187 9367
rect 21281 9333 21315 9367
rect 23857 9333 23891 9367
rect 25237 9333 25271 9367
rect 31769 9333 31803 9367
rect 33793 9333 33827 9367
rect 35909 9333 35943 9367
rect 36737 9333 36771 9367
rect 37657 9333 37691 9367
rect 38669 9333 38703 9367
rect 41337 9333 41371 9367
rect 46581 9333 46615 9367
rect 47593 9333 47627 9367
rect 51089 9333 51123 9367
rect 51641 9333 51675 9367
rect 53481 9333 53515 9367
rect 55137 9333 55171 9367
rect 56885 9333 56919 9367
rect 6469 9129 6503 9163
rect 6929 9129 6963 9163
rect 7205 9129 7239 9163
rect 8769 9129 8803 9163
rect 10425 9129 10459 9163
rect 15945 9129 15979 9163
rect 18061 9129 18095 9163
rect 19625 9129 19659 9163
rect 23305 9129 23339 9163
rect 26525 9129 26559 9163
rect 29837 9129 29871 9163
rect 33149 9129 33183 9163
rect 34529 9129 34563 9163
rect 36461 9129 36495 9163
rect 37565 9129 37599 9163
rect 38945 9129 38979 9163
rect 39313 9129 39347 9163
rect 42257 9129 42291 9163
rect 44005 9129 44039 9163
rect 45845 9129 45879 9163
rect 49341 9129 49375 9163
rect 49709 9129 49743 9163
rect 50353 9129 50387 9163
rect 52193 9129 52227 9163
rect 52653 9129 52687 9163
rect 53665 9129 53699 9163
rect 55137 9129 55171 9163
rect 56241 9129 56275 9163
rect 57621 9129 57655 9163
rect 11621 9061 11655 9095
rect 26433 9061 26467 9095
rect 40417 9061 40451 9095
rect 46397 9061 46431 9095
rect 48329 9061 48363 9095
rect 54033 9061 54067 9095
rect 54677 9061 54711 9095
rect 55965 9061 55999 9095
rect 4353 8993 4387 9027
rect 10885 8993 10919 9027
rect 10977 8993 11011 9027
rect 16589 8993 16623 9027
rect 16773 8993 16807 9027
rect 16957 8993 16991 9027
rect 18613 8993 18647 9027
rect 19533 8993 19567 9027
rect 20177 8993 20211 9027
rect 23857 8993 23891 9027
rect 25053 8993 25087 9027
rect 25789 8993 25823 9027
rect 27077 8993 27111 9027
rect 28181 8993 28215 9027
rect 29193 8993 29227 9027
rect 30665 8993 30699 9027
rect 33701 8993 33735 9027
rect 33885 8993 33919 9027
rect 35173 8993 35207 9027
rect 35909 8993 35943 9027
rect 38117 8993 38151 9027
rect 38393 8993 38427 9027
rect 47409 8993 47443 9027
rect 47685 8993 47719 9027
rect 47869 8993 47903 9027
rect 48697 8993 48731 9027
rect 50813 8993 50847 9027
rect 55321 8993 55355 9027
rect 56793 8993 56827 9027
rect 56977 8993 57011 9027
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 4445 8925 4479 8959
rect 7389 8925 7423 8959
rect 7656 8925 7690 8959
rect 9781 8925 9815 8959
rect 10333 8925 10367 8959
rect 20085 8925 20119 8959
rect 22845 8925 22879 8959
rect 25605 8925 25639 8959
rect 26065 8925 26099 8959
rect 28457 8925 28491 8959
rect 31493 8925 31527 8959
rect 35265 8925 35299 8959
rect 43453 8925 43487 8959
rect 45293 8925 45327 8959
rect 47961 8925 47995 8959
rect 51080 8925 51114 8959
rect 58265 8925 58299 8959
rect 9137 8857 9171 8891
rect 11437 8857 11471 8891
rect 11897 8857 11931 8891
rect 15761 8857 15795 8891
rect 19073 8857 19107 8891
rect 29009 8857 29043 8891
rect 35357 8857 35391 8891
rect 42165 8857 42199 8891
rect 52929 8857 52963 8891
rect 10793 8789 10827 8823
rect 12357 8789 12391 8823
rect 17049 8789 17083 8823
rect 17417 8789 17451 8823
rect 17969 8789 18003 8823
rect 19993 8789 20027 8823
rect 23121 8789 23155 8823
rect 24869 8789 24903 8823
rect 25973 8789 26007 8823
rect 27445 8789 27479 8823
rect 28641 8789 28675 8823
rect 29101 8789 29135 8823
rect 30113 8789 30147 8823
rect 30481 8789 30515 8823
rect 30573 8789 30607 8823
rect 30941 8789 30975 8823
rect 31953 8789 31987 8823
rect 35725 8789 35759 8823
rect 42901 8789 42935 8823
rect 44649 8789 44683 8823
rect 57713 8789 57747 8823
rect 5457 8585 5491 8619
rect 7573 8585 7607 8619
rect 8033 8585 8067 8619
rect 9505 8585 9539 8619
rect 11805 8585 11839 8619
rect 18337 8585 18371 8619
rect 25237 8585 25271 8619
rect 28457 8585 28491 8619
rect 29929 8585 29963 8619
rect 30757 8585 30791 8619
rect 30849 8585 30883 8619
rect 34897 8585 34931 8619
rect 35909 8585 35943 8619
rect 48513 8585 48547 8619
rect 50169 8585 50203 8619
rect 51549 8585 51583 8619
rect 52377 8585 52411 8619
rect 55873 8585 55907 8619
rect 6193 8517 6227 8551
rect 6561 8517 6595 8551
rect 7941 8517 7975 8551
rect 16497 8517 16531 8551
rect 18889 8517 18923 8551
rect 26556 8517 26590 8551
rect 26985 8517 27019 8551
rect 42800 8517 42834 8551
rect 50077 8517 50111 8551
rect 50537 8517 50571 8551
rect 57345 8517 57379 8551
rect 7205 8449 7239 8483
rect 8493 8449 8527 8483
rect 10149 8449 10183 8483
rect 11161 8449 11195 8483
rect 11897 8449 11931 8483
rect 12357 8449 12391 8483
rect 17693 8449 17727 8483
rect 18797 8449 18831 8483
rect 19901 8449 19935 8483
rect 26801 8449 26835 8483
rect 27905 8449 27939 8483
rect 29009 8449 29043 8483
rect 29377 8449 29411 8483
rect 30205 8449 30239 8483
rect 35541 8449 35575 8483
rect 38669 8449 38703 8483
rect 42533 8449 42567 8483
rect 50629 8449 50663 8483
rect 53481 8449 53515 8483
rect 55965 8449 55999 8483
rect 57253 8449 57287 8483
rect 57897 8449 57931 8483
rect 4997 8381 5031 8415
rect 8125 8381 8159 8415
rect 8769 8381 8803 8415
rect 10287 8381 10321 8415
rect 10425 8381 10459 8415
rect 10701 8381 10735 8415
rect 11345 8381 11379 8415
rect 11621 8381 11655 8415
rect 12909 8381 12943 8415
rect 17049 8381 17083 8415
rect 19073 8381 19107 8415
rect 19257 8381 19291 8415
rect 19993 8381 20027 8415
rect 24041 8381 24075 8415
rect 27537 8381 27571 8415
rect 31401 8381 31435 8415
rect 36645 8381 36679 8415
rect 41429 8381 41463 8415
rect 41613 8381 41647 8415
rect 44557 8381 44591 8415
rect 47593 8381 47627 8415
rect 50721 8381 50755 8415
rect 54585 8381 54619 8415
rect 54769 8381 54803 8415
rect 56241 8381 56275 8415
rect 57437 8381 57471 8415
rect 58449 8381 58483 8415
rect 12265 8313 12299 8347
rect 17601 8313 17635 8347
rect 18429 8313 18463 8347
rect 36093 8313 36127 8347
rect 43913 8313 43947 8347
rect 52009 8313 52043 8347
rect 52929 8313 52963 8347
rect 53849 8313 53883 8347
rect 55321 8313 55355 8347
rect 56885 8313 56919 8347
rect 4629 8245 4663 8279
rect 5825 8245 5859 8279
rect 14105 8245 14139 8279
rect 20637 8245 20671 8279
rect 23489 8245 23523 8279
rect 25421 8245 25455 8279
rect 34529 8245 34563 8279
rect 38393 8245 38427 8279
rect 40785 8245 40819 8279
rect 42165 8245 42199 8279
rect 44005 8245 44039 8279
rect 48237 8245 48271 8279
rect 53941 8245 53975 8279
rect 55597 8245 55631 8279
rect 56793 8245 56827 8279
rect 8033 8041 8067 8075
rect 11897 8041 11931 8075
rect 13921 8041 13955 8075
rect 19073 8041 19107 8075
rect 24133 8041 24167 8075
rect 29745 8041 29779 8075
rect 33609 8041 33643 8075
rect 35265 8041 35299 8075
rect 40877 8041 40911 8075
rect 42809 8041 42843 8075
rect 42993 8041 43027 8075
rect 45293 8041 45327 8075
rect 46949 8041 46983 8075
rect 50445 8041 50479 8075
rect 52745 8041 52779 8075
rect 53205 8041 53239 8075
rect 53573 8041 53607 8075
rect 56609 8041 56643 8075
rect 58081 8041 58115 8075
rect 3801 7973 3835 8007
rect 5733 7973 5767 8007
rect 17325 7973 17359 8007
rect 20453 7973 20487 8007
rect 23121 7973 23155 8007
rect 27905 7973 27939 8007
rect 40785 7973 40819 8007
rect 3617 7905 3651 7939
rect 4445 7905 4479 7939
rect 4813 7905 4847 7939
rect 5641 7905 5675 7939
rect 6377 7905 6411 7939
rect 6837 7905 6871 7939
rect 12541 7905 12575 7939
rect 19257 7905 19291 7939
rect 20060 7905 20094 7939
rect 20177 7905 20211 7939
rect 21097 7905 21131 7939
rect 22661 7905 22695 7939
rect 23673 7905 23707 7939
rect 25145 7905 25179 7939
rect 25789 7905 25823 7939
rect 31125 7905 31159 7939
rect 41521 7905 41555 7939
rect 42257 7905 42291 7939
rect 43545 7905 43579 7939
rect 48329 7905 48363 7939
rect 50813 7905 50847 7939
rect 53757 7905 53791 7939
rect 7389 7837 7423 7871
rect 8217 7837 8251 7871
rect 8953 7837 8987 7871
rect 10517 7837 10551 7871
rect 13461 7837 13495 7871
rect 14749 7837 14783 7871
rect 17233 7837 17267 7871
rect 17693 7837 17727 7871
rect 19901 7837 19935 7871
rect 20913 7837 20947 7871
rect 23029 7837 23063 7871
rect 24409 7837 24443 7871
rect 25881 7837 25915 7871
rect 31769 7837 31803 7871
rect 33149 7837 33183 7871
rect 36093 7837 36127 7871
rect 36829 7837 36863 7871
rect 37565 7837 37599 7871
rect 38117 7837 38151 7871
rect 39405 7837 39439 7871
rect 41245 7837 41279 7871
rect 41337 7837 41371 7871
rect 42073 7837 42107 7871
rect 42165 7837 42199 7871
rect 43453 7837 43487 7871
rect 44557 7837 44591 7871
rect 48973 7837 49007 7871
rect 50997 7837 51031 7871
rect 52285 7837 52319 7871
rect 55965 7837 55999 7871
rect 56701 7837 56735 7871
rect 56957 7837 56991 7871
rect 58357 7837 58391 7871
rect 6101 7769 6135 7803
rect 8769 7769 8803 7803
rect 9198 7769 9232 7803
rect 10784 7769 10818 7803
rect 11989 7769 12023 7803
rect 17509 7769 17543 7803
rect 17960 7769 17994 7803
rect 23489 7769 23523 7803
rect 25053 7769 25087 7803
rect 30880 7769 30914 7803
rect 31217 7769 31251 7803
rect 35357 7769 35391 7803
rect 48084 7769 48118 7803
rect 48421 7769 48455 7803
rect 51733 7769 51767 7803
rect 54024 7769 54058 7803
rect 55321 7769 55355 7803
rect 2973 7701 3007 7735
rect 4169 7701 4203 7735
rect 4261 7701 4295 7735
rect 4997 7701 5031 7735
rect 6193 7701 6227 7735
rect 10333 7701 10367 7735
rect 12909 7701 12943 7735
rect 14105 7701 14139 7735
rect 15117 7701 15151 7735
rect 15853 7701 15887 7735
rect 21465 7701 21499 7735
rect 23581 7701 23615 7735
rect 27169 7701 27203 7735
rect 32597 7701 32631 7735
rect 35541 7701 35575 7735
rect 36277 7701 36311 7735
rect 37013 7701 37047 7735
rect 38761 7701 38795 7735
rect 38853 7701 38887 7735
rect 41705 7701 41739 7735
rect 43361 7701 43395 7735
rect 43913 7701 43947 7735
rect 51641 7701 51675 7735
rect 55137 7701 55171 7735
rect 4261 7497 4295 7531
rect 6837 7497 6871 7531
rect 8861 7497 8895 7531
rect 9229 7497 9263 7531
rect 9321 7497 9355 7531
rect 9873 7497 9907 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 18889 7497 18923 7531
rect 19441 7497 19475 7531
rect 23949 7497 23983 7531
rect 24041 7497 24075 7531
rect 24501 7497 24535 7531
rect 30481 7497 30515 7531
rect 30573 7497 30607 7531
rect 30941 7497 30975 7531
rect 32781 7497 32815 7531
rect 35909 7497 35943 7531
rect 38945 7497 38979 7531
rect 41705 7497 41739 7531
rect 41981 7497 42015 7531
rect 44373 7497 44407 7531
rect 47869 7497 47903 7531
rect 48329 7497 48363 7531
rect 51733 7497 51767 7531
rect 52193 7497 52227 7531
rect 54861 7497 54895 7531
rect 8493 7429 8527 7463
rect 11805 7429 11839 7463
rect 12624 7429 12658 7463
rect 14473 7429 14507 7463
rect 15669 7429 15703 7463
rect 34796 7429 34830 7463
rect 36461 7429 36495 7463
rect 40592 7429 40626 7463
rect 44833 7429 44867 7463
rect 47961 7429 47995 7463
rect 48789 7429 48823 7463
rect 58265 7429 58299 7463
rect 2412 7361 2446 7395
rect 4997 7361 5031 7395
rect 6009 7361 6043 7395
rect 8125 7361 8159 7395
rect 12357 7361 12391 7395
rect 17509 7361 17543 7395
rect 17776 7361 17810 7395
rect 19349 7361 19383 7395
rect 20260 7361 20294 7395
rect 22569 7361 22603 7395
rect 22836 7361 22870 7395
rect 24409 7361 24443 7395
rect 25605 7361 25639 7395
rect 25881 7361 25915 7395
rect 26617 7361 26651 7395
rect 27353 7361 27387 7395
rect 27813 7361 27847 7395
rect 33149 7361 33183 7395
rect 33241 7361 33275 7395
rect 34253 7361 34287 7395
rect 36369 7361 36403 7395
rect 37565 7361 37599 7395
rect 37832 7361 37866 7395
rect 39037 7361 39071 7395
rect 40325 7361 40359 7395
rect 43085 7361 43119 7395
rect 43223 7361 43257 7395
rect 43361 7361 43395 7395
rect 44097 7361 44131 7395
rect 44741 7361 44775 7395
rect 45201 7361 45235 7395
rect 48973 7361 49007 7395
rect 49893 7361 49927 7395
rect 51109 7361 51143 7395
rect 51365 7361 51399 7395
rect 51825 7361 51859 7395
rect 53481 7361 53515 7395
rect 53748 7361 53782 7395
rect 56241 7361 56275 7395
rect 56379 7361 56413 7395
rect 56517 7361 56551 7395
rect 57253 7361 57287 7395
rect 58449 7361 58483 7395
rect 2145 7293 2179 7327
rect 3617 7293 3651 7327
rect 5156 7293 5190 7327
rect 5273 7293 5307 7327
rect 5549 7293 5583 7327
rect 6193 7293 6227 7327
rect 9413 7293 9447 7327
rect 10425 7293 10459 7327
rect 14289 7293 14323 7327
rect 15025 7293 15059 7327
rect 17325 7293 17359 7327
rect 19625 7293 19659 7327
rect 19993 7293 20027 7327
rect 22385 7293 22419 7327
rect 24685 7293 24719 7327
rect 25743 7293 25777 7327
rect 26801 7293 26835 7327
rect 27445 7293 27479 7327
rect 27537 7293 27571 7327
rect 28365 7293 28399 7327
rect 29377 7293 29411 7327
rect 30113 7293 30147 7327
rect 30389 7293 30423 7327
rect 32597 7293 32631 7327
rect 33333 7293 33367 7327
rect 33609 7293 33643 7327
rect 34529 7293 34563 7327
rect 36553 7293 36587 7327
rect 37013 7293 37047 7327
rect 39589 7293 39623 7327
rect 44281 7293 44315 7327
rect 44925 7293 44959 7327
rect 45753 7293 45787 7327
rect 46489 7293 46523 7327
rect 46673 7293 46707 7327
rect 47685 7293 47719 7327
rect 48697 7293 48731 7327
rect 51641 7293 51675 7327
rect 53297 7293 53331 7327
rect 56793 7293 56827 7327
rect 57437 7293 57471 7327
rect 14013 7225 14047 7259
rect 16037 7225 16071 7259
rect 21373 7225 21407 7259
rect 26157 7225 26191 7259
rect 31217 7225 31251 7259
rect 43637 7225 43671 7259
rect 52561 7225 52595 7259
rect 3525 7157 3559 7191
rect 4353 7157 4387 7191
rect 11069 7157 11103 7191
rect 12081 7157 12115 7191
rect 13737 7157 13771 7191
rect 16405 7157 16439 7191
rect 16681 7157 16715 7191
rect 18981 7157 19015 7191
rect 21833 7157 21867 7191
rect 24961 7157 24995 7191
rect 26985 7157 27019 7191
rect 28733 7157 28767 7191
rect 29469 7157 29503 7191
rect 36001 7157 36035 7191
rect 42441 7157 42475 7191
rect 45937 7157 45971 7191
rect 47317 7157 47351 7191
rect 49433 7157 49467 7191
rect 49985 7157 50019 7191
rect 52745 7157 52779 7191
rect 55229 7157 55263 7191
rect 55597 7157 55631 7191
rect 58081 7157 58115 7191
rect 3433 6953 3467 6987
rect 9137 6953 9171 6987
rect 13921 6953 13955 6987
rect 17509 6953 17543 6987
rect 18429 6953 18463 6987
rect 19533 6953 19567 6987
rect 21005 6953 21039 6987
rect 25053 6953 25087 6987
rect 27813 6953 27847 6987
rect 29377 6953 29411 6987
rect 33425 6953 33459 6987
rect 36185 6953 36219 6987
rect 37105 6953 37139 6987
rect 46397 6953 46431 6987
rect 52561 6953 52595 6987
rect 56057 6953 56091 6987
rect 15393 6885 15427 6919
rect 41705 6885 41739 6919
rect 51273 6885 51307 6919
rect 4445 6817 4479 6851
rect 10057 6817 10091 6851
rect 11897 6817 11931 6851
rect 15117 6817 15151 6851
rect 16037 6817 16071 6851
rect 18981 6817 19015 6851
rect 20269 6817 20303 6851
rect 21741 6817 21775 6851
rect 22477 6817 22511 6851
rect 25513 6817 25547 6851
rect 25962 6817 25996 6851
rect 27997 6817 28031 6851
rect 33977 6817 34011 6851
rect 34161 6817 34195 6851
rect 36829 6817 36863 6851
rect 38669 6817 38703 6851
rect 38853 6817 38887 6851
rect 43177 6817 43211 6851
rect 46581 6817 46615 6851
rect 47225 6817 47259 6851
rect 47501 6817 47535 6851
rect 47618 6817 47652 6851
rect 48973 6817 49007 6851
rect 49065 6817 49099 6851
rect 50675 6817 50709 6851
rect 51549 6817 51583 6851
rect 51825 6817 51859 6851
rect 54125 6817 54159 6851
rect 55045 6817 55079 6851
rect 55505 6817 55539 6851
rect 2053 6749 2087 6783
rect 4905 6749 4939 6783
rect 5172 6749 5206 6783
rect 6377 6749 6411 6783
rect 8401 6749 8435 6783
rect 10793 6749 10827 6783
rect 11437 6749 11471 6783
rect 12541 6749 12575 6783
rect 14841 6749 14875 6783
rect 14979 6749 15013 6783
rect 15853 6749 15887 6783
rect 16129 6749 16163 6783
rect 18153 6749 18187 6783
rect 20545 6749 20579 6783
rect 21557 6749 21591 6783
rect 24409 6749 24443 6783
rect 29561 6749 29595 6783
rect 31585 6749 31619 6783
rect 32045 6749 32079 6783
rect 34713 6749 34747 6783
rect 38485 6749 38519 6783
rect 40049 6749 40083 6783
rect 40325 6749 40359 6783
rect 42349 6749 42383 6783
rect 45017 6749 45051 6783
rect 45284 6749 45318 6783
rect 46765 6749 46799 6783
rect 47777 6749 47811 6783
rect 49985 6749 50019 6783
rect 50813 6749 50847 6783
rect 51687 6749 51721 6783
rect 53941 6749 53975 6783
rect 54309 6749 54343 6783
rect 56425 6749 56459 6783
rect 58449 6749 58483 6783
rect 2320 6681 2354 6715
rect 6644 6681 6678 6715
rect 7849 6681 7883 6715
rect 9597 6681 9631 6715
rect 12808 6681 12842 6715
rect 16396 6681 16430 6715
rect 17601 6681 17635 6715
rect 20453 6681 20487 6715
rect 21925 6681 21959 6715
rect 22744 6681 22778 6715
rect 25329 6681 25363 6715
rect 26240 6681 26274 6715
rect 28264 6681 28298 6715
rect 29806 6681 29840 6715
rect 32312 6681 32346 6715
rect 34980 6681 35014 6715
rect 38240 6681 38274 6715
rect 40592 6681 40626 6715
rect 41797 6681 41831 6715
rect 43444 6681 43478 6715
rect 48421 6681 48455 6715
rect 48881 6681 48915 6715
rect 53696 6681 53730 6715
rect 55597 6681 55631 6715
rect 56692 6681 56726 6715
rect 57897 6681 57931 6715
rect 3801 6613 3835 6647
rect 4169 6613 4203 6647
rect 4261 6613 4295 6647
rect 6285 6613 6319 6647
rect 7757 6613 7791 6647
rect 10149 6613 10183 6647
rect 10885 6613 10919 6647
rect 12449 6613 12483 6647
rect 14197 6613 14231 6647
rect 19809 6613 19843 6647
rect 20913 6613 20947 6647
rect 23857 6613 23891 6647
rect 24225 6613 24259 6647
rect 27353 6613 27387 6647
rect 30941 6613 30975 6647
rect 31033 6613 31067 6647
rect 33517 6613 33551 6647
rect 33885 6613 33919 6647
rect 36093 6613 36127 6647
rect 36553 6613 36587 6647
rect 36645 6613 36679 6647
rect 38945 6613 38979 6647
rect 39313 6613 39347 6647
rect 39681 6613 39715 6647
rect 44557 6613 44591 6647
rect 48513 6613 48547 6647
rect 49341 6613 49375 6647
rect 50445 6613 50479 6647
rect 52469 6613 52503 6647
rect 54401 6613 54435 6647
rect 54769 6613 54803 6647
rect 55689 6613 55723 6647
rect 57805 6613 57839 6647
rect 3157 6409 3191 6443
rect 4537 6409 4571 6443
rect 6193 6409 6227 6443
rect 7297 6409 7331 6443
rect 7665 6409 7699 6443
rect 11069 6409 11103 6443
rect 12633 6409 12667 6443
rect 13185 6409 13219 6443
rect 16129 6409 16163 6443
rect 16957 6409 16991 6443
rect 17049 6409 17083 6443
rect 17417 6409 17451 6443
rect 20453 6409 20487 6443
rect 22937 6409 22971 6443
rect 24869 6409 24903 6443
rect 25881 6409 25915 6443
rect 26249 6409 26283 6443
rect 26709 6409 26743 6443
rect 26985 6409 27019 6443
rect 27905 6409 27939 6443
rect 28181 6409 28215 6443
rect 30021 6409 30055 6443
rect 33793 6409 33827 6443
rect 35725 6409 35759 6443
rect 36829 6409 36863 6443
rect 40049 6409 40083 6443
rect 43085 6409 43119 6443
rect 44281 6409 44315 6443
rect 45385 6409 45419 6443
rect 45845 6409 45879 6443
rect 47593 6409 47627 6443
rect 48053 6409 48087 6443
rect 48421 6409 48455 6443
rect 52101 6409 52135 6443
rect 53113 6409 53147 6443
rect 54217 6409 54251 6443
rect 54677 6409 54711 6443
rect 56149 6409 56183 6443
rect 57069 6409 57103 6443
rect 57437 6409 57471 6443
rect 2697 6341 2731 6375
rect 9956 6341 9990 6375
rect 13093 6341 13127 6375
rect 13820 6341 13854 6375
rect 16221 6341 16255 6375
rect 17969 6341 18003 6375
rect 30389 6341 30423 6375
rect 36185 6341 36219 6375
rect 47961 6341 47995 6375
rect 49586 6341 49620 6375
rect 52193 6341 52227 6375
rect 56517 6341 56551 6375
rect 3801 6273 3835 6307
rect 3893 6273 3927 6307
rect 7205 6273 7239 6307
rect 8309 6273 8343 6307
rect 9689 6273 9723 6307
rect 12081 6273 12115 6307
rect 15209 6273 15243 6307
rect 20821 6273 20855 6307
rect 23489 6273 23523 6307
rect 26341 6273 26375 6307
rect 27629 6273 27663 6307
rect 29285 6273 29319 6307
rect 32137 6273 32171 6307
rect 32404 6273 32438 6307
rect 34713 6273 34747 6307
rect 35449 6273 35483 6307
rect 36093 6273 36127 6307
rect 37657 6273 37691 6307
rect 39497 6273 39531 6307
rect 39957 6273 39991 6307
rect 42441 6273 42475 6307
rect 45477 6273 45511 6307
rect 46029 6273 46063 6307
rect 46296 6273 46330 6307
rect 49341 6273 49375 6307
rect 51181 6273 51215 6307
rect 53205 6273 53239 6307
rect 55321 6273 55355 6307
rect 55505 6273 55539 6307
rect 58449 6273 58483 6307
rect 2329 6205 2363 6239
rect 7113 6205 7147 6239
rect 7757 6205 7791 6239
rect 9229 6205 9263 6239
rect 13277 6205 13311 6239
rect 13553 6205 13587 6239
rect 16313 6205 16347 6239
rect 16773 6205 16807 6239
rect 18061 6205 18095 6239
rect 18797 6205 18831 6239
rect 20085 6205 20119 6239
rect 24225 6205 24259 6239
rect 26065 6205 26099 6239
rect 28825 6205 28859 6239
rect 29377 6205 29411 6239
rect 29561 6205 29595 6239
rect 30481 6205 30515 6239
rect 30573 6205 30607 6239
rect 31033 6205 31067 6239
rect 34437 6205 34471 6239
rect 34596 6205 34630 6239
rect 35633 6205 35667 6239
rect 36277 6205 36311 6239
rect 37841 6205 37875 6239
rect 38577 6205 38611 6239
rect 38715 6205 38749 6239
rect 38853 6205 38887 6239
rect 40141 6205 40175 6239
rect 45293 6205 45327 6239
rect 48145 6205 48179 6239
rect 48973 6205 49007 6239
rect 51273 6205 51307 6239
rect 51457 6205 51491 6239
rect 51917 6205 51951 6239
rect 53389 6205 53423 6239
rect 53573 6205 53607 6239
rect 56885 6205 56919 6239
rect 56977 6205 57011 6239
rect 57897 6205 57931 6239
rect 1961 6137 1995 6171
rect 4997 6137 5031 6171
rect 5365 6137 5399 6171
rect 6745 6137 6779 6171
rect 14933 6137 14967 6171
rect 19533 6137 19567 6171
rect 21281 6137 21315 6171
rect 25421 6137 25455 6171
rect 28917 6137 28951 6171
rect 31401 6137 31435 6171
rect 34989 6137 35023 6171
rect 38301 6137 38335 6171
rect 47409 6137 47443 6171
rect 50813 6137 50847 6171
rect 52561 6137 52595 6171
rect 2973 6069 3007 6103
rect 5825 6069 5859 6103
rect 8677 6069 8711 6103
rect 11897 6069 11931 6103
rect 12725 6069 12759 6103
rect 15577 6069 15611 6103
rect 15761 6069 15795 6103
rect 18705 6069 18739 6103
rect 19441 6069 19475 6103
rect 21557 6069 21591 6103
rect 22017 6069 22051 6103
rect 22661 6069 22695 6103
rect 23673 6069 23707 6103
rect 33517 6069 33551 6103
rect 37473 6069 37507 6103
rect 39589 6069 39623 6103
rect 44649 6069 44683 6103
rect 45017 6069 45051 6103
rect 50721 6069 50755 6103
rect 52745 6069 52779 6103
rect 54585 6069 54619 6103
rect 1869 5865 1903 5899
rect 8953 5865 8987 5899
rect 10977 5865 11011 5899
rect 13001 5865 13035 5899
rect 13093 5865 13127 5899
rect 14749 5865 14783 5899
rect 15209 5865 15243 5899
rect 19257 5865 19291 5899
rect 22017 5865 22051 5899
rect 24041 5865 24075 5899
rect 29745 5865 29779 5899
rect 30389 5865 30423 5899
rect 31125 5865 31159 5899
rect 32965 5865 32999 5899
rect 34437 5865 34471 5899
rect 35357 5865 35391 5899
rect 38853 5865 38887 5899
rect 46397 5865 46431 5899
rect 46949 5865 46983 5899
rect 47869 5865 47903 5899
rect 48237 5865 48271 5899
rect 48697 5865 48731 5899
rect 51641 5865 51675 5899
rect 52009 5865 52043 5899
rect 3341 5797 3375 5831
rect 6101 5797 6135 5831
rect 8769 5797 8803 5831
rect 12173 5797 12207 5831
rect 22845 5797 22879 5831
rect 26801 5797 26835 5831
rect 38761 5797 38795 5831
rect 45201 5797 45235 5831
rect 1961 5729 1995 5763
rect 4445 5729 4479 5763
rect 4629 5729 4663 5763
rect 6837 5729 6871 5763
rect 9413 5729 9447 5763
rect 9505 5729 9539 5763
rect 10333 5729 10367 5763
rect 13737 5729 13771 5763
rect 14105 5729 14139 5763
rect 18429 5729 18463 5763
rect 20637 5729 20671 5763
rect 22753 5729 22787 5763
rect 23397 5729 23431 5763
rect 26157 5729 26191 5763
rect 26341 5729 26375 5763
rect 27445 5729 27479 5763
rect 33517 5729 33551 5763
rect 33793 5729 33827 5763
rect 37565 5729 37599 5763
rect 38117 5729 38151 5763
rect 44741 5729 44775 5763
rect 47593 5729 47627 5763
rect 50997 5729 51031 5763
rect 6285 5661 6319 5695
rect 7573 5661 7607 5695
rect 8309 5661 8343 5695
rect 10517 5661 10551 5695
rect 10609 5661 10643 5695
rect 11621 5661 11655 5695
rect 15669 5661 15703 5695
rect 16773 5661 16807 5695
rect 17601 5661 17635 5695
rect 18337 5661 18371 5695
rect 21281 5661 21315 5695
rect 24961 5661 24995 5695
rect 25881 5661 25915 5695
rect 35449 5661 35483 5695
rect 37841 5661 37875 5695
rect 39405 5661 39439 5695
rect 40141 5661 40175 5695
rect 41429 5661 41463 5695
rect 41797 5661 41831 5695
rect 42441 5661 42475 5695
rect 42993 5661 43027 5695
rect 44373 5661 44407 5695
rect 49709 5661 49743 5695
rect 50721 5661 50755 5695
rect 52837 5661 52871 5695
rect 54125 5661 54159 5695
rect 54861 5661 54895 5695
rect 55873 5661 55907 5695
rect 56609 5661 56643 5695
rect 57345 5661 57379 5695
rect 57897 5661 57931 5695
rect 2228 5593 2262 5627
rect 4169 5593 4203 5627
rect 5273 5593 5307 5627
rect 5825 5593 5859 5627
rect 9321 5593 9355 5627
rect 11069 5593 11103 5627
rect 13461 5593 13495 5627
rect 20392 5593 20426 5627
rect 20729 5593 20763 5627
rect 23213 5593 23247 5627
rect 26433 5593 26467 5627
rect 30297 5593 30331 5627
rect 37197 5593 37231 5627
rect 38393 5593 38427 5627
rect 39957 5593 39991 5627
rect 47777 5593 47811 5627
rect 53297 5593 53331 5627
rect 57713 5593 57747 5627
rect 3801 5525 3835 5559
rect 4261 5525 4295 5559
rect 7021 5525 7055 5559
rect 7757 5525 7791 5559
rect 10057 5525 10091 5559
rect 12633 5525 12667 5559
rect 13553 5525 13587 5559
rect 15577 5525 15611 5559
rect 16313 5525 16347 5559
rect 16957 5525 16991 5559
rect 17693 5525 17727 5559
rect 19073 5525 19107 5559
rect 22109 5525 22143 5559
rect 23305 5525 23339 5559
rect 24409 5525 24443 5559
rect 25329 5525 25363 5559
rect 26893 5525 26927 5559
rect 30757 5525 30791 5559
rect 38301 5525 38335 5559
rect 40877 5525 40911 5559
rect 42349 5525 42383 5559
rect 43821 5525 43855 5559
rect 49065 5525 49099 5559
rect 50169 5525 50203 5559
rect 52285 5525 52319 5559
rect 53573 5525 53607 5559
rect 54309 5525 54343 5559
rect 55321 5525 55355 5559
rect 56057 5525 56091 5559
rect 56793 5525 56827 5559
rect 58541 5525 58575 5559
rect 3065 5321 3099 5355
rect 5733 5321 5767 5355
rect 9413 5321 9447 5355
rect 11989 5321 12023 5355
rect 15393 5321 15427 5355
rect 18245 5321 18279 5355
rect 18337 5321 18371 5355
rect 20085 5321 20119 5355
rect 22385 5321 22419 5355
rect 23949 5321 23983 5355
rect 24317 5321 24351 5355
rect 24409 5321 24443 5355
rect 25421 5321 25455 5355
rect 27261 5321 27295 5355
rect 27997 5321 28031 5355
rect 28733 5321 28767 5355
rect 36921 5321 36955 5355
rect 40877 5321 40911 5355
rect 41061 5321 41095 5355
rect 41521 5321 41555 5355
rect 43913 5321 43947 5355
rect 46765 5321 46799 5355
rect 53205 5321 53239 5355
rect 54677 5321 54711 5355
rect 55045 5321 55079 5355
rect 55137 5321 55171 5355
rect 57529 5321 57563 5355
rect 4537 5253 4571 5287
rect 8300 5253 8334 5287
rect 13829 5253 13863 5287
rect 17132 5253 17166 5287
rect 19625 5253 19659 5287
rect 20453 5253 20487 5287
rect 22744 5253 22778 5287
rect 26556 5253 26590 5287
rect 29469 5253 29503 5287
rect 37565 5253 37599 5287
rect 42073 5253 42107 5287
rect 44373 5253 44407 5287
rect 45109 5253 45143 5287
rect 45477 5253 45511 5287
rect 49249 5253 49283 5287
rect 50997 5253 51031 5287
rect 56250 5253 56284 5287
rect 1869 5185 1903 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 6644 5185 6678 5219
rect 8033 5185 8067 5219
rect 9505 5185 9539 5219
rect 10542 5185 10576 5219
rect 11345 5185 11379 5219
rect 11897 5185 11931 5219
rect 16865 5185 16899 5219
rect 18705 5185 18739 5219
rect 19717 5185 19751 5219
rect 20545 5185 20579 5219
rect 25053 5185 25087 5219
rect 26801 5185 26835 5219
rect 27353 5185 27387 5219
rect 30205 5185 30239 5219
rect 41429 5185 41463 5219
rect 43085 5185 43119 5219
rect 44281 5185 44315 5219
rect 45293 5185 45327 5219
rect 48717 5185 48751 5219
rect 48973 5185 49007 5219
rect 51825 5185 51859 5219
rect 53297 5185 53331 5219
rect 54585 5185 54619 5219
rect 56517 5185 56551 5219
rect 57713 5185 57747 5219
rect 2973 5117 3007 5151
rect 3709 5117 3743 5151
rect 3801 5117 3835 5151
rect 5089 5117 5123 5151
rect 5641 5117 5675 5151
rect 9689 5117 9723 5151
rect 10425 5117 10459 5151
rect 10701 5117 10735 5151
rect 12081 5117 12115 5151
rect 12909 5117 12943 5151
rect 14289 5117 14323 5151
rect 15669 5117 15703 5151
rect 16497 5117 16531 5151
rect 18797 5117 18831 5151
rect 18889 5117 18923 5151
rect 19533 5117 19567 5151
rect 20361 5117 20395 5151
rect 21097 5117 21131 5151
rect 22477 5117 22511 5151
rect 24501 5117 24535 5151
rect 27169 5117 27203 5151
rect 28365 5117 28399 5151
rect 30389 5117 30423 5151
rect 31309 5117 31343 5151
rect 36369 5117 36403 5151
rect 38301 5117 38335 5151
rect 39221 5117 39255 5151
rect 39865 5117 39899 5151
rect 41705 5117 41739 5151
rect 42441 5117 42475 5151
rect 43729 5117 43763 5151
rect 44557 5117 44591 5151
rect 46029 5117 46063 5151
rect 47409 5117 47443 5151
rect 51641 5117 51675 5151
rect 52377 5117 52411 5151
rect 53481 5117 53515 5151
rect 54493 5117 54527 5151
rect 57161 5117 57195 5151
rect 58449 5117 58483 5151
rect 4445 5049 4479 5083
rect 10149 5049 10183 5083
rect 23857 5049 23891 5083
rect 33793 5049 33827 5083
rect 35725 5049 35759 5083
rect 47593 5049 47627 5083
rect 2237 4981 2271 5015
rect 2329 4981 2363 5015
rect 6193 4981 6227 5015
rect 7757 4981 7791 5015
rect 11529 4981 11563 5015
rect 12357 4981 12391 5015
rect 13461 4981 13495 5015
rect 14105 4981 14139 5015
rect 14933 4981 14967 5015
rect 15853 4981 15887 5015
rect 20913 4981 20947 5015
rect 21649 4981 21683 5015
rect 27721 4981 27755 5015
rect 29561 4981 29595 5015
rect 31033 4981 31067 5015
rect 31677 4981 31711 5015
rect 33425 4981 33459 5015
rect 35817 4981 35851 5015
rect 37749 4981 37783 5015
rect 38577 4981 38611 5015
rect 39313 4981 39347 5015
rect 40509 4981 40543 5015
rect 43177 4981 43211 5015
rect 45017 4981 45051 5015
rect 46581 4981 46615 5015
rect 51089 4981 51123 5015
rect 52929 4981 52963 5015
rect 54125 4981 54159 5015
rect 56609 4981 56643 5015
rect 57897 4981 57931 5015
rect 3249 4777 3283 4811
rect 7021 4777 7055 4811
rect 14933 4777 14967 4811
rect 15761 4777 15795 4811
rect 17601 4777 17635 4811
rect 19809 4777 19843 4811
rect 24225 4777 24259 4811
rect 26249 4777 26283 4811
rect 28457 4777 28491 4811
rect 33701 4777 33735 4811
rect 34437 4777 34471 4811
rect 37841 4777 37875 4811
rect 38761 4777 38795 4811
rect 41797 4777 41831 4811
rect 48329 4777 48363 4811
rect 51549 4777 51583 4811
rect 53297 4777 53331 4811
rect 55873 4777 55907 4811
rect 4445 4709 4479 4743
rect 11253 4709 11287 4743
rect 14657 4709 14691 4743
rect 23489 4709 23523 4743
rect 30205 4709 30239 4743
rect 32505 4709 32539 4743
rect 33057 4709 33091 4743
rect 33609 4709 33643 4743
rect 38669 4709 38703 4743
rect 44833 4709 44867 4743
rect 47961 4709 47995 4743
rect 49065 4709 49099 4743
rect 55137 4709 55171 4743
rect 1869 4641 1903 4675
rect 3801 4641 3835 4675
rect 4838 4641 4872 4675
rect 4997 4641 5031 4675
rect 6377 4641 6411 4675
rect 7481 4641 7515 4675
rect 9137 4641 9171 4675
rect 10609 4641 10643 4675
rect 11897 4641 11931 4675
rect 12541 4641 12575 4675
rect 18245 4641 18279 4675
rect 23581 4641 23615 4675
rect 24409 4641 24443 4675
rect 24593 4641 24627 4675
rect 25053 4641 25087 4675
rect 25329 4641 25363 4675
rect 25467 4641 25501 4675
rect 26709 4641 26743 4675
rect 29745 4641 29779 4675
rect 30598 4641 30632 4675
rect 30757 4641 30791 4675
rect 32045 4641 32079 4675
rect 37197 4641 37231 4675
rect 38117 4641 38151 4675
rect 40049 4641 40083 4675
rect 42625 4641 42659 4675
rect 43269 4641 43303 4675
rect 43683 4641 43717 4675
rect 43821 4641 43855 4675
rect 45569 4641 45603 4675
rect 47133 4641 47167 4675
rect 47409 4641 47443 4675
rect 48421 4641 48455 4675
rect 50169 4641 50203 4675
rect 55597 4641 55631 4675
rect 56241 4641 56275 4675
rect 56425 4641 56459 4675
rect 1777 4573 1811 4607
rect 3985 4573 4019 4607
rect 4721 4573 4755 4607
rect 5641 4573 5675 4607
rect 6561 4573 6595 4607
rect 6653 4573 6687 4607
rect 8125 4573 8159 4607
rect 9781 4573 9815 4607
rect 10885 4573 10919 4607
rect 13185 4573 13219 4607
rect 13921 4573 13955 4607
rect 15117 4573 15151 4607
rect 17233 4573 17267 4607
rect 18429 4573 18463 4607
rect 20453 4573 20487 4607
rect 21189 4573 21223 4607
rect 21465 4573 21499 4607
rect 22109 4573 22143 4607
rect 22365 4573 22399 4607
rect 25605 4573 25639 4607
rect 27445 4573 27479 4607
rect 28089 4573 28123 4607
rect 29377 4573 29411 4607
rect 29561 4573 29595 4607
rect 30481 4573 30515 4607
rect 31953 4573 31987 4607
rect 33885 4573 33919 4607
rect 34253 4573 34287 4607
rect 35541 4573 35575 4607
rect 36277 4573 36311 4607
rect 37473 4573 37507 4607
rect 38209 4573 38243 4607
rect 39313 4573 39347 4607
rect 40417 4573 40451 4607
rect 42441 4573 42475 4607
rect 42809 4573 42843 4607
rect 43545 4573 43579 4607
rect 45845 4573 45879 4607
rect 46397 4573 46431 4607
rect 47593 4573 47627 4607
rect 49709 4573 49743 4607
rect 50436 4573 50470 4607
rect 52193 4573 52227 4607
rect 52929 4573 52963 4607
rect 53113 4573 53147 4607
rect 53757 4573 53791 4607
rect 54024 4573 54058 4607
rect 58265 4573 58299 4607
rect 2136 4505 2170 4539
rect 3433 4505 3467 4539
rect 6101 4505 6135 4539
rect 8769 4505 8803 4539
rect 15301 4505 15335 4539
rect 31401 4505 31435 4539
rect 31861 4505 31895 4539
rect 40684 4505 40718 4539
rect 44465 4505 44499 4539
rect 45385 4505 45419 4539
rect 55413 4505 55447 4539
rect 56517 4505 56551 4539
rect 57161 4505 57195 4539
rect 3525 4437 3559 4471
rect 8033 4437 8067 4471
rect 9689 4437 9723 4471
rect 10425 4437 10459 4471
rect 10793 4437 10827 4471
rect 11345 4437 11379 4471
rect 12449 4437 12483 4471
rect 13277 4437 13311 4471
rect 17969 4437 18003 4471
rect 18061 4437 18095 4471
rect 19073 4437 19107 4471
rect 19901 4437 19935 4471
rect 20637 4437 20671 4471
rect 22017 4437 22051 4471
rect 26801 4437 26835 4471
rect 27537 4437 27571 4471
rect 28733 4437 28767 4471
rect 31493 4437 31527 4471
rect 34989 4437 35023 4471
rect 35725 4437 35759 4471
rect 36645 4437 36679 4471
rect 37381 4437 37415 4471
rect 38301 4437 38335 4471
rect 41889 4437 41923 4471
rect 45017 4437 45051 4471
rect 45477 4437 45511 4471
rect 47501 4437 47535 4471
rect 49157 4437 49191 4471
rect 51641 4437 51675 4471
rect 52377 4437 52411 4471
rect 53573 4437 53607 4471
rect 56885 4437 56919 4471
rect 2973 4233 3007 4267
rect 3341 4233 3375 4267
rect 8033 4233 8067 4267
rect 8861 4233 8895 4267
rect 9229 4233 9263 4267
rect 9321 4233 9355 4267
rect 9781 4233 9815 4267
rect 10241 4233 10275 4267
rect 10701 4233 10735 4267
rect 13921 4233 13955 4267
rect 15945 4233 15979 4267
rect 18245 4233 18279 4267
rect 20177 4233 20211 4267
rect 20269 4233 20303 4267
rect 20729 4233 20763 4267
rect 21557 4233 21591 4267
rect 24041 4233 24075 4267
rect 25789 4233 25823 4267
rect 27261 4233 27295 4267
rect 27721 4233 27755 4267
rect 29745 4233 29779 4267
rect 31033 4233 31067 4267
rect 35081 4233 35115 4267
rect 35909 4233 35943 4267
rect 38669 4233 38703 4267
rect 39037 4233 39071 4267
rect 39497 4233 39531 4267
rect 41429 4233 41463 4267
rect 41889 4233 41923 4267
rect 42809 4233 42843 4267
rect 43269 4233 43303 4267
rect 44741 4233 44775 4267
rect 45201 4233 45235 4267
rect 45569 4233 45603 4267
rect 48697 4233 48731 4267
rect 49065 4233 49099 4267
rect 49525 4233 49559 4267
rect 50445 4233 50479 4267
rect 52285 4233 52319 4267
rect 53113 4233 53147 4267
rect 56149 4233 56183 4267
rect 6561 4165 6595 4199
rect 6837 4165 6871 4199
rect 8677 4165 8711 4199
rect 10609 4165 10643 4199
rect 25881 4165 25915 4199
rect 27353 4165 27387 4199
rect 30113 4165 30147 4199
rect 30941 4165 30975 4199
rect 35449 4165 35483 4199
rect 37556 4165 37590 4199
rect 39129 4165 39163 4199
rect 51917 4165 51951 4199
rect 3433 4097 3467 4131
rect 4813 4097 4847 4131
rect 6377 4097 6411 4131
rect 7389 4097 7423 4131
rect 8493 4097 8527 4131
rect 9965 4097 9999 4131
rect 13461 4097 13495 4131
rect 16865 4097 16899 4131
rect 17132 4097 17166 4131
rect 19257 4097 19291 4131
rect 19533 4097 19567 4131
rect 20637 4097 20671 4131
rect 28089 4097 28123 4131
rect 28273 4097 28307 4131
rect 28540 4097 28574 4131
rect 30205 4097 30239 4131
rect 31677 4097 31711 4131
rect 35541 4097 35575 4131
rect 36277 4097 36311 4131
rect 37013 4097 37047 4131
rect 40141 4097 40175 4131
rect 41521 4097 41555 4131
rect 41981 4097 42015 4131
rect 42901 4097 42935 4131
rect 43361 4097 43395 4131
rect 43628 4097 43662 4131
rect 45109 4097 45143 4131
rect 46397 4097 46431 4131
rect 48605 4097 48639 4131
rect 50353 4097 50387 4131
rect 54493 4097 54527 4131
rect 55346 4097 55380 4131
rect 57713 4097 57747 4131
rect 58449 4097 58483 4131
rect 2145 4029 2179 4063
rect 2329 4029 2363 4063
rect 3617 4029 3651 4063
rect 4169 4029 4203 4063
rect 5457 4029 5491 4063
rect 5641 4029 5675 4063
rect 6193 4029 6227 4063
rect 8309 4029 8343 4063
rect 9505 4029 9539 4063
rect 10885 4029 10919 4063
rect 12081 4029 12115 4063
rect 12449 4029 12483 4063
rect 14197 4029 14231 4063
rect 14933 4029 14967 4063
rect 15485 4029 15519 4063
rect 16037 4029 16071 4063
rect 16129 4029 16163 4063
rect 18337 4029 18371 4063
rect 18521 4029 18555 4063
rect 18981 4029 19015 4063
rect 19374 4029 19408 4063
rect 20821 4029 20855 4063
rect 22293 4029 22327 4063
rect 23029 4029 23063 4063
rect 23581 4029 23615 4063
rect 24133 4029 24167 4063
rect 24225 4029 24259 4063
rect 25237 4029 25271 4063
rect 26617 4029 26651 4063
rect 27169 4029 27203 4063
rect 30297 4029 30331 4063
rect 31125 4029 31159 4063
rect 32689 4029 32723 4063
rect 33425 4029 33459 4063
rect 34161 4029 34195 4063
rect 34897 4029 34931 4063
rect 35725 4029 35759 4063
rect 36369 4029 36403 4063
rect 36553 4029 36587 4063
rect 37289 4029 37323 4063
rect 38945 4029 38979 4063
rect 40877 4029 40911 4063
rect 41337 4029 41371 4063
rect 42717 4029 42751 4063
rect 44925 4029 44959 4063
rect 46213 4029 46247 4063
rect 46949 4029 46983 4063
rect 48145 4029 48179 4063
rect 48421 4029 48455 4063
rect 49249 4029 49283 4063
rect 49433 4029 49467 4063
rect 50261 4029 50295 4063
rect 51733 4029 51767 4063
rect 51825 4029 51859 4063
rect 52837 4029 52871 4063
rect 53021 4029 53055 4063
rect 54125 4029 54159 4063
rect 54309 4029 54343 4063
rect 55229 4029 55263 4063
rect 55505 4029 55539 4063
rect 57253 4029 57287 4063
rect 4721 3961 4755 3995
rect 11253 3961 11287 3995
rect 15577 3961 15611 3995
rect 23673 3961 23707 3995
rect 27905 3961 27939 3995
rect 29653 3961 29687 3995
rect 30573 3961 30607 3995
rect 32137 3961 32171 3995
rect 40325 3961 40359 3995
rect 47317 3961 47351 3995
rect 49893 3961 49927 3995
rect 50813 3961 50847 3995
rect 53481 3961 53515 3995
rect 54953 3961 54987 3995
rect 1501 3893 1535 3927
rect 2881 3893 2915 3927
rect 11529 3893 11563 3927
rect 14749 3893 14783 3927
rect 22109 3893 22143 3927
rect 22845 3893 22879 3927
rect 24593 3893 24627 3927
rect 25513 3893 25547 3927
rect 26065 3893 26099 3927
rect 31493 3893 31527 3927
rect 32873 3893 32907 3927
rect 33609 3893 33643 3927
rect 34345 3893 34379 3927
rect 36829 3893 36863 3927
rect 39589 3893 39623 3927
rect 42165 3893 42199 3927
rect 45661 3893 45695 3927
rect 47593 3893 47627 3927
rect 51181 3893 51215 3927
rect 53573 3893 53607 3927
rect 57897 3893 57931 3927
rect 3249 3689 3283 3723
rect 3893 3689 3927 3723
rect 4997 3689 5031 3723
rect 9781 3689 9815 3723
rect 11437 3689 11471 3723
rect 14105 3689 14139 3723
rect 16405 3689 16439 3723
rect 16497 3689 16531 3723
rect 19349 3689 19383 3723
rect 21005 3689 21039 3723
rect 24225 3689 24259 3723
rect 27629 3689 27663 3723
rect 29745 3689 29779 3723
rect 32965 3689 32999 3723
rect 34437 3689 34471 3723
rect 39037 3689 39071 3723
rect 39313 3689 39347 3723
rect 40049 3689 40083 3723
rect 41797 3689 41831 3723
rect 42901 3689 42935 3723
rect 44557 3689 44591 3723
rect 46397 3689 46431 3723
rect 49341 3689 49375 3723
rect 53205 3689 53239 3723
rect 57713 3689 57747 3723
rect 9689 3621 9723 3655
rect 12449 3621 12483 3655
rect 17509 3621 17543 3655
rect 17693 3621 17727 3655
rect 49617 3621 49651 3655
rect 54677 3621 54711 3655
rect 54953 3621 54987 3655
rect 57621 3621 57655 3655
rect 3617 3553 3651 3587
rect 4537 3553 4571 3587
rect 5457 3553 5491 3587
rect 5641 3553 5675 3587
rect 7757 3553 7791 3587
rect 11805 3553 11839 3587
rect 11989 3553 12023 3587
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 15025 3553 15059 3587
rect 16957 3553 16991 3587
rect 17141 3553 17175 3587
rect 19073 3553 19107 3587
rect 39681 3553 39715 3587
rect 42349 3553 42383 3587
rect 42533 3553 42567 3587
rect 44281 3553 44315 3587
rect 45017 3553 45051 3587
rect 50813 3553 50847 3587
rect 53297 3553 53331 3587
rect 55413 3553 55447 3587
rect 56241 3553 56275 3587
rect 58173 3553 58207 3587
rect 58265 3553 58299 3587
rect 1593 3485 1627 3519
rect 1860 3485 1894 3519
rect 3433 3485 3467 3519
rect 4353 3485 4387 3519
rect 5365 3485 5399 3519
rect 5825 3485 5859 3519
rect 7297 3485 7331 3519
rect 9137 3485 9171 3519
rect 10894 3485 10928 3519
rect 11161 3485 11195 3519
rect 11621 3485 11655 3519
rect 12541 3485 12575 3519
rect 12808 3485 12842 3519
rect 14473 3485 14507 3519
rect 16865 3485 16899 3519
rect 18806 3485 18840 3519
rect 19533 3485 19567 3519
rect 19625 3485 19659 3519
rect 19892 3485 19926 3519
rect 22210 3485 22244 3519
rect 22477 3485 22511 3519
rect 22845 3485 22879 3519
rect 23112 3485 23146 3519
rect 24777 3485 24811 3519
rect 26249 3485 26283 3519
rect 26516 3485 26550 3519
rect 28457 3485 28491 3519
rect 28825 3485 28859 3519
rect 29561 3485 29595 3519
rect 29929 3485 29963 3519
rect 31585 3485 31619 3519
rect 33057 3485 33091 3519
rect 34713 3485 34747 3519
rect 36369 3485 36403 3519
rect 37657 3485 37691 3519
rect 37924 3485 37958 3519
rect 39129 3485 39163 3519
rect 39865 3485 39899 3519
rect 40417 3485 40451 3519
rect 40684 3485 40718 3519
rect 42257 3485 42291 3519
rect 44025 3485 44059 3519
rect 46489 3485 46523 3519
rect 47961 3485 47995 3519
rect 49801 3485 49835 3519
rect 50537 3485 50571 3519
rect 51825 3485 51859 3519
rect 53564 3485 53598 3519
rect 54769 3485 54803 3519
rect 55597 3485 55631 3519
rect 56508 3485 56542 3519
rect 58081 3485 58115 3519
rect 6070 3417 6104 3451
rect 15270 3417 15304 3451
rect 25022 3417 25056 3451
rect 29377 3417 29411 3451
rect 30174 3417 30208 3451
rect 31852 3417 31886 3451
rect 33324 3417 33358 3451
rect 34980 3417 35014 3451
rect 37105 3417 37139 3451
rect 45284 3417 45318 3451
rect 46756 3417 46790 3451
rect 48228 3417 48262 3451
rect 52092 3417 52126 3451
rect 2973 3349 3007 3383
rect 4261 3349 4295 3383
rect 7205 3349 7239 3383
rect 12081 3349 12115 3383
rect 13921 3349 13955 3383
rect 21097 3349 21131 3383
rect 24685 3349 24719 3383
rect 26157 3349 26191 3383
rect 27905 3349 27939 3383
rect 31309 3349 31343 3383
rect 36093 3349 36127 3383
rect 41889 3349 41923 3383
rect 47869 3349 47903 3383
rect 55689 3349 55723 3383
rect 56057 3349 56091 3383
rect 2789 3145 2823 3179
rect 4261 3145 4295 3179
rect 5457 3145 5491 3179
rect 7757 3145 7791 3179
rect 8217 3145 8251 3179
rect 11989 3145 12023 3179
rect 12173 3145 12207 3179
rect 14289 3145 14323 3179
rect 16405 3145 16439 3179
rect 16773 3145 16807 3179
rect 18061 3145 18095 3179
rect 20821 3145 20855 3179
rect 21833 3145 21867 3179
rect 22201 3145 22235 3179
rect 22937 3145 22971 3179
rect 25513 3145 25547 3179
rect 25973 3145 26007 3179
rect 26709 3145 26743 3179
rect 30389 3145 30423 3179
rect 30757 3145 30791 3179
rect 32505 3145 32539 3179
rect 32873 3145 32907 3179
rect 33333 3145 33367 3179
rect 36001 3145 36035 3179
rect 36277 3145 36311 3179
rect 37289 3145 37323 3179
rect 39405 3145 39439 3179
rect 40141 3145 40175 3179
rect 41797 3145 41831 3179
rect 42073 3145 42107 3179
rect 45385 3145 45419 3179
rect 47041 3145 47075 3179
rect 47409 3145 47443 3179
rect 49893 3145 49927 3179
rect 50997 3145 51031 3179
rect 56149 3145 56183 3179
rect 57897 3145 57931 3179
rect 1593 3077 1627 3111
rect 3126 3077 3160 3111
rect 5825 3077 5859 3111
rect 15516 3077 15550 3111
rect 18429 3077 18463 3111
rect 25881 3077 25915 3111
rect 29162 3077 29196 3111
rect 32413 3077 32447 3111
rect 33425 3077 33459 3111
rect 33885 3077 33919 3111
rect 34888 3077 34922 3111
rect 47593 3077 47627 3111
rect 48780 3077 48814 3111
rect 55137 3077 55171 3111
rect 56600 3077 56634 3111
rect 1961 3009 1995 3043
rect 2881 3009 2915 3043
rect 4445 3009 4479 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 6377 3009 6411 3043
rect 6644 3009 6678 3043
rect 8125 3009 8159 3043
rect 9330 3009 9364 3043
rect 9597 3009 9631 3043
rect 11089 3009 11123 3043
rect 11345 3009 11379 3043
rect 11805 3009 11839 3043
rect 13286 3009 13320 3043
rect 13553 3009 13587 3043
rect 15754 3009 15788 3043
rect 15945 3009 15979 3043
rect 16129 3009 16163 3043
rect 16957 3009 16991 3043
rect 17417 3009 17451 3043
rect 20085 3009 20119 3043
rect 22753 3009 22787 3043
rect 25053 3009 25087 3043
rect 26525 3009 26559 3043
rect 27353 3009 27387 3043
rect 28917 3009 28951 3043
rect 30849 3009 30883 3043
rect 31217 3009 31251 3043
rect 34621 3009 34655 3043
rect 36829 3009 36863 3043
rect 38025 3009 38059 3043
rect 38292 3009 38326 3043
rect 40417 3009 40451 3043
rect 40684 3009 40718 3043
rect 41889 3009 41923 3043
rect 42625 3009 42659 3043
rect 45109 3009 45143 3043
rect 46305 3009 46339 3043
rect 48520 3009 48554 3043
rect 50537 3009 50571 3043
rect 50813 3009 50847 3043
rect 51096 3009 51130 3043
rect 51356 3009 51390 3043
rect 53113 3009 53147 3043
rect 53205 3009 53239 3043
rect 53665 3009 53699 3043
rect 55965 3009 55999 3043
rect 56333 3009 56367 3043
rect 2145 2941 2179 2975
rect 4905 2941 4939 2975
rect 13737 2941 13771 2975
rect 17969 2941 18003 2975
rect 18521 2941 18555 2975
rect 18705 2941 18739 2975
rect 19073 2941 19107 2975
rect 21097 2941 21131 2975
rect 21649 2941 21683 2975
rect 22293 2941 22327 2975
rect 22477 2941 22511 2975
rect 23213 2941 23247 2975
rect 24041 2941 24075 2975
rect 26157 2941 26191 2975
rect 27629 2941 27663 2975
rect 30941 2941 30975 2975
rect 31861 2941 31895 2975
rect 32321 2941 32355 2975
rect 33149 2941 33183 2975
rect 34437 2941 34471 2975
rect 37841 2941 37875 2975
rect 39497 2941 39531 2975
rect 42901 2941 42935 2975
rect 44097 2941 44131 2975
rect 45937 2941 45971 2975
rect 46765 2941 46799 2975
rect 46949 2941 46983 2975
rect 48145 2941 48179 2975
rect 53021 2941 53055 2975
rect 54125 2941 54159 2975
rect 55689 2941 55723 2975
rect 58449 2941 58483 2975
rect 7941 2873 7975 2907
rect 14381 2873 14415 2907
rect 30297 2873 30331 2907
rect 33793 2873 33827 2907
rect 57713 2873 57747 2907
rect 4629 2805 4663 2839
rect 9965 2805 9999 2839
rect 23765 2805 23799 2839
rect 46489 2805 46523 2839
rect 49985 2805 50019 2839
rect 52469 2805 52503 2839
rect 53573 2805 53607 2839
rect 2145 2601 2179 2635
rect 2881 2601 2915 2635
rect 5273 2601 5307 2635
rect 6193 2601 6227 2635
rect 9873 2601 9907 2635
rect 12449 2601 12483 2635
rect 18889 2601 18923 2635
rect 20177 2601 20211 2635
rect 22109 2601 22143 2635
rect 24133 2601 24167 2635
rect 25329 2601 25363 2635
rect 27905 2601 27939 2635
rect 30389 2601 30423 2635
rect 34253 2601 34287 2635
rect 36185 2601 36219 2635
rect 39405 2601 39439 2635
rect 41337 2601 41371 2635
rect 43913 2601 43947 2635
rect 45201 2601 45235 2635
rect 47041 2601 47075 2635
rect 47409 2601 47443 2635
rect 49065 2601 49099 2635
rect 51641 2601 51675 2635
rect 54217 2601 54251 2635
rect 56885 2601 56919 2635
rect 6377 2533 6411 2567
rect 16773 2533 16807 2567
rect 3065 2465 3099 2499
rect 4261 2465 4295 2499
rect 6837 2465 6871 2499
rect 6929 2465 6963 2499
rect 13461 2465 13495 2499
rect 15577 2465 15611 2499
rect 17693 2465 17727 2499
rect 22661 2465 22695 2499
rect 28733 2465 28767 2499
rect 35173 2465 35207 2499
rect 37749 2465 37783 2499
rect 40325 2465 40359 2499
rect 41981 2465 42015 2499
rect 42901 2465 42935 2499
rect 50629 2465 50663 2499
rect 57437 2465 57471 2499
rect 58449 2465 58483 2499
rect 1593 2397 1627 2431
rect 2329 2397 2363 2431
rect 3801 2397 3835 2431
rect 5457 2397 5491 2431
rect 5641 2397 5675 2431
rect 7389 2397 7423 2431
rect 9321 2397 9355 2431
rect 11161 2397 11195 2431
rect 11897 2397 11931 2431
rect 13921 2397 13955 2431
rect 14473 2397 14507 2431
rect 15209 2397 15243 2431
rect 16957 2397 16991 2431
rect 17233 2397 17267 2431
rect 19073 2397 19107 2431
rect 19625 2397 19659 2431
rect 21465 2397 21499 2431
rect 21925 2397 21959 2431
rect 22201 2397 22235 2431
rect 23949 2397 23983 2431
rect 24777 2397 24811 2431
rect 26617 2397 26651 2431
rect 27353 2397 27387 2431
rect 28181 2397 28215 2431
rect 29837 2397 29871 2431
rect 31861 2397 31895 2431
rect 33333 2397 33367 2431
rect 33609 2397 33643 2431
rect 34805 2397 34839 2431
rect 36737 2397 36771 2431
rect 37289 2397 37323 2431
rect 38761 2397 38795 2431
rect 39865 2397 39899 2431
rect 42441 2397 42475 2431
rect 44465 2397 44499 2431
rect 45017 2397 45051 2431
rect 46673 2397 46707 2431
rect 46857 2397 46891 2431
rect 48789 2397 48823 2431
rect 49617 2397 49651 2431
rect 50169 2397 50203 2431
rect 52193 2397 52227 2431
rect 53941 2397 53975 2431
rect 54769 2397 54803 2431
rect 56701 2397 56735 2431
rect 57253 2397 57287 2431
rect 57345 2397 57379 2431
rect 6745 2329 6779 2363
rect 8585 2329 8619 2363
rect 10425 2329 10459 2363
rect 15025 2329 15059 2363
rect 20453 2329 20487 2363
rect 25605 2329 25639 2363
rect 30665 2329 30699 2363
rect 32321 2329 32355 2363
rect 45569 2329 45603 2363
rect 47777 2329 47811 2363
rect 52929 2329 52963 2363
rect 55505 2329 55539 2363
rect 3617 2261 3651 2295
rect 57897 2261 57931 2295
<< metal1 >>
rect 1104 27770 58880 27792
rect 1104 27718 8172 27770
rect 8224 27718 8236 27770
rect 8288 27718 8300 27770
rect 8352 27718 8364 27770
rect 8416 27718 8428 27770
rect 8480 27718 22616 27770
rect 22668 27718 22680 27770
rect 22732 27718 22744 27770
rect 22796 27718 22808 27770
rect 22860 27718 22872 27770
rect 22924 27718 37060 27770
rect 37112 27718 37124 27770
rect 37176 27718 37188 27770
rect 37240 27718 37252 27770
rect 37304 27718 37316 27770
rect 37368 27718 51504 27770
rect 51556 27718 51568 27770
rect 51620 27718 51632 27770
rect 51684 27718 51696 27770
rect 51748 27718 51760 27770
rect 51812 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 59040 27248
rect 1104 27174 15394 27226
rect 15446 27174 15458 27226
rect 15510 27174 15522 27226
rect 15574 27174 15586 27226
rect 15638 27174 15650 27226
rect 15702 27174 29838 27226
rect 29890 27174 29902 27226
rect 29954 27174 29966 27226
rect 30018 27174 30030 27226
rect 30082 27174 30094 27226
rect 30146 27174 44282 27226
rect 44334 27174 44346 27226
rect 44398 27174 44410 27226
rect 44462 27174 44474 27226
rect 44526 27174 44538 27226
rect 44590 27174 58726 27226
rect 58778 27174 58790 27226
rect 58842 27174 58854 27226
rect 58906 27174 58918 27226
rect 58970 27174 58982 27226
rect 59034 27174 59040 27226
rect 1104 27152 59040 27174
rect 1104 26682 58880 26704
rect 1104 26630 8172 26682
rect 8224 26630 8236 26682
rect 8288 26630 8300 26682
rect 8352 26630 8364 26682
rect 8416 26630 8428 26682
rect 8480 26630 22616 26682
rect 22668 26630 22680 26682
rect 22732 26630 22744 26682
rect 22796 26630 22808 26682
rect 22860 26630 22872 26682
rect 22924 26630 37060 26682
rect 37112 26630 37124 26682
rect 37176 26630 37188 26682
rect 37240 26630 37252 26682
rect 37304 26630 37316 26682
rect 37368 26630 51504 26682
rect 51556 26630 51568 26682
rect 51620 26630 51632 26682
rect 51684 26630 51696 26682
rect 51748 26630 51760 26682
rect 51812 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 59040 26160
rect 1104 26086 15394 26138
rect 15446 26086 15458 26138
rect 15510 26086 15522 26138
rect 15574 26086 15586 26138
rect 15638 26086 15650 26138
rect 15702 26086 29838 26138
rect 29890 26086 29902 26138
rect 29954 26086 29966 26138
rect 30018 26086 30030 26138
rect 30082 26086 30094 26138
rect 30146 26086 44282 26138
rect 44334 26086 44346 26138
rect 44398 26086 44410 26138
rect 44462 26086 44474 26138
rect 44526 26086 44538 26138
rect 44590 26086 58726 26138
rect 58778 26086 58790 26138
rect 58842 26086 58854 26138
rect 58906 26086 58918 26138
rect 58970 26086 58982 26138
rect 59034 26086 59040 26138
rect 1104 26064 59040 26086
rect 1104 25594 58880 25616
rect 1104 25542 8172 25594
rect 8224 25542 8236 25594
rect 8288 25542 8300 25594
rect 8352 25542 8364 25594
rect 8416 25542 8428 25594
rect 8480 25542 22616 25594
rect 22668 25542 22680 25594
rect 22732 25542 22744 25594
rect 22796 25542 22808 25594
rect 22860 25542 22872 25594
rect 22924 25542 37060 25594
rect 37112 25542 37124 25594
rect 37176 25542 37188 25594
rect 37240 25542 37252 25594
rect 37304 25542 37316 25594
rect 37368 25542 51504 25594
rect 51556 25542 51568 25594
rect 51620 25542 51632 25594
rect 51684 25542 51696 25594
rect 51748 25542 51760 25594
rect 51812 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 59040 25072
rect 1104 24998 15394 25050
rect 15446 24998 15458 25050
rect 15510 24998 15522 25050
rect 15574 24998 15586 25050
rect 15638 24998 15650 25050
rect 15702 24998 29838 25050
rect 29890 24998 29902 25050
rect 29954 24998 29966 25050
rect 30018 24998 30030 25050
rect 30082 24998 30094 25050
rect 30146 24998 44282 25050
rect 44334 24998 44346 25050
rect 44398 24998 44410 25050
rect 44462 24998 44474 25050
rect 44526 24998 44538 25050
rect 44590 24998 58726 25050
rect 58778 24998 58790 25050
rect 58842 24998 58854 25050
rect 58906 24998 58918 25050
rect 58970 24998 58982 25050
rect 59034 24998 59040 25050
rect 1104 24976 59040 24998
rect 1104 24506 58880 24528
rect 1104 24454 8172 24506
rect 8224 24454 8236 24506
rect 8288 24454 8300 24506
rect 8352 24454 8364 24506
rect 8416 24454 8428 24506
rect 8480 24454 22616 24506
rect 22668 24454 22680 24506
rect 22732 24454 22744 24506
rect 22796 24454 22808 24506
rect 22860 24454 22872 24506
rect 22924 24454 37060 24506
rect 37112 24454 37124 24506
rect 37176 24454 37188 24506
rect 37240 24454 37252 24506
rect 37304 24454 37316 24506
rect 37368 24454 51504 24506
rect 51556 24454 51568 24506
rect 51620 24454 51632 24506
rect 51684 24454 51696 24506
rect 51748 24454 51760 24506
rect 51812 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 59040 23984
rect 1104 23910 15394 23962
rect 15446 23910 15458 23962
rect 15510 23910 15522 23962
rect 15574 23910 15586 23962
rect 15638 23910 15650 23962
rect 15702 23910 29838 23962
rect 29890 23910 29902 23962
rect 29954 23910 29966 23962
rect 30018 23910 30030 23962
rect 30082 23910 30094 23962
rect 30146 23910 44282 23962
rect 44334 23910 44346 23962
rect 44398 23910 44410 23962
rect 44462 23910 44474 23962
rect 44526 23910 44538 23962
rect 44590 23910 58726 23962
rect 58778 23910 58790 23962
rect 58842 23910 58854 23962
rect 58906 23910 58918 23962
rect 58970 23910 58982 23962
rect 59034 23910 59040 23962
rect 1104 23888 59040 23910
rect 15194 23604 15200 23656
rect 15252 23604 15258 23656
rect 15286 23604 15292 23656
rect 15344 23604 15350 23656
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 18138 23644 18144 23656
rect 18095 23616 18144 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 18230 23604 18236 23656
rect 18288 23604 18294 23656
rect 47578 23604 47584 23656
rect 47636 23604 47642 23656
rect 53282 23604 53288 23656
rect 53340 23604 53346 23656
rect 54018 23604 54024 23656
rect 54076 23604 54082 23656
rect 54478 23576 54484 23588
rect 52472 23548 54484 23576
rect 14550 23468 14556 23520
rect 14608 23468 14614 23520
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 16206 23508 16212 23520
rect 15979 23480 16212 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 17402 23468 17408 23520
rect 17460 23468 17466 23520
rect 18874 23468 18880 23520
rect 18932 23468 18938 23520
rect 46842 23468 46848 23520
rect 46900 23468 46906 23520
rect 47397 23511 47455 23517
rect 47397 23477 47409 23511
rect 47443 23508 47455 23511
rect 48130 23508 48136 23520
rect 47443 23480 48136 23508
rect 47443 23477 47455 23480
rect 47397 23471 47455 23477
rect 48130 23468 48136 23480
rect 48188 23468 48194 23520
rect 48222 23468 48228 23520
rect 48280 23468 48286 23520
rect 49326 23468 49332 23520
rect 49384 23508 49390 23520
rect 52472 23517 52500 23548
rect 54478 23536 54484 23548
rect 54536 23536 54542 23588
rect 52457 23511 52515 23517
rect 52457 23508 52469 23511
rect 49384 23480 52469 23508
rect 49384 23468 49390 23480
rect 52457 23477 52469 23480
rect 52503 23477 52515 23511
rect 52457 23471 52515 23477
rect 52730 23468 52736 23520
rect 52788 23468 52794 23520
rect 53466 23468 53472 23520
rect 53524 23468 53530 23520
rect 1104 23418 58880 23440
rect 1104 23366 8172 23418
rect 8224 23366 8236 23418
rect 8288 23366 8300 23418
rect 8352 23366 8364 23418
rect 8416 23366 8428 23418
rect 8480 23366 22616 23418
rect 22668 23366 22680 23418
rect 22732 23366 22744 23418
rect 22796 23366 22808 23418
rect 22860 23366 22872 23418
rect 22924 23366 37060 23418
rect 37112 23366 37124 23418
rect 37176 23366 37188 23418
rect 37240 23366 37252 23418
rect 37304 23366 37316 23418
rect 37368 23366 51504 23418
rect 51556 23366 51568 23418
rect 51620 23366 51632 23418
rect 51684 23366 51696 23418
rect 51748 23366 51760 23418
rect 51812 23366 58880 23418
rect 1104 23344 58880 23366
rect 17773 23307 17831 23313
rect 15120 23276 17724 23304
rect 15120 23180 15148 23276
rect 15473 23239 15531 23245
rect 15473 23205 15485 23239
rect 15519 23236 15531 23239
rect 17696 23236 17724 23276
rect 17773 23273 17785 23307
rect 17819 23304 17831 23307
rect 18230 23304 18236 23316
rect 17819 23276 18236 23304
rect 17819 23273 17831 23276
rect 17773 23267 17831 23273
rect 18230 23264 18236 23276
rect 18288 23264 18294 23316
rect 42518 23264 42524 23316
rect 42576 23304 42582 23316
rect 46842 23304 46848 23316
rect 42576 23276 46848 23304
rect 42576 23264 42582 23276
rect 46842 23264 46848 23276
rect 46900 23304 46906 23316
rect 52546 23304 52552 23316
rect 46900 23276 52552 23304
rect 46900 23264 46906 23276
rect 19613 23239 19671 23245
rect 19613 23236 19625 23239
rect 15519 23208 15608 23236
rect 17696 23208 19625 23236
rect 15519 23205 15531 23208
rect 15473 23199 15531 23205
rect 15102 23128 15108 23180
rect 15160 23128 15166 23180
rect 15580 23177 15608 23208
rect 19613 23205 19625 23208
rect 19659 23236 19671 23239
rect 20438 23236 20444 23248
rect 19659 23208 20444 23236
rect 19659 23205 19671 23208
rect 19613 23199 19671 23205
rect 20438 23196 20444 23208
rect 20496 23196 20502 23248
rect 46937 23239 46995 23245
rect 46937 23205 46949 23239
rect 46983 23205 46995 23239
rect 46937 23199 46995 23205
rect 15565 23171 15623 23177
rect 15565 23137 15577 23171
rect 15611 23137 15623 23171
rect 15565 23131 15623 23137
rect 46845 23171 46903 23177
rect 46845 23137 46857 23171
rect 46891 23168 46903 23171
rect 46952 23168 46980 23199
rect 46891 23140 46980 23168
rect 47581 23171 47639 23177
rect 46891 23137 46903 23140
rect 46845 23131 46903 23137
rect 47581 23137 47593 23171
rect 47627 23168 47639 23171
rect 47688 23168 47716 23276
rect 52546 23264 52552 23276
rect 52604 23264 52610 23316
rect 53285 23307 53343 23313
rect 53285 23273 53297 23307
rect 53331 23304 53343 23307
rect 54018 23304 54024 23316
rect 53331 23276 54024 23304
rect 53331 23273 53343 23276
rect 53285 23267 53343 23273
rect 54018 23264 54024 23276
rect 54076 23264 54082 23316
rect 47765 23239 47823 23245
rect 47765 23205 47777 23239
rect 47811 23236 47823 23239
rect 48590 23236 48596 23248
rect 47811 23208 48596 23236
rect 47811 23205 47823 23208
rect 47765 23199 47823 23205
rect 48590 23196 48596 23208
rect 48648 23196 48654 23248
rect 49973 23239 50031 23245
rect 49973 23205 49985 23239
rect 50019 23236 50031 23239
rect 55033 23239 55091 23245
rect 50019 23208 50752 23236
rect 50019 23205 50031 23208
rect 49973 23199 50031 23205
rect 47627 23140 47716 23168
rect 47627 23137 47639 23140
rect 47581 23131 47639 23137
rect 48130 23128 48136 23180
rect 48188 23168 48194 23180
rect 50724 23177 50752 23208
rect 55033 23205 55045 23239
rect 55079 23236 55091 23239
rect 55079 23208 55214 23236
rect 55079 23205 55091 23208
rect 55033 23199 55091 23205
rect 48317 23171 48375 23177
rect 48317 23168 48329 23171
rect 48188 23140 48329 23168
rect 48188 23128 48194 23140
rect 48317 23137 48329 23140
rect 48363 23137 48375 23171
rect 50709 23171 50767 23177
rect 48317 23131 48375 23137
rect 48516 23140 48728 23168
rect 6638 23060 6644 23112
rect 6696 23060 6702 23112
rect 12066 23060 12072 23112
rect 12124 23060 12130 23112
rect 14090 23060 14096 23112
rect 14148 23100 14154 23112
rect 16393 23103 16451 23109
rect 16393 23100 16405 23103
rect 14148 23072 16405 23100
rect 14148 23060 14154 23072
rect 16393 23069 16405 23072
rect 16439 23069 16451 23103
rect 16393 23063 16451 23069
rect 16660 23103 16718 23109
rect 16660 23069 16672 23103
rect 16706 23100 16718 23103
rect 17402 23100 17408 23112
rect 16706 23072 17408 23100
rect 16706 23069 16718 23072
rect 16660 23063 16718 23069
rect 14366 23041 14372 23044
rect 14360 22995 14372 23041
rect 14366 22992 14372 22995
rect 14424 22992 14430 23044
rect 16408 23032 16436 23063
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 17954 23060 17960 23112
rect 18012 23100 18018 23112
rect 18601 23103 18659 23109
rect 18601 23100 18613 23103
rect 18012 23072 18613 23100
rect 18012 23060 18018 23072
rect 18601 23069 18613 23072
rect 18647 23069 18659 23103
rect 18601 23063 18659 23069
rect 20346 23060 20352 23112
rect 20404 23060 20410 23112
rect 22278 23060 22284 23112
rect 22336 23100 22342 23112
rect 22741 23103 22799 23109
rect 22741 23100 22753 23103
rect 22336 23072 22753 23100
rect 22336 23060 22342 23072
rect 22741 23069 22753 23072
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 23566 23060 23572 23112
rect 23624 23060 23630 23112
rect 34054 23060 34060 23112
rect 34112 23060 34118 23112
rect 36446 23060 36452 23112
rect 36504 23060 36510 23112
rect 40402 23060 40408 23112
rect 40460 23060 40466 23112
rect 45554 23060 45560 23112
rect 45612 23060 45618 23112
rect 48148 23100 48176 23128
rect 45664 23072 48176 23100
rect 48225 23103 48283 23109
rect 16758 23032 16764 23044
rect 16408 23004 16764 23032
rect 16758 22992 16764 23004
rect 16816 23032 16822 23044
rect 16816 23004 19288 23032
rect 16816 22992 16822 23004
rect 19260 22976 19288 23004
rect 35802 22992 35808 23044
rect 35860 23032 35866 23044
rect 36817 23035 36875 23041
rect 36817 23032 36829 23035
rect 35860 23004 36829 23032
rect 35860 22992 35866 23004
rect 36817 23001 36829 23004
rect 36863 23001 36875 23035
rect 36817 22995 36875 23001
rect 42702 22992 42708 23044
rect 42760 23032 42766 23044
rect 45664 23032 45692 23072
rect 48225 23069 48237 23103
rect 48271 23100 48283 23103
rect 48516 23100 48544 23140
rect 48271 23072 48544 23100
rect 48593 23103 48651 23109
rect 48271 23069 48283 23072
rect 48225 23063 48283 23069
rect 48593 23069 48605 23103
rect 48639 23069 48651 23103
rect 48700 23100 48728 23140
rect 50709 23137 50721 23171
rect 50755 23137 50767 23171
rect 55186 23168 55214 23208
rect 55861 23171 55919 23177
rect 55861 23168 55873 23171
rect 55186 23140 55873 23168
rect 50709 23131 50767 23137
rect 55861 23137 55873 23140
rect 55907 23137 55919 23171
rect 55861 23131 55919 23137
rect 49142 23100 49148 23112
rect 48700 23072 49148 23100
rect 48593 23063 48651 23069
rect 42760 23004 45692 23032
rect 47305 23035 47363 23041
rect 42760 22992 42766 23004
rect 47305 23001 47317 23035
rect 47351 23032 47363 23035
rect 47351 23004 48268 23032
rect 47351 23001 47363 23004
rect 47305 22995 47363 23001
rect 48240 22976 48268 23004
rect 6086 22924 6092 22976
rect 6144 22924 6150 22976
rect 11054 22924 11060 22976
rect 11112 22964 11118 22976
rect 11517 22967 11575 22973
rect 11517 22964 11529 22967
rect 11112 22936 11529 22964
rect 11112 22924 11118 22936
rect 11517 22933 11529 22936
rect 11563 22933 11575 22967
rect 11517 22927 11575 22933
rect 16209 22967 16267 22973
rect 16209 22933 16221 22967
rect 16255 22964 16267 22967
rect 16298 22964 16304 22976
rect 16255 22936 16304 22964
rect 16255 22933 16267 22936
rect 16209 22927 16267 22933
rect 16298 22924 16304 22936
rect 16356 22924 16362 22976
rect 18046 22924 18052 22976
rect 18104 22924 18110 22976
rect 19242 22924 19248 22976
rect 19300 22924 19306 22976
rect 19794 22924 19800 22976
rect 19852 22924 19858 22976
rect 22186 22924 22192 22976
rect 22244 22924 22250 22976
rect 23017 22967 23075 22973
rect 23017 22933 23029 22967
rect 23063 22964 23075 22967
rect 23198 22964 23204 22976
rect 23063 22936 23204 22964
rect 23063 22933 23075 22936
rect 23017 22927 23075 22933
rect 23198 22924 23204 22936
rect 23256 22924 23262 22976
rect 33410 22924 33416 22976
rect 33468 22924 33474 22976
rect 34238 22924 34244 22976
rect 34296 22964 34302 22976
rect 34333 22967 34391 22973
rect 34333 22964 34345 22967
rect 34296 22936 34345 22964
rect 34296 22924 34302 22936
rect 34333 22933 34345 22936
rect 34379 22933 34391 22967
rect 34333 22927 34391 22933
rect 35897 22967 35955 22973
rect 35897 22933 35909 22967
rect 35943 22964 35955 22967
rect 35986 22964 35992 22976
rect 35943 22936 35992 22964
rect 35943 22933 35955 22936
rect 35897 22927 35955 22933
rect 35986 22924 35992 22936
rect 36044 22924 36050 22976
rect 39850 22924 39856 22976
rect 39908 22924 39914 22976
rect 45002 22924 45008 22976
rect 45060 22924 45066 22976
rect 46198 22924 46204 22976
rect 46256 22924 46262 22976
rect 47397 22967 47455 22973
rect 47397 22933 47409 22967
rect 47443 22964 47455 22967
rect 48038 22964 48044 22976
rect 47443 22936 48044 22964
rect 47443 22933 47455 22936
rect 47397 22927 47455 22933
rect 48038 22924 48044 22936
rect 48096 22964 48102 22976
rect 48133 22967 48191 22973
rect 48133 22964 48145 22967
rect 48096 22936 48145 22964
rect 48096 22924 48102 22936
rect 48133 22933 48145 22936
rect 48179 22933 48191 22967
rect 48133 22927 48191 22933
rect 48222 22924 48228 22976
rect 48280 22924 48286 22976
rect 48608 22964 48636 23063
rect 49142 23060 49148 23072
rect 49200 23060 49206 23112
rect 51534 23060 51540 23112
rect 51592 23060 51598 23112
rect 51902 23060 51908 23112
rect 51960 23100 51966 23112
rect 53653 23103 53711 23109
rect 53653 23100 53665 23103
rect 51960 23072 53665 23100
rect 51960 23060 51966 23072
rect 53653 23069 53665 23072
rect 53699 23100 53711 23103
rect 55214 23100 55220 23112
rect 53699 23072 55220 23100
rect 53699 23069 53711 23072
rect 53653 23063 53711 23069
rect 55214 23060 55220 23072
rect 55272 23060 55278 23112
rect 56594 23060 56600 23112
rect 56652 23060 56658 23112
rect 48860 23035 48918 23041
rect 48860 23001 48872 23035
rect 48906 23032 48918 23035
rect 49050 23032 49056 23044
rect 48906 23004 49056 23032
rect 48906 23001 48918 23004
rect 48860 22995 48918 23001
rect 49050 22992 49056 23004
rect 49108 22992 49114 23044
rect 52172 23035 52230 23041
rect 52172 23001 52184 23035
rect 52218 23032 52230 23035
rect 52730 23032 52736 23044
rect 52218 23004 52736 23032
rect 52218 23001 52230 23004
rect 52172 22995 52230 23001
rect 52730 22992 52736 23004
rect 52788 22992 52794 23044
rect 53920 23035 53978 23041
rect 53920 23001 53932 23035
rect 53966 23032 53978 23035
rect 54202 23032 54208 23044
rect 53966 23004 54208 23032
rect 53966 23001 53978 23004
rect 53920 22995 53978 23001
rect 54202 22992 54208 23004
rect 54260 22992 54266 23044
rect 49970 22964 49976 22976
rect 48608 22936 49976 22964
rect 49970 22924 49976 22936
rect 50028 22924 50034 22976
rect 50062 22924 50068 22976
rect 50120 22964 50126 22976
rect 50157 22967 50215 22973
rect 50157 22964 50169 22967
rect 50120 22936 50169 22964
rect 50120 22924 50126 22936
rect 50157 22933 50169 22936
rect 50203 22933 50215 22967
rect 50157 22927 50215 22933
rect 50246 22924 50252 22976
rect 50304 22964 50310 22976
rect 50893 22967 50951 22973
rect 50893 22964 50905 22967
rect 50304 22936 50905 22964
rect 50304 22924 50310 22936
rect 50893 22933 50905 22936
rect 50939 22933 50951 22967
rect 50893 22927 50951 22933
rect 55122 22924 55128 22976
rect 55180 22964 55186 22976
rect 55309 22967 55367 22973
rect 55309 22964 55321 22967
rect 55180 22936 55321 22964
rect 55180 22924 55186 22936
rect 55309 22933 55321 22936
rect 55355 22933 55367 22967
rect 55309 22927 55367 22933
rect 56042 22924 56048 22976
rect 56100 22924 56106 22976
rect 1104 22874 59040 22896
rect 1104 22822 15394 22874
rect 15446 22822 15458 22874
rect 15510 22822 15522 22874
rect 15574 22822 15586 22874
rect 15638 22822 15650 22874
rect 15702 22822 29838 22874
rect 29890 22822 29902 22874
rect 29954 22822 29966 22874
rect 30018 22822 30030 22874
rect 30082 22822 30094 22874
rect 30146 22822 44282 22874
rect 44334 22822 44346 22874
rect 44398 22822 44410 22874
rect 44462 22822 44474 22874
rect 44526 22822 44538 22874
rect 44590 22822 58726 22874
rect 58778 22822 58790 22874
rect 58842 22822 58854 22874
rect 58906 22822 58918 22874
rect 58970 22822 58982 22874
rect 59034 22822 59040 22874
rect 1104 22800 59040 22822
rect 12158 22720 12164 22772
rect 12216 22760 12222 22772
rect 12989 22763 13047 22769
rect 12989 22760 13001 22763
rect 12216 22732 13001 22760
rect 12216 22720 12222 22732
rect 12989 22729 13001 22732
rect 13035 22760 13047 22763
rect 15105 22763 15163 22769
rect 13035 22732 14688 22760
rect 13035 22729 13047 22732
rect 12989 22723 13047 22729
rect 14090 22692 14096 22704
rect 13648 22664 14096 22692
rect 13648 22636 13676 22664
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 14550 22652 14556 22704
rect 14608 22652 14614 22704
rect 14660 22692 14688 22732
rect 15105 22729 15117 22763
rect 15151 22760 15163 22763
rect 15194 22760 15200 22772
rect 15151 22732 15200 22760
rect 15151 22729 15163 22732
rect 15105 22723 15163 22729
rect 15194 22720 15200 22732
rect 15252 22720 15258 22772
rect 15565 22763 15623 22769
rect 15565 22729 15577 22763
rect 15611 22760 15623 22763
rect 17126 22760 17132 22772
rect 15611 22732 17132 22760
rect 15611 22729 15623 22732
rect 15565 22723 15623 22729
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18049 22763 18107 22769
rect 18049 22760 18061 22763
rect 18012 22732 18061 22760
rect 18012 22720 18018 22732
rect 18049 22729 18061 22732
rect 18095 22729 18107 22763
rect 18049 22723 18107 22729
rect 18138 22720 18144 22772
rect 18196 22720 18202 22772
rect 18601 22763 18659 22769
rect 18601 22729 18613 22763
rect 18647 22760 18659 22763
rect 18874 22760 18880 22772
rect 18647 22732 18880 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 19889 22763 19947 22769
rect 19889 22729 19901 22763
rect 19935 22760 19947 22763
rect 20346 22760 20352 22772
rect 19935 22732 20352 22760
rect 19935 22729 19947 22732
rect 19889 22723 19947 22729
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 22186 22720 22192 22772
rect 22244 22720 22250 22772
rect 23201 22763 23259 22769
rect 23201 22729 23213 22763
rect 23247 22760 23259 22763
rect 23566 22760 23572 22772
rect 23247 22732 23572 22760
rect 23247 22729 23259 22732
rect 23201 22723 23259 22729
rect 23566 22720 23572 22732
rect 23624 22720 23630 22772
rect 36081 22763 36139 22769
rect 36081 22729 36093 22763
rect 36127 22760 36139 22763
rect 36446 22760 36452 22772
rect 36127 22732 36452 22760
rect 36127 22729 36139 22732
rect 36081 22723 36139 22729
rect 36446 22720 36452 22732
rect 36504 22720 36510 22772
rect 36541 22763 36599 22769
rect 36541 22729 36553 22763
rect 36587 22760 36599 22763
rect 37921 22763 37979 22769
rect 37921 22760 37933 22763
rect 36587 22732 37933 22760
rect 36587 22729 36599 22732
rect 36541 22723 36599 22729
rect 37921 22729 37933 22732
rect 37967 22760 37979 22763
rect 38654 22760 38660 22772
rect 37967 22732 38660 22760
rect 37967 22729 37979 22732
rect 37921 22723 37979 22729
rect 38654 22720 38660 22732
rect 38712 22720 38718 22772
rect 39850 22720 39856 22772
rect 39908 22720 39914 22772
rect 46198 22720 46204 22772
rect 46256 22720 46262 22772
rect 47397 22763 47455 22769
rect 47397 22729 47409 22763
rect 47443 22760 47455 22763
rect 47578 22760 47584 22772
rect 47443 22732 47584 22760
rect 47443 22729 47455 22732
rect 47397 22723 47455 22729
rect 47578 22720 47584 22732
rect 47636 22720 47642 22772
rect 48130 22720 48136 22772
rect 48188 22760 48194 22772
rect 48188 22732 51304 22760
rect 48188 22720 48194 22732
rect 14660 22664 15608 22692
rect 13630 22584 13636 22636
rect 13688 22584 13694 22636
rect 13900 22627 13958 22633
rect 13900 22593 13912 22627
rect 13946 22624 13958 22627
rect 14568 22624 14596 22652
rect 13946 22596 14596 22624
rect 13946 22593 13958 22596
rect 13900 22587 13958 22593
rect 15470 22584 15476 22636
rect 15528 22584 15534 22636
rect 15580 22624 15608 22664
rect 16758 22652 16764 22704
rect 16816 22652 16822 22704
rect 21361 22695 21419 22701
rect 21361 22692 21373 22695
rect 20180 22664 21373 22692
rect 16669 22627 16727 22633
rect 15580 22596 16620 22624
rect 3694 22516 3700 22568
rect 3752 22516 3758 22568
rect 4430 22516 4436 22568
rect 4488 22516 4494 22568
rect 7098 22516 7104 22568
rect 7156 22516 7162 22568
rect 9766 22516 9772 22568
rect 9824 22516 9830 22568
rect 10042 22516 10048 22568
rect 10100 22516 10106 22568
rect 10686 22516 10692 22568
rect 10744 22516 10750 22568
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 15286 22516 15292 22568
rect 15344 22516 15350 22568
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22556 15807 22559
rect 16114 22556 16120 22568
rect 15795 22528 16120 22556
rect 15795 22525 15807 22528
rect 15749 22519 15807 22525
rect 16114 22516 16120 22528
rect 16172 22516 16178 22568
rect 4890 22448 4896 22500
rect 4948 22488 4954 22500
rect 9950 22488 9956 22500
rect 4948 22460 9956 22488
rect 4948 22448 4954 22460
rect 9950 22448 9956 22460
rect 10008 22448 10014 22500
rect 15013 22491 15071 22497
rect 10152 22460 13676 22488
rect 10152 22432 10180 22460
rect 3050 22380 3056 22432
rect 3108 22380 3114 22432
rect 3878 22380 3884 22432
rect 3936 22380 3942 22432
rect 5718 22380 5724 22432
rect 5776 22420 5782 22432
rect 6457 22423 6515 22429
rect 6457 22420 6469 22423
rect 5776 22392 6469 22420
rect 5776 22380 5782 22392
rect 6457 22389 6469 22392
rect 6503 22389 6515 22423
rect 6457 22383 6515 22389
rect 9214 22380 9220 22432
rect 9272 22380 9278 22432
rect 10134 22380 10140 22432
rect 10192 22380 10198 22432
rect 10597 22423 10655 22429
rect 10597 22389 10609 22423
rect 10643 22420 10655 22423
rect 10870 22420 10876 22432
rect 10643 22392 10876 22420
rect 10643 22389 10655 22392
rect 10597 22383 10655 22389
rect 10870 22380 10876 22392
rect 10928 22380 10934 22432
rect 11330 22380 11336 22432
rect 11388 22380 11394 22432
rect 12618 22380 12624 22432
rect 12676 22380 12682 22432
rect 13648 22420 13676 22460
rect 15013 22457 15025 22491
rect 15059 22488 15071 22491
rect 15304 22488 15332 22516
rect 16592 22500 16620 22596
rect 16669 22593 16681 22627
rect 16715 22624 16727 22627
rect 16776 22624 16804 22652
rect 16715 22596 16804 22624
rect 16936 22627 16994 22633
rect 16715 22593 16727 22596
rect 16669 22587 16727 22593
rect 16936 22593 16948 22627
rect 16982 22624 16994 22627
rect 16982 22596 17908 22624
rect 16982 22593 16994 22596
rect 16936 22587 16994 22593
rect 15059 22460 15332 22488
rect 15059 22457 15071 22460
rect 15013 22451 15071 22457
rect 16574 22448 16580 22500
rect 16632 22448 16638 22500
rect 17880 22488 17908 22596
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18012 22596 18521 22624
rect 18012 22584 18018 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 18690 22516 18696 22568
rect 18748 22516 18754 22568
rect 19518 22516 19524 22568
rect 19576 22516 19582 22568
rect 20180 22556 20208 22664
rect 21361 22661 21373 22664
rect 21407 22661 21419 22695
rect 21361 22655 21419 22661
rect 22088 22695 22146 22701
rect 22088 22661 22100 22695
rect 22134 22692 22146 22695
rect 22204 22692 22232 22720
rect 22134 22664 22232 22692
rect 22134 22661 22146 22664
rect 22088 22655 22146 22661
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22624 20315 22627
rect 20622 22624 20628 22636
rect 20303 22596 20628 22624
rect 20303 22593 20315 22596
rect 20257 22587 20315 22593
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 21376 22624 21404 22655
rect 32030 22652 32036 22704
rect 32088 22692 32094 22704
rect 35989 22695 36047 22701
rect 35989 22692 36001 22695
rect 32088 22664 36001 22692
rect 32088 22652 32094 22664
rect 35989 22661 36001 22664
rect 36035 22692 36047 22695
rect 38832 22695 38890 22701
rect 36035 22664 36768 22692
rect 36035 22661 36047 22664
rect 35989 22655 36047 22661
rect 22370 22624 22376 22636
rect 21376 22596 22376 22624
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 33413 22627 33471 22633
rect 33413 22593 33425 22627
rect 33459 22624 33471 22627
rect 33778 22624 33784 22636
rect 33459 22596 33784 22624
rect 33459 22593 33471 22596
rect 33413 22587 33471 22593
rect 33778 22584 33784 22596
rect 33836 22624 33842 22636
rect 33873 22627 33931 22633
rect 33873 22624 33885 22627
rect 33836 22596 33885 22624
rect 33836 22584 33842 22596
rect 33873 22593 33885 22596
rect 33919 22593 33931 22627
rect 33873 22587 33931 22593
rect 34330 22584 34336 22636
rect 34388 22624 34394 22636
rect 35161 22627 35219 22633
rect 35161 22624 35173 22627
rect 34388 22596 35173 22624
rect 34388 22584 34394 22596
rect 35161 22593 35173 22596
rect 35207 22593 35219 22627
rect 35161 22587 35219 22593
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 36740 22624 36768 22664
rect 38832 22661 38844 22695
rect 38878 22692 38890 22695
rect 39868 22692 39896 22720
rect 38878 22664 39896 22692
rect 43824 22664 46060 22692
rect 38878 22661 38890 22664
rect 38832 22655 38890 22661
rect 36740 22596 42748 22624
rect 20349 22559 20407 22565
rect 20349 22556 20361 22559
rect 20180 22528 20361 22556
rect 20349 22525 20361 22528
rect 20395 22525 20407 22559
rect 20349 22519 20407 22525
rect 20438 22516 20444 22568
rect 20496 22556 20502 22568
rect 20496 22528 20576 22556
rect 20496 22516 20502 22528
rect 18969 22491 19027 22497
rect 18969 22488 18981 22491
rect 17880 22460 18981 22488
rect 18969 22457 18981 22460
rect 19015 22457 19027 22491
rect 18969 22451 19027 22457
rect 13814 22420 13820 22432
rect 13648 22392 13820 22420
rect 13814 22380 13820 22392
rect 13872 22380 13878 22432
rect 20548 22420 20576 22528
rect 20714 22516 20720 22568
rect 20772 22516 20778 22568
rect 21821 22559 21879 22565
rect 21821 22525 21833 22559
rect 21867 22525 21879 22559
rect 21821 22519 21879 22525
rect 20806 22448 20812 22500
rect 20864 22488 20870 22500
rect 21836 22488 21864 22519
rect 23382 22516 23388 22568
rect 23440 22556 23446 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23440 22528 23857 22556
rect 23440 22516 23446 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 23845 22519 23903 22525
rect 26326 22516 26332 22568
rect 26384 22516 26390 22568
rect 27890 22516 27896 22568
rect 27948 22556 27954 22568
rect 28445 22559 28503 22565
rect 28445 22556 28457 22559
rect 27948 22528 28457 22556
rect 27948 22516 27954 22528
rect 28445 22525 28457 22528
rect 28491 22525 28503 22559
rect 28445 22519 28503 22525
rect 29178 22516 29184 22568
rect 29236 22516 29242 22568
rect 31570 22516 31576 22568
rect 31628 22516 31634 22568
rect 31662 22516 31668 22568
rect 31720 22556 31726 22568
rect 32125 22559 32183 22565
rect 32125 22556 32137 22559
rect 31720 22528 32137 22556
rect 31720 22516 31726 22528
rect 32125 22525 32137 22528
rect 32171 22525 32183 22559
rect 32125 22519 32183 22525
rect 33229 22559 33287 22565
rect 33229 22525 33241 22559
rect 33275 22525 33287 22559
rect 33229 22519 33287 22525
rect 24854 22488 24860 22500
rect 20864 22460 21864 22488
rect 23216 22460 24860 22488
rect 20864 22448 20870 22460
rect 23216 22420 23244 22460
rect 24854 22448 24860 22460
rect 24912 22448 24918 22500
rect 26786 22448 26792 22500
rect 26844 22488 26850 22500
rect 26844 22460 28212 22488
rect 26844 22448 26850 22460
rect 28184 22432 28212 22460
rect 20548 22392 23244 22420
rect 23290 22380 23296 22432
rect 23348 22380 23354 22432
rect 25590 22380 25596 22432
rect 25648 22420 25654 22432
rect 25777 22423 25835 22429
rect 25777 22420 25789 22423
rect 25648 22392 25789 22420
rect 25648 22380 25654 22392
rect 25777 22389 25789 22392
rect 25823 22389 25835 22423
rect 25777 22383 25835 22389
rect 27249 22423 27307 22429
rect 27249 22389 27261 22423
rect 27295 22420 27307 22423
rect 27706 22420 27712 22432
rect 27295 22392 27712 22420
rect 27295 22389 27307 22392
rect 27249 22383 27307 22389
rect 27706 22380 27712 22392
rect 27764 22380 27770 22432
rect 27798 22380 27804 22432
rect 27856 22420 27862 22432
rect 27893 22423 27951 22429
rect 27893 22420 27905 22423
rect 27856 22392 27905 22420
rect 27856 22380 27862 22392
rect 27893 22389 27905 22392
rect 27939 22389 27951 22423
rect 27893 22383 27951 22389
rect 28166 22380 28172 22432
rect 28224 22380 28230 22432
rect 28626 22380 28632 22432
rect 28684 22380 28690 22432
rect 30558 22380 30564 22432
rect 30616 22380 30622 22432
rect 31018 22380 31024 22432
rect 31076 22380 31082 22432
rect 32769 22423 32827 22429
rect 32769 22389 32781 22423
rect 32815 22420 32827 22423
rect 33042 22420 33048 22432
rect 32815 22392 33048 22420
rect 32815 22389 32827 22392
rect 32769 22383 32827 22389
rect 33042 22380 33048 22392
rect 33100 22380 33106 22432
rect 33244 22420 33272 22519
rect 33318 22516 33324 22568
rect 33376 22516 33382 22568
rect 33962 22516 33968 22568
rect 34020 22556 34026 22568
rect 34425 22559 34483 22565
rect 34425 22556 34437 22559
rect 34020 22528 34437 22556
rect 34020 22516 34026 22528
rect 34425 22525 34437 22528
rect 34471 22525 34483 22559
rect 34425 22519 34483 22525
rect 33781 22491 33839 22497
rect 33781 22457 33793 22491
rect 33827 22488 33839 22491
rect 35250 22488 35256 22500
rect 33827 22460 35256 22488
rect 33827 22457 33839 22460
rect 33781 22451 33839 22457
rect 35250 22448 35256 22460
rect 35308 22448 35314 22500
rect 36464 22488 36492 22587
rect 36740 22565 36768 22596
rect 42720 22568 42748 22596
rect 36725 22559 36783 22565
rect 36725 22525 36737 22559
rect 36771 22525 36783 22559
rect 36725 22519 36783 22525
rect 37369 22559 37427 22565
rect 37369 22525 37381 22559
rect 37415 22556 37427 22559
rect 37458 22556 37464 22568
rect 37415 22528 37464 22556
rect 37415 22525 37427 22528
rect 37369 22519 37427 22525
rect 37458 22516 37464 22528
rect 37516 22516 37522 22568
rect 38562 22516 38568 22568
rect 38620 22516 38626 22568
rect 40586 22516 40592 22568
rect 40644 22516 40650 22568
rect 41417 22559 41475 22565
rect 41417 22525 41429 22559
rect 41463 22525 41475 22559
rect 41417 22519 41475 22525
rect 39945 22491 40003 22497
rect 36464 22460 37596 22488
rect 37568 22432 37596 22460
rect 39945 22457 39957 22491
rect 39991 22488 40003 22491
rect 41432 22488 41460 22519
rect 42058 22516 42064 22568
rect 42116 22516 42122 22568
rect 42426 22516 42432 22568
rect 42484 22516 42490 22568
rect 42702 22516 42708 22568
rect 42760 22516 42766 22568
rect 43438 22516 43444 22568
rect 43496 22556 43502 22568
rect 43824 22565 43852 22664
rect 44076 22627 44134 22633
rect 44076 22593 44088 22627
rect 44122 22624 44134 22627
rect 45002 22624 45008 22636
rect 44122 22596 45008 22624
rect 44122 22593 44134 22596
rect 44076 22587 44134 22593
rect 45002 22584 45008 22596
rect 45060 22584 45066 22636
rect 46032 22565 46060 22664
rect 46216 22624 46244 22720
rect 49970 22652 49976 22704
rect 50028 22692 50034 22704
rect 51074 22692 51080 22704
rect 50028 22664 51080 22692
rect 50028 22652 50034 22664
rect 46273 22627 46331 22633
rect 46273 22624 46285 22627
rect 46216 22596 46285 22624
rect 46273 22593 46285 22596
rect 46319 22593 46331 22627
rect 46273 22587 46331 22593
rect 48866 22584 48872 22636
rect 48924 22584 48930 22636
rect 49142 22584 49148 22636
rect 49200 22584 49206 22636
rect 50062 22584 50068 22636
rect 50120 22584 50126 22636
rect 50172 22633 50200 22664
rect 51074 22652 51080 22664
rect 51132 22652 51138 22704
rect 50157 22627 50215 22633
rect 50157 22593 50169 22627
rect 50203 22593 50215 22627
rect 50157 22587 50215 22593
rect 50246 22584 50252 22636
rect 50304 22584 50310 22636
rect 50424 22627 50482 22633
rect 50424 22593 50436 22627
rect 50470 22624 50482 22627
rect 51166 22624 51172 22636
rect 50470 22596 51172 22624
rect 50470 22593 50482 22596
rect 50424 22587 50482 22593
rect 51166 22584 51172 22596
rect 51224 22584 51230 22636
rect 43809 22559 43867 22565
rect 43809 22556 43821 22559
rect 43496 22528 43821 22556
rect 43496 22516 43502 22528
rect 43809 22525 43821 22528
rect 43855 22525 43867 22559
rect 45833 22559 45891 22565
rect 45833 22556 45845 22559
rect 43809 22519 43867 22525
rect 45526 22528 45845 22556
rect 39991 22460 41460 22488
rect 45189 22491 45247 22497
rect 39991 22457 40003 22460
rect 39945 22451 40003 22457
rect 45189 22457 45201 22491
rect 45235 22488 45247 22491
rect 45526 22488 45554 22528
rect 45833 22525 45845 22528
rect 45879 22525 45891 22559
rect 45833 22519 45891 22525
rect 46017 22559 46075 22565
rect 46017 22525 46029 22559
rect 46063 22525 46075 22559
rect 46017 22519 46075 22525
rect 45235 22460 45554 22488
rect 45235 22457 45247 22460
rect 45189 22451 45247 22457
rect 34238 22420 34244 22432
rect 33244 22392 34244 22420
rect 34238 22380 34244 22392
rect 34296 22380 34302 22432
rect 34422 22380 34428 22432
rect 34480 22420 34486 22432
rect 34609 22423 34667 22429
rect 34609 22420 34621 22423
rect 34480 22392 34621 22420
rect 34480 22380 34486 22392
rect 34609 22389 34621 22392
rect 34655 22389 34667 22423
rect 34609 22383 34667 22389
rect 37550 22380 37556 22432
rect 37608 22380 37614 22432
rect 38289 22423 38347 22429
rect 38289 22389 38301 22423
rect 38335 22420 38347 22423
rect 38930 22420 38936 22432
rect 38335 22392 38936 22420
rect 38335 22389 38347 22392
rect 38289 22383 38347 22389
rect 38930 22380 38936 22392
rect 38988 22380 38994 22432
rect 39206 22380 39212 22432
rect 39264 22420 39270 22432
rect 40037 22423 40095 22429
rect 40037 22420 40049 22423
rect 39264 22392 40049 22420
rect 39264 22380 39270 22392
rect 40037 22389 40049 22392
rect 40083 22389 40095 22423
rect 40037 22383 40095 22389
rect 40770 22380 40776 22432
rect 40828 22380 40834 22432
rect 41506 22380 41512 22432
rect 41564 22380 41570 22432
rect 43073 22423 43131 22429
rect 43073 22389 43085 22423
rect 43119 22420 43131 22423
rect 43622 22420 43628 22432
rect 43119 22392 43628 22420
rect 43119 22389 43131 22392
rect 43073 22383 43131 22389
rect 43622 22380 43628 22392
rect 43680 22380 43686 22432
rect 45278 22380 45284 22432
rect 45336 22380 45342 22432
rect 46032 22420 46060 22519
rect 48222 22516 48228 22568
rect 48280 22556 48286 22568
rect 49007 22559 49065 22565
rect 49007 22556 49019 22559
rect 48280 22528 49019 22556
rect 48280 22516 48286 22528
rect 49007 22525 49019 22528
rect 49053 22525 49065 22559
rect 49007 22519 49065 22525
rect 49881 22559 49939 22565
rect 49881 22525 49893 22559
rect 49927 22556 49939 22559
rect 50264 22556 50292 22584
rect 49927 22528 50292 22556
rect 51276 22556 51304 22732
rect 51534 22720 51540 22772
rect 51592 22720 51598 22772
rect 52549 22763 52607 22769
rect 52549 22729 52561 22763
rect 52595 22760 52607 22763
rect 53282 22760 53288 22772
rect 52595 22732 53288 22760
rect 52595 22729 52607 22732
rect 52549 22723 52607 22729
rect 53282 22720 53288 22732
rect 53340 22720 53346 22772
rect 53466 22720 53472 22772
rect 53524 22720 53530 22772
rect 56594 22720 56600 22772
rect 56652 22720 56658 22772
rect 52089 22695 52147 22701
rect 52089 22661 52101 22695
rect 52135 22692 52147 22695
rect 53484 22692 53512 22720
rect 56042 22692 56048 22704
rect 52135 22664 53512 22692
rect 54956 22664 56048 22692
rect 52135 22661 52147 22664
rect 52089 22655 52147 22661
rect 52181 22627 52239 22633
rect 52181 22593 52193 22627
rect 52227 22624 52239 22627
rect 53282 22624 53288 22636
rect 52227 22596 53288 22624
rect 52227 22593 52239 22596
rect 52181 22587 52239 22593
rect 53282 22584 53288 22596
rect 53340 22584 53346 22636
rect 54956 22633 54984 22664
rect 56042 22652 56048 22664
rect 56100 22652 56106 22704
rect 54941 22627 54999 22633
rect 54941 22593 54953 22627
rect 54987 22593 54999 22627
rect 54941 22587 54999 22593
rect 55214 22584 55220 22636
rect 55272 22584 55278 22636
rect 55484 22627 55542 22633
rect 55484 22593 55496 22627
rect 55530 22624 55542 22627
rect 56689 22627 56747 22633
rect 56689 22624 56701 22627
rect 55530 22596 56701 22624
rect 55530 22593 55542 22596
rect 55484 22587 55542 22593
rect 56689 22593 56701 22596
rect 56735 22593 56747 22627
rect 56689 22587 56747 22593
rect 51997 22559 52055 22565
rect 51997 22556 52009 22559
rect 51276 22528 52009 22556
rect 49927 22525 49939 22528
rect 49881 22519 49939 22525
rect 51997 22525 52009 22528
rect 52043 22556 52055 22559
rect 52917 22559 52975 22565
rect 52917 22556 52929 22559
rect 52043 22528 52929 22556
rect 52043 22525 52055 22528
rect 51997 22519 52055 22525
rect 52917 22525 52929 22528
rect 52963 22525 52975 22559
rect 52917 22519 52975 22525
rect 53926 22516 53932 22568
rect 53984 22516 53990 22568
rect 54018 22516 54024 22568
rect 54076 22565 54082 22568
rect 54076 22559 54125 22565
rect 54076 22525 54079 22559
rect 54113 22525 54125 22559
rect 54076 22519 54125 22525
rect 54205 22559 54263 22565
rect 54205 22525 54217 22559
rect 54251 22556 54263 22559
rect 54251 22528 54432 22556
rect 54251 22525 54263 22528
rect 54205 22519 54263 22525
rect 54076 22516 54082 22519
rect 49418 22448 49424 22500
rect 49476 22448 49482 22500
rect 46658 22420 46664 22432
rect 46032 22392 46664 22420
rect 46658 22380 46664 22392
rect 46716 22380 46722 22432
rect 47946 22380 47952 22432
rect 48004 22380 48010 22432
rect 48225 22423 48283 22429
rect 48225 22389 48237 22423
rect 48271 22420 48283 22423
rect 49602 22420 49608 22432
rect 48271 22392 49608 22420
rect 48271 22389 48283 22392
rect 48225 22383 48283 22389
rect 49602 22380 49608 22392
rect 49660 22380 49666 22432
rect 53285 22423 53343 22429
rect 53285 22389 53297 22423
rect 53331 22420 53343 22423
rect 53926 22420 53932 22432
rect 53331 22392 53932 22420
rect 53331 22389 53343 22392
rect 53285 22383 53343 22389
rect 53926 22380 53932 22392
rect 53984 22380 53990 22432
rect 54110 22380 54116 22432
rect 54168 22420 54174 22432
rect 54404 22420 54432 22528
rect 54478 22516 54484 22568
rect 54536 22516 54542 22568
rect 54570 22516 54576 22568
rect 54628 22556 54634 22568
rect 55122 22556 55128 22568
rect 54628 22528 55128 22556
rect 54628 22516 54634 22528
rect 55122 22516 55128 22528
rect 55180 22516 55186 22568
rect 57238 22516 57244 22568
rect 57296 22516 57302 22568
rect 54168 22392 54432 22420
rect 54168 22380 54174 22392
rect 1104 22330 58880 22352
rect 1104 22278 8172 22330
rect 8224 22278 8236 22330
rect 8288 22278 8300 22330
rect 8352 22278 8364 22330
rect 8416 22278 8428 22330
rect 8480 22278 22616 22330
rect 22668 22278 22680 22330
rect 22732 22278 22744 22330
rect 22796 22278 22808 22330
rect 22860 22278 22872 22330
rect 22924 22278 37060 22330
rect 37112 22278 37124 22330
rect 37176 22278 37188 22330
rect 37240 22278 37252 22330
rect 37304 22278 37316 22330
rect 37368 22278 51504 22330
rect 51556 22278 51568 22330
rect 51620 22278 51632 22330
rect 51684 22278 51696 22330
rect 51748 22278 51760 22330
rect 51812 22278 58880 22330
rect 1104 22256 58880 22278
rect 3694 22176 3700 22228
rect 3752 22216 3758 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3752 22188 3801 22216
rect 3752 22176 3758 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 3789 22179 3847 22185
rect 4890 22176 4896 22228
rect 4948 22176 4954 22228
rect 7098 22176 7104 22228
rect 7156 22176 7162 22228
rect 9585 22219 9643 22225
rect 9585 22185 9597 22219
rect 9631 22216 9643 22219
rect 9766 22216 9772 22228
rect 9631 22188 9772 22216
rect 9631 22185 9643 22188
rect 9585 22179 9643 22185
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 10505 22219 10563 22225
rect 10505 22185 10517 22219
rect 10551 22216 10563 22219
rect 11146 22216 11152 22228
rect 10551 22188 11152 22216
rect 10551 22185 10563 22188
rect 10505 22179 10563 22185
rect 11146 22176 11152 22188
rect 11204 22216 11210 22228
rect 12066 22216 12072 22228
rect 11204 22188 12072 22216
rect 11204 22176 11210 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 13814 22216 13820 22228
rect 13775 22188 13820 22216
rect 13814 22176 13820 22188
rect 13872 22176 13878 22228
rect 16390 22216 16396 22228
rect 15212 22188 16396 22216
rect 4908 22148 4936 22176
rect 4448 22120 4936 22148
rect 4448 22089 4476 22120
rect 4433 22083 4491 22089
rect 4433 22049 4445 22083
rect 4479 22080 4491 22083
rect 4479 22052 4513 22080
rect 4479 22049 4491 22052
rect 4433 22043 4491 22049
rect 10134 22040 10140 22092
rect 10192 22040 10198 22092
rect 12158 22040 12164 22092
rect 12216 22040 12222 22092
rect 2958 21972 2964 22024
rect 3016 21972 3022 22024
rect 4706 21972 4712 22024
rect 4764 21972 4770 22024
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 22012 5779 22015
rect 6454 22012 6460 22024
rect 5767 21984 6460 22012
rect 5767 21981 5779 21984
rect 5721 21975 5779 21981
rect 6454 21972 6460 21984
rect 6512 21972 6518 22024
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 9030 21972 9036 22024
rect 9088 22012 9094 22024
rect 11885 22015 11943 22021
rect 11885 22012 11897 22015
rect 9088 21984 11897 22012
rect 9088 21972 9094 21984
rect 11885 21981 11897 21984
rect 11931 21981 11943 22015
rect 11885 21975 11943 21981
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 21981 13415 22015
rect 13832 22012 13860 22176
rect 15212 22148 15240 22188
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 20714 22176 20720 22228
rect 20772 22176 20778 22228
rect 23382 22176 23388 22228
rect 23440 22176 23446 22228
rect 25961 22219 26019 22225
rect 25961 22185 25973 22219
rect 26007 22216 26019 22219
rect 26326 22216 26332 22228
rect 26007 22188 26332 22216
rect 26007 22185 26019 22188
rect 25961 22179 26019 22185
rect 26326 22176 26332 22188
rect 26384 22176 26390 22228
rect 26786 22176 26792 22228
rect 26844 22176 26850 22228
rect 28905 22219 28963 22225
rect 28905 22185 28917 22219
rect 28951 22216 28963 22219
rect 29178 22216 29184 22228
rect 28951 22188 29184 22216
rect 28951 22185 28963 22188
rect 28905 22179 28963 22185
rect 29178 22176 29184 22188
rect 29236 22176 29242 22228
rect 31481 22219 31539 22225
rect 31481 22185 31493 22219
rect 31527 22216 31539 22219
rect 31570 22216 31576 22228
rect 31527 22188 31576 22216
rect 31527 22185 31539 22188
rect 31481 22179 31539 22185
rect 31570 22176 31576 22188
rect 31628 22176 31634 22228
rect 33873 22219 33931 22225
rect 31680 22188 33456 22216
rect 15028 22120 15240 22148
rect 15028 22089 15056 22120
rect 17126 22108 17132 22160
rect 17184 22148 17190 22160
rect 17862 22148 17868 22160
rect 17184 22120 17868 22148
rect 17184 22108 17190 22120
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 15197 22083 15255 22089
rect 15059 22052 15093 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15197 22049 15209 22083
rect 15243 22049 15255 22083
rect 15197 22043 15255 22049
rect 15102 22012 15108 22024
rect 13832 21984 15108 22012
rect 13357 21975 13415 21981
rect 3605 21947 3663 21953
rect 3605 21913 3617 21947
rect 3651 21944 3663 21947
rect 4157 21947 4215 21953
rect 4157 21944 4169 21947
rect 3651 21916 4169 21944
rect 3651 21913 3663 21916
rect 3605 21907 3663 21913
rect 4157 21913 4169 21916
rect 4203 21944 4215 21947
rect 5988 21947 6046 21953
rect 4203 21916 4660 21944
rect 4203 21913 4215 21916
rect 4157 21907 4215 21913
rect 4632 21888 4660 21916
rect 5000 21916 5948 21944
rect 5000 21888 5028 21916
rect 4246 21836 4252 21888
rect 4304 21836 4310 21888
rect 4614 21836 4620 21888
rect 4672 21836 4678 21888
rect 4982 21836 4988 21888
rect 5040 21836 5046 21888
rect 5258 21836 5264 21888
rect 5316 21836 5322 21888
rect 5920 21876 5948 21916
rect 5988 21913 6000 21947
rect 6034 21944 6046 21947
rect 6086 21944 6092 21956
rect 6034 21916 6092 21944
rect 6034 21913 6046 21916
rect 5988 21907 6046 21913
rect 6086 21904 6092 21916
rect 6144 21904 6150 21956
rect 9401 21947 9459 21953
rect 9401 21944 9413 21947
rect 7116 21916 9413 21944
rect 7116 21876 7144 21916
rect 9401 21913 9413 21916
rect 9447 21944 9459 21947
rect 10134 21944 10140 21956
rect 9447 21916 10140 21944
rect 9447 21913 9459 21916
rect 9401 21907 9459 21913
rect 10134 21904 10140 21916
rect 10192 21904 10198 21956
rect 11330 21904 11336 21956
rect 11388 21944 11394 21956
rect 11618 21947 11676 21953
rect 11618 21944 11630 21947
rect 11388 21916 11630 21944
rect 11388 21904 11394 21916
rect 11618 21913 11630 21916
rect 11664 21913 11676 21947
rect 13372 21944 13400 21975
rect 15102 21972 15108 21984
rect 15160 22012 15166 22024
rect 15212 22012 15240 22043
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 16298 22080 16304 22092
rect 15436 22052 16304 22080
rect 15436 22040 15442 22052
rect 16298 22040 16304 22052
rect 16356 22089 16362 22092
rect 16356 22083 16405 22089
rect 16356 22049 16359 22083
rect 16393 22080 16405 22083
rect 16393 22052 16449 22080
rect 16393 22049 16405 22052
rect 16356 22043 16405 22049
rect 16356 22040 16362 22043
rect 16482 22040 16488 22092
rect 16540 22040 16546 22092
rect 16666 22040 16672 22092
rect 16724 22080 16730 22092
rect 16761 22083 16819 22089
rect 16761 22080 16773 22083
rect 16724 22052 16773 22080
rect 16724 22040 16730 22052
rect 16761 22049 16773 22052
rect 16807 22049 16819 22083
rect 16761 22043 16819 22049
rect 17405 22083 17463 22089
rect 17405 22049 17417 22083
rect 17451 22049 17463 22083
rect 17405 22043 17463 22049
rect 15160 21984 15240 22012
rect 15160 21972 15166 21984
rect 16206 21972 16212 22024
rect 16264 21972 16270 22024
rect 17221 22015 17279 22021
rect 17221 21981 17233 22015
rect 17267 21981 17279 22015
rect 17420 22012 17448 22043
rect 17678 22040 17684 22092
rect 17736 22040 17742 22092
rect 17788 22089 17816 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 26804 22148 26832 22176
rect 23768 22120 26832 22148
rect 17773 22083 17831 22089
rect 17773 22049 17785 22083
rect 17819 22080 17831 22083
rect 21361 22083 21419 22089
rect 17819 22052 17853 22080
rect 17819 22049 17831 22052
rect 17773 22043 17831 22049
rect 21361 22049 21373 22083
rect 21407 22080 21419 22083
rect 21726 22080 21732 22092
rect 21407 22052 21732 22080
rect 21407 22049 21419 22052
rect 21361 22043 21419 22049
rect 21726 22040 21732 22052
rect 21784 22080 21790 22092
rect 22097 22083 22155 22089
rect 22097 22080 22109 22083
rect 21784 22052 22109 22080
rect 21784 22040 21790 22052
rect 22097 22049 22109 22052
rect 22143 22049 22155 22083
rect 22097 22043 22155 22049
rect 22370 22040 22376 22092
rect 22428 22040 22434 22092
rect 22554 22040 22560 22092
rect 22612 22080 22618 22092
rect 22649 22083 22707 22089
rect 22649 22080 22661 22083
rect 22612 22052 22661 22080
rect 22612 22040 22618 22052
rect 22649 22049 22661 22052
rect 22695 22080 22707 22083
rect 23768 22080 23796 22120
rect 30558 22108 30564 22160
rect 30616 22148 30622 22160
rect 31680 22148 31708 22188
rect 30616 22120 31708 22148
rect 33428 22148 33456 22188
rect 33873 22185 33885 22219
rect 33919 22216 33931 22219
rect 34330 22216 34336 22228
rect 33919 22188 34336 22216
rect 33919 22185 33931 22188
rect 33873 22179 33931 22185
rect 34330 22176 34336 22188
rect 34388 22176 34394 22228
rect 35066 22176 35072 22228
rect 35124 22216 35130 22228
rect 35802 22216 35808 22228
rect 35124 22188 35808 22216
rect 35124 22176 35130 22188
rect 35802 22176 35808 22188
rect 35860 22216 35866 22228
rect 39853 22219 39911 22225
rect 35860 22188 39252 22216
rect 35860 22176 35866 22188
rect 35084 22148 35112 22176
rect 33428 22120 35112 22148
rect 30616 22108 30622 22120
rect 22695 22052 23796 22080
rect 22695 22049 22707 22052
rect 22649 22043 22707 22049
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 24084 22052 24808 22080
rect 24084 22040 24090 22052
rect 18874 22012 18880 22024
rect 17420 21984 18880 22012
rect 17221 21975 17279 21981
rect 11618 21907 11676 21913
rect 12728 21916 13400 21944
rect 17236 21944 17264 21975
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 19242 21972 19248 22024
rect 19300 22012 19306 22024
rect 19337 22015 19395 22021
rect 19337 22012 19349 22015
rect 19300 21984 19349 22012
rect 19300 21972 19306 21984
rect 19337 21981 19349 21984
rect 19383 22012 19395 22015
rect 20806 22012 20812 22024
rect 19383 21984 20812 22012
rect 19383 21981 19395 21984
rect 19337 21975 19395 21981
rect 20806 21972 20812 21984
rect 20864 21972 20870 22024
rect 22186 21972 22192 22024
rect 22244 22021 22250 22024
rect 22244 22015 22293 22021
rect 22244 21981 22247 22015
rect 22281 21981 22293 22015
rect 22244 21975 22293 21981
rect 23109 22015 23167 22021
rect 23109 21981 23121 22015
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 22244 21972 22250 21975
rect 17865 21947 17923 21953
rect 17865 21944 17877 21947
rect 17236 21916 17877 21944
rect 5920 21848 7144 21876
rect 7190 21836 7196 21888
rect 7248 21836 7254 21888
rect 9858 21836 9864 21888
rect 9916 21876 9922 21888
rect 9953 21879 10011 21885
rect 9953 21876 9965 21879
rect 9916 21848 9965 21876
rect 9916 21836 9922 21848
rect 9953 21845 9965 21848
rect 9999 21845 10011 21879
rect 9953 21839 10011 21845
rect 10045 21879 10103 21885
rect 10045 21845 10057 21879
rect 10091 21876 10103 21879
rect 10870 21876 10876 21888
rect 10091 21848 10876 21876
rect 10091 21845 10103 21848
rect 10045 21839 10103 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 10962 21836 10968 21888
rect 11020 21876 11026 21888
rect 12253 21879 12311 21885
rect 12253 21876 12265 21879
rect 11020 21848 12265 21876
rect 11020 21836 11026 21848
rect 12253 21845 12265 21848
rect 12299 21845 12311 21879
rect 12253 21839 12311 21845
rect 12345 21879 12403 21885
rect 12345 21845 12357 21879
rect 12391 21876 12403 21879
rect 12434 21876 12440 21888
rect 12391 21848 12440 21876
rect 12391 21845 12403 21848
rect 12345 21839 12403 21845
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 12728 21885 12756 21916
rect 17865 21913 17877 21916
rect 17911 21944 17923 21947
rect 17954 21944 17960 21956
rect 17911 21916 17960 21944
rect 17911 21913 17923 21916
rect 17865 21907 17923 21913
rect 17954 21904 17960 21916
rect 18012 21904 18018 21956
rect 19604 21947 19662 21953
rect 18248 21916 19472 21944
rect 12713 21879 12771 21885
rect 12713 21845 12725 21879
rect 12759 21845 12771 21879
rect 12713 21839 12771 21845
rect 12802 21836 12808 21888
rect 12860 21836 12866 21888
rect 14274 21836 14280 21888
rect 14332 21876 14338 21888
rect 14369 21879 14427 21885
rect 14369 21876 14381 21879
rect 14332 21848 14381 21876
rect 14332 21836 14338 21848
rect 14369 21845 14381 21848
rect 14415 21845 14427 21879
rect 14369 21839 14427 21845
rect 14550 21836 14556 21888
rect 14608 21836 14614 21888
rect 14918 21836 14924 21888
rect 14976 21836 14982 21888
rect 15565 21879 15623 21885
rect 15565 21845 15577 21879
rect 15611 21876 15623 21879
rect 16850 21876 16856 21888
rect 15611 21848 16856 21876
rect 15611 21845 15623 21848
rect 15565 21839 15623 21845
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 18248 21885 18276 21916
rect 19444 21888 19472 21916
rect 19604 21913 19616 21947
rect 19650 21944 19662 21947
rect 19794 21944 19800 21956
rect 19650 21916 19800 21944
rect 19650 21913 19662 21916
rect 19604 21907 19662 21913
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 23124 21944 23152 21975
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 23256 21984 23305 22012
rect 23256 21972 23262 21984
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 23753 21947 23811 21953
rect 23753 21944 23765 21947
rect 23124 21916 23765 21944
rect 23753 21913 23765 21916
rect 23799 21944 23811 21947
rect 24397 21947 24455 21953
rect 24397 21944 24409 21947
rect 23799 21916 24409 21944
rect 23799 21913 23811 21916
rect 23753 21907 23811 21913
rect 24397 21913 24409 21916
rect 24443 21913 24455 21947
rect 24780 21944 24808 22052
rect 24854 22040 24860 22092
rect 24912 22080 24918 22092
rect 31312 22089 31340 22120
rect 25777 22083 25835 22089
rect 25777 22080 25789 22083
rect 24912 22052 25789 22080
rect 24912 22040 24918 22052
rect 25777 22049 25789 22052
rect 25823 22080 25835 22083
rect 26513 22083 26571 22089
rect 26513 22080 26525 22083
rect 25823 22052 26525 22080
rect 25823 22049 25835 22052
rect 25777 22043 25835 22049
rect 26513 22049 26525 22052
rect 26559 22049 26571 22083
rect 31297 22083 31355 22089
rect 26513 22043 26571 22049
rect 26620 22052 27016 22080
rect 24946 21972 24952 22024
rect 25004 21972 25010 22024
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 22012 26387 22015
rect 26620 22012 26648 22052
rect 26988 22024 27016 22052
rect 31297 22049 31309 22083
rect 31343 22080 31355 22083
rect 32030 22080 32036 22092
rect 31343 22052 31377 22080
rect 31726 22052 32036 22080
rect 31343 22049 31355 22052
rect 31297 22043 31355 22049
rect 26375 21984 26648 22012
rect 26375 21981 26387 21984
rect 26329 21975 26387 21981
rect 26694 21972 26700 22024
rect 26752 22012 26758 22024
rect 26789 22015 26847 22021
rect 26789 22012 26801 22015
rect 26752 21984 26801 22012
rect 26752 21972 26758 21984
rect 26789 21981 26801 21984
rect 26835 21981 26847 22015
rect 26789 21975 26847 21981
rect 26970 21972 26976 22024
rect 27028 21972 27034 22024
rect 27525 22015 27583 22021
rect 27525 21981 27537 22015
rect 27571 22012 27583 22015
rect 27571 21984 28028 22012
rect 27571 21981 27583 21984
rect 27525 21975 27583 21981
rect 28000 21956 28028 21984
rect 29362 21972 29368 22024
rect 29420 22012 29426 22024
rect 30101 22015 30159 22021
rect 30101 22012 30113 22015
rect 29420 21984 30113 22012
rect 29420 21972 29426 21984
rect 30101 21981 30113 21984
rect 30147 21981 30159 22015
rect 30101 21975 30159 21981
rect 30561 22015 30619 22021
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 31570 22012 31576 22024
rect 30607 21984 31576 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 31570 21972 31576 21984
rect 31628 22012 31634 22024
rect 31726 22012 31754 22052
rect 32030 22040 32036 22052
rect 32088 22040 32094 22092
rect 35434 22080 35440 22092
rect 35176 22052 35440 22080
rect 31628 21984 31754 22012
rect 32493 22015 32551 22021
rect 31628 21972 31634 21984
rect 32493 21981 32505 22015
rect 32539 22012 32551 22015
rect 32582 22012 32588 22024
rect 32539 21984 32588 22012
rect 32539 21981 32551 21984
rect 32493 21975 32551 21981
rect 32582 21972 32588 21984
rect 32640 22012 32646 22024
rect 35176 22012 35204 22052
rect 35434 22040 35440 22052
rect 35492 22040 35498 22092
rect 37476 22089 37504 22188
rect 39114 22108 39120 22160
rect 39172 22108 39178 22160
rect 39224 22148 39252 22188
rect 39853 22185 39865 22219
rect 39899 22216 39911 22219
rect 40586 22216 40592 22228
rect 39899 22188 40592 22216
rect 39899 22185 39911 22188
rect 39853 22179 39911 22185
rect 40586 22176 40592 22188
rect 40644 22176 40650 22228
rect 41785 22219 41843 22225
rect 41785 22185 41797 22219
rect 41831 22216 41843 22219
rect 42058 22216 42064 22228
rect 41831 22188 42064 22216
rect 41831 22185 41843 22188
rect 41785 22179 41843 22185
rect 42058 22176 42064 22188
rect 42116 22176 42122 22228
rect 42610 22176 42616 22228
rect 42668 22176 42674 22228
rect 43456 22188 45048 22216
rect 41138 22148 41144 22160
rect 39224 22120 41144 22148
rect 41138 22108 41144 22120
rect 41196 22108 41202 22160
rect 43456 22148 43484 22188
rect 41340 22120 43484 22148
rect 45020 22148 45048 22188
rect 48866 22176 48872 22228
rect 48924 22216 48930 22228
rect 48961 22219 49019 22225
rect 48961 22216 48973 22219
rect 48924 22188 48973 22216
rect 48924 22176 48930 22188
rect 48961 22185 48973 22188
rect 49007 22185 49019 22219
rect 48961 22179 49019 22185
rect 49418 22176 49424 22228
rect 49476 22176 49482 22228
rect 50062 22216 50068 22228
rect 49712 22188 50068 22216
rect 46566 22148 46572 22160
rect 45020 22120 46572 22148
rect 37461 22083 37519 22089
rect 37461 22049 37473 22083
rect 37507 22049 37519 22083
rect 37826 22080 37832 22092
rect 37461 22043 37519 22049
rect 37568 22052 37832 22080
rect 32640 21984 35204 22012
rect 32640 21972 32646 21984
rect 35250 21972 35256 22024
rect 35308 21972 35314 22024
rect 37277 22015 37335 22021
rect 37277 21981 37289 22015
rect 37323 22012 37335 22015
rect 37568 22012 37596 22052
rect 37826 22040 37832 22052
rect 37884 22080 37890 22092
rect 38519 22083 38577 22089
rect 38519 22080 38531 22083
rect 37884 22052 38531 22080
rect 37884 22040 37890 22052
rect 38519 22049 38531 22052
rect 38565 22049 38577 22083
rect 38519 22043 38577 22049
rect 38654 22040 38660 22092
rect 38712 22040 38718 22092
rect 38930 22080 38936 22092
rect 38891 22052 38936 22080
rect 38930 22040 38936 22052
rect 38988 22080 38994 22092
rect 39132 22080 39160 22108
rect 38988 22052 39160 22080
rect 39393 22083 39451 22089
rect 38988 22040 38994 22052
rect 39393 22049 39405 22083
rect 39439 22080 39451 22083
rect 40034 22080 40040 22092
rect 39439 22052 40040 22080
rect 39439 22049 39451 22052
rect 39393 22043 39451 22049
rect 40034 22040 40040 22052
rect 40092 22040 40098 22092
rect 40494 22040 40500 22092
rect 40552 22080 40558 22092
rect 41340 22080 41368 22120
rect 40552 22052 41368 22080
rect 41693 22083 41751 22089
rect 40552 22040 40558 22052
rect 41693 22049 41705 22083
rect 41739 22080 41751 22083
rect 42429 22083 42487 22089
rect 42429 22080 42441 22083
rect 41739 22052 42441 22080
rect 41739 22049 41751 22052
rect 41693 22043 41751 22049
rect 42429 22049 42441 22052
rect 42475 22080 42487 22083
rect 42518 22080 42524 22092
rect 42475 22052 42524 22080
rect 42475 22049 42487 22052
rect 42429 22043 42487 22049
rect 37323 21984 37596 22012
rect 37323 21981 37335 21984
rect 37277 21975 37335 21981
rect 38378 21972 38384 22024
rect 38436 21972 38442 22024
rect 39577 22015 39635 22021
rect 39577 21981 39589 22015
rect 39623 22012 39635 22015
rect 40313 22015 40371 22021
rect 40313 22012 40325 22015
rect 39623 21984 40325 22012
rect 39623 21981 39635 21984
rect 39577 21975 39635 21981
rect 40313 21981 40325 21984
rect 40359 22012 40371 22015
rect 40681 22015 40739 22021
rect 40681 22012 40693 22015
rect 40359 21984 40693 22012
rect 40359 21981 40371 21984
rect 40313 21975 40371 21981
rect 40681 21981 40693 21984
rect 40727 21981 40739 22015
rect 40681 21975 40739 21981
rect 41233 22015 41291 22021
rect 41233 21981 41245 22015
rect 41279 21981 41291 22015
rect 41233 21975 41291 21981
rect 27798 21953 27804 21956
rect 24780 21916 27568 21944
rect 24397 21907 24455 21913
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21845 18291 21879
rect 18233 21839 18291 21845
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 19058 21876 19064 21888
rect 18656 21848 19064 21876
rect 18656 21836 18662 21848
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19426 21836 19432 21888
rect 19484 21836 19490 21888
rect 21453 21879 21511 21885
rect 21453 21845 21465 21879
rect 21499 21876 21511 21879
rect 22462 21876 22468 21888
rect 21499 21848 22468 21876
rect 21499 21845 21511 21848
rect 21453 21839 21511 21845
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 23106 21836 23112 21888
rect 23164 21876 23170 21888
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23164 21848 23857 21876
rect 23164 21836 23170 21848
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 23845 21839 23903 21845
rect 26421 21879 26479 21885
rect 26421 21845 26433 21879
rect 26467 21876 26479 21879
rect 27430 21876 27436 21888
rect 26467 21848 27436 21876
rect 26467 21845 26479 21848
rect 26421 21839 26479 21845
rect 27430 21836 27436 21848
rect 27488 21836 27494 21888
rect 27540 21876 27568 21916
rect 27792 21907 27804 21953
rect 27798 21904 27804 21907
rect 27856 21904 27862 21956
rect 27982 21904 27988 21956
rect 28040 21904 28046 21956
rect 31021 21947 31079 21953
rect 31021 21913 31033 21947
rect 31067 21944 31079 21947
rect 32214 21944 32220 21956
rect 31067 21916 32220 21944
rect 31067 21913 31079 21916
rect 31021 21907 31079 21913
rect 32214 21904 32220 21916
rect 32272 21904 32278 21956
rect 32760 21947 32818 21953
rect 32760 21913 32772 21947
rect 32806 21944 32818 21947
rect 33410 21944 33416 21956
rect 32806 21916 33416 21944
rect 32806 21913 32818 21916
rect 32760 21907 32818 21913
rect 33410 21904 33416 21916
rect 33468 21904 33474 21956
rect 35704 21947 35762 21953
rect 35704 21913 35716 21947
rect 35750 21944 35762 21947
rect 36354 21944 36360 21956
rect 35750 21916 36360 21944
rect 35750 21913 35762 21916
rect 35704 21907 35762 21913
rect 36354 21904 36360 21916
rect 36412 21904 36418 21956
rect 41248 21944 41276 21975
rect 41414 21972 41420 22024
rect 41472 22012 41478 22024
rect 41708 22012 41736 22043
rect 42518 22040 42524 22052
rect 42576 22040 42582 22092
rect 42702 22040 42708 22092
rect 42760 22080 42766 22092
rect 45112 22089 45140 22120
rect 46566 22108 46572 22120
rect 46624 22108 46630 22160
rect 47946 22108 47952 22160
rect 48004 22148 48010 22160
rect 49436 22148 49464 22176
rect 48004 22120 49464 22148
rect 48004 22108 48010 22120
rect 43165 22083 43223 22089
rect 43165 22080 43177 22083
rect 42760 22052 43177 22080
rect 42760 22040 42766 22052
rect 43165 22049 43177 22052
rect 43211 22049 43223 22083
rect 43165 22043 43223 22049
rect 45097 22083 45155 22089
rect 45097 22049 45109 22083
rect 45143 22080 45155 22083
rect 45143 22052 45177 22080
rect 45143 22049 45155 22052
rect 45097 22043 45155 22049
rect 48590 22040 48596 22092
rect 48648 22040 48654 22092
rect 49712 22089 49740 22188
rect 50062 22176 50068 22188
rect 50120 22176 50126 22228
rect 51074 22176 51080 22228
rect 51132 22216 51138 22228
rect 51902 22216 51908 22228
rect 51132 22188 51908 22216
rect 51132 22176 51138 22188
rect 49697 22083 49755 22089
rect 49697 22049 49709 22083
rect 49743 22049 49755 22083
rect 49697 22043 49755 22049
rect 49881 22083 49939 22089
rect 49881 22049 49893 22083
rect 49927 22049 49939 22083
rect 49881 22043 49939 22049
rect 41472 21984 41736 22012
rect 41472 21972 41478 21984
rect 43438 21972 43444 22024
rect 43496 21972 43502 22024
rect 43708 22015 43766 22021
rect 43708 21981 43720 22015
rect 43754 22012 43766 22015
rect 45833 22015 45891 22021
rect 45833 22012 45845 22015
rect 43754 21984 45845 22012
rect 43754 21981 43766 21984
rect 43708 21975 43766 21981
rect 45833 21981 45845 21984
rect 45879 21981 45891 22015
rect 45833 21975 45891 21981
rect 46385 22015 46443 22021
rect 46385 21981 46397 22015
rect 46431 21981 46443 22015
rect 46385 21975 46443 21981
rect 46569 22015 46627 22021
rect 46569 21981 46581 22015
rect 46615 22012 46627 22015
rect 46658 22012 46664 22024
rect 46615 21984 46664 22012
rect 46615 21981 46627 21984
rect 46569 21975 46627 21981
rect 39684 21916 41276 21944
rect 42153 21947 42211 21953
rect 29273 21879 29331 21885
rect 29273 21876 29285 21879
rect 27540 21848 29285 21876
rect 29273 21845 29285 21848
rect 29319 21876 29331 21879
rect 29454 21876 29460 21888
rect 29319 21848 29460 21876
rect 29319 21845 29331 21848
rect 29273 21839 29331 21845
rect 29454 21836 29460 21848
rect 29512 21836 29518 21888
rect 29546 21836 29552 21888
rect 29604 21836 29610 21888
rect 30650 21836 30656 21888
rect 30708 21836 30714 21888
rect 31113 21879 31171 21885
rect 31113 21845 31125 21879
rect 31159 21876 31171 21879
rect 31478 21876 31484 21888
rect 31159 21848 31484 21876
rect 31159 21845 31171 21848
rect 31113 21839 31171 21845
rect 31478 21836 31484 21848
rect 31536 21876 31542 21888
rect 31849 21879 31907 21885
rect 31849 21876 31861 21879
rect 31536 21848 31861 21876
rect 31536 21836 31542 21848
rect 31849 21845 31861 21848
rect 31895 21845 31907 21879
rect 31849 21839 31907 21845
rect 31941 21879 31999 21885
rect 31941 21845 31953 21879
rect 31987 21876 31999 21879
rect 33042 21876 33048 21888
rect 31987 21848 33048 21876
rect 31987 21845 31999 21848
rect 31941 21839 31999 21845
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 34146 21836 34152 21888
rect 34204 21836 34210 21888
rect 34698 21836 34704 21888
rect 34756 21836 34762 21888
rect 36814 21836 36820 21888
rect 36872 21836 36878 21888
rect 36906 21836 36912 21888
rect 36964 21836 36970 21888
rect 37369 21879 37427 21885
rect 37369 21845 37381 21879
rect 37415 21876 37427 21879
rect 37550 21876 37556 21888
rect 37415 21848 37556 21876
rect 37415 21845 37427 21848
rect 37369 21839 37427 21845
rect 37550 21836 37556 21848
rect 37608 21836 37614 21888
rect 37737 21879 37795 21885
rect 37737 21845 37749 21879
rect 37783 21876 37795 21879
rect 39022 21876 39028 21888
rect 37783 21848 39028 21876
rect 37783 21845 37795 21848
rect 37737 21839 37795 21845
rect 39022 21836 39028 21848
rect 39080 21836 39086 21888
rect 39574 21836 39580 21888
rect 39632 21876 39638 21888
rect 39684 21876 39712 21916
rect 42153 21913 42165 21947
rect 42199 21944 42211 21947
rect 43622 21944 43628 21956
rect 42199 21916 43628 21944
rect 42199 21913 42211 21916
rect 42153 21907 42211 21913
rect 43622 21904 43628 21916
rect 43680 21904 43686 21956
rect 46400 21944 46428 21975
rect 46658 21972 46664 21984
rect 46716 21972 46722 22024
rect 44836 21916 45508 21944
rect 39632 21848 39712 21876
rect 39632 21836 39638 21848
rect 40126 21836 40132 21888
rect 40184 21876 40190 21888
rect 40221 21879 40279 21885
rect 40221 21876 40233 21879
rect 40184 21848 40233 21876
rect 40184 21836 40190 21848
rect 40221 21845 40233 21848
rect 40267 21845 40279 21879
rect 40221 21839 40279 21845
rect 42245 21879 42303 21885
rect 42245 21845 42257 21879
rect 42291 21876 42303 21879
rect 42518 21876 42524 21888
rect 42291 21848 42524 21876
rect 42291 21845 42303 21848
rect 42245 21839 42303 21845
rect 42518 21836 42524 21848
rect 42576 21876 42582 21888
rect 42981 21879 43039 21885
rect 42981 21876 42993 21879
rect 42576 21848 42993 21876
rect 42576 21836 42582 21848
rect 42981 21845 42993 21848
rect 43027 21845 43039 21879
rect 42981 21839 43039 21845
rect 43073 21879 43131 21885
rect 43073 21845 43085 21879
rect 43119 21876 43131 21879
rect 43806 21876 43812 21888
rect 43119 21848 43812 21876
rect 43119 21845 43131 21848
rect 43073 21839 43131 21845
rect 43806 21836 43812 21848
rect 43864 21836 43870 21888
rect 44836 21885 44864 21916
rect 45480 21888 45508 21916
rect 45756 21916 46428 21944
rect 46836 21947 46894 21953
rect 44821 21879 44879 21885
rect 44821 21845 44833 21879
rect 44867 21845 44879 21879
rect 44821 21839 44879 21845
rect 45278 21836 45284 21888
rect 45336 21836 45342 21888
rect 45370 21836 45376 21888
rect 45428 21836 45434 21888
rect 45462 21836 45468 21888
rect 45520 21836 45526 21888
rect 45756 21885 45784 21916
rect 46836 21913 46848 21947
rect 46882 21944 46894 21947
rect 48041 21947 48099 21953
rect 48041 21944 48053 21947
rect 46882 21916 48053 21944
rect 46882 21913 46894 21916
rect 46836 21907 46894 21913
rect 48041 21913 48053 21916
rect 48087 21913 48099 21947
rect 48041 21907 48099 21913
rect 48130 21904 48136 21956
rect 48188 21944 48194 21956
rect 48188 21916 49464 21944
rect 48188 21904 48194 21916
rect 49436 21888 49464 21916
rect 49510 21904 49516 21956
rect 49568 21944 49574 21956
rect 49896 21944 49924 22043
rect 50154 22040 50160 22092
rect 50212 22080 50218 22092
rect 51552 22089 51580 22188
rect 51902 22176 51908 22188
rect 51960 22176 51966 22228
rect 52546 22108 52552 22160
rect 52604 22148 52610 22160
rect 52604 22120 53604 22148
rect 52604 22108 52610 22120
rect 53576 22094 53604 22120
rect 53576 22089 53641 22094
rect 50249 22083 50307 22089
rect 50249 22080 50261 22083
rect 50212 22052 50261 22080
rect 50212 22040 50218 22052
rect 50249 22049 50261 22052
rect 50295 22049 50307 22083
rect 50249 22043 50307 22049
rect 51537 22083 51595 22089
rect 51537 22049 51549 22083
rect 51583 22049 51595 22083
rect 51537 22043 51595 22049
rect 53561 22083 53641 22089
rect 53561 22049 53573 22083
rect 53607 22066 53641 22083
rect 53607 22049 53619 22066
rect 53561 22043 53619 22049
rect 54570 22040 54576 22092
rect 54628 22040 54634 22092
rect 54662 22040 54668 22092
rect 54720 22040 54726 22092
rect 55214 22040 55220 22092
rect 55272 22080 55278 22092
rect 55401 22083 55459 22089
rect 55401 22080 55413 22083
rect 55272 22052 55413 22080
rect 55272 22040 55278 22052
rect 55401 22049 55413 22052
rect 55447 22049 55459 22083
rect 55401 22043 55459 22049
rect 53377 22015 53435 22021
rect 53377 21981 53389 22015
rect 53423 22012 53435 22015
rect 54018 22012 54024 22024
rect 53423 21984 54024 22012
rect 53423 21981 53435 21984
rect 53377 21975 53435 21981
rect 54018 21972 54024 21984
rect 54076 21972 54082 22024
rect 55677 22015 55735 22021
rect 55677 21981 55689 22015
rect 55723 22012 55735 22015
rect 56042 22012 56048 22024
rect 55723 21984 56048 22012
rect 55723 21981 55735 21984
rect 55677 21975 55735 21981
rect 56042 21972 56048 21984
rect 56100 21972 56106 22024
rect 49568 21916 49924 21944
rect 49568 21904 49574 21916
rect 50246 21904 50252 21956
rect 50304 21944 50310 21956
rect 50525 21947 50583 21953
rect 50525 21944 50537 21947
rect 50304 21916 50537 21944
rect 50304 21904 50310 21916
rect 50525 21913 50537 21916
rect 50571 21913 50583 21947
rect 50525 21907 50583 21913
rect 51804 21947 51862 21953
rect 51804 21913 51816 21947
rect 51850 21944 51862 21947
rect 52730 21944 52736 21956
rect 51850 21916 52736 21944
rect 51850 21913 51862 21916
rect 51804 21907 51862 21913
rect 52730 21904 52736 21916
rect 52788 21904 52794 21956
rect 53466 21904 53472 21956
rect 53524 21944 53530 21956
rect 53524 21916 54524 21944
rect 53524 21904 53530 21916
rect 45741 21879 45799 21885
rect 45741 21845 45753 21879
rect 45787 21845 45799 21879
rect 45741 21839 45799 21845
rect 47946 21836 47952 21888
rect 48004 21836 48010 21888
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 49418 21836 49424 21888
rect 49476 21876 49482 21888
rect 49605 21879 49663 21885
rect 49605 21876 49617 21879
rect 49476 21848 49617 21876
rect 49476 21836 49482 21848
rect 49605 21845 49617 21848
rect 49651 21876 49663 21879
rect 50433 21879 50491 21885
rect 50433 21876 50445 21879
rect 49651 21848 50445 21876
rect 49651 21845 49663 21848
rect 49605 21839 49663 21845
rect 50433 21845 50445 21848
rect 50479 21845 50491 21879
rect 50433 21839 50491 21845
rect 50890 21836 50896 21888
rect 50948 21836 50954 21888
rect 52914 21836 52920 21888
rect 52972 21836 52978 21888
rect 53009 21879 53067 21885
rect 53009 21845 53021 21879
rect 53055 21876 53067 21879
rect 53282 21876 53288 21888
rect 53055 21848 53288 21876
rect 53055 21845 53067 21848
rect 53009 21839 53067 21845
rect 53282 21836 53288 21848
rect 53340 21836 53346 21888
rect 54110 21836 54116 21888
rect 54168 21836 54174 21888
rect 54496 21885 54524 21916
rect 54481 21879 54539 21885
rect 54481 21845 54493 21879
rect 54527 21876 54539 21879
rect 54570 21876 54576 21888
rect 54527 21848 54576 21876
rect 54527 21845 54539 21848
rect 54481 21839 54539 21845
rect 54570 21836 54576 21848
rect 54628 21876 54634 21888
rect 55585 21879 55643 21885
rect 55585 21876 55597 21879
rect 54628 21848 55597 21876
rect 54628 21836 54634 21848
rect 55585 21845 55597 21848
rect 55631 21845 55643 21879
rect 55585 21839 55643 21845
rect 56045 21879 56103 21885
rect 56045 21845 56057 21879
rect 56091 21876 56103 21879
rect 57238 21876 57244 21888
rect 56091 21848 57244 21876
rect 56091 21845 56103 21848
rect 56045 21839 56103 21845
rect 57238 21836 57244 21848
rect 57296 21836 57302 21888
rect 1104 21786 59040 21808
rect 1104 21734 15394 21786
rect 15446 21734 15458 21786
rect 15510 21734 15522 21786
rect 15574 21734 15586 21786
rect 15638 21734 15650 21786
rect 15702 21734 29838 21786
rect 29890 21734 29902 21786
rect 29954 21734 29966 21786
rect 30018 21734 30030 21786
rect 30082 21734 30094 21786
rect 30146 21734 44282 21786
rect 44334 21734 44346 21786
rect 44398 21734 44410 21786
rect 44462 21734 44474 21786
rect 44526 21734 44538 21786
rect 44590 21734 58726 21786
rect 58778 21734 58790 21786
rect 58842 21734 58854 21786
rect 58906 21734 58918 21786
rect 58970 21734 58982 21786
rect 59034 21734 59040 21786
rect 1104 21712 59040 21734
rect 1949 21675 2007 21681
rect 1949 21641 1961 21675
rect 1995 21672 2007 21675
rect 2958 21672 2964 21684
rect 1995 21644 2964 21672
rect 1995 21641 2007 21644
rect 1949 21635 2007 21641
rect 2958 21632 2964 21644
rect 3016 21632 3022 21684
rect 4706 21632 4712 21684
rect 4764 21672 4770 21684
rect 4801 21675 4859 21681
rect 4801 21672 4813 21675
rect 4764 21644 4813 21672
rect 4764 21632 4770 21644
rect 4801 21641 4813 21644
rect 4847 21641 4859 21675
rect 4801 21635 4859 21641
rect 5718 21632 5724 21684
rect 5776 21632 5782 21684
rect 6181 21675 6239 21681
rect 6181 21641 6193 21675
rect 6227 21672 6239 21675
rect 6638 21672 6644 21684
rect 6227 21644 6644 21672
rect 6227 21641 6239 21644
rect 6181 21635 6239 21641
rect 6638 21632 6644 21644
rect 6696 21632 6702 21684
rect 7190 21632 7196 21684
rect 7248 21632 7254 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 10100 21644 10241 21672
rect 10100 21632 10106 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 10229 21635 10287 21641
rect 10597 21675 10655 21681
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10686 21672 10692 21684
rect 10643 21644 10692 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11054 21632 11060 21684
rect 11112 21632 11118 21684
rect 11517 21675 11575 21681
rect 11517 21641 11529 21675
rect 11563 21672 11575 21675
rect 11974 21672 11980 21684
rect 11563 21644 11980 21672
rect 11563 21641 11575 21644
rect 11517 21635 11575 21641
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 14461 21675 14519 21681
rect 14461 21672 14473 21675
rect 14424 21644 14473 21672
rect 14424 21632 14430 21644
rect 14461 21641 14473 21644
rect 14507 21641 14519 21675
rect 14461 21635 14519 21641
rect 16114 21632 16120 21684
rect 16172 21672 16178 21684
rect 21082 21672 21088 21684
rect 16172 21644 21088 21672
rect 16172 21632 16178 21644
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 21361 21675 21419 21681
rect 21361 21641 21373 21675
rect 21407 21672 21419 21675
rect 22370 21672 22376 21684
rect 21407 21644 22376 21672
rect 21407 21641 21419 21644
rect 21361 21635 21419 21641
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 23845 21675 23903 21681
rect 23845 21641 23857 21675
rect 23891 21672 23903 21675
rect 24946 21672 24952 21684
rect 23891 21644 24952 21672
rect 23891 21641 23903 21644
rect 23845 21635 23903 21641
rect 24946 21632 24952 21644
rect 25004 21632 25010 21684
rect 27982 21672 27988 21684
rect 25332 21644 27988 21672
rect 3050 21564 3056 21616
rect 3108 21613 3114 21616
rect 3108 21604 3120 21613
rect 6724 21607 6782 21613
rect 3108 21576 3153 21604
rect 3436 21576 6500 21604
rect 3108 21567 3120 21576
rect 3108 21564 3114 21567
rect 3436 21545 3464 21576
rect 3694 21545 3700 21548
rect 3329 21539 3387 21545
rect 3329 21505 3341 21539
rect 3375 21536 3387 21539
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 3375 21508 3433 21536
rect 3375 21505 3387 21508
rect 3329 21499 3387 21505
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3688 21536 3700 21545
rect 3655 21508 3700 21536
rect 3421 21499 3479 21505
rect 3688 21499 3700 21508
rect 3694 21496 3700 21499
rect 3752 21496 3758 21548
rect 4246 21496 4252 21548
rect 4304 21536 4310 21548
rect 5813 21539 5871 21545
rect 5813 21536 5825 21539
rect 4304 21508 5825 21536
rect 4304 21496 4310 21508
rect 5813 21505 5825 21508
rect 5859 21536 5871 21539
rect 6178 21536 6184 21548
rect 5859 21508 6184 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 6472 21480 6500 21576
rect 6724 21573 6736 21607
rect 6770 21604 6782 21607
rect 7208 21604 7236 21632
rect 6770 21576 7236 21604
rect 9116 21607 9174 21613
rect 6770 21573 6782 21576
rect 6724 21567 6782 21573
rect 9116 21573 9128 21607
rect 9162 21604 9174 21607
rect 9214 21604 9220 21616
rect 9162 21576 9220 21604
rect 9162 21573 9174 21576
rect 9116 21567 9174 21573
rect 9214 21564 9220 21576
rect 9272 21564 9278 21616
rect 9858 21564 9864 21616
rect 9916 21604 9922 21616
rect 12652 21607 12710 21613
rect 9916 21576 10180 21604
rect 9916 21564 9922 21576
rect 10152 21548 10180 21576
rect 12652 21573 12664 21607
rect 12698 21604 12710 21607
rect 12820 21604 12848 21632
rect 12698 21576 12848 21604
rect 12698 21573 12710 21576
rect 12652 21567 12710 21573
rect 20806 21564 20812 21616
rect 20864 21604 20870 21616
rect 25332 21604 25360 21644
rect 27982 21632 27988 21644
rect 28040 21632 28046 21684
rect 29273 21675 29331 21681
rect 29273 21641 29285 21675
rect 29319 21672 29331 21675
rect 29546 21672 29552 21684
rect 29319 21644 29552 21672
rect 29319 21641 29331 21644
rect 29273 21635 29331 21641
rect 25590 21613 25596 21616
rect 25584 21604 25596 21613
rect 20864 21576 25360 21604
rect 25551 21576 25596 21604
rect 20864 21564 20870 21576
rect 7484 21508 9904 21536
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5399 21440 5641 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5629 21437 5641 21440
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 5644 21332 5672 21431
rect 6454 21428 6460 21480
rect 6512 21428 6518 21480
rect 7484 21332 7512 21508
rect 8481 21471 8539 21477
rect 8481 21468 8493 21471
rect 7852 21440 8493 21468
rect 7852 21409 7880 21440
rect 8481 21437 8493 21440
rect 8527 21437 8539 21471
rect 8481 21431 8539 21437
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21437 8907 21471
rect 9876 21468 9904 21508
rect 10134 21496 10140 21548
rect 10192 21536 10198 21548
rect 10962 21536 10968 21548
rect 10192 21508 10968 21536
rect 10192 21496 10198 21508
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 12897 21539 12955 21545
rect 11256 21508 12848 21536
rect 11256 21477 11284 21508
rect 11241 21471 11299 21477
rect 11241 21468 11253 21471
rect 9876 21440 11253 21468
rect 8849 21431 8907 21437
rect 11241 21437 11253 21440
rect 11287 21437 11299 21471
rect 12820 21468 12848 21508
rect 12897 21505 12909 21539
rect 12943 21536 12955 21539
rect 13630 21536 13636 21548
rect 12943 21508 13636 21536
rect 12943 21505 12955 21508
rect 12897 21499 12955 21505
rect 13630 21496 13636 21508
rect 13688 21496 13694 21548
rect 14550 21496 14556 21548
rect 14608 21536 14614 21548
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 14608 21508 15025 21536
rect 14608 21496 14614 21508
rect 15013 21505 15025 21508
rect 15059 21505 15071 21539
rect 15013 21499 15071 21505
rect 18782 21496 18788 21548
rect 18840 21536 18846 21548
rect 22480 21545 22508 21576
rect 25332 21548 25360 21576
rect 25584 21567 25596 21576
rect 25590 21564 25596 21567
rect 25648 21564 25654 21616
rect 19153 21539 19211 21545
rect 19153 21536 19165 21539
rect 18840 21508 19165 21536
rect 18840 21496 18846 21508
rect 19153 21505 19165 21508
rect 19199 21536 19211 21539
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 19199 21508 21005 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 20993 21505 21005 21508
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 22732 21539 22790 21545
rect 22732 21505 22744 21539
rect 22778 21536 22790 21539
rect 23290 21536 23296 21548
rect 22778 21508 23296 21536
rect 22778 21505 22790 21508
rect 22732 21499 22790 21505
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 25314 21496 25320 21548
rect 25372 21496 25378 21548
rect 27893 21539 27951 21545
rect 27893 21505 27905 21539
rect 27939 21505 27951 21539
rect 27893 21499 27951 21505
rect 12820 21440 13308 21468
rect 11241 21431 11299 21437
rect 7837 21403 7895 21409
rect 7837 21369 7849 21403
rect 7883 21369 7895 21403
rect 7837 21363 7895 21369
rect 5644 21304 7512 21332
rect 7926 21292 7932 21344
rect 7984 21292 7990 21344
rect 8864 21332 8892 21431
rect 9030 21332 9036 21344
rect 8864 21304 9036 21332
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 13280 21341 13308 21440
rect 18432 21440 22508 21468
rect 18432 21344 18460 21440
rect 22094 21400 22100 21412
rect 19076 21372 22100 21400
rect 19076 21344 19104 21372
rect 22094 21360 22100 21372
rect 22152 21360 22158 21412
rect 13265 21335 13323 21341
rect 13265 21301 13277 21335
rect 13311 21332 13323 21335
rect 13538 21332 13544 21344
rect 13311 21304 13544 21332
rect 13311 21301 13323 21304
rect 13265 21295 13323 21301
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 15378 21292 15384 21344
rect 15436 21332 15442 21344
rect 16206 21332 16212 21344
rect 15436 21304 16212 21332
rect 15436 21292 15442 21304
rect 16206 21292 16212 21304
rect 16264 21292 16270 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 16632 21304 17417 21332
rect 16632 21292 16638 21304
rect 17405 21301 17417 21304
rect 17451 21332 17463 21335
rect 17678 21332 17684 21344
rect 17451 21304 17684 21332
rect 17451 21301 17463 21304
rect 17405 21295 17463 21301
rect 17678 21292 17684 21304
rect 17736 21332 17742 21344
rect 18414 21332 18420 21344
rect 17736 21304 18420 21332
rect 17736 21292 17742 21304
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 19058 21292 19064 21344
rect 19116 21292 19122 21344
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19300 21304 19533 21332
rect 19300 21292 19306 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 22480 21332 22508 21440
rect 27430 21428 27436 21480
rect 27488 21468 27494 21480
rect 27798 21477 27804 21480
rect 27607 21471 27665 21477
rect 27607 21468 27619 21471
rect 27488 21440 27619 21468
rect 27488 21428 27494 21440
rect 27607 21437 27619 21440
rect 27653 21437 27665 21471
rect 27607 21431 27665 21437
rect 27755 21471 27804 21477
rect 27755 21437 27767 21471
rect 27801 21437 27804 21471
rect 27755 21431 27804 21437
rect 27798 21428 27804 21431
rect 27856 21428 27862 21480
rect 27908 21468 27936 21499
rect 28442 21496 28448 21548
rect 28500 21536 28506 21548
rect 28813 21539 28871 21545
rect 28813 21536 28825 21539
rect 28500 21508 28825 21536
rect 28500 21496 28506 21508
rect 28813 21505 28825 21508
rect 28859 21505 28871 21539
rect 28813 21499 28871 21505
rect 28074 21468 28080 21480
rect 27908 21440 28080 21468
rect 28074 21428 28080 21440
rect 28132 21428 28138 21480
rect 28629 21471 28687 21477
rect 28629 21437 28641 21471
rect 28675 21468 28687 21471
rect 29288 21468 29316 21635
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 31573 21675 31631 21681
rect 31573 21641 31585 21675
rect 31619 21672 31631 21675
rect 31662 21672 31668 21684
rect 31619 21644 31668 21672
rect 31619 21641 31631 21644
rect 31573 21635 31631 21641
rect 31662 21632 31668 21644
rect 31720 21632 31726 21684
rect 33318 21672 33324 21684
rect 32324 21644 33324 21672
rect 29454 21564 29460 21616
rect 29512 21564 29518 21616
rect 30460 21607 30518 21613
rect 30460 21573 30472 21607
rect 30506 21604 30518 21607
rect 31018 21604 31024 21616
rect 30506 21576 31024 21604
rect 30506 21573 30518 21576
rect 30460 21567 30518 21573
rect 31018 21564 31024 21576
rect 31076 21564 31082 21616
rect 31478 21564 31484 21616
rect 31536 21604 31542 21616
rect 32324 21604 32352 21644
rect 33318 21632 33324 21644
rect 33376 21632 33382 21684
rect 34054 21632 34060 21684
rect 34112 21632 34118 21684
rect 34422 21632 34428 21684
rect 34480 21672 34486 21684
rect 34517 21675 34575 21681
rect 34517 21672 34529 21675
rect 34480 21644 34529 21672
rect 34480 21632 34486 21644
rect 34517 21641 34529 21644
rect 34563 21641 34575 21675
rect 34517 21635 34575 21641
rect 36817 21675 36875 21681
rect 36817 21641 36829 21675
rect 36863 21672 36875 21675
rect 37458 21672 37464 21684
rect 36863 21644 37464 21672
rect 36863 21641 36875 21644
rect 36817 21635 36875 21641
rect 37458 21632 37464 21644
rect 37516 21632 37522 21684
rect 37826 21632 37832 21684
rect 37884 21672 37890 21684
rect 37921 21675 37979 21681
rect 37921 21672 37933 21675
rect 37884 21644 37933 21672
rect 37884 21632 37890 21644
rect 37921 21641 37933 21644
rect 37967 21641 37979 21675
rect 37921 21635 37979 21641
rect 39574 21632 39580 21684
rect 39632 21632 39638 21684
rect 39669 21675 39727 21681
rect 39669 21641 39681 21675
rect 39715 21672 39727 21675
rect 40402 21672 40408 21684
rect 39715 21644 40408 21672
rect 39715 21641 39727 21644
rect 39669 21635 39727 21641
rect 40402 21632 40408 21644
rect 40460 21632 40466 21684
rect 43438 21672 43444 21684
rect 41386 21644 43444 21672
rect 34440 21604 34468 21632
rect 38562 21604 38568 21616
rect 31536 21576 32352 21604
rect 33980 21576 34468 21604
rect 35452 21576 36768 21604
rect 31536 21564 31542 21576
rect 29472 21477 29500 21564
rect 32950 21545 32956 21548
rect 32769 21539 32827 21545
rect 32769 21505 32781 21539
rect 32815 21536 32827 21539
rect 32928 21539 32956 21545
rect 32815 21508 32895 21536
rect 32815 21505 32827 21508
rect 32769 21499 32827 21505
rect 28675 21440 29316 21468
rect 29365 21471 29423 21477
rect 28675 21437 28687 21440
rect 28629 21431 28687 21437
rect 29365 21437 29377 21471
rect 29411 21437 29423 21471
rect 29365 21431 29423 21437
rect 29457 21471 29515 21477
rect 29457 21437 29469 21471
rect 29503 21437 29515 21471
rect 29457 21431 29515 21437
rect 26694 21360 26700 21412
rect 26752 21360 26758 21412
rect 28169 21403 28227 21409
rect 28169 21369 28181 21403
rect 28215 21400 28227 21403
rect 28350 21400 28356 21412
rect 28215 21372 28356 21400
rect 28215 21369 28227 21372
rect 28169 21363 28227 21369
rect 28350 21360 28356 21372
rect 28408 21360 28414 21412
rect 29380 21400 29408 21431
rect 30098 21428 30104 21480
rect 30156 21468 30162 21480
rect 30193 21471 30251 21477
rect 30193 21468 30205 21471
rect 30156 21440 30205 21468
rect 30156 21428 30162 21440
rect 30193 21437 30205 21440
rect 30239 21437 30251 21471
rect 32867 21468 32895 21508
rect 32928 21505 32940 21539
rect 32928 21499 32956 21505
rect 32950 21496 32956 21499
rect 33008 21496 33014 21548
rect 33042 21496 33048 21548
rect 33100 21496 33106 21548
rect 33778 21496 33784 21548
rect 33836 21496 33842 21548
rect 33980 21545 34008 21576
rect 35452 21548 35480 21576
rect 33965 21539 34023 21545
rect 33965 21505 33977 21539
rect 34011 21505 34023 21539
rect 33965 21499 34023 21505
rect 34425 21539 34483 21545
rect 34425 21505 34437 21539
rect 34471 21505 34483 21539
rect 34425 21499 34483 21505
rect 32867 21440 33456 21468
rect 30193 21431 30251 21437
rect 28828 21372 29408 21400
rect 24026 21332 24032 21344
rect 22480 21304 24032 21332
rect 19521 21295 19579 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 26973 21335 27031 21341
rect 26973 21301 26985 21335
rect 27019 21332 27031 21335
rect 27614 21332 27620 21344
rect 27019 21304 27620 21332
rect 27019 21301 27031 21304
rect 26973 21295 27031 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 28258 21292 28264 21344
rect 28316 21332 28322 21344
rect 28828 21332 28856 21372
rect 33318 21360 33324 21412
rect 33376 21360 33382 21412
rect 33428 21400 33456 21440
rect 33594 21428 33600 21480
rect 33652 21468 33658 21480
rect 34440 21468 34468 21499
rect 35434 21496 35440 21548
rect 35492 21496 35498 21548
rect 35704 21539 35762 21545
rect 35704 21505 35716 21539
rect 35750 21536 35762 21539
rect 35986 21536 35992 21548
rect 35750 21508 35992 21536
rect 35750 21505 35762 21508
rect 35704 21499 35762 21505
rect 35986 21496 35992 21508
rect 36044 21496 36050 21548
rect 33652 21440 34468 21468
rect 34609 21471 34667 21477
rect 33652 21428 33658 21440
rect 34609 21437 34621 21471
rect 34655 21437 34667 21471
rect 36740 21468 36768 21576
rect 38304 21576 38568 21604
rect 36814 21496 36820 21548
rect 36872 21536 36878 21548
rect 37277 21539 37335 21545
rect 37277 21536 37289 21539
rect 36872 21508 37289 21536
rect 36872 21496 36878 21508
rect 37277 21505 37289 21508
rect 37323 21505 37335 21539
rect 37277 21499 37335 21505
rect 38197 21471 38255 21477
rect 38197 21468 38209 21471
rect 36740 21440 38209 21468
rect 34609 21431 34667 21437
rect 38197 21437 38209 21440
rect 38243 21468 38255 21471
rect 38304 21468 38332 21576
rect 38562 21564 38568 21576
rect 38620 21604 38626 21616
rect 41386 21604 41414 21644
rect 43438 21632 43444 21644
rect 43496 21632 43502 21684
rect 45186 21672 45192 21684
rect 44560 21644 45192 21672
rect 38620 21576 41414 21604
rect 38620 21564 38626 21576
rect 38464 21539 38522 21545
rect 38464 21505 38476 21539
rect 38510 21536 38522 21539
rect 39206 21536 39212 21548
rect 38510 21508 39212 21536
rect 38510 21505 38522 21508
rect 38464 21499 38522 21505
rect 39206 21496 39212 21508
rect 39264 21496 39270 21548
rect 40034 21496 40040 21548
rect 40092 21536 40098 21548
rect 40770 21536 40776 21548
rect 40092 21508 40776 21536
rect 40092 21496 40098 21508
rect 40770 21496 40776 21508
rect 40828 21496 40834 21548
rect 40880 21545 40908 21576
rect 42702 21564 42708 21616
rect 42760 21564 42766 21616
rect 40865 21539 40923 21545
rect 40865 21505 40877 21539
rect 40911 21505 40923 21539
rect 40865 21499 40923 21505
rect 41132 21539 41190 21545
rect 41132 21505 41144 21539
rect 41178 21536 41190 21539
rect 41506 21536 41512 21548
rect 41178 21508 41512 21536
rect 41178 21505 41190 21508
rect 41132 21499 41190 21505
rect 41506 21496 41512 21508
rect 41564 21496 41570 21548
rect 43622 21496 43628 21548
rect 43680 21545 43686 21548
rect 43680 21539 43729 21545
rect 43680 21505 43683 21539
rect 43717 21505 43729 21539
rect 43680 21499 43729 21505
rect 43680 21496 43686 21499
rect 43806 21496 43812 21548
rect 43864 21496 43870 21548
rect 44560 21545 44588 21644
rect 45186 21632 45192 21644
rect 45244 21632 45250 21684
rect 45554 21632 45560 21684
rect 45612 21632 45618 21684
rect 49050 21632 49056 21684
rect 49108 21632 49114 21684
rect 49142 21632 49148 21684
rect 49200 21632 49206 21684
rect 51166 21632 51172 21684
rect 51224 21632 51230 21684
rect 52546 21632 52552 21684
rect 52604 21632 52610 21684
rect 52730 21632 52736 21684
rect 52788 21632 52794 21684
rect 54018 21632 54024 21684
rect 54076 21672 54082 21684
rect 54113 21675 54171 21681
rect 54113 21672 54125 21675
rect 54076 21644 54125 21672
rect 54076 21632 54082 21644
rect 54113 21641 54125 21644
rect 54159 21641 54171 21675
rect 54113 21635 54171 21641
rect 54202 21632 54208 21684
rect 54260 21632 54266 21684
rect 45278 21604 45284 21616
rect 44744 21576 45284 21604
rect 44744 21545 44772 21576
rect 45278 21564 45284 21576
rect 45336 21604 45342 21616
rect 45649 21607 45707 21613
rect 45649 21604 45661 21607
rect 45336 21576 45661 21604
rect 45336 21564 45342 21576
rect 45649 21573 45661 21576
rect 45695 21573 45707 21607
rect 45649 21567 45707 21573
rect 48777 21607 48835 21613
rect 48777 21573 48789 21607
rect 48823 21604 48835 21607
rect 49160 21604 49188 21632
rect 48823 21576 49188 21604
rect 48823 21573 48835 21576
rect 48777 21567 48835 21573
rect 52914 21564 52920 21616
rect 52972 21604 52978 21616
rect 52972 21576 53512 21604
rect 52972 21564 52978 21576
rect 44545 21539 44603 21545
rect 44545 21505 44557 21539
rect 44591 21505 44603 21539
rect 44545 21499 44603 21505
rect 44729 21539 44787 21545
rect 44729 21505 44741 21539
rect 44775 21505 44787 21539
rect 44729 21499 44787 21505
rect 44928 21508 45508 21536
rect 44928 21480 44956 21508
rect 38243 21440 38332 21468
rect 38243 21437 38255 21440
rect 38197 21431 38255 21437
rect 34624 21400 34652 21431
rect 40126 21428 40132 21480
rect 40184 21428 40190 21480
rect 40313 21471 40371 21477
rect 40313 21437 40325 21471
rect 40359 21468 40371 21471
rect 43533 21471 43591 21477
rect 40359 21440 40816 21468
rect 40359 21437 40371 21440
rect 40313 21431 40371 21437
rect 33428 21372 33824 21400
rect 33796 21344 33824 21372
rect 34072 21372 34652 21400
rect 34072 21344 34100 21372
rect 28316 21304 28856 21332
rect 28905 21335 28963 21341
rect 28316 21292 28322 21304
rect 28905 21301 28917 21335
rect 28951 21332 28963 21335
rect 29270 21332 29276 21344
rect 28951 21304 29276 21332
rect 28951 21301 28963 21304
rect 28905 21295 28963 21301
rect 29270 21292 29276 21304
rect 29328 21292 29334 21344
rect 31846 21292 31852 21344
rect 31904 21292 31910 21344
rect 32125 21335 32183 21341
rect 32125 21301 32137 21335
rect 32171 21332 32183 21335
rect 33502 21332 33508 21344
rect 32171 21304 33508 21332
rect 32171 21301 32183 21304
rect 32125 21295 32183 21301
rect 33502 21292 33508 21304
rect 33560 21292 33566 21344
rect 33778 21292 33784 21344
rect 33836 21292 33842 21344
rect 34054 21292 34060 21344
rect 34112 21292 34118 21344
rect 34624 21332 34652 21372
rect 40788 21344 40816 21440
rect 43533 21437 43545 21471
rect 43579 21468 43591 21471
rect 44818 21468 44824 21480
rect 43579 21440 44824 21468
rect 43579 21437 43591 21440
rect 43533 21431 43591 21437
rect 44818 21428 44824 21440
rect 44876 21428 44882 21480
rect 44910 21428 44916 21480
rect 44968 21428 44974 21480
rect 45002 21428 45008 21480
rect 45060 21468 45066 21480
rect 45097 21471 45155 21477
rect 45097 21468 45109 21471
rect 45060 21440 45109 21468
rect 45060 21428 45066 21440
rect 45097 21437 45109 21440
rect 45143 21468 45155 21471
rect 45370 21468 45376 21480
rect 45143 21440 45376 21468
rect 45143 21437 45155 21440
rect 45097 21431 45155 21437
rect 45370 21428 45376 21440
rect 45428 21428 45434 21480
rect 45480 21468 45508 21508
rect 45554 21496 45560 21548
rect 45612 21536 45618 21548
rect 46201 21539 46259 21545
rect 46201 21536 46213 21539
rect 45612 21508 46213 21536
rect 45612 21496 45618 21508
rect 46201 21505 46213 21508
rect 46247 21505 46259 21539
rect 46201 21499 46259 21505
rect 47946 21496 47952 21548
rect 48004 21536 48010 21548
rect 48133 21539 48191 21545
rect 48133 21536 48145 21539
rect 48004 21508 48145 21536
rect 48004 21496 48010 21508
rect 48133 21505 48145 21508
rect 48179 21505 48191 21539
rect 48133 21499 48191 21505
rect 49234 21496 49240 21548
rect 49292 21536 49298 21548
rect 49605 21539 49663 21545
rect 49605 21536 49617 21539
rect 49292 21508 49617 21536
rect 49292 21496 49298 21508
rect 49605 21505 49617 21508
rect 49651 21505 49663 21539
rect 49605 21499 49663 21505
rect 50890 21496 50896 21548
rect 50948 21536 50954 21548
rect 51721 21539 51779 21545
rect 51721 21536 51733 21539
rect 50948 21508 51733 21536
rect 50948 21496 50954 21508
rect 51721 21505 51733 21508
rect 51767 21505 51779 21539
rect 51721 21499 51779 21505
rect 53282 21496 53288 21548
rect 53340 21496 53346 21548
rect 53484 21545 53512 21576
rect 53469 21539 53527 21545
rect 53469 21505 53481 21539
rect 53515 21505 53527 21539
rect 53469 21499 53527 21505
rect 54110 21496 54116 21548
rect 54168 21536 54174 21548
rect 54757 21539 54815 21545
rect 54757 21536 54769 21539
rect 54168 21508 54769 21536
rect 54168 21496 54174 21508
rect 54757 21505 54769 21508
rect 54803 21505 54815 21539
rect 54757 21499 54815 21505
rect 45480 21440 50108 21468
rect 42245 21403 42303 21409
rect 42245 21369 42257 21403
rect 42291 21400 42303 21403
rect 42426 21400 42432 21412
rect 42291 21372 42432 21400
rect 42291 21369 42303 21372
rect 42245 21363 42303 21369
rect 42426 21360 42432 21372
rect 42484 21360 42490 21412
rect 44085 21403 44143 21409
rect 44085 21369 44097 21403
rect 44131 21400 44143 21403
rect 45554 21400 45560 21412
rect 44131 21372 45560 21400
rect 44131 21369 44143 21372
rect 44085 21363 44143 21369
rect 45554 21360 45560 21372
rect 45612 21400 45618 21412
rect 48958 21400 48964 21412
rect 45612 21372 48964 21400
rect 45612 21360 45618 21372
rect 48958 21360 48964 21372
rect 49016 21400 49022 21412
rect 49326 21400 49332 21412
rect 49016 21372 49332 21400
rect 49016 21360 49022 21372
rect 49326 21360 49332 21372
rect 49384 21360 49390 21412
rect 40402 21332 40408 21344
rect 34624 21304 40408 21332
rect 40402 21292 40408 21304
rect 40460 21292 40466 21344
rect 40770 21292 40776 21344
rect 40828 21292 40834 21344
rect 42889 21335 42947 21341
rect 42889 21301 42901 21335
rect 42935 21332 42947 21335
rect 44726 21332 44732 21344
rect 42935 21304 44732 21332
rect 42935 21301 42947 21304
rect 42889 21295 42947 21301
rect 44726 21292 44732 21304
rect 44784 21292 44790 21344
rect 46566 21292 46572 21344
rect 46624 21332 46630 21344
rect 46661 21335 46719 21341
rect 46661 21332 46673 21335
rect 46624 21304 46673 21332
rect 46624 21292 46630 21304
rect 46661 21301 46673 21304
rect 46707 21332 46719 21335
rect 48590 21332 48596 21344
rect 46707 21304 48596 21332
rect 46707 21301 46719 21304
rect 46661 21295 46719 21301
rect 48590 21292 48596 21304
rect 48648 21292 48654 21344
rect 50080 21341 50108 21440
rect 55214 21400 55220 21412
rect 51046 21372 55220 21400
rect 50065 21335 50123 21341
rect 50065 21301 50077 21335
rect 50111 21332 50123 21335
rect 50154 21332 50160 21344
rect 50111 21304 50160 21332
rect 50111 21301 50123 21304
rect 50065 21295 50123 21301
rect 50154 21292 50160 21304
rect 50212 21332 50218 21344
rect 51046 21332 51074 21372
rect 55214 21360 55220 21372
rect 55272 21360 55278 21412
rect 50212 21304 51074 21332
rect 50212 21292 50218 21304
rect 1104 21242 58880 21264
rect 1104 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 22616 21242
rect 22668 21190 22680 21242
rect 22732 21190 22744 21242
rect 22796 21190 22808 21242
rect 22860 21190 22872 21242
rect 22924 21190 37060 21242
rect 37112 21190 37124 21242
rect 37176 21190 37188 21242
rect 37240 21190 37252 21242
rect 37304 21190 37316 21242
rect 37368 21190 51504 21242
rect 51556 21190 51568 21242
rect 51620 21190 51632 21242
rect 51684 21190 51696 21242
rect 51748 21190 51760 21242
rect 51812 21190 58880 21242
rect 1104 21168 58880 21190
rect 3973 21131 4031 21137
rect 3973 21097 3985 21131
rect 4019 21128 4031 21131
rect 4430 21128 4436 21140
rect 4019 21100 4436 21128
rect 4019 21097 4031 21100
rect 3973 21091 4031 21097
rect 4430 21088 4436 21100
rect 4488 21088 4494 21140
rect 7193 21131 7251 21137
rect 5276 21100 6408 21128
rect 5276 21072 5304 21100
rect 5258 21060 5264 21072
rect 4448 21032 5264 21060
rect 4448 21001 4476 21032
rect 5258 21020 5264 21032
rect 5316 21020 5322 21072
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 4525 20995 4583 21001
rect 4525 20961 4537 20995
rect 4571 20961 4583 20995
rect 4525 20955 4583 20961
rect 4540 20924 4568 20955
rect 4614 20952 4620 21004
rect 4672 20992 4678 21004
rect 6043 20995 6101 21001
rect 6043 20992 6055 20995
rect 4672 20964 6055 20992
rect 4672 20952 4678 20964
rect 6043 20961 6055 20964
rect 6089 20961 6101 20995
rect 6043 20955 6101 20961
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20992 6239 20995
rect 6380 20992 6408 21100
rect 7193 21097 7205 21131
rect 7239 21128 7251 21131
rect 7742 21128 7748 21140
rect 7239 21100 7748 21128
rect 7239 21097 7251 21100
rect 7193 21091 7251 21097
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 7926 21088 7932 21140
rect 7984 21088 7990 21140
rect 12434 21128 12440 21140
rect 10796 21100 12440 21128
rect 7944 21060 7972 21088
rect 7668 21032 7972 21060
rect 6227 20964 6408 20992
rect 6457 20995 6515 21001
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 6457 20961 6469 20995
rect 6503 20992 6515 20995
rect 7006 20992 7012 21004
rect 6503 20964 7012 20992
rect 6503 20961 6515 20964
rect 6457 20955 6515 20961
rect 7006 20952 7012 20964
rect 7064 20952 7070 21004
rect 7098 20952 7104 21004
rect 7156 20952 7162 21004
rect 4982 20924 4988 20936
rect 4540 20896 4988 20924
rect 4982 20884 4988 20896
rect 5040 20884 5046 20936
rect 5902 20884 5908 20936
rect 5960 20884 5966 20936
rect 6917 20927 6975 20933
rect 6917 20893 6929 20927
rect 6963 20924 6975 20927
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 6963 20896 7573 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 7561 20893 7573 20896
rect 7607 20924 7619 20927
rect 7668 20924 7696 21032
rect 10796 21001 10824 21100
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 16850 21088 16856 21140
rect 16908 21088 16914 21140
rect 22186 21128 22192 21140
rect 22066 21100 22192 21128
rect 10870 21020 10876 21072
rect 10928 21060 10934 21072
rect 10928 21032 11376 21060
rect 10928 21020 10934 21032
rect 7837 20995 7895 21001
rect 7837 20961 7849 20995
rect 7883 20961 7895 20995
rect 7837 20955 7895 20961
rect 10781 20995 10839 21001
rect 10781 20961 10793 20995
rect 10827 20961 10839 20995
rect 11146 20992 11152 21004
rect 10781 20955 10839 20961
rect 10888 20964 11152 20992
rect 7607 20896 7696 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 7852 20856 7880 20955
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9030 20924 9036 20936
rect 8987 20896 9036 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9030 20884 9036 20896
rect 9088 20884 9094 20936
rect 10597 20927 10655 20933
rect 9140 20896 10456 20924
rect 8297 20859 8355 20865
rect 8297 20856 8309 20859
rect 7852 20828 8309 20856
rect 8297 20825 8309 20828
rect 8343 20856 8355 20859
rect 9140 20856 9168 20896
rect 8343 20828 9168 20856
rect 9208 20859 9266 20865
rect 8343 20825 8355 20828
rect 8297 20819 8355 20825
rect 9208 20825 9220 20859
rect 9254 20856 9266 20859
rect 9306 20856 9312 20868
rect 9254 20828 9312 20856
rect 9254 20825 9266 20828
rect 9208 20819 9266 20825
rect 9306 20816 9312 20828
rect 9364 20816 9370 20868
rect 4246 20748 4252 20800
rect 4304 20788 4310 20800
rect 4341 20791 4399 20797
rect 4341 20788 4353 20791
rect 4304 20760 4353 20788
rect 4304 20748 4310 20760
rect 4341 20757 4353 20760
rect 4387 20757 4399 20791
rect 4341 20751 4399 20757
rect 5261 20791 5319 20797
rect 5261 20757 5273 20791
rect 5307 20788 5319 20791
rect 6086 20788 6092 20800
rect 5307 20760 6092 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 6178 20748 6184 20800
rect 6236 20788 6242 20800
rect 7653 20791 7711 20797
rect 7653 20788 7665 20791
rect 6236 20760 7665 20788
rect 6236 20748 6242 20760
rect 7653 20757 7665 20760
rect 7699 20757 7711 20791
rect 7653 20751 7711 20757
rect 8665 20791 8723 20797
rect 8665 20757 8677 20791
rect 8711 20788 8723 20791
rect 8754 20788 8760 20800
rect 8711 20760 8760 20788
rect 8711 20757 8723 20760
rect 8665 20751 8723 20757
rect 8754 20748 8760 20760
rect 8812 20748 8818 20800
rect 10318 20748 10324 20800
rect 10376 20748 10382 20800
rect 10428 20788 10456 20896
rect 10597 20893 10609 20927
rect 10643 20924 10655 20927
rect 10888 20924 10916 20964
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 11238 20952 11244 21004
rect 11296 20952 11302 21004
rect 11348 20992 11376 21032
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 16666 21060 16672 21072
rect 14332 21032 16672 21060
rect 14332 21020 14338 21032
rect 16666 21020 16672 21032
rect 16724 21020 16730 21072
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 11348 20964 11529 20992
rect 11517 20961 11529 20964
rect 11563 20961 11575 20995
rect 11517 20955 11575 20961
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 15378 20992 15384 21004
rect 11848 20964 15384 20992
rect 11848 20952 11854 20964
rect 15378 20952 15384 20964
rect 15436 20952 15442 21004
rect 16390 20952 16396 21004
rect 16448 20952 16454 21004
rect 10643 20896 10916 20924
rect 10643 20893 10655 20896
rect 10597 20887 10655 20893
rect 11606 20884 11612 20936
rect 11664 20933 11670 20936
rect 11664 20927 11692 20933
rect 11680 20893 11692 20927
rect 11664 20887 11692 20893
rect 11664 20884 11670 20887
rect 15010 20884 15016 20936
rect 15068 20884 15074 20936
rect 15286 20884 15292 20936
rect 15344 20884 15350 20936
rect 16408 20856 16436 20952
rect 16868 20933 16896 21088
rect 20625 21063 20683 21069
rect 20625 21029 20637 21063
rect 20671 21060 20683 21063
rect 20671 21032 21588 21060
rect 20671 21029 20683 21032
rect 20625 21023 20683 21029
rect 17037 20995 17095 21001
rect 17037 20961 17049 20995
rect 17083 20961 17095 20995
rect 17037 20955 17095 20961
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 17052 20856 17080 20955
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 21177 20995 21235 21001
rect 21177 20992 21189 20995
rect 20772 20964 21189 20992
rect 20772 20952 20778 20964
rect 17954 20884 17960 20936
rect 18012 20884 18018 20936
rect 18874 20884 18880 20936
rect 18932 20924 18938 20936
rect 19242 20924 19248 20936
rect 18932 20896 19248 20924
rect 18932 20884 18938 20896
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 16408 20828 17080 20856
rect 19512 20859 19570 20865
rect 19512 20825 19524 20859
rect 19558 20856 19570 20859
rect 20162 20856 20168 20868
rect 19558 20828 20168 20856
rect 19558 20825 19570 20828
rect 19512 20819 19570 20825
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 12066 20788 12072 20800
rect 10428 20760 12072 20788
rect 12066 20748 12072 20760
rect 12124 20748 12130 20800
rect 12437 20791 12495 20797
rect 12437 20757 12449 20791
rect 12483 20788 12495 20791
rect 13906 20788 13912 20800
rect 12483 20760 13912 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 14461 20791 14519 20797
rect 14461 20788 14473 20791
rect 14424 20760 14473 20788
rect 14424 20748 14430 20760
rect 14461 20757 14473 20760
rect 14507 20757 14519 20791
rect 14461 20751 14519 20757
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 16482 20748 16488 20800
rect 16540 20748 16546 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17402 20748 17408 20800
rect 17460 20748 17466 20800
rect 20714 20748 20720 20800
rect 20772 20748 20778 20800
rect 21008 20788 21036 20964
rect 21177 20961 21189 20964
rect 21223 20961 21235 20995
rect 21177 20955 21235 20961
rect 21266 20952 21272 21004
rect 21324 20952 21330 21004
rect 21560 21001 21588 21032
rect 21545 20995 21603 21001
rect 21545 20961 21557 20995
rect 21591 20961 21603 20995
rect 21545 20955 21603 20961
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20924 21143 20927
rect 22066 20924 22094 21100
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 22278 21088 22284 21140
rect 22336 21088 22342 21140
rect 23385 21131 23443 21137
rect 23385 21097 23397 21131
rect 23431 21128 23443 21131
rect 24026 21128 24032 21140
rect 23431 21100 24032 21128
rect 23431 21097 23443 21100
rect 23385 21091 23443 21097
rect 24026 21088 24032 21100
rect 24084 21088 24090 21140
rect 25314 21128 25320 21140
rect 25056 21100 25320 21128
rect 22925 20995 22983 21001
rect 22925 20961 22937 20995
rect 22971 20992 22983 20995
rect 23382 20992 23388 21004
rect 22971 20964 23388 20992
rect 22971 20961 22983 20964
rect 22925 20955 22983 20961
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 25056 21001 25084 21100
rect 25314 21088 25320 21100
rect 25372 21088 25378 21140
rect 29362 21088 29368 21140
rect 29420 21088 29426 21140
rect 31846 21088 31852 21140
rect 31904 21088 31910 21140
rect 32214 21088 32220 21140
rect 32272 21088 32278 21140
rect 33318 21128 33324 21140
rect 32600 21100 33324 21128
rect 31864 21060 31892 21088
rect 32600 21060 32628 21100
rect 33318 21088 33324 21100
rect 33376 21088 33382 21140
rect 33962 21088 33968 21140
rect 34020 21088 34026 21140
rect 34698 21088 34704 21140
rect 34756 21088 34762 21140
rect 36354 21088 36360 21140
rect 36412 21088 36418 21140
rect 38562 21088 38568 21140
rect 38620 21128 38626 21140
rect 39209 21131 39267 21137
rect 39209 21128 39221 21131
rect 38620 21100 39221 21128
rect 38620 21088 38626 21100
rect 39209 21097 39221 21100
rect 39255 21097 39267 21131
rect 39209 21091 39267 21097
rect 31864 21032 32628 21060
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 27065 20995 27123 21001
rect 27065 20961 27077 20995
rect 27111 20961 27123 20995
rect 27065 20955 27123 20961
rect 21131 20896 22094 20924
rect 22741 20927 22799 20933
rect 21131 20893 21143 20896
rect 21085 20887 21143 20893
rect 22741 20893 22753 20927
rect 22787 20924 22799 20927
rect 23198 20924 23204 20936
rect 22787 20896 23204 20924
rect 22787 20893 22799 20896
rect 22741 20887 22799 20893
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 27080 20924 27108 20955
rect 27982 20952 27988 21004
rect 28040 20952 28046 21004
rect 32582 20992 32588 21004
rect 31404 20964 32588 20992
rect 27525 20927 27583 20933
rect 27525 20924 27537 20927
rect 25240 20896 27537 20924
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 25240 20856 25268 20896
rect 27525 20893 27537 20896
rect 27571 20893 27583 20927
rect 27525 20887 27583 20893
rect 29638 20884 29644 20936
rect 29696 20924 29702 20936
rect 30098 20924 30104 20936
rect 29696 20896 30104 20924
rect 29696 20884 29702 20896
rect 30098 20884 30104 20896
rect 30156 20924 30162 20936
rect 31404 20924 31432 20964
rect 32582 20952 32588 20964
rect 32640 20952 32646 21004
rect 31573 20927 31631 20933
rect 31573 20924 31585 20927
rect 30156 20896 31432 20924
rect 31496 20896 31585 20924
rect 30156 20884 30162 20896
rect 21324 20828 25268 20856
rect 25308 20859 25366 20865
rect 21324 20816 21330 20828
rect 25308 20825 25320 20859
rect 25354 20856 25366 20859
rect 25958 20856 25964 20868
rect 25354 20828 25964 20856
rect 25354 20825 25366 20828
rect 25308 20819 25366 20825
rect 25958 20816 25964 20828
rect 26016 20816 26022 20868
rect 26881 20859 26939 20865
rect 26881 20825 26893 20859
rect 26927 20856 26939 20859
rect 27798 20856 27804 20868
rect 26927 20828 27804 20856
rect 26927 20825 26939 20828
rect 26881 20819 26939 20825
rect 27798 20816 27804 20828
rect 27856 20816 27862 20868
rect 28252 20859 28310 20865
rect 28252 20825 28264 20859
rect 28298 20856 28310 20859
rect 28718 20856 28724 20868
rect 28298 20828 28724 20856
rect 28298 20825 28310 20828
rect 28252 20819 28310 20825
rect 28718 20816 28724 20828
rect 28776 20816 28782 20868
rect 30368 20859 30426 20865
rect 30368 20825 30380 20859
rect 30414 20856 30426 20859
rect 30558 20856 30564 20868
rect 30414 20828 30564 20856
rect 30414 20825 30426 20828
rect 30368 20819 30426 20825
rect 30558 20816 30564 20828
rect 30616 20816 30622 20868
rect 22649 20791 22707 20797
rect 22649 20788 22661 20791
rect 21008 20760 22661 20788
rect 22649 20757 22661 20760
rect 22695 20788 22707 20791
rect 23106 20788 23112 20800
rect 22695 20760 23112 20788
rect 22695 20757 22707 20760
rect 22649 20751 22707 20757
rect 23106 20748 23112 20760
rect 23164 20748 23170 20800
rect 26418 20748 26424 20800
rect 26476 20748 26482 20800
rect 26510 20748 26516 20800
rect 26568 20748 26574 20800
rect 26970 20748 26976 20800
rect 27028 20748 27034 20800
rect 31496 20797 31524 20896
rect 31573 20893 31585 20896
rect 31619 20893 31631 20927
rect 31573 20887 31631 20893
rect 32852 20927 32910 20933
rect 32852 20893 32864 20927
rect 32898 20924 32910 20927
rect 34716 20924 34744 21088
rect 37642 21020 37648 21072
rect 37700 21060 37706 21072
rect 38378 21060 38384 21072
rect 37700 21032 38384 21060
rect 37700 21020 37706 21032
rect 38378 21020 38384 21032
rect 38436 21020 38442 21072
rect 36906 20952 36912 21004
rect 36964 20952 36970 21004
rect 39224 20992 39252 21091
rect 40402 21088 40408 21140
rect 40460 21088 40466 21140
rect 43806 21088 43812 21140
rect 43864 21128 43870 21140
rect 44177 21131 44235 21137
rect 44177 21128 44189 21131
rect 43864 21100 44189 21128
rect 43864 21088 43870 21100
rect 44177 21097 44189 21100
rect 44223 21097 44235 21131
rect 44177 21091 44235 21097
rect 44818 21088 44824 21140
rect 44876 21128 44882 21140
rect 45186 21128 45192 21140
rect 44876 21100 45192 21128
rect 44876 21088 44882 21100
rect 45186 21088 45192 21100
rect 45244 21088 45250 21140
rect 45554 21088 45560 21140
rect 45612 21088 45618 21140
rect 49050 21088 49056 21140
rect 49108 21128 49114 21140
rect 49510 21128 49516 21140
rect 49108 21100 49516 21128
rect 49108 21088 49114 21100
rect 49510 21088 49516 21100
rect 49568 21128 49574 21140
rect 53929 21131 53987 21137
rect 53929 21128 53941 21131
rect 49568 21100 53941 21128
rect 49568 21088 49574 21100
rect 53929 21097 53941 21100
rect 53975 21128 53987 21131
rect 54662 21128 54668 21140
rect 53975 21100 54668 21128
rect 53975 21097 53987 21100
rect 53929 21091 53987 21097
rect 54662 21088 54668 21100
rect 54720 21088 54726 21140
rect 42705 21063 42763 21069
rect 42705 21029 42717 21063
rect 42751 21060 42763 21063
rect 44729 21063 44787 21069
rect 42751 21032 43576 21060
rect 42751 21029 42763 21032
rect 42705 21023 42763 21029
rect 41325 20995 41383 21001
rect 41325 20992 41337 20995
rect 39224 20964 41337 20992
rect 41325 20961 41337 20964
rect 41371 20961 41383 20995
rect 41325 20955 41383 20961
rect 42610 20952 42616 21004
rect 42668 20992 42674 21004
rect 43548 21001 43576 21032
rect 44729 21029 44741 21063
rect 44775 21060 44787 21063
rect 44910 21060 44916 21072
rect 44775 21032 44916 21060
rect 44775 21029 44787 21032
rect 44729 21023 44787 21029
rect 43349 20995 43407 21001
rect 43349 20992 43361 20995
rect 42668 20964 43361 20992
rect 42668 20952 42674 20964
rect 43349 20961 43361 20964
rect 43395 20961 43407 20995
rect 43349 20955 43407 20961
rect 43533 20995 43591 21001
rect 43533 20961 43545 20995
rect 43579 20961 43591 20995
rect 43533 20955 43591 20961
rect 32898 20896 34744 20924
rect 32898 20893 32910 20896
rect 32852 20887 32910 20893
rect 40770 20884 40776 20936
rect 40828 20924 40834 20936
rect 44744 20924 44772 21023
rect 44910 21020 44916 21032
rect 44968 21020 44974 21072
rect 54478 21020 54484 21072
rect 54536 21060 54542 21072
rect 54941 21063 54999 21069
rect 54941 21060 54953 21063
rect 54536 21032 54953 21060
rect 54536 21020 54542 21032
rect 54941 21029 54953 21032
rect 54987 21060 54999 21063
rect 56502 21060 56508 21072
rect 54987 21032 56508 21060
rect 54987 21029 54999 21032
rect 54941 21023 54999 21029
rect 56502 21020 56508 21032
rect 56560 21020 56566 21072
rect 48130 20952 48136 21004
rect 48188 20992 48194 21004
rect 48774 20992 48780 21004
rect 48188 20964 48780 20992
rect 48188 20952 48194 20964
rect 48774 20952 48780 20964
rect 48832 20992 48838 21004
rect 54573 20995 54631 21001
rect 54573 20992 54585 20995
rect 48832 20964 54585 20992
rect 48832 20952 48838 20964
rect 54573 20961 54585 20964
rect 54619 20992 54631 20995
rect 55214 20992 55220 21004
rect 54619 20964 55220 20992
rect 54619 20961 54631 20964
rect 54573 20955 54631 20961
rect 55214 20952 55220 20964
rect 55272 20952 55278 21004
rect 40828 20896 44772 20924
rect 40828 20884 40834 20896
rect 55858 20884 55864 20936
rect 55916 20884 55922 20936
rect 56042 20884 56048 20936
rect 56100 20884 56106 20936
rect 57330 20884 57336 20936
rect 57388 20884 57394 20936
rect 37921 20859 37979 20865
rect 37921 20856 37933 20859
rect 37844 20828 37933 20856
rect 37844 20800 37872 20828
rect 37921 20825 37933 20828
rect 37967 20856 37979 20859
rect 40037 20859 40095 20865
rect 40037 20856 40049 20859
rect 37967 20828 40049 20856
rect 37967 20825 37979 20828
rect 37921 20819 37979 20825
rect 40037 20825 40049 20828
rect 40083 20825 40095 20859
rect 40037 20819 40095 20825
rect 41592 20859 41650 20865
rect 41592 20825 41604 20859
rect 41638 20856 41650 20859
rect 42797 20859 42855 20865
rect 42797 20856 42809 20859
rect 41638 20828 42809 20856
rect 41638 20825 41650 20828
rect 41592 20819 41650 20825
rect 42797 20825 42809 20828
rect 42843 20825 42855 20859
rect 55398 20856 55404 20868
rect 42797 20819 42855 20825
rect 53852 20828 55404 20856
rect 53852 20800 53880 20828
rect 55398 20816 55404 20828
rect 55456 20816 55462 20868
rect 31481 20791 31539 20797
rect 31481 20757 31493 20791
rect 31527 20757 31539 20791
rect 31481 20751 31539 20757
rect 33778 20748 33784 20800
rect 33836 20788 33842 20800
rect 34241 20791 34299 20797
rect 34241 20788 34253 20791
rect 33836 20760 34253 20788
rect 33836 20748 33842 20760
rect 34241 20757 34253 20760
rect 34287 20757 34299 20791
rect 34241 20751 34299 20757
rect 37826 20748 37832 20800
rect 37884 20748 37890 20800
rect 48590 20748 48596 20800
rect 48648 20788 48654 20800
rect 49050 20788 49056 20800
rect 48648 20760 49056 20788
rect 48648 20748 48654 20760
rect 49050 20748 49056 20760
rect 49108 20748 49114 20800
rect 52454 20748 52460 20800
rect 52512 20788 52518 20800
rect 53101 20791 53159 20797
rect 53101 20788 53113 20791
rect 52512 20760 53113 20788
rect 52512 20748 52518 20760
rect 53101 20757 53113 20760
rect 53147 20788 53159 20791
rect 53834 20788 53840 20800
rect 53147 20760 53840 20788
rect 53147 20757 53159 20760
rect 53101 20751 53159 20757
rect 53834 20748 53840 20760
rect 53892 20748 53898 20800
rect 55306 20748 55312 20800
rect 55364 20748 55370 20800
rect 56686 20748 56692 20800
rect 56744 20748 56750 20800
rect 56778 20748 56784 20800
rect 56836 20748 56842 20800
rect 1104 20698 59040 20720
rect 1104 20646 15394 20698
rect 15446 20646 15458 20698
rect 15510 20646 15522 20698
rect 15574 20646 15586 20698
rect 15638 20646 15650 20698
rect 15702 20646 29838 20698
rect 29890 20646 29902 20698
rect 29954 20646 29966 20698
rect 30018 20646 30030 20698
rect 30082 20646 30094 20698
rect 30146 20646 44282 20698
rect 44334 20646 44346 20698
rect 44398 20646 44410 20698
rect 44462 20646 44474 20698
rect 44526 20646 44538 20698
rect 44590 20646 58726 20698
rect 58778 20646 58790 20698
rect 58842 20646 58854 20698
rect 58906 20646 58918 20698
rect 58970 20646 58982 20698
rect 59034 20646 59040 20698
rect 1104 20624 59040 20646
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 6917 20587 6975 20593
rect 6917 20584 6929 20587
rect 6144 20556 6929 20584
rect 6144 20544 6150 20556
rect 6917 20553 6929 20556
rect 6963 20553 6975 20587
rect 6917 20547 6975 20553
rect 7006 20544 7012 20596
rect 7064 20584 7070 20596
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 7064 20556 7941 20584
rect 7064 20544 7070 20556
rect 7929 20553 7941 20556
rect 7975 20553 7987 20587
rect 7929 20547 7987 20553
rect 9769 20587 9827 20593
rect 9769 20553 9781 20587
rect 9815 20584 9827 20587
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 9815 20556 10885 20584
rect 9815 20553 9827 20556
rect 9769 20547 9827 20553
rect 10873 20553 10885 20556
rect 10919 20584 10931 20587
rect 11606 20584 11612 20596
rect 10919 20556 11612 20584
rect 10919 20553 10931 20556
rect 10873 20547 10931 20553
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 11790 20544 11796 20596
rect 11848 20544 11854 20596
rect 14461 20587 14519 20593
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 15010 20584 15016 20596
rect 14507 20556 15016 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 17313 20587 17371 20593
rect 17313 20553 17325 20587
rect 17359 20584 17371 20587
rect 17402 20584 17408 20596
rect 17359 20556 17408 20584
rect 17359 20553 17371 20556
rect 17313 20547 17371 20553
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 20162 20544 20168 20596
rect 20220 20544 20226 20596
rect 21082 20544 21088 20596
rect 21140 20544 21146 20596
rect 22462 20544 22468 20596
rect 22520 20584 22526 20596
rect 23290 20584 23296 20596
rect 22520 20556 23296 20584
rect 22520 20544 22526 20556
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 25958 20544 25964 20596
rect 26016 20544 26022 20596
rect 27617 20587 27675 20593
rect 27617 20553 27629 20587
rect 27663 20584 27675 20587
rect 27798 20584 27804 20596
rect 27663 20556 27804 20584
rect 27663 20553 27675 20556
rect 27617 20547 27675 20553
rect 27798 20544 27804 20556
rect 27856 20544 27862 20596
rect 27890 20544 27896 20596
rect 27948 20544 27954 20596
rect 28353 20587 28411 20593
rect 28353 20553 28365 20587
rect 28399 20584 28411 20587
rect 28442 20584 28448 20596
rect 28399 20556 28448 20584
rect 28399 20553 28411 20556
rect 28353 20547 28411 20553
rect 28442 20544 28448 20556
rect 28500 20544 28506 20596
rect 28718 20544 28724 20596
rect 28776 20544 28782 20596
rect 30558 20544 30564 20596
rect 30616 20544 30622 20596
rect 37642 20544 37648 20596
rect 37700 20544 37706 20596
rect 54662 20544 54668 20596
rect 54720 20584 54726 20596
rect 55309 20587 55367 20593
rect 55309 20584 55321 20587
rect 54720 20556 55321 20584
rect 54720 20544 54726 20556
rect 55309 20553 55321 20556
rect 55355 20553 55367 20587
rect 55309 20547 55367 20553
rect 55677 20587 55735 20593
rect 55677 20553 55689 20587
rect 55723 20584 55735 20587
rect 55858 20584 55864 20596
rect 55723 20556 55864 20584
rect 55723 20553 55735 20556
rect 55677 20547 55735 20553
rect 55858 20544 55864 20556
rect 55916 20544 55922 20596
rect 11241 20519 11299 20525
rect 11241 20485 11253 20519
rect 11287 20516 11299 20519
rect 11808 20516 11836 20544
rect 11287 20488 11836 20516
rect 11287 20485 11299 20488
rect 11241 20479 11299 20485
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 22189 20519 22247 20525
rect 22189 20516 22201 20519
rect 22152 20488 22201 20516
rect 22152 20476 22158 20488
rect 22189 20485 22201 20488
rect 22235 20516 22247 20519
rect 23382 20516 23388 20528
rect 22235 20488 23388 20516
rect 22235 20485 22247 20488
rect 22189 20479 22247 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 26970 20476 26976 20528
rect 27028 20516 27034 20528
rect 28258 20516 28264 20528
rect 27028 20488 28264 20516
rect 27028 20476 27034 20488
rect 28258 20476 28264 20488
rect 28316 20476 28322 20528
rect 44634 20476 44640 20528
rect 44692 20516 44698 20528
rect 50246 20516 50252 20528
rect 44692 20488 50252 20516
rect 44692 20476 44698 20488
rect 50246 20476 50252 20488
rect 50304 20476 50310 20528
rect 56588 20519 56646 20525
rect 54680 20488 56548 20516
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 9907 20420 10180 20448
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10152 20392 10180 20420
rect 10318 20408 10324 20460
rect 10376 20408 10382 20460
rect 14829 20451 14887 20457
rect 14829 20417 14841 20451
rect 14875 20448 14887 20451
rect 15838 20448 15844 20460
rect 14875 20420 15844 20448
rect 14875 20417 14887 20420
rect 14829 20411 14887 20417
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 17052 20420 18368 20448
rect 4522 20340 4528 20392
rect 4580 20340 4586 20392
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5960 20352 7021 20380
rect 5960 20340 5966 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20380 7251 20383
rect 7239 20352 7328 20380
rect 7239 20349 7251 20352
rect 7193 20343 7251 20349
rect 7300 20256 7328 20352
rect 10042 20340 10048 20392
rect 10100 20340 10106 20392
rect 10134 20340 10140 20392
rect 10192 20340 10198 20392
rect 14918 20340 14924 20392
rect 14976 20340 14982 20392
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 15028 20312 15056 20343
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 15252 20352 15485 20380
rect 15252 20340 15258 20352
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 15473 20343 15531 20349
rect 16022 20340 16028 20392
rect 16080 20380 16086 20392
rect 17052 20389 17080 20420
rect 16485 20383 16543 20389
rect 16485 20380 16497 20383
rect 16080 20352 16497 20380
rect 16080 20340 16086 20352
rect 16485 20349 16497 20352
rect 16531 20380 16543 20383
rect 17037 20383 17095 20389
rect 17037 20380 17049 20383
rect 16531 20352 17049 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 17037 20349 17049 20352
rect 17083 20349 17095 20383
rect 17037 20343 17095 20349
rect 17126 20340 17132 20392
rect 17184 20380 17190 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 17184 20352 17233 20380
rect 17184 20340 17190 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 18233 20383 18291 20389
rect 18233 20380 18245 20383
rect 17221 20343 17279 20349
rect 17696 20352 18245 20380
rect 17696 20321 17724 20352
rect 18233 20349 18245 20352
rect 18279 20349 18291 20383
rect 18340 20380 18368 20420
rect 20714 20408 20720 20460
rect 20772 20408 20778 20460
rect 26418 20408 26424 20460
rect 26476 20408 26482 20460
rect 26510 20408 26516 20460
rect 26568 20408 26574 20460
rect 29270 20408 29276 20460
rect 29328 20408 29334 20460
rect 30650 20408 30656 20460
rect 30708 20448 30714 20460
rect 31113 20451 31171 20457
rect 31113 20448 31125 20451
rect 30708 20420 31125 20448
rect 30708 20408 30714 20420
rect 31113 20417 31125 20420
rect 31159 20417 31171 20451
rect 54570 20448 54576 20460
rect 31113 20411 31171 20417
rect 49344 20420 54576 20448
rect 22462 20380 22468 20392
rect 18340 20352 22468 20380
rect 18233 20343 18291 20349
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 23474 20340 23480 20392
rect 23532 20340 23538 20392
rect 26436 20380 26464 20408
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26436 20352 26985 20380
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 28442 20340 28448 20392
rect 28500 20340 28506 20392
rect 45554 20340 45560 20392
rect 45612 20340 45618 20392
rect 48222 20340 48228 20392
rect 48280 20340 48286 20392
rect 48406 20340 48412 20392
rect 48464 20340 48470 20392
rect 49344 20324 49372 20420
rect 54570 20408 54576 20420
rect 54628 20408 54634 20460
rect 54202 20340 54208 20392
rect 54260 20340 54266 20392
rect 14292 20284 15056 20312
rect 16117 20315 16175 20321
rect 5074 20204 5080 20256
rect 5132 20204 5138 20256
rect 6546 20204 6552 20256
rect 6604 20204 6610 20256
rect 7282 20204 7288 20256
rect 7340 20244 7346 20256
rect 7561 20247 7619 20253
rect 7561 20244 7573 20247
rect 7340 20216 7573 20244
rect 7340 20204 7346 20216
rect 7561 20213 7573 20216
rect 7607 20213 7619 20247
rect 7561 20207 7619 20213
rect 9398 20204 9404 20256
rect 9456 20204 9462 20256
rect 14090 20204 14096 20256
rect 14148 20244 14154 20256
rect 14292 20253 14320 20284
rect 16117 20281 16129 20315
rect 16163 20312 16175 20315
rect 17681 20315 17739 20321
rect 16163 20284 16528 20312
rect 16163 20281 16175 20284
rect 16117 20275 16175 20281
rect 16500 20256 16528 20284
rect 17681 20281 17693 20315
rect 17727 20281 17739 20315
rect 49326 20312 49332 20324
rect 17681 20275 17739 20281
rect 44560 20284 49332 20312
rect 44560 20256 44588 20284
rect 49326 20272 49332 20284
rect 49384 20272 49390 20324
rect 50065 20315 50123 20321
rect 50065 20281 50077 20315
rect 50111 20312 50123 20315
rect 50246 20312 50252 20324
rect 50111 20284 50252 20312
rect 50111 20281 50123 20284
rect 50065 20275 50123 20281
rect 50246 20272 50252 20284
rect 50304 20312 50310 20324
rect 54680 20312 54708 20488
rect 55122 20448 55128 20460
rect 55048 20420 55128 20448
rect 55048 20389 55076 20420
rect 55122 20408 55128 20420
rect 55180 20408 55186 20460
rect 55398 20408 55404 20460
rect 55456 20448 55462 20460
rect 55953 20451 56011 20457
rect 55953 20448 55965 20451
rect 55456 20420 55965 20448
rect 55456 20408 55462 20420
rect 55953 20417 55965 20420
rect 55999 20417 56011 20451
rect 56520 20448 56548 20488
rect 56588 20485 56600 20519
rect 56634 20516 56646 20519
rect 56778 20516 56784 20528
rect 56634 20488 56784 20516
rect 56634 20485 56646 20488
rect 56588 20479 56646 20485
rect 56778 20476 56784 20488
rect 56836 20476 56842 20528
rect 56870 20448 56876 20460
rect 56520 20420 56876 20448
rect 55953 20411 56011 20417
rect 56870 20408 56876 20420
rect 56928 20408 56934 20460
rect 55033 20383 55091 20389
rect 55033 20349 55045 20383
rect 55079 20349 55091 20383
rect 55033 20343 55091 20349
rect 55217 20383 55275 20389
rect 55217 20349 55229 20383
rect 55263 20349 55275 20383
rect 55217 20343 55275 20349
rect 50304 20284 54708 20312
rect 50304 20272 50310 20284
rect 14277 20247 14335 20253
rect 14277 20244 14289 20247
rect 14148 20216 14289 20244
rect 14148 20204 14154 20216
rect 14277 20213 14289 20216
rect 14323 20213 14335 20247
rect 14277 20207 14335 20213
rect 16482 20204 16488 20256
rect 16540 20204 16546 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18656 20216 18889 20244
rect 18656 20204 18662 20216
rect 18877 20213 18889 20216
rect 18923 20213 18935 20247
rect 18877 20207 18935 20213
rect 22833 20247 22891 20253
rect 22833 20213 22845 20247
rect 22879 20244 22891 20247
rect 23014 20244 23020 20256
rect 22879 20216 23020 20244
rect 22879 20213 22891 20216
rect 22833 20207 22891 20213
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 38102 20204 38108 20256
rect 38160 20244 38166 20256
rect 38381 20247 38439 20253
rect 38381 20244 38393 20247
rect 38160 20216 38393 20244
rect 38160 20204 38166 20216
rect 38381 20213 38393 20216
rect 38427 20213 38439 20247
rect 38381 20207 38439 20213
rect 39758 20204 39764 20256
rect 39816 20204 39822 20256
rect 44542 20204 44548 20256
rect 44600 20204 44606 20256
rect 44818 20204 44824 20256
rect 44876 20204 44882 20256
rect 44913 20247 44971 20253
rect 44913 20213 44925 20247
rect 44959 20244 44971 20247
rect 45370 20244 45376 20256
rect 44959 20216 45376 20244
rect 44959 20213 44971 20216
rect 44913 20207 44971 20213
rect 45370 20204 45376 20216
rect 45428 20204 45434 20256
rect 47302 20204 47308 20256
rect 47360 20244 47366 20256
rect 47673 20247 47731 20253
rect 47673 20244 47685 20247
rect 47360 20216 47685 20244
rect 47360 20204 47366 20216
rect 47673 20213 47685 20216
rect 47719 20213 47731 20247
rect 47673 20207 47731 20213
rect 48682 20204 48688 20256
rect 48740 20244 48746 20256
rect 49053 20247 49111 20253
rect 49053 20244 49065 20247
rect 48740 20216 49065 20244
rect 48740 20204 48746 20216
rect 49053 20213 49065 20216
rect 49099 20213 49111 20247
rect 49053 20207 49111 20213
rect 53650 20204 53656 20256
rect 53708 20204 53714 20256
rect 55232 20244 55260 20343
rect 56318 20340 56324 20392
rect 56376 20340 56382 20392
rect 58437 20383 58495 20389
rect 58437 20380 58449 20383
rect 57716 20352 58449 20380
rect 57716 20321 57744 20352
rect 58437 20349 58449 20352
rect 58483 20349 58495 20383
rect 58437 20343 58495 20349
rect 57701 20315 57759 20321
rect 57701 20281 57713 20315
rect 57747 20281 57759 20315
rect 57701 20275 57759 20281
rect 56686 20244 56692 20256
rect 55232 20216 56692 20244
rect 56686 20204 56692 20216
rect 56744 20204 56750 20256
rect 57238 20204 57244 20256
rect 57296 20244 57302 20256
rect 57885 20247 57943 20253
rect 57885 20244 57897 20247
rect 57296 20216 57897 20244
rect 57296 20204 57302 20216
rect 57885 20213 57897 20216
rect 57931 20213 57943 20247
rect 57885 20207 57943 20213
rect 1104 20154 58880 20176
rect 1104 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 22616 20154
rect 22668 20102 22680 20154
rect 22732 20102 22744 20154
rect 22796 20102 22808 20154
rect 22860 20102 22872 20154
rect 22924 20102 37060 20154
rect 37112 20102 37124 20154
rect 37176 20102 37188 20154
rect 37240 20102 37252 20154
rect 37304 20102 37316 20154
rect 37368 20102 51504 20154
rect 51556 20102 51568 20154
rect 51620 20102 51632 20154
rect 51684 20102 51696 20154
rect 51748 20102 51760 20154
rect 51812 20102 58880 20154
rect 1104 20080 58880 20102
rect 4522 20000 4528 20052
rect 4580 20000 4586 20052
rect 8665 20043 8723 20049
rect 8665 20009 8677 20043
rect 8711 20040 8723 20043
rect 18690 20040 18696 20052
rect 8711 20012 18696 20040
rect 8711 20009 8723 20012
rect 8665 20003 8723 20009
rect 3973 19907 4031 19913
rect 3973 19873 3985 19907
rect 4019 19904 4031 19907
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 4019 19876 5733 19904
rect 4019 19873 4031 19876
rect 3973 19867 4031 19873
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 4798 19796 4804 19848
rect 4856 19796 4862 19848
rect 5736 19836 5764 19867
rect 6549 19839 6607 19845
rect 5736 19808 6500 19836
rect 4065 19771 4123 19777
rect 4065 19737 4077 19771
rect 4111 19768 4123 19771
rect 5445 19771 5503 19777
rect 5445 19768 5457 19771
rect 4111 19740 5457 19768
rect 4111 19737 4123 19740
rect 4065 19731 4123 19737
rect 5445 19737 5457 19740
rect 5491 19768 5503 19771
rect 6086 19768 6092 19780
rect 5491 19740 6092 19768
rect 5491 19737 5503 19740
rect 5445 19731 5503 19737
rect 6086 19728 6092 19740
rect 6144 19728 6150 19780
rect 6472 19768 6500 19808
rect 6549 19805 6561 19839
rect 6595 19836 6607 19839
rect 8680 19836 8708 20003
rect 18690 20000 18696 20012
rect 18748 20000 18754 20052
rect 21726 20000 21732 20052
rect 21784 20000 21790 20052
rect 23474 20000 23480 20052
rect 23532 20040 23538 20052
rect 23569 20043 23627 20049
rect 23569 20040 23581 20043
rect 23532 20012 23581 20040
rect 23532 20000 23538 20012
rect 23569 20009 23581 20012
rect 23615 20009 23627 20043
rect 23569 20003 23627 20009
rect 27801 20043 27859 20049
rect 27801 20009 27813 20043
rect 27847 20040 27859 20043
rect 28442 20040 28448 20052
rect 27847 20012 28448 20040
rect 27847 20009 27859 20012
rect 27801 20003 27859 20009
rect 9306 19932 9312 19984
rect 9364 19932 9370 19984
rect 9398 19932 9404 19984
rect 9456 19932 9462 19984
rect 10689 19975 10747 19981
rect 10689 19941 10701 19975
rect 10735 19972 10747 19975
rect 11238 19972 11244 19984
rect 10735 19944 11244 19972
rect 10735 19941 10747 19944
rect 10689 19935 10747 19941
rect 11238 19932 11244 19944
rect 11296 19932 11302 19984
rect 15286 19932 15292 19984
rect 15344 19972 15350 19984
rect 15473 19975 15531 19981
rect 15473 19972 15485 19975
rect 15344 19944 15485 19972
rect 15344 19932 15350 19944
rect 15473 19941 15485 19944
rect 15519 19941 15531 19975
rect 15473 19935 15531 19941
rect 16666 19932 16672 19984
rect 16724 19972 16730 19984
rect 16761 19975 16819 19981
rect 16761 19972 16773 19975
rect 16724 19944 16773 19972
rect 16724 19932 16730 19944
rect 16761 19941 16773 19944
rect 16807 19941 16819 19975
rect 16761 19935 16819 19941
rect 17402 19932 17408 19984
rect 17460 19932 17466 19984
rect 9416 19904 9444 19932
rect 9861 19907 9919 19913
rect 9861 19904 9873 19907
rect 9416 19876 9873 19904
rect 9861 19873 9873 19876
rect 9907 19873 9919 19907
rect 9861 19867 9919 19873
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13872 19876 14105 19904
rect 13872 19864 13878 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 16347 19907 16405 19913
rect 16347 19904 16359 19907
rect 15896 19876 16359 19904
rect 15896 19864 15902 19876
rect 16347 19873 16359 19876
rect 16393 19873 16405 19907
rect 16347 19867 16405 19873
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 17420 19904 17448 19932
rect 17267 19876 17448 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 14366 19845 14372 19848
rect 14360 19836 14372 19845
rect 6595 19808 8708 19836
rect 14327 19808 14372 19836
rect 6595 19805 6607 19808
rect 6549 19799 6607 19805
rect 14360 19799 14372 19808
rect 14366 19796 14372 19799
rect 14424 19796 14430 19848
rect 16206 19796 16212 19848
rect 16264 19796 16270 19848
rect 16482 19796 16488 19848
rect 16540 19796 16546 19848
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19836 17463 19839
rect 17451 19808 17908 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 17880 19780 17908 19808
rect 18046 19796 18052 19848
rect 18104 19836 18110 19848
rect 18874 19836 18880 19848
rect 18104 19808 18880 19836
rect 18104 19796 18110 19808
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 20254 19796 20260 19848
rect 20312 19796 20318 19848
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 21744 19836 21772 20000
rect 23032 19944 23336 19972
rect 22462 19864 22468 19916
rect 22520 19904 22526 19916
rect 23032 19913 23060 19944
rect 22741 19907 22799 19913
rect 22741 19904 22753 19907
rect 22520 19876 22753 19904
rect 22520 19864 22526 19876
rect 22741 19873 22753 19876
rect 22787 19904 22799 19907
rect 23017 19907 23075 19913
rect 23017 19904 23029 19907
rect 22787 19876 23029 19904
rect 22787 19873 22799 19876
rect 22741 19867 22799 19873
rect 23017 19873 23029 19876
rect 23063 19873 23075 19907
rect 23017 19867 23075 19873
rect 23106 19864 23112 19916
rect 23164 19864 23170 19916
rect 23198 19864 23204 19916
rect 23256 19864 23262 19916
rect 23308 19904 23336 19944
rect 23382 19932 23388 19984
rect 23440 19972 23446 19984
rect 27816 19972 27844 20003
rect 28442 20000 28448 20012
rect 28500 20000 28506 20052
rect 39132 20012 41414 20040
rect 23440 19944 27844 19972
rect 38565 19975 38623 19981
rect 23440 19932 23446 19944
rect 38565 19941 38577 19975
rect 38611 19972 38623 19975
rect 38838 19972 38844 19984
rect 38611 19944 38844 19972
rect 38611 19941 38623 19944
rect 38565 19935 38623 19941
rect 38838 19932 38844 19944
rect 38896 19932 38902 19984
rect 23308 19876 27476 19904
rect 23216 19836 23244 19864
rect 21744 19808 23244 19836
rect 24946 19796 24952 19848
rect 25004 19796 25010 19848
rect 26234 19796 26240 19848
rect 26292 19796 26298 19848
rect 26510 19796 26516 19848
rect 26568 19796 26574 19848
rect 9674 19768 9680 19780
rect 6472 19740 9680 19768
rect 9674 19728 9680 19740
rect 9732 19728 9738 19780
rect 10042 19728 10048 19780
rect 10100 19768 10106 19780
rect 10321 19771 10379 19777
rect 10321 19768 10333 19771
rect 10100 19740 10333 19768
rect 10100 19728 10106 19740
rect 10321 19737 10333 19740
rect 10367 19768 10379 19771
rect 10367 19740 10824 19768
rect 10367 19737 10379 19740
rect 10321 19731 10379 19737
rect 10796 19712 10824 19740
rect 17862 19728 17868 19780
rect 17920 19728 17926 19780
rect 17954 19728 17960 19780
rect 18012 19728 18018 19780
rect 18598 19728 18604 19780
rect 18656 19777 18662 19780
rect 18656 19768 18668 19777
rect 18656 19740 18701 19768
rect 18656 19731 18668 19740
rect 18656 19728 18662 19731
rect 21082 19728 21088 19780
rect 21140 19768 21146 19780
rect 21140 19740 22876 19768
rect 21140 19728 21146 19740
rect 4157 19703 4215 19709
rect 4157 19669 4169 19703
rect 4203 19700 4215 19703
rect 4246 19700 4252 19712
rect 4203 19672 4252 19700
rect 4203 19669 4215 19672
rect 4157 19663 4215 19669
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 6454 19660 6460 19712
rect 6512 19700 6518 19712
rect 8021 19703 8079 19709
rect 8021 19700 8033 19703
rect 6512 19672 8033 19700
rect 6512 19660 6518 19672
rect 8021 19669 8033 19672
rect 8067 19700 8079 19703
rect 9122 19700 9128 19712
rect 8067 19672 9128 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 10778 19660 10784 19712
rect 10836 19660 10842 19712
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 12250 19700 12256 19712
rect 11296 19672 12256 19700
rect 11296 19660 11302 19672
rect 12250 19660 12256 19672
rect 12308 19700 12314 19712
rect 13817 19703 13875 19709
rect 13817 19700 13829 19703
rect 12308 19672 13829 19700
rect 12308 19660 12314 19672
rect 13817 19669 13829 19672
rect 13863 19700 13875 19703
rect 14274 19700 14280 19712
rect 13863 19672 14280 19700
rect 13863 19669 13875 19672
rect 13817 19663 13875 19669
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 15565 19703 15623 19709
rect 15565 19669 15577 19703
rect 15611 19700 15623 19703
rect 16942 19700 16948 19712
rect 15611 19672 16948 19700
rect 15611 19669 15623 19672
rect 15565 19663 15623 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 17972 19700 18000 19728
rect 22848 19712 22876 19740
rect 22922 19728 22928 19780
rect 22980 19768 22986 19780
rect 23201 19771 23259 19777
rect 23201 19768 23213 19771
rect 22980 19740 23213 19768
rect 22980 19728 22986 19740
rect 23201 19737 23213 19740
rect 23247 19768 23259 19771
rect 24397 19771 24455 19777
rect 24397 19768 24409 19771
rect 23247 19740 24409 19768
rect 23247 19737 23259 19740
rect 23201 19731 23259 19737
rect 24397 19737 24409 19740
rect 24443 19737 24455 19771
rect 24397 19731 24455 19737
rect 27448 19712 27476 19876
rect 36906 19864 36912 19916
rect 36964 19904 36970 19916
rect 37461 19907 37519 19913
rect 37461 19904 37473 19907
rect 36964 19876 37473 19904
rect 36964 19864 36970 19876
rect 37461 19873 37473 19876
rect 37507 19873 37519 19907
rect 37461 19867 37519 19873
rect 38102 19864 38108 19916
rect 38160 19904 38166 19916
rect 39132 19913 39160 20012
rect 41386 19972 41414 20012
rect 48222 20000 48228 20052
rect 48280 20000 48286 20052
rect 48406 20000 48412 20052
rect 48464 20000 48470 20052
rect 49326 20000 49332 20052
rect 49384 20000 49390 20052
rect 50246 20000 50252 20052
rect 50304 20000 50310 20052
rect 54570 20000 54576 20052
rect 54628 20000 54634 20052
rect 56686 20000 56692 20052
rect 56744 20000 56750 20052
rect 56870 20000 56876 20052
rect 56928 20040 56934 20052
rect 56928 20012 57468 20040
rect 56928 20000 56934 20012
rect 43993 19975 44051 19981
rect 43993 19972 44005 19975
rect 41386 19944 44005 19972
rect 43993 19941 44005 19944
rect 44039 19972 44051 19975
rect 44910 19972 44916 19984
rect 44039 19944 44916 19972
rect 44039 19941 44051 19944
rect 43993 19935 44051 19941
rect 44652 19916 44680 19944
rect 44910 19932 44916 19944
rect 44968 19932 44974 19984
rect 45741 19975 45799 19981
rect 45741 19941 45753 19975
rect 45787 19972 45799 19975
rect 48133 19975 48191 19981
rect 45787 19944 46428 19972
rect 45787 19941 45799 19944
rect 45741 19935 45799 19941
rect 39117 19907 39175 19913
rect 39117 19904 39129 19907
rect 38160 19876 39129 19904
rect 38160 19864 38166 19876
rect 39117 19873 39129 19876
rect 39163 19873 39175 19907
rect 39117 19867 39175 19873
rect 39758 19864 39764 19916
rect 39816 19904 39822 19916
rect 40037 19907 40095 19913
rect 40037 19904 40049 19907
rect 39816 19876 40049 19904
rect 39816 19864 39822 19876
rect 40037 19873 40049 19876
rect 40083 19904 40095 19907
rect 44542 19904 44548 19916
rect 40083 19876 44548 19904
rect 40083 19873 40095 19876
rect 40037 19867 40095 19873
rect 44542 19864 44548 19876
rect 44600 19864 44606 19916
rect 44634 19864 44640 19916
rect 44692 19864 44698 19916
rect 44818 19864 44824 19916
rect 44876 19904 44882 19916
rect 46400 19913 46428 19944
rect 48133 19941 48145 19975
rect 48179 19972 48191 19975
rect 48424 19972 48452 20000
rect 48179 19944 48452 19972
rect 48608 19944 49280 19972
rect 48179 19941 48191 19944
rect 48133 19935 48191 19941
rect 45097 19907 45155 19913
rect 45097 19904 45109 19907
rect 44876 19876 45109 19904
rect 44876 19864 44882 19876
rect 45097 19873 45109 19876
rect 45143 19873 45155 19907
rect 45097 19867 45155 19873
rect 46385 19907 46443 19913
rect 46385 19873 46397 19907
rect 46431 19873 46443 19907
rect 46385 19867 46443 19873
rect 46658 19864 46664 19916
rect 46716 19904 46722 19916
rect 46753 19907 46811 19913
rect 46753 19904 46765 19907
rect 46716 19876 46765 19904
rect 46716 19864 46722 19876
rect 46753 19873 46765 19876
rect 46799 19873 46811 19907
rect 46753 19867 46811 19873
rect 30650 19796 30656 19848
rect 30708 19796 30714 19848
rect 31386 19796 31392 19848
rect 31444 19796 31450 19848
rect 35437 19839 35495 19845
rect 35437 19836 35449 19839
rect 35360 19808 35449 19836
rect 33778 19768 33784 19780
rect 32324 19740 33784 19768
rect 32324 19712 32352 19740
rect 33778 19728 33784 19740
rect 33836 19728 33842 19780
rect 35360 19712 35388 19808
rect 35437 19805 35449 19808
rect 35483 19805 35495 19839
rect 35437 19799 35495 19805
rect 37642 19796 37648 19848
rect 37700 19796 37706 19848
rect 39022 19796 39028 19848
rect 39080 19836 39086 19848
rect 40221 19839 40279 19845
rect 40221 19836 40233 19839
rect 39080 19808 40233 19836
rect 39080 19796 39086 19808
rect 40221 19805 40233 19808
rect 40267 19805 40279 19839
rect 40221 19799 40279 19805
rect 41966 19796 41972 19848
rect 42024 19796 42030 19848
rect 42702 19796 42708 19848
rect 42760 19836 42766 19848
rect 44453 19839 44511 19845
rect 44453 19836 44465 19839
rect 42760 19808 44465 19836
rect 42760 19796 42766 19808
rect 44453 19805 44465 19808
rect 44499 19836 44511 19839
rect 45002 19836 45008 19848
rect 44499 19808 45008 19836
rect 44499 19805 44511 19808
rect 44453 19799 44511 19805
rect 45002 19796 45008 19808
rect 45060 19836 45066 19848
rect 45281 19839 45339 19845
rect 45281 19836 45293 19839
rect 45060 19808 45293 19836
rect 45060 19796 45066 19808
rect 45281 19805 45293 19808
rect 45327 19805 45339 19839
rect 45281 19799 45339 19805
rect 47020 19839 47078 19845
rect 47020 19805 47032 19839
rect 47066 19836 47078 19839
rect 47302 19836 47308 19848
rect 47066 19808 47308 19836
rect 47066 19805 47078 19808
rect 47020 19799 47078 19805
rect 47302 19796 47308 19808
rect 47360 19796 47366 19848
rect 47854 19796 47860 19848
rect 47912 19836 47918 19848
rect 48608 19845 48636 19944
rect 49252 19916 49280 19944
rect 48682 19864 48688 19916
rect 48740 19864 48746 19916
rect 48774 19864 48780 19916
rect 48832 19864 48838 19916
rect 49234 19864 49240 19916
rect 49292 19864 49298 19916
rect 49344 19904 49372 20000
rect 50264 19913 50292 20000
rect 49789 19907 49847 19913
rect 49789 19904 49801 19907
rect 49344 19876 49801 19904
rect 49789 19873 49801 19876
rect 49835 19873 49847 19907
rect 49789 19867 49847 19873
rect 50249 19907 50307 19913
rect 50249 19873 50261 19907
rect 50295 19873 50307 19907
rect 50249 19867 50307 19873
rect 50433 19907 50491 19913
rect 50433 19873 50445 19907
rect 50479 19904 50491 19907
rect 50985 19907 51043 19913
rect 50985 19904 50997 19907
rect 50479 19876 50997 19904
rect 50479 19873 50491 19876
rect 50433 19867 50491 19873
rect 50985 19873 50997 19876
rect 51031 19873 51043 19907
rect 52917 19907 52975 19913
rect 52917 19904 52929 19907
rect 50985 19867 51043 19873
rect 51920 19876 52929 19904
rect 48593 19839 48651 19845
rect 48593 19836 48605 19839
rect 47912 19808 48605 19836
rect 47912 19796 47918 19808
rect 48593 19805 48605 19808
rect 48639 19805 48651 19839
rect 48700 19836 48728 19864
rect 51920 19848 51948 19876
rect 52917 19873 52929 19876
rect 52963 19873 52975 19907
rect 54588 19904 54616 20000
rect 56502 19932 56508 19984
rect 56560 19932 56566 19984
rect 54941 19907 54999 19913
rect 54941 19904 54953 19907
rect 54588 19876 54953 19904
rect 52917 19867 52975 19873
rect 54941 19873 54953 19876
rect 54987 19873 54999 19907
rect 54941 19867 54999 19873
rect 55398 19864 55404 19916
rect 55456 19904 55462 19916
rect 55953 19907 56011 19913
rect 55953 19904 55965 19907
rect 55456 19876 55965 19904
rect 55456 19864 55462 19876
rect 55953 19873 55965 19876
rect 55999 19873 56011 19907
rect 55953 19867 56011 19873
rect 56229 19907 56287 19913
rect 56229 19873 56241 19907
rect 56275 19904 56287 19907
rect 56704 19904 56732 20000
rect 57440 19916 57468 20012
rect 57238 19904 57244 19916
rect 56275 19876 56732 19904
rect 57072 19876 57244 19904
rect 56275 19873 56287 19876
rect 56229 19867 56287 19873
rect 49326 19836 49332 19848
rect 48700 19808 49332 19836
rect 48593 19799 48651 19805
rect 49326 19796 49332 19808
rect 49384 19796 49390 19848
rect 49602 19796 49608 19848
rect 49660 19796 49666 19848
rect 50338 19796 50344 19848
rect 50396 19836 50402 19848
rect 51537 19839 51595 19845
rect 51537 19836 51549 19839
rect 50396 19808 51549 19836
rect 50396 19796 50402 19808
rect 51537 19805 51549 19808
rect 51583 19805 51595 19839
rect 51537 19799 51595 19805
rect 51902 19796 51908 19848
rect 51960 19796 51966 19848
rect 52273 19839 52331 19845
rect 52273 19805 52285 19839
rect 52319 19805 52331 19839
rect 52273 19799 52331 19805
rect 53184 19839 53242 19845
rect 53184 19805 53196 19839
rect 53230 19836 53242 19839
rect 53650 19836 53656 19848
rect 53230 19808 53656 19836
rect 53230 19805 53242 19808
rect 53184 19799 53242 19805
rect 35704 19771 35762 19777
rect 35704 19737 35716 19771
rect 35750 19768 35762 19771
rect 36909 19771 36967 19777
rect 36909 19768 36921 19771
rect 35750 19740 36921 19768
rect 35750 19737 35762 19740
rect 35704 19731 35762 19737
rect 36909 19737 36921 19740
rect 36955 19737 36967 19771
rect 39574 19768 39580 19780
rect 36909 19731 36967 19737
rect 38672 19740 39580 19768
rect 38672 19712 38700 19740
rect 39574 19728 39580 19740
rect 39632 19728 39638 19780
rect 48406 19728 48412 19780
rect 48464 19768 48470 19780
rect 49697 19771 49755 19777
rect 49697 19768 49709 19771
rect 48464 19740 49709 19768
rect 48464 19728 48470 19740
rect 49697 19737 49709 19740
rect 49743 19737 49755 19771
rect 52288 19768 52316 19799
rect 53650 19796 53656 19808
rect 53708 19796 53714 19848
rect 53926 19796 53932 19848
rect 53984 19836 53990 19848
rect 56134 19845 56140 19848
rect 54757 19839 54815 19845
rect 54757 19836 54769 19839
rect 53984 19808 54769 19836
rect 53984 19796 53990 19808
rect 54757 19805 54769 19808
rect 54803 19805 54815 19839
rect 54757 19799 54815 19805
rect 56112 19839 56140 19845
rect 56112 19805 56124 19839
rect 56112 19799 56140 19805
rect 56134 19796 56140 19799
rect 56192 19796 56198 19848
rect 56965 19839 57023 19845
rect 56965 19805 56977 19839
rect 57011 19836 57023 19839
rect 57072 19836 57100 19876
rect 57238 19864 57244 19876
rect 57296 19864 57302 19916
rect 57422 19864 57428 19916
rect 57480 19904 57486 19916
rect 58253 19907 58311 19913
rect 58253 19904 58265 19907
rect 57480 19876 58265 19904
rect 57480 19864 57486 19876
rect 58253 19873 58265 19876
rect 58299 19873 58311 19907
rect 58253 19867 58311 19873
rect 57011 19808 57100 19836
rect 57149 19839 57207 19845
rect 57011 19805 57023 19808
rect 56965 19799 57023 19805
rect 57149 19805 57161 19839
rect 57195 19836 57207 19839
rect 57195 19808 57560 19836
rect 57195 19805 57207 19808
rect 57149 19799 57207 19805
rect 55214 19768 55220 19780
rect 49697 19731 49755 19737
rect 50908 19740 51074 19768
rect 17543 19672 18000 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 19702 19660 19708 19712
rect 19760 19660 19766 19712
rect 22097 19703 22155 19709
rect 22097 19669 22109 19703
rect 22143 19700 22155 19703
rect 22278 19700 22284 19712
rect 22143 19672 22284 19700
rect 22143 19669 22155 19672
rect 22097 19663 22155 19669
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 22830 19660 22836 19712
rect 22888 19660 22894 19712
rect 23842 19660 23848 19712
rect 23900 19660 23906 19712
rect 25590 19660 25596 19712
rect 25648 19660 25654 19712
rect 27062 19660 27068 19712
rect 27120 19660 27126 19712
rect 27430 19660 27436 19712
rect 27488 19660 27494 19712
rect 29730 19660 29736 19712
rect 29788 19700 29794 19712
rect 30101 19703 30159 19709
rect 30101 19700 30113 19703
rect 29788 19672 30113 19700
rect 29788 19660 29794 19672
rect 30101 19669 30113 19672
rect 30147 19669 30159 19703
rect 30101 19663 30159 19669
rect 30834 19660 30840 19712
rect 30892 19660 30898 19712
rect 31754 19660 31760 19712
rect 31812 19660 31818 19712
rect 32306 19660 32312 19712
rect 32364 19660 32370 19712
rect 33505 19703 33563 19709
rect 33505 19669 33517 19703
rect 33551 19700 33563 19703
rect 33686 19700 33692 19712
rect 33551 19672 33692 19700
rect 33551 19669 33563 19672
rect 33505 19663 33563 19669
rect 33686 19660 33692 19672
rect 33744 19660 33750 19712
rect 35342 19660 35348 19712
rect 35400 19660 35406 19712
rect 36817 19703 36875 19709
rect 36817 19669 36829 19703
rect 36863 19700 36875 19703
rect 37550 19700 37556 19712
rect 36863 19672 37556 19700
rect 36863 19669 36875 19672
rect 36817 19663 36875 19669
rect 37550 19660 37556 19672
rect 37608 19660 37614 19712
rect 37734 19660 37740 19712
rect 37792 19700 37798 19712
rect 38289 19703 38347 19709
rect 38289 19700 38301 19703
rect 37792 19672 38301 19700
rect 37792 19660 37798 19672
rect 38289 19669 38301 19672
rect 38335 19700 38347 19703
rect 38470 19700 38476 19712
rect 38335 19672 38476 19700
rect 38335 19669 38347 19672
rect 38289 19663 38347 19669
rect 38470 19660 38476 19672
rect 38528 19660 38534 19712
rect 38654 19660 38660 19712
rect 38712 19660 38718 19712
rect 38930 19660 38936 19712
rect 38988 19660 38994 19712
rect 39022 19660 39028 19712
rect 39080 19660 39086 19712
rect 39114 19660 39120 19712
rect 39172 19700 39178 19712
rect 40129 19703 40187 19709
rect 40129 19700 40141 19703
rect 39172 19672 40141 19700
rect 39172 19660 39178 19672
rect 40129 19669 40141 19672
rect 40175 19669 40187 19703
rect 40129 19663 40187 19669
rect 40586 19660 40592 19712
rect 40644 19660 40650 19712
rect 41414 19660 41420 19712
rect 41472 19660 41478 19712
rect 44085 19703 44143 19709
rect 44085 19669 44097 19703
rect 44131 19700 44143 19703
rect 44174 19700 44180 19712
rect 44131 19672 44180 19700
rect 44131 19669 44143 19672
rect 44085 19663 44143 19669
rect 44174 19660 44180 19672
rect 44232 19660 44238 19712
rect 44545 19703 44603 19709
rect 44545 19669 44557 19703
rect 44591 19700 44603 19703
rect 44634 19700 44640 19712
rect 44591 19672 44640 19700
rect 44591 19669 44603 19672
rect 44545 19663 44603 19669
rect 44634 19660 44640 19672
rect 44692 19660 44698 19712
rect 45370 19660 45376 19712
rect 45428 19660 45434 19712
rect 45830 19660 45836 19712
rect 45888 19660 45894 19712
rect 48774 19660 48780 19712
rect 48832 19700 48838 19712
rect 49237 19703 49295 19709
rect 49237 19700 49249 19703
rect 48832 19672 49249 19700
rect 48832 19660 48838 19672
rect 49237 19669 49249 19672
rect 49283 19669 49295 19703
rect 49237 19663 49295 19669
rect 49418 19660 49424 19712
rect 49476 19700 49482 19712
rect 49878 19700 49884 19712
rect 49476 19672 49884 19700
rect 49476 19660 49482 19672
rect 49878 19660 49884 19672
rect 49936 19700 49942 19712
rect 50908 19709 50936 19740
rect 50525 19703 50583 19709
rect 50525 19700 50537 19703
rect 49936 19672 50537 19700
rect 49936 19660 49942 19672
rect 50525 19669 50537 19672
rect 50571 19669 50583 19703
rect 50525 19663 50583 19669
rect 50893 19703 50951 19709
rect 50893 19669 50905 19703
rect 50939 19669 50951 19703
rect 51046 19700 51074 19740
rect 51644 19740 52316 19768
rect 54312 19740 55220 19768
rect 51644 19700 51672 19740
rect 51046 19672 51672 19700
rect 50893 19663 50951 19669
rect 51718 19660 51724 19712
rect 51776 19660 51782 19712
rect 54312 19709 54340 19740
rect 55214 19728 55220 19740
rect 55272 19728 55278 19780
rect 57532 19712 57560 19808
rect 54297 19703 54355 19709
rect 54297 19669 54309 19703
rect 54343 19669 54355 19703
rect 54297 19663 54355 19669
rect 54386 19660 54392 19712
rect 54444 19660 54450 19712
rect 54849 19703 54907 19709
rect 54849 19669 54861 19703
rect 54895 19700 54907 19703
rect 55309 19703 55367 19709
rect 55309 19700 55321 19703
rect 54895 19672 55321 19700
rect 54895 19669 54907 19672
rect 54849 19663 54907 19669
rect 55309 19669 55321 19672
rect 55355 19669 55367 19703
rect 55309 19663 55367 19669
rect 57514 19660 57520 19712
rect 57572 19660 57578 19712
rect 57606 19660 57612 19712
rect 57664 19660 57670 19712
rect 57974 19660 57980 19712
rect 58032 19660 58038 19712
rect 1104 19610 59040 19632
rect 1104 19558 15394 19610
rect 15446 19558 15458 19610
rect 15510 19558 15522 19610
rect 15574 19558 15586 19610
rect 15638 19558 15650 19610
rect 15702 19558 29838 19610
rect 29890 19558 29902 19610
rect 29954 19558 29966 19610
rect 30018 19558 30030 19610
rect 30082 19558 30094 19610
rect 30146 19558 44282 19610
rect 44334 19558 44346 19610
rect 44398 19558 44410 19610
rect 44462 19558 44474 19610
rect 44526 19558 44538 19610
rect 44590 19558 58726 19610
rect 58778 19558 58790 19610
rect 58842 19558 58854 19610
rect 58906 19558 58918 19610
rect 58970 19558 58982 19610
rect 59034 19558 59040 19610
rect 1104 19536 59040 19558
rect 3973 19499 4031 19505
rect 3973 19465 3985 19499
rect 4019 19496 4031 19499
rect 4798 19496 4804 19508
rect 4019 19468 4804 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19465 7803 19499
rect 7745 19459 7803 19465
rect 7760 19428 7788 19459
rect 11238 19456 11244 19508
rect 11296 19496 11302 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11296 19468 11713 19496
rect 11296 19456 11302 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 15194 19456 15200 19508
rect 15252 19456 15258 19508
rect 15749 19499 15807 19505
rect 15749 19465 15761 19499
rect 15795 19496 15807 19499
rect 16482 19496 16488 19508
rect 15795 19468 16488 19496
rect 15795 19465 15807 19468
rect 15749 19459 15807 19465
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 17954 19496 17960 19508
rect 16715 19468 17960 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 17954 19456 17960 19468
rect 18012 19496 18018 19508
rect 19797 19499 19855 19505
rect 18012 19468 18736 19496
rect 18012 19456 18018 19468
rect 2516 19400 5396 19428
rect 7760 19400 8524 19428
rect 2406 19320 2412 19372
rect 2464 19360 2470 19372
rect 2516 19369 2544 19400
rect 2774 19369 2780 19372
rect 2501 19363 2559 19369
rect 2501 19360 2513 19363
rect 2464 19332 2513 19360
rect 2464 19320 2470 19332
rect 2501 19329 2513 19332
rect 2547 19329 2559 19363
rect 2501 19323 2559 19329
rect 2768 19323 2780 19369
rect 2774 19320 2780 19323
rect 2832 19320 2838 19372
rect 5074 19320 5080 19372
rect 5132 19369 5138 19372
rect 5368 19369 5396 19400
rect 5132 19360 5144 19369
rect 5353 19363 5411 19369
rect 5132 19332 5177 19360
rect 5132 19323 5144 19332
rect 5353 19329 5365 19363
rect 5399 19360 5411 19363
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 5399 19332 6377 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 6365 19329 6377 19332
rect 6411 19360 6423 19363
rect 6454 19360 6460 19372
rect 6411 19332 6460 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 5132 19320 5138 19323
rect 6454 19320 6460 19332
rect 6512 19320 6518 19372
rect 6632 19363 6690 19369
rect 6632 19329 6644 19363
rect 6678 19360 6690 19363
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 6678 19332 7849 19360
rect 6678 19329 6690 19332
rect 6632 19323 6690 19329
rect 7837 19329 7849 19332
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 5445 19295 5503 19301
rect 5445 19292 5457 19295
rect 5368 19264 5457 19292
rect 3881 19227 3939 19233
rect 3881 19193 3893 19227
rect 3927 19224 3939 19227
rect 3927 19196 4476 19224
rect 3927 19193 3939 19196
rect 3881 19187 3939 19193
rect 4448 19156 4476 19196
rect 5368 19156 5396 19264
rect 5445 19261 5457 19264
rect 5491 19261 5503 19295
rect 5445 19255 5503 19261
rect 7926 19252 7932 19304
rect 7984 19292 7990 19304
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 7984 19264 8401 19292
rect 7984 19252 7990 19264
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8496 19292 8524 19400
rect 14918 19388 14924 19440
rect 14976 19428 14982 19440
rect 15657 19431 15715 19437
rect 15657 19428 15669 19431
rect 14976 19400 15669 19428
rect 14976 19388 14982 19400
rect 15657 19397 15669 19400
rect 15703 19428 15715 19431
rect 17126 19428 17132 19440
rect 15703 19400 17132 19428
rect 15703 19397 15715 19400
rect 15657 19391 15715 19397
rect 17126 19388 17132 19400
rect 17184 19388 17190 19440
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11149 19363 11207 19369
rect 11149 19360 11161 19363
rect 11112 19332 11161 19360
rect 11112 19320 11118 19332
rect 11149 19329 11161 19332
rect 11195 19360 11207 19363
rect 11195 19332 12112 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 12084 19304 12112 19332
rect 13814 19320 13820 19372
rect 13872 19320 13878 19372
rect 14084 19363 14142 19369
rect 14084 19329 14096 19363
rect 14130 19360 14142 19363
rect 14366 19360 14372 19372
rect 14130 19332 14372 19360
rect 14130 19329 14142 19332
rect 14084 19323 14142 19329
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 16022 19320 16028 19372
rect 16080 19320 16086 19372
rect 17793 19363 17851 19369
rect 17793 19329 17805 19363
rect 17839 19360 17851 19363
rect 17954 19360 17960 19372
rect 17839 19332 17960 19360
rect 17839 19329 17851 19332
rect 17793 19323 17851 19329
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18046 19320 18052 19372
rect 18104 19320 18110 19372
rect 18708 19369 18736 19468
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20254 19496 20260 19508
rect 19843 19468 20260 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 21082 19456 21088 19508
rect 21140 19456 21146 19508
rect 22922 19496 22928 19508
rect 22020 19468 22928 19496
rect 20165 19431 20223 19437
rect 20165 19397 20177 19431
rect 20211 19428 20223 19431
rect 21100 19428 21128 19456
rect 20211 19400 21128 19428
rect 20211 19397 20223 19400
rect 20165 19391 20223 19397
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 20622 19360 20628 19372
rect 20303 19332 20628 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19360 21879 19363
rect 21910 19360 21916 19372
rect 21867 19332 21916 19360
rect 21867 19329 21879 19332
rect 21821 19323 21879 19329
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22020 19369 22048 19468
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 24121 19499 24179 19505
rect 24121 19496 24133 19499
rect 23348 19468 24133 19496
rect 23348 19456 23354 19468
rect 24121 19465 24133 19468
rect 24167 19465 24179 19499
rect 24121 19459 24179 19465
rect 25590 19456 25596 19508
rect 25648 19456 25654 19508
rect 26510 19456 26516 19508
rect 26568 19456 26574 19508
rect 30285 19499 30343 19505
rect 30285 19465 30297 19499
rect 30331 19496 30343 19499
rect 30650 19496 30656 19508
rect 30331 19468 30656 19496
rect 30331 19465 30343 19468
rect 30285 19459 30343 19465
rect 30650 19456 30656 19468
rect 30708 19456 30714 19508
rect 30745 19499 30803 19505
rect 30745 19465 30757 19499
rect 30791 19496 30803 19499
rect 30834 19496 30840 19508
rect 30791 19468 30840 19496
rect 30791 19465 30803 19468
rect 30745 19459 30803 19465
rect 30834 19456 30840 19468
rect 30892 19456 30898 19508
rect 34057 19499 34115 19505
rect 34057 19465 34069 19499
rect 34103 19496 34115 19499
rect 35250 19496 35256 19508
rect 34103 19468 35256 19496
rect 34103 19465 34115 19468
rect 34057 19459 34115 19465
rect 35250 19456 35256 19468
rect 35308 19456 35314 19508
rect 36909 19499 36967 19505
rect 36909 19465 36921 19499
rect 36955 19496 36967 19499
rect 37642 19496 37648 19508
rect 36955 19468 37648 19496
rect 36955 19465 36967 19468
rect 36909 19459 36967 19465
rect 37642 19456 37648 19468
rect 37700 19456 37706 19508
rect 37737 19499 37795 19505
rect 37737 19465 37749 19499
rect 37783 19496 37795 19499
rect 39114 19496 39120 19508
rect 37783 19468 39120 19496
rect 37783 19465 37795 19468
rect 37737 19459 37795 19465
rect 39114 19456 39120 19468
rect 39172 19456 39178 19508
rect 40218 19496 40224 19508
rect 39408 19468 40224 19496
rect 25400 19431 25458 19437
rect 25400 19397 25412 19431
rect 25446 19428 25458 19431
rect 25608 19428 25636 19456
rect 25446 19400 25636 19428
rect 35796 19431 35854 19437
rect 25446 19397 25458 19400
rect 25400 19391 25458 19397
rect 35796 19397 35808 19431
rect 35842 19428 35854 19431
rect 35986 19428 35992 19440
rect 35842 19400 35992 19428
rect 35842 19397 35854 19400
rect 35796 19391 35854 19397
rect 35986 19388 35992 19400
rect 36044 19388 36050 19440
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19329 22063 19363
rect 23661 19363 23719 19369
rect 22005 19323 22063 19329
rect 9125 19295 9183 19301
rect 9125 19292 9137 19295
rect 8496 19264 9137 19292
rect 8389 19255 8447 19261
rect 9125 19261 9137 19264
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 10226 19252 10232 19304
rect 10284 19252 10290 19304
rect 10594 19252 10600 19304
rect 10652 19252 10658 19304
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12618 19252 12624 19304
rect 12676 19252 12682 19304
rect 15838 19252 15844 19304
rect 15896 19252 15902 19304
rect 16040 19224 16068 19320
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 19392 19264 20361 19292
rect 19392 19252 19398 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20349 19255 20407 19261
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 21928 19264 22753 19292
rect 21174 19224 21180 19236
rect 15212 19196 16068 19224
rect 18064 19196 21180 19224
rect 4448 19128 5396 19156
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6089 19159 6147 19165
rect 6089 19156 6101 19159
rect 6052 19128 6101 19156
rect 6052 19116 6058 19128
rect 6089 19125 6101 19128
rect 6135 19125 6147 19159
rect 6089 19119 6147 19125
rect 8570 19116 8576 19168
rect 8628 19116 8634 19168
rect 9677 19159 9735 19165
rect 9677 19125 9689 19159
rect 9723 19156 9735 19159
rect 9766 19156 9772 19168
rect 9723 19128 9772 19156
rect 9723 19125 9735 19128
rect 9677 19119 9735 19125
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12069 19159 12127 19165
rect 12069 19156 12081 19159
rect 11940 19128 12081 19156
rect 11940 19116 11946 19128
rect 12069 19125 12081 19128
rect 12115 19125 12127 19159
rect 12069 19119 12127 19125
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 15212 19156 15240 19196
rect 13136 19128 15240 19156
rect 13136 19116 13142 19128
rect 15286 19116 15292 19168
rect 15344 19116 15350 19168
rect 16206 19116 16212 19168
rect 16264 19156 16270 19168
rect 16393 19159 16451 19165
rect 16393 19156 16405 19159
rect 16264 19128 16405 19156
rect 16264 19116 16270 19128
rect 16393 19125 16405 19128
rect 16439 19156 16451 19159
rect 18064 19156 18092 19196
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 21928 19224 21956 19264
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22830 19294 22836 19346
rect 22888 19301 22894 19346
rect 23661 19329 23673 19363
rect 23707 19360 23719 19363
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23707 19332 24041 19360
rect 23707 19329 23719 19332
rect 23661 19323 23719 19329
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 25133 19363 25191 19369
rect 25133 19360 25145 19363
rect 24029 19323 24087 19329
rect 24872 19332 25145 19360
rect 24872 19304 24900 19332
rect 25133 19329 25145 19332
rect 25179 19329 25191 19363
rect 25133 19323 25191 19329
rect 27522 19320 27528 19372
rect 27580 19360 27586 19372
rect 27801 19363 27859 19369
rect 27801 19360 27813 19363
rect 27580 19332 27813 19360
rect 27580 19320 27586 19332
rect 27801 19329 27813 19332
rect 27847 19329 27859 19363
rect 27801 19323 27859 19329
rect 30653 19363 30711 19369
rect 30653 19329 30665 19363
rect 30699 19360 30711 19363
rect 31478 19360 31484 19372
rect 30699 19332 31484 19360
rect 30699 19329 30711 19332
rect 30653 19323 30711 19329
rect 31478 19320 31484 19332
rect 31536 19320 31542 19372
rect 32944 19363 33002 19369
rect 32944 19329 32956 19363
rect 32990 19360 33002 19363
rect 34149 19363 34207 19369
rect 34149 19360 34161 19363
rect 32990 19332 34161 19360
rect 32990 19329 33002 19332
rect 32944 19323 33002 19329
rect 34149 19329 34161 19332
rect 34195 19329 34207 19363
rect 34149 19323 34207 19329
rect 35434 19320 35440 19372
rect 35492 19360 35498 19372
rect 35529 19363 35587 19369
rect 35529 19360 35541 19363
rect 35492 19332 35541 19360
rect 35492 19320 35498 19332
rect 35529 19329 35541 19332
rect 35575 19329 35587 19363
rect 35529 19323 35587 19329
rect 38470 19320 38476 19372
rect 38528 19369 38534 19372
rect 39408 19369 39436 19468
rect 40218 19456 40224 19468
rect 40276 19456 40282 19508
rect 45554 19456 45560 19508
rect 45612 19496 45618 19508
rect 45649 19499 45707 19505
rect 45649 19496 45661 19499
rect 45612 19468 45661 19496
rect 45612 19456 45618 19468
rect 45649 19465 45661 19468
rect 45695 19465 45707 19499
rect 45649 19459 45707 19465
rect 45830 19456 45836 19508
rect 45888 19456 45894 19508
rect 47397 19499 47455 19505
rect 47397 19465 47409 19499
rect 47443 19496 47455 19499
rect 47949 19499 48007 19505
rect 47949 19496 47961 19499
rect 47443 19468 47961 19496
rect 47443 19465 47455 19468
rect 47397 19459 47455 19465
rect 47949 19465 47961 19468
rect 47995 19496 48007 19499
rect 49142 19496 49148 19508
rect 47995 19468 49148 19496
rect 47995 19465 48007 19468
rect 47949 19459 48007 19465
rect 49142 19456 49148 19468
rect 49200 19456 49206 19508
rect 50338 19456 50344 19508
rect 50396 19456 50402 19508
rect 51718 19456 51724 19508
rect 51776 19456 51782 19508
rect 54021 19499 54079 19505
rect 54021 19496 54033 19499
rect 51920 19468 54033 19496
rect 39574 19388 39580 19440
rect 39632 19428 39638 19440
rect 44536 19431 44594 19437
rect 39632 19400 39712 19428
rect 39632 19388 39638 19400
rect 39684 19369 39712 19400
rect 44536 19397 44548 19431
rect 44582 19428 44594 19431
rect 45848 19428 45876 19456
rect 44582 19400 45876 19428
rect 44582 19397 44594 19400
rect 44536 19391 44594 19397
rect 47854 19388 47860 19440
rect 47912 19388 47918 19440
rect 48406 19388 48412 19440
rect 48464 19388 48470 19440
rect 38528 19363 38577 19369
rect 38528 19329 38531 19363
rect 38565 19329 38577 19363
rect 38528 19323 38577 19329
rect 39393 19363 39451 19369
rect 39393 19329 39405 19363
rect 39439 19329 39451 19363
rect 39393 19323 39451 19329
rect 39669 19363 39727 19369
rect 39669 19329 39681 19363
rect 39715 19329 39727 19363
rect 39669 19323 39727 19329
rect 39936 19363 39994 19369
rect 39936 19329 39948 19363
rect 39982 19360 39994 19363
rect 41141 19363 41199 19369
rect 41141 19360 41153 19363
rect 39982 19332 41153 19360
rect 39982 19329 39994 19332
rect 39936 19323 39994 19329
rect 41141 19329 41153 19332
rect 41187 19329 41199 19363
rect 44269 19363 44327 19369
rect 44269 19360 44281 19363
rect 41141 19323 41199 19329
rect 44008 19332 44281 19360
rect 38528 19320 38534 19323
rect 22888 19295 22916 19301
rect 22848 19264 22870 19294
rect 22741 19255 22799 19261
rect 22858 19261 22870 19264
rect 22904 19261 22916 19295
rect 22858 19255 22916 19261
rect 23017 19295 23075 19301
rect 23017 19261 23029 19295
rect 23063 19292 23075 19295
rect 23198 19292 23204 19304
rect 23063 19264 23204 19292
rect 23063 19261 23075 19264
rect 23017 19255 23075 19261
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 23842 19292 23848 19304
rect 23400 19264 23848 19292
rect 21468 19196 21956 19224
rect 16439 19128 18092 19156
rect 16439 19125 16451 19128
rect 16393 19119 16451 19125
rect 18138 19116 18144 19168
rect 18196 19116 18202 19168
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 19392 19128 19625 19156
rect 19392 19116 19398 19128
rect 19613 19125 19625 19128
rect 19659 19125 19671 19159
rect 19613 19119 19671 19125
rect 21082 19116 21088 19168
rect 21140 19156 21146 19168
rect 21468 19165 21496 19196
rect 22278 19184 22284 19236
rect 22336 19224 22342 19236
rect 22462 19224 22468 19236
rect 22336 19196 22468 19224
rect 22336 19184 22342 19196
rect 22462 19184 22468 19196
rect 22520 19184 22526 19236
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 21140 19128 21465 19156
rect 21140 19116 21146 19128
rect 21453 19125 21465 19128
rect 21499 19125 21511 19159
rect 21453 19119 21511 19125
rect 21542 19116 21548 19168
rect 21600 19156 21606 19168
rect 23400 19156 23428 19264
rect 23842 19252 23848 19264
rect 23900 19252 23906 19304
rect 24854 19252 24860 19304
rect 24912 19252 24918 19304
rect 27154 19252 27160 19304
rect 27212 19252 27218 19304
rect 30190 19252 30196 19304
rect 30248 19252 30254 19304
rect 30929 19295 30987 19301
rect 30929 19261 30941 19295
rect 30975 19261 30987 19295
rect 30929 19255 30987 19261
rect 29270 19184 29276 19236
rect 29328 19224 29334 19236
rect 30944 19224 30972 19255
rect 31294 19252 31300 19304
rect 31352 19252 31358 19304
rect 32122 19252 32128 19304
rect 32180 19292 32186 19304
rect 32582 19292 32588 19304
rect 32180 19264 32588 19292
rect 32180 19252 32186 19264
rect 32582 19252 32588 19264
rect 32640 19292 32646 19304
rect 32677 19295 32735 19301
rect 32677 19292 32689 19295
rect 32640 19264 32689 19292
rect 32640 19252 32646 19264
rect 32677 19261 32689 19264
rect 32723 19261 32735 19295
rect 32677 19255 32735 19261
rect 34698 19252 34704 19304
rect 34756 19252 34762 19304
rect 38378 19252 38384 19304
rect 38436 19252 38442 19304
rect 38657 19295 38715 19301
rect 38657 19261 38669 19295
rect 38703 19292 38715 19295
rect 38933 19295 38991 19301
rect 38703 19264 38884 19292
rect 38703 19261 38715 19264
rect 38657 19255 38715 19261
rect 31754 19224 31760 19236
rect 29328 19196 31760 19224
rect 29328 19184 29334 19196
rect 31754 19184 31760 19196
rect 31812 19224 31818 19236
rect 31812 19196 32536 19224
rect 31812 19184 31818 19196
rect 21600 19128 23428 19156
rect 21600 19116 21606 19128
rect 24486 19116 24492 19168
rect 24544 19116 24550 19168
rect 27890 19116 27896 19168
rect 27948 19156 27954 19168
rect 28077 19159 28135 19165
rect 28077 19156 28089 19159
rect 27948 19128 28089 19156
rect 27948 19116 27954 19128
rect 28077 19125 28089 19128
rect 28123 19125 28135 19159
rect 28077 19119 28135 19125
rect 29546 19116 29552 19168
rect 29604 19116 29610 19168
rect 31938 19116 31944 19168
rect 31996 19116 32002 19168
rect 32398 19116 32404 19168
rect 32456 19116 32462 19168
rect 32508 19156 32536 19196
rect 36722 19156 36728 19168
rect 32508 19128 36728 19156
rect 36722 19116 36728 19128
rect 36780 19116 36786 19168
rect 37553 19159 37611 19165
rect 37553 19125 37565 19159
rect 37599 19156 37611 19159
rect 37642 19156 37648 19168
rect 37599 19128 37648 19156
rect 37599 19125 37611 19128
rect 37553 19119 37611 19125
rect 37642 19116 37648 19128
rect 37700 19116 37706 19168
rect 37918 19116 37924 19168
rect 37976 19156 37982 19168
rect 38856 19156 38884 19264
rect 38933 19261 38945 19295
rect 38979 19292 38991 19295
rect 39206 19292 39212 19304
rect 38979 19264 39212 19292
rect 38979 19261 38991 19264
rect 38933 19255 38991 19261
rect 39206 19252 39212 19264
rect 39264 19252 39270 19304
rect 39577 19295 39635 19301
rect 39577 19261 39589 19295
rect 39623 19261 39635 19295
rect 39577 19255 39635 19261
rect 37976 19128 38884 19156
rect 39592 19156 39620 19255
rect 40954 19252 40960 19304
rect 41012 19292 41018 19304
rect 41693 19295 41751 19301
rect 41693 19292 41705 19295
rect 41012 19264 41705 19292
rect 41012 19252 41018 19264
rect 41693 19261 41705 19264
rect 41739 19261 41751 19295
rect 41693 19255 41751 19261
rect 42426 19252 42432 19304
rect 42484 19252 42490 19304
rect 43438 19252 43444 19304
rect 43496 19292 43502 19304
rect 44008 19292 44036 19332
rect 44269 19329 44281 19332
rect 44315 19329 44327 19363
rect 44269 19323 44327 19329
rect 49142 19320 49148 19372
rect 49200 19369 49206 19372
rect 49200 19363 49249 19369
rect 49200 19329 49203 19363
rect 49237 19329 49249 19363
rect 49200 19323 49249 19329
rect 49200 19320 49206 19323
rect 49326 19320 49332 19372
rect 49384 19320 49390 19372
rect 50249 19363 50307 19369
rect 50249 19329 50261 19363
rect 50295 19360 50307 19363
rect 50356 19360 50384 19456
rect 51476 19431 51534 19437
rect 51476 19397 51488 19431
rect 51522 19428 51534 19431
rect 51736 19428 51764 19456
rect 51522 19400 51764 19428
rect 51522 19397 51534 19400
rect 51476 19391 51534 19397
rect 51920 19372 51948 19468
rect 54021 19465 54033 19468
rect 54067 19465 54079 19499
rect 54021 19459 54079 19465
rect 55953 19499 56011 19505
rect 55953 19465 55965 19499
rect 55999 19496 56011 19499
rect 56042 19496 56048 19508
rect 55999 19468 56048 19496
rect 55999 19465 56011 19468
rect 55953 19459 56011 19465
rect 50295 19332 50384 19360
rect 51721 19363 51779 19369
rect 50295 19329 50307 19332
rect 50249 19323 50307 19329
rect 51721 19329 51733 19363
rect 51767 19360 51779 19363
rect 51902 19360 51908 19372
rect 51767 19332 51908 19360
rect 51767 19329 51779 19332
rect 51721 19323 51779 19329
rect 51902 19320 51908 19332
rect 51960 19320 51966 19372
rect 52733 19363 52791 19369
rect 52733 19360 52745 19363
rect 52472 19332 52745 19360
rect 43496 19264 44036 19292
rect 43496 19252 43502 19264
rect 44174 19252 44180 19304
rect 44232 19252 44238 19304
rect 46290 19252 46296 19304
rect 46348 19252 46354 19304
rect 46750 19252 46756 19304
rect 46808 19252 46814 19304
rect 47762 19252 47768 19304
rect 47820 19252 47826 19304
rect 49050 19252 49056 19304
rect 49108 19292 49114 19304
rect 49108 19264 49556 19292
rect 49108 19252 49114 19264
rect 44082 19224 44088 19236
rect 43364 19196 44088 19224
rect 39850 19156 39856 19168
rect 39592 19128 39856 19156
rect 37976 19116 37982 19128
rect 39850 19116 39856 19128
rect 39908 19116 39914 19168
rect 41046 19116 41052 19168
rect 41104 19116 41110 19168
rect 41874 19116 41880 19168
rect 41932 19156 41938 19168
rect 42061 19159 42119 19165
rect 42061 19156 42073 19159
rect 41932 19128 42073 19156
rect 41932 19116 41938 19128
rect 42061 19125 42073 19128
rect 42107 19125 42119 19159
rect 42061 19119 42119 19125
rect 42886 19116 42892 19168
rect 42944 19156 42950 19168
rect 43073 19159 43131 19165
rect 43073 19156 43085 19159
rect 42944 19128 43085 19156
rect 42944 19116 42950 19128
rect 43073 19125 43085 19128
rect 43119 19125 43131 19159
rect 43073 19119 43131 19125
rect 43254 19116 43260 19168
rect 43312 19156 43318 19168
rect 43364 19165 43392 19196
rect 44082 19184 44088 19196
rect 44140 19184 44146 19236
rect 43349 19159 43407 19165
rect 43349 19156 43361 19159
rect 43312 19128 43361 19156
rect 43312 19116 43318 19128
rect 43349 19125 43361 19128
rect 43395 19125 43407 19159
rect 43349 19119 43407 19125
rect 43530 19116 43536 19168
rect 43588 19116 43594 19168
rect 44634 19116 44640 19168
rect 44692 19156 44698 19168
rect 45741 19159 45799 19165
rect 45741 19156 45753 19159
rect 44692 19128 45753 19156
rect 44692 19116 44698 19128
rect 45741 19125 45753 19128
rect 45787 19125 45799 19159
rect 45741 19119 45799 19125
rect 45830 19116 45836 19168
rect 45888 19156 45894 19168
rect 46934 19156 46940 19168
rect 45888 19128 46940 19156
rect 45888 19116 45894 19128
rect 46934 19116 46940 19128
rect 46992 19156 46998 19168
rect 48130 19156 48136 19168
rect 46992 19128 48136 19156
rect 46992 19116 46998 19128
rect 48130 19116 48136 19128
rect 48188 19116 48194 19168
rect 48314 19116 48320 19168
rect 48372 19116 48378 19168
rect 49528 19156 49556 19264
rect 50062 19252 50068 19304
rect 50120 19252 50126 19304
rect 49602 19184 49608 19236
rect 49660 19184 49666 19236
rect 52472 19168 52500 19332
rect 52733 19329 52745 19332
rect 52779 19329 52791 19363
rect 54036 19360 54064 19459
rect 56042 19456 56048 19468
rect 56100 19456 56106 19508
rect 57701 19499 57759 19505
rect 57701 19465 57713 19499
rect 57747 19496 57759 19499
rect 58250 19496 58256 19508
rect 57747 19468 58256 19496
rect 57747 19465 57759 19468
rect 57701 19459 57759 19465
rect 58250 19456 58256 19468
rect 58308 19456 58314 19508
rect 54588 19400 55444 19428
rect 54588 19372 54616 19400
rect 54570 19360 54576 19372
rect 54036 19332 54576 19360
rect 52733 19323 52791 19329
rect 54570 19320 54576 19332
rect 54628 19320 54634 19372
rect 54840 19363 54898 19369
rect 54840 19329 54852 19363
rect 54886 19360 54898 19363
rect 55306 19360 55312 19372
rect 54886 19332 55312 19360
rect 54886 19329 54898 19332
rect 54840 19323 54898 19329
rect 55306 19320 55312 19332
rect 55364 19320 55370 19372
rect 55416 19360 55444 19400
rect 56318 19360 56324 19372
rect 55416 19332 56324 19360
rect 56318 19320 56324 19332
rect 56376 19320 56382 19372
rect 56588 19363 56646 19369
rect 56588 19329 56600 19363
rect 56634 19360 56646 19363
rect 57885 19363 57943 19369
rect 57885 19360 57897 19363
rect 56634 19332 57897 19360
rect 56634 19329 56646 19332
rect 56588 19323 56646 19329
rect 57885 19329 57897 19332
rect 57931 19329 57943 19363
rect 57885 19323 57943 19329
rect 57974 19320 57980 19372
rect 58032 19360 58038 19372
rect 58437 19363 58495 19369
rect 58437 19360 58449 19363
rect 58032 19332 58449 19360
rect 58032 19320 58038 19332
rect 58437 19329 58449 19332
rect 58483 19329 58495 19363
rect 58437 19323 58495 19329
rect 52362 19156 52368 19168
rect 49528 19128 52368 19156
rect 52362 19116 52368 19128
rect 52420 19116 52426 19168
rect 52454 19116 52460 19168
rect 52512 19116 52518 19168
rect 1104 19066 58880 19088
rect 1104 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 22616 19066
rect 22668 19014 22680 19066
rect 22732 19014 22744 19066
rect 22796 19014 22808 19066
rect 22860 19014 22872 19066
rect 22924 19014 37060 19066
rect 37112 19014 37124 19066
rect 37176 19014 37188 19066
rect 37240 19014 37252 19066
rect 37304 19014 37316 19066
rect 37368 19014 51504 19066
rect 51556 19014 51568 19066
rect 51620 19014 51632 19066
rect 51684 19014 51696 19066
rect 51748 19014 51760 19066
rect 51812 19014 58880 19066
rect 1104 18992 58880 19014
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2832 18924 2973 18952
rect 2832 18912 2838 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 2961 18915 3019 18921
rect 5169 18955 5227 18961
rect 5169 18921 5181 18955
rect 5215 18952 5227 18955
rect 5902 18952 5908 18964
rect 5215 18924 5908 18952
rect 5215 18921 5227 18924
rect 5169 18915 5227 18921
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 7926 18912 7932 18964
rect 7984 18912 7990 18964
rect 9674 18912 9680 18964
rect 9732 18912 9738 18964
rect 9861 18955 9919 18961
rect 9861 18921 9873 18955
rect 9907 18952 9919 18955
rect 10226 18952 10232 18964
rect 9907 18924 10232 18952
rect 9907 18921 9919 18924
rect 9861 18915 9919 18921
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 12345 18955 12403 18961
rect 12345 18921 12357 18955
rect 12391 18952 12403 18955
rect 12618 18952 12624 18964
rect 12391 18924 12624 18952
rect 12391 18921 12403 18924
rect 12345 18915 12403 18921
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 13078 18912 13084 18964
rect 13136 18912 13142 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14424 18924 14749 18952
rect 14424 18912 14430 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 16390 18912 16396 18964
rect 16448 18952 16454 18964
rect 16448 18924 17632 18952
rect 16448 18912 16454 18924
rect 3789 18887 3847 18893
rect 3789 18853 3801 18887
rect 3835 18853 3847 18887
rect 3789 18847 3847 18853
rect 6365 18887 6423 18893
rect 6365 18853 6377 18887
rect 6411 18884 6423 18887
rect 6822 18884 6828 18896
rect 6411 18856 6828 18884
rect 6411 18853 6423 18856
rect 6365 18847 6423 18853
rect 3605 18819 3663 18825
rect 3605 18785 3617 18819
rect 3651 18816 3663 18819
rect 3804 18816 3832 18847
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 9125 18887 9183 18893
rect 9125 18884 9137 18887
rect 8496 18856 9137 18884
rect 3651 18788 3832 18816
rect 4433 18819 4491 18825
rect 3651 18785 3663 18788
rect 3605 18779 3663 18785
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4798 18816 4804 18828
rect 4479 18788 4804 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 5994 18825 6000 18828
rect 5951 18819 6000 18825
rect 5951 18816 5963 18819
rect 5276 18788 5963 18816
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 5276 18748 5304 18788
rect 5951 18785 5963 18788
rect 5997 18785 6000 18819
rect 5951 18779 6000 18785
rect 5994 18776 6000 18779
rect 6052 18776 6058 18828
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7742 18816 7748 18828
rect 7331 18788 7748 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8496 18825 8524 18856
rect 9125 18853 9137 18856
rect 9171 18853 9183 18887
rect 9692 18884 9720 18912
rect 9692 18856 10456 18884
rect 9125 18847 9183 18853
rect 8481 18819 8539 18825
rect 8481 18785 8493 18819
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 8570 18776 8576 18828
rect 8628 18776 8634 18828
rect 4203 18720 5304 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18748 7067 18751
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7055 18720 8401 18748
rect 7055 18717 7067 18720
rect 7009 18711 7067 18717
rect 8389 18717 8401 18720
rect 8435 18748 8447 18751
rect 8588 18748 8616 18776
rect 8435 18720 8616 18748
rect 9140 18748 9168 18847
rect 10428 18828 10456 18856
rect 10410 18776 10416 18828
rect 10468 18776 10474 18828
rect 13096 18825 13124 18912
rect 17405 18887 17463 18893
rect 17405 18853 17417 18887
rect 17451 18884 17463 18887
rect 17604 18884 17632 18924
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18141 18955 18199 18961
rect 18141 18952 18153 18955
rect 18012 18924 18153 18952
rect 18012 18912 18018 18924
rect 18141 18921 18153 18924
rect 18187 18921 18199 18955
rect 18141 18915 18199 18921
rect 18248 18924 20208 18952
rect 18248 18884 18276 18924
rect 17451 18856 17540 18884
rect 17604 18856 18276 18884
rect 20180 18884 20208 18924
rect 20530 18912 20536 18964
rect 20588 18952 20594 18964
rect 20625 18955 20683 18961
rect 20625 18952 20637 18955
rect 20588 18924 20637 18952
rect 20588 18912 20594 18924
rect 20625 18921 20637 18924
rect 20671 18921 20683 18955
rect 20625 18915 20683 18921
rect 21450 18912 21456 18964
rect 21508 18912 21514 18964
rect 23937 18955 23995 18961
rect 23937 18921 23949 18955
rect 23983 18952 23995 18955
rect 24946 18952 24952 18964
rect 23983 18924 24952 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 25777 18955 25835 18961
rect 25777 18921 25789 18955
rect 25823 18952 25835 18955
rect 26234 18952 26240 18964
rect 25823 18924 26240 18952
rect 25823 18921 25835 18924
rect 25777 18915 25835 18921
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 26973 18955 27031 18961
rect 26973 18921 26985 18955
rect 27019 18952 27031 18955
rect 27154 18952 27160 18964
rect 27019 18924 27160 18952
rect 27019 18921 27031 18924
rect 26973 18915 27031 18921
rect 27154 18912 27160 18924
rect 27212 18912 27218 18964
rect 27430 18912 27436 18964
rect 27488 18952 27494 18964
rect 31021 18955 31079 18961
rect 27488 18924 30696 18952
rect 27488 18912 27494 18924
rect 21468 18884 21496 18912
rect 20180 18856 21496 18884
rect 17451 18853 17463 18856
rect 17405 18847 17463 18853
rect 13081 18819 13139 18825
rect 10888 18788 11100 18816
rect 10888 18748 10916 18788
rect 9140 18720 10916 18748
rect 10965 18751 11023 18757
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 10965 18717 10977 18751
rect 11011 18717 11023 18751
rect 11072 18748 11100 18788
rect 13081 18785 13093 18819
rect 13127 18785 13139 18819
rect 13081 18779 13139 18785
rect 15286 18776 15292 18828
rect 15344 18776 15350 18828
rect 16577 18819 16635 18825
rect 16577 18785 16589 18819
rect 16623 18816 16635 18819
rect 16758 18816 16764 18828
rect 16623 18788 16764 18816
rect 16623 18785 16635 18788
rect 16577 18779 16635 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 17512 18825 17540 18856
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18138 18776 18144 18828
rect 18196 18776 18202 18828
rect 26329 18819 26387 18825
rect 26329 18816 26341 18819
rect 24872 18788 26341 18816
rect 11072 18720 11376 18748
rect 10965 18711 11023 18717
rect 4246 18640 4252 18692
rect 4304 18680 4310 18692
rect 6840 18680 6868 18711
rect 7466 18680 7472 18692
rect 4304 18652 5396 18680
rect 6840 18652 7472 18680
rect 4304 18640 4310 18652
rect 5368 18612 5396 18652
rect 7466 18640 7472 18652
rect 7524 18640 7530 18692
rect 8297 18683 8355 18689
rect 8297 18680 8309 18683
rect 7760 18652 8309 18680
rect 5810 18612 5816 18624
rect 5368 18584 5816 18612
rect 5810 18572 5816 18584
rect 5868 18612 5874 18624
rect 7377 18615 7435 18621
rect 7377 18612 7389 18615
rect 5868 18584 7389 18612
rect 5868 18572 5874 18584
rect 7377 18581 7389 18584
rect 7423 18612 7435 18615
rect 7760 18612 7788 18652
rect 8297 18649 8309 18652
rect 8343 18649 8355 18683
rect 8297 18643 8355 18649
rect 10321 18683 10379 18689
rect 10321 18649 10333 18683
rect 10367 18680 10379 18683
rect 10870 18680 10876 18692
rect 10367 18652 10876 18680
rect 10367 18649 10379 18652
rect 10321 18643 10379 18649
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 10980 18624 11008 18711
rect 11348 18692 11376 18720
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 12216 18720 12909 18748
rect 12216 18708 12222 18720
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 13814 18708 13820 18760
rect 13872 18708 13878 18760
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18748 17003 18751
rect 18156 18748 18184 18776
rect 16991 18720 18184 18748
rect 19061 18751 19119 18757
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 19061 18717 19073 18751
rect 19107 18748 19119 18751
rect 19150 18748 19156 18760
rect 19107 18720 19156 18748
rect 19107 18717 19119 18720
rect 19061 18711 19119 18717
rect 19150 18708 19156 18720
rect 19208 18748 19214 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19208 18720 19257 18748
rect 19208 18708 19214 18720
rect 19245 18717 19257 18720
rect 19291 18748 19303 18751
rect 20993 18751 21051 18757
rect 20993 18748 21005 18751
rect 19291 18720 21005 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 20993 18717 21005 18720
rect 21039 18748 21051 18751
rect 22462 18748 22468 18760
rect 21039 18720 22468 18748
rect 21039 18717 21051 18720
rect 20993 18711 21051 18717
rect 22462 18708 22468 18720
rect 22520 18748 22526 18760
rect 22557 18751 22615 18757
rect 22557 18748 22569 18751
rect 22520 18720 22569 18748
rect 22520 18708 22526 18720
rect 22557 18717 22569 18720
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 11210 18683 11268 18689
rect 11210 18680 11222 18683
rect 11112 18652 11222 18680
rect 11112 18640 11118 18652
rect 11210 18649 11222 18652
rect 11256 18649 11268 18683
rect 11210 18643 11268 18649
rect 11330 18640 11336 18692
rect 11388 18640 11394 18692
rect 12805 18683 12863 18689
rect 12805 18680 12817 18683
rect 11716 18652 12817 18680
rect 11716 18624 11744 18652
rect 12805 18649 12817 18652
rect 12851 18680 12863 18683
rect 13265 18683 13323 18689
rect 13265 18680 13277 18683
rect 12851 18652 13277 18680
rect 12851 18649 12863 18652
rect 12805 18643 12863 18649
rect 13265 18649 13277 18652
rect 13311 18649 13323 18683
rect 13265 18643 13323 18649
rect 14090 18640 14096 18692
rect 14148 18680 14154 18692
rect 19334 18680 19340 18692
rect 14148 18652 19340 18680
rect 14148 18640 14154 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 19512 18683 19570 18689
rect 19512 18649 19524 18683
rect 19558 18680 19570 18683
rect 19702 18680 19708 18692
rect 19558 18652 19708 18680
rect 19558 18649 19570 18652
rect 19512 18643 19570 18649
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 21910 18640 21916 18692
rect 21968 18640 21974 18692
rect 22186 18640 22192 18692
rect 22244 18689 22250 18692
rect 22244 18643 22256 18689
rect 22824 18683 22882 18689
rect 22824 18649 22836 18683
rect 22870 18680 22882 18683
rect 23014 18680 23020 18692
rect 22870 18652 23020 18680
rect 22870 18649 22882 18652
rect 22824 18643 22882 18649
rect 22244 18640 22250 18643
rect 23014 18640 23020 18652
rect 23072 18640 23078 18692
rect 7423 18584 7788 18612
rect 7423 18581 7435 18584
rect 7377 18575 7435 18581
rect 7834 18572 7840 18624
rect 7892 18572 7898 18624
rect 10226 18572 10232 18624
rect 10284 18572 10290 18624
rect 10962 18572 10968 18624
rect 11020 18572 11026 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12437 18615 12495 18621
rect 12437 18581 12449 18615
rect 12483 18612 12495 18615
rect 12986 18612 12992 18624
rect 12483 18584 12992 18612
rect 12483 18581 12495 18584
rect 12437 18575 12495 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 15657 18615 15715 18621
rect 15657 18612 15669 18615
rect 15252 18584 15669 18612
rect 15252 18572 15258 18584
rect 15657 18581 15669 18584
rect 15703 18612 15715 18615
rect 15838 18612 15844 18624
rect 15703 18584 15844 18612
rect 15703 18581 15715 18584
rect 15657 18575 15715 18581
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 17037 18615 17095 18621
rect 17037 18581 17049 18615
rect 17083 18612 17095 18615
rect 17126 18612 17132 18624
rect 17083 18584 17132 18612
rect 17083 18581 17095 18584
rect 17037 18575 17095 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 21928 18612 21956 18640
rect 21131 18584 21956 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 22002 18572 22008 18624
rect 22060 18612 22066 18624
rect 24872 18621 24900 18788
rect 26329 18785 26341 18788
rect 26375 18785 26387 18819
rect 27448 18816 27476 18912
rect 27525 18819 27583 18825
rect 27525 18816 27537 18819
rect 27448 18788 27537 18816
rect 26329 18779 26387 18785
rect 27525 18785 27537 18788
rect 27571 18785 27583 18819
rect 28353 18819 28411 18825
rect 28353 18816 28365 18819
rect 27525 18779 27583 18785
rect 27632 18788 28365 18816
rect 25590 18708 25596 18760
rect 25648 18708 25654 18760
rect 26970 18748 26976 18760
rect 26436 18720 26976 18748
rect 26145 18683 26203 18689
rect 26145 18649 26157 18683
rect 26191 18680 26203 18683
rect 26436 18680 26464 18720
rect 26970 18708 26976 18720
rect 27028 18748 27034 18760
rect 27433 18751 27491 18757
rect 27433 18748 27445 18751
rect 27028 18720 27445 18748
rect 27028 18708 27034 18720
rect 27433 18717 27445 18720
rect 27479 18717 27491 18751
rect 27433 18711 27491 18717
rect 26191 18652 26464 18680
rect 26191 18649 26203 18652
rect 26145 18643 26203 18649
rect 26436 18624 26464 18652
rect 27154 18640 27160 18692
rect 27212 18680 27218 18692
rect 27341 18683 27399 18689
rect 27341 18680 27353 18683
rect 27212 18652 27353 18680
rect 27212 18640 27218 18652
rect 27341 18649 27353 18652
rect 27387 18649 27399 18683
rect 27341 18643 27399 18649
rect 24857 18615 24915 18621
rect 24857 18612 24869 18615
rect 22060 18584 24869 18612
rect 22060 18572 22066 18584
rect 24857 18581 24869 18584
rect 24903 18581 24915 18615
rect 24857 18575 24915 18581
rect 25038 18572 25044 18624
rect 25096 18572 25102 18624
rect 26234 18572 26240 18624
rect 26292 18572 26298 18624
rect 26418 18572 26424 18624
rect 26476 18572 26482 18624
rect 26510 18572 26516 18624
rect 26568 18612 26574 18624
rect 26789 18615 26847 18621
rect 26789 18612 26801 18615
rect 26568 18584 26801 18612
rect 26568 18572 26574 18584
rect 26789 18581 26801 18584
rect 26835 18612 26847 18615
rect 27632 18612 27660 18788
rect 28353 18785 28365 18788
rect 28399 18785 28411 18819
rect 28353 18779 28411 18785
rect 27706 18708 27712 18760
rect 27764 18748 27770 18760
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 27764 18720 28181 18748
rect 27764 18708 27770 18720
rect 28169 18717 28181 18720
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 28368 18680 28396 18779
rect 29638 18776 29644 18828
rect 29696 18776 29702 18828
rect 29546 18708 29552 18760
rect 29604 18748 29610 18760
rect 29897 18751 29955 18757
rect 29897 18748 29909 18751
rect 29604 18720 29909 18748
rect 29604 18708 29610 18720
rect 29897 18717 29909 18720
rect 29943 18717 29955 18751
rect 30668 18748 30696 18924
rect 31021 18921 31033 18955
rect 31067 18952 31079 18955
rect 31294 18952 31300 18964
rect 31067 18924 31300 18952
rect 31067 18921 31079 18924
rect 31021 18915 31079 18921
rect 31294 18912 31300 18924
rect 31352 18912 31358 18964
rect 32398 18952 32404 18964
rect 31864 18924 32404 18952
rect 31864 18896 31892 18924
rect 32398 18912 32404 18924
rect 32456 18952 32462 18964
rect 34333 18955 34391 18961
rect 32456 18924 32904 18952
rect 32456 18912 32462 18924
rect 31846 18844 31852 18896
rect 31904 18844 31910 18896
rect 32876 18893 32904 18924
rect 34333 18921 34345 18955
rect 34379 18952 34391 18955
rect 34698 18952 34704 18964
rect 34379 18924 34704 18952
rect 34379 18921 34391 18924
rect 34333 18915 34391 18921
rect 34698 18912 34704 18924
rect 34756 18912 34762 18964
rect 36906 18912 36912 18964
rect 36964 18912 36970 18964
rect 37642 18912 37648 18964
rect 37700 18952 37706 18964
rect 39206 18952 39212 18964
rect 37700 18924 39212 18952
rect 37700 18912 37706 18924
rect 39206 18912 39212 18924
rect 39264 18912 39270 18964
rect 40589 18955 40647 18961
rect 40589 18921 40601 18955
rect 40635 18952 40647 18955
rect 40954 18952 40960 18964
rect 40635 18924 40960 18952
rect 40635 18921 40647 18924
rect 40589 18915 40647 18921
rect 40954 18912 40960 18924
rect 41012 18912 41018 18964
rect 41693 18955 41751 18961
rect 41693 18921 41705 18955
rect 41739 18952 41751 18955
rect 41966 18952 41972 18964
rect 41739 18924 41972 18952
rect 41739 18921 41751 18924
rect 41693 18915 41751 18921
rect 41966 18912 41972 18924
rect 42024 18912 42030 18964
rect 42518 18912 42524 18964
rect 42576 18952 42582 18964
rect 42797 18955 42855 18961
rect 42797 18952 42809 18955
rect 42576 18924 42809 18952
rect 42576 18912 42582 18924
rect 42797 18921 42809 18924
rect 42843 18952 42855 18955
rect 45830 18952 45836 18964
rect 42843 18924 45836 18952
rect 42843 18921 42855 18924
rect 42797 18915 42855 18921
rect 45830 18912 45836 18924
rect 45888 18912 45894 18964
rect 46661 18955 46719 18961
rect 46661 18921 46673 18955
rect 46707 18952 46719 18955
rect 46750 18952 46756 18964
rect 46707 18924 46756 18952
rect 46707 18921 46719 18924
rect 46661 18915 46719 18921
rect 46750 18912 46756 18924
rect 46808 18912 46814 18964
rect 48222 18952 48228 18964
rect 46952 18924 48228 18952
rect 32861 18887 32919 18893
rect 32861 18853 32873 18887
rect 32907 18853 32919 18887
rect 46293 18887 46351 18893
rect 46293 18884 46305 18887
rect 32861 18847 32919 18853
rect 45664 18856 46305 18884
rect 31938 18776 31944 18828
rect 31996 18816 32002 18828
rect 31996 18788 32435 18816
rect 31996 18776 32002 18788
rect 30668 18720 31754 18748
rect 29897 18711 29955 18717
rect 31726 18692 31754 18720
rect 32306 18708 32312 18760
rect 32364 18708 32370 18760
rect 32407 18748 32435 18788
rect 32766 18776 32772 18828
rect 32824 18816 32830 18828
rect 32824 18788 33640 18816
rect 32824 18776 32830 18788
rect 32468 18751 32526 18757
rect 32468 18748 32480 18751
rect 32407 18720 32480 18748
rect 32468 18717 32480 18720
rect 32514 18717 32526 18751
rect 32468 18711 32526 18717
rect 32582 18708 32588 18760
rect 32640 18708 32646 18760
rect 33321 18751 33379 18757
rect 33321 18717 33333 18751
rect 33367 18717 33379 18751
rect 33321 18711 33379 18717
rect 29638 18680 29644 18692
rect 28368 18652 29644 18680
rect 29638 18640 29644 18652
rect 29696 18640 29702 18692
rect 31726 18652 31760 18692
rect 31754 18640 31760 18652
rect 31812 18640 31818 18692
rect 33336 18680 33364 18711
rect 33410 18708 33416 18760
rect 33468 18748 33474 18760
rect 33505 18751 33563 18757
rect 33505 18748 33517 18751
rect 33468 18720 33517 18748
rect 33468 18708 33474 18720
rect 33505 18717 33517 18720
rect 33551 18717 33563 18751
rect 33612 18748 33640 18788
rect 33686 18776 33692 18828
rect 33744 18776 33750 18828
rect 35250 18776 35256 18828
rect 35308 18776 35314 18828
rect 35434 18776 35440 18828
rect 35492 18816 35498 18828
rect 35989 18819 36047 18825
rect 35989 18816 36001 18819
rect 35492 18788 36001 18816
rect 35492 18776 35498 18788
rect 35989 18785 36001 18788
rect 36035 18816 36047 18819
rect 36633 18819 36691 18825
rect 36633 18816 36645 18819
rect 36035 18788 36645 18816
rect 36035 18785 36047 18788
rect 35989 18779 36047 18785
rect 36633 18785 36645 18788
rect 36679 18785 36691 18819
rect 36633 18779 36691 18785
rect 36722 18776 36728 18828
rect 36780 18816 36786 18828
rect 37461 18819 37519 18825
rect 37461 18816 37473 18819
rect 36780 18788 37473 18816
rect 36780 18776 36786 18788
rect 37461 18785 37473 18788
rect 37507 18785 37519 18819
rect 37918 18816 37924 18828
rect 37461 18779 37519 18785
rect 37844 18788 37924 18816
rect 33873 18751 33931 18757
rect 33873 18748 33885 18751
rect 33612 18720 33885 18748
rect 33505 18711 33563 18717
rect 33873 18717 33885 18720
rect 33919 18717 33931 18751
rect 33873 18711 33931 18717
rect 37369 18751 37427 18757
rect 37369 18717 37381 18751
rect 37415 18748 37427 18751
rect 37844 18748 37872 18788
rect 37918 18776 37924 18788
rect 37976 18776 37982 18828
rect 40037 18819 40095 18825
rect 40037 18785 40049 18819
rect 40083 18785 40095 18819
rect 40037 18779 40095 18785
rect 38105 18751 38163 18757
rect 38105 18748 38117 18751
rect 37415 18720 37872 18748
rect 37936 18720 38117 18748
rect 37415 18717 37427 18720
rect 37369 18711 37427 18717
rect 33965 18683 34023 18689
rect 33965 18680 33977 18683
rect 33336 18652 33977 18680
rect 33965 18649 33977 18652
rect 34011 18680 34023 18683
rect 34701 18683 34759 18689
rect 34701 18680 34713 18683
rect 34011 18652 34713 18680
rect 34011 18649 34023 18652
rect 33965 18643 34023 18649
rect 34701 18649 34713 18652
rect 34747 18649 34759 18683
rect 34701 18643 34759 18649
rect 36449 18683 36507 18689
rect 36449 18649 36461 18683
rect 36495 18680 36507 18683
rect 37734 18680 37740 18692
rect 36495 18652 37740 18680
rect 36495 18649 36507 18652
rect 36449 18643 36507 18649
rect 37734 18640 37740 18652
rect 37792 18640 37798 18692
rect 26835 18584 27660 18612
rect 26835 18581 26847 18584
rect 26789 18575 26847 18581
rect 27798 18572 27804 18624
rect 27856 18572 27862 18624
rect 28261 18615 28319 18621
rect 28261 18581 28273 18615
rect 28307 18612 28319 18615
rect 28810 18612 28816 18624
rect 28307 18584 28816 18612
rect 28307 18581 28319 18584
rect 28261 18575 28319 18581
rect 28810 18572 28816 18584
rect 28868 18572 28874 18624
rect 30374 18572 30380 18624
rect 30432 18612 30438 18624
rect 31389 18615 31447 18621
rect 31389 18612 31401 18615
rect 30432 18584 31401 18612
rect 30432 18572 30438 18584
rect 31389 18581 31401 18584
rect 31435 18581 31447 18615
rect 31389 18575 31447 18581
rect 31665 18615 31723 18621
rect 31665 18581 31677 18615
rect 31711 18612 31723 18615
rect 32858 18612 32864 18624
rect 31711 18584 32864 18612
rect 31711 18581 31723 18584
rect 31665 18575 31723 18581
rect 32858 18572 32864 18584
rect 32916 18572 32922 18624
rect 36078 18572 36084 18624
rect 36136 18572 36142 18624
rect 36541 18615 36599 18621
rect 36541 18581 36553 18615
rect 36587 18612 36599 18615
rect 37274 18612 37280 18624
rect 36587 18584 37280 18612
rect 36587 18581 36599 18584
rect 36541 18575 36599 18581
rect 37274 18572 37280 18584
rect 37332 18572 37338 18624
rect 37458 18572 37464 18624
rect 37516 18612 37522 18624
rect 37936 18621 37964 18720
rect 38105 18717 38117 18720
rect 38151 18748 38163 18751
rect 38654 18748 38660 18760
rect 38151 18720 38660 18748
rect 38151 18717 38163 18720
rect 38105 18711 38163 18717
rect 38654 18708 38660 18720
rect 38712 18708 38718 18760
rect 39942 18708 39948 18760
rect 40000 18748 40006 18760
rect 40052 18748 40080 18779
rect 41046 18776 41052 18828
rect 41104 18816 41110 18828
rect 41233 18819 41291 18825
rect 41233 18816 41245 18819
rect 41104 18788 41245 18816
rect 41104 18776 41110 18788
rect 41233 18785 41245 18788
rect 41279 18785 41291 18819
rect 41233 18779 41291 18785
rect 41874 18776 41880 18828
rect 41932 18816 41938 18828
rect 42245 18819 42303 18825
rect 42245 18816 42257 18819
rect 41932 18788 42257 18816
rect 41932 18776 41938 18788
rect 42245 18785 42257 18788
rect 42291 18785 42303 18819
rect 42245 18779 42303 18785
rect 43346 18776 43352 18828
rect 43404 18816 43410 18828
rect 43404 18788 43567 18816
rect 43404 18776 43410 18788
rect 40000 18720 40080 18748
rect 40000 18708 40006 18720
rect 40218 18708 40224 18760
rect 40276 18748 40282 18760
rect 40681 18751 40739 18757
rect 40681 18748 40693 18751
rect 40276 18720 40693 18748
rect 40276 18708 40282 18720
rect 40681 18717 40693 18720
rect 40727 18717 40739 18751
rect 40681 18711 40739 18717
rect 42061 18751 42119 18757
rect 42061 18717 42073 18751
rect 42107 18748 42119 18751
rect 42886 18748 42892 18760
rect 42107 18720 42892 18748
rect 42107 18717 42119 18720
rect 42061 18711 42119 18717
rect 42886 18708 42892 18720
rect 42944 18708 42950 18760
rect 43539 18757 43567 18788
rect 44082 18776 44088 18828
rect 44140 18776 44146 18828
rect 44634 18776 44640 18828
rect 44692 18816 44698 18828
rect 44729 18819 44787 18825
rect 44729 18816 44741 18819
rect 44692 18788 44741 18816
rect 44692 18776 44698 18788
rect 44729 18785 44741 18788
rect 44775 18785 44787 18819
rect 44729 18779 44787 18785
rect 43714 18757 43720 18760
rect 43533 18751 43591 18757
rect 43533 18717 43545 18751
rect 43579 18717 43591 18751
rect 43533 18711 43591 18717
rect 43692 18751 43720 18757
rect 43692 18717 43704 18751
rect 43692 18711 43720 18717
rect 43714 18708 43720 18711
rect 43772 18708 43778 18760
rect 43806 18708 43812 18760
rect 43864 18708 43870 18760
rect 44545 18751 44603 18757
rect 44545 18717 44557 18751
rect 44591 18748 44603 18751
rect 45370 18748 45376 18760
rect 44591 18720 45376 18748
rect 44591 18717 44603 18720
rect 44545 18711 44603 18717
rect 45370 18708 45376 18720
rect 45428 18708 45434 18760
rect 38372 18683 38430 18689
rect 38372 18649 38384 18683
rect 38418 18680 38430 18683
rect 38470 18680 38476 18692
rect 38418 18652 38476 18680
rect 38418 18649 38430 18652
rect 38372 18643 38430 18649
rect 38470 18640 38476 18652
rect 38528 18640 38534 18692
rect 38930 18640 38936 18692
rect 38988 18680 38994 18692
rect 38988 18652 40172 18680
rect 38988 18640 38994 18652
rect 40144 18624 40172 18652
rect 45002 18640 45008 18692
rect 45060 18680 45066 18692
rect 45664 18680 45692 18856
rect 46293 18853 46305 18856
rect 46339 18884 46351 18887
rect 46952 18884 46980 18924
rect 48222 18912 48228 18924
rect 48280 18952 48286 18964
rect 48866 18952 48872 18964
rect 48280 18924 48872 18952
rect 48280 18912 48286 18924
rect 48866 18912 48872 18924
rect 48924 18912 48930 18964
rect 49694 18912 49700 18964
rect 49752 18912 49758 18964
rect 49973 18955 50031 18961
rect 49973 18921 49985 18955
rect 50019 18952 50031 18955
rect 50062 18952 50068 18964
rect 50019 18924 50068 18952
rect 50019 18921 50031 18924
rect 49973 18915 50031 18921
rect 50062 18912 50068 18924
rect 50120 18912 50126 18964
rect 54113 18955 54171 18961
rect 50172 18924 53604 18952
rect 46339 18856 46980 18884
rect 49712 18884 49740 18912
rect 50172 18884 50200 18924
rect 49712 18856 50200 18884
rect 46339 18853 46351 18856
rect 46293 18847 46351 18853
rect 48041 18819 48099 18825
rect 48041 18785 48053 18819
rect 48087 18816 48099 18819
rect 48130 18816 48136 18828
rect 48087 18788 48136 18816
rect 48087 18785 48099 18788
rect 48041 18779 48099 18785
rect 48130 18776 48136 18788
rect 48188 18816 48194 18828
rect 48188 18788 49464 18816
rect 48188 18776 48194 18788
rect 48314 18708 48320 18760
rect 48372 18748 48378 18760
rect 48685 18751 48743 18757
rect 48685 18748 48697 18751
rect 48372 18720 48697 18748
rect 48372 18708 48378 18720
rect 48685 18717 48697 18720
rect 48731 18717 48743 18751
rect 48685 18711 48743 18717
rect 49329 18751 49387 18757
rect 49329 18717 49341 18751
rect 49375 18717 49387 18751
rect 49436 18748 49464 18788
rect 51537 18751 51595 18757
rect 51537 18748 51549 18751
rect 49436 18720 51549 18748
rect 49329 18711 49387 18717
rect 45060 18652 45692 18680
rect 45741 18683 45799 18689
rect 45060 18640 45066 18652
rect 45741 18649 45753 18683
rect 45787 18649 45799 18683
rect 45741 18643 45799 18649
rect 47796 18683 47854 18689
rect 47796 18649 47808 18683
rect 47842 18680 47854 18683
rect 48133 18683 48191 18689
rect 48133 18680 48145 18683
rect 47842 18652 48145 18680
rect 47842 18649 47854 18652
rect 47796 18643 47854 18649
rect 48133 18649 48145 18652
rect 48179 18649 48191 18683
rect 48133 18643 48191 18649
rect 37921 18615 37979 18621
rect 37921 18612 37933 18615
rect 37516 18584 37933 18612
rect 37516 18572 37522 18584
rect 37921 18581 37933 18584
rect 37967 18581 37979 18615
rect 37921 18575 37979 18581
rect 39485 18615 39543 18621
rect 39485 18581 39497 18615
rect 39531 18612 39543 18615
rect 39850 18612 39856 18624
rect 39531 18584 39856 18612
rect 39531 18581 39543 18584
rect 39485 18575 39543 18581
rect 39850 18572 39856 18584
rect 39908 18572 39914 18624
rect 40126 18572 40132 18624
rect 40184 18572 40190 18624
rect 42153 18615 42211 18621
rect 42153 18581 42165 18615
rect 42199 18612 42211 18615
rect 42610 18612 42616 18624
rect 42199 18584 42616 18612
rect 42199 18581 42211 18584
rect 42153 18575 42211 18581
rect 42610 18572 42616 18584
rect 42668 18572 42674 18624
rect 42889 18615 42947 18621
rect 42889 18581 42901 18615
rect 42935 18612 42947 18615
rect 44174 18612 44180 18624
rect 42935 18584 44180 18612
rect 42935 18581 42947 18584
rect 42889 18575 42947 18581
rect 44174 18572 44180 18584
rect 44232 18572 44238 18624
rect 45278 18572 45284 18624
rect 45336 18612 45342 18624
rect 45756 18612 45784 18643
rect 49050 18640 49056 18692
rect 49108 18640 49114 18692
rect 49344 18680 49372 18711
rect 51184 18692 51212 18720
rect 51537 18717 51549 18720
rect 51583 18748 51595 18751
rect 51813 18751 51871 18757
rect 51813 18748 51825 18751
rect 51583 18720 51825 18748
rect 51583 18717 51595 18720
rect 51537 18711 51595 18717
rect 51813 18717 51825 18720
rect 51859 18748 51871 18751
rect 51902 18748 51908 18760
rect 51859 18720 51908 18748
rect 51859 18717 51871 18720
rect 51813 18711 51871 18717
rect 51902 18708 51908 18720
rect 51960 18708 51966 18760
rect 49344 18652 50200 18680
rect 47394 18612 47400 18624
rect 45336 18584 47400 18612
rect 45336 18572 45342 18584
rect 47394 18572 47400 18584
rect 47452 18612 47458 18624
rect 49068 18612 49096 18640
rect 50172 18621 50200 18652
rect 51166 18640 51172 18692
rect 51224 18640 51230 18692
rect 51292 18683 51350 18689
rect 51292 18649 51304 18683
rect 51338 18680 51350 18683
rect 51626 18680 51632 18692
rect 51338 18652 51632 18680
rect 51338 18649 51350 18652
rect 51292 18643 51350 18649
rect 51626 18640 51632 18652
rect 51684 18640 51690 18692
rect 52080 18683 52138 18689
rect 52080 18649 52092 18683
rect 52126 18680 52138 18683
rect 52730 18680 52736 18692
rect 52126 18652 52736 18680
rect 52126 18649 52138 18652
rect 52080 18643 52138 18649
rect 52730 18640 52736 18652
rect 52788 18640 52794 18692
rect 53576 18680 53604 18924
rect 54113 18921 54125 18955
rect 54159 18952 54171 18955
rect 54202 18952 54208 18964
rect 54159 18924 54208 18952
rect 54159 18921 54171 18924
rect 54113 18915 54171 18921
rect 54202 18912 54208 18924
rect 54260 18912 54266 18964
rect 55953 18955 56011 18961
rect 55953 18921 55965 18955
rect 55999 18952 56011 18955
rect 56134 18952 56140 18964
rect 55999 18924 56140 18952
rect 55999 18921 56011 18924
rect 55953 18915 56011 18921
rect 53650 18844 53656 18896
rect 53708 18844 53714 18896
rect 54478 18844 54484 18896
rect 54536 18884 54542 18896
rect 54536 18856 54708 18884
rect 54536 18844 54542 18856
rect 53668 18816 53696 18844
rect 54680 18825 54708 18856
rect 53837 18819 53895 18825
rect 53837 18816 53849 18819
rect 53668 18788 53849 18816
rect 53837 18785 53849 18788
rect 53883 18785 53895 18819
rect 53837 18779 53895 18785
rect 54665 18819 54723 18825
rect 54665 18785 54677 18819
rect 54711 18785 54723 18819
rect 54665 18779 54723 18785
rect 55214 18776 55220 18828
rect 55272 18816 55278 18828
rect 55309 18819 55367 18825
rect 55309 18816 55321 18819
rect 55272 18788 55321 18816
rect 55272 18776 55278 18788
rect 55309 18785 55321 18788
rect 55355 18785 55367 18819
rect 55309 18779 55367 18785
rect 53653 18751 53711 18757
rect 53653 18717 53665 18751
rect 53699 18748 53711 18751
rect 54386 18748 54392 18760
rect 53699 18720 54392 18748
rect 53699 18717 53711 18720
rect 53653 18711 53711 18717
rect 54386 18708 54392 18720
rect 54444 18708 54450 18760
rect 54481 18751 54539 18757
rect 54481 18717 54493 18751
rect 54527 18748 54539 18751
rect 55968 18748 55996 18915
rect 56134 18912 56140 18924
rect 56192 18912 56198 18964
rect 56781 18955 56839 18961
rect 56781 18921 56793 18955
rect 56827 18952 56839 18955
rect 57330 18952 57336 18964
rect 56827 18924 57336 18952
rect 56827 18921 56839 18924
rect 56781 18915 56839 18921
rect 57330 18912 57336 18924
rect 57388 18912 57394 18964
rect 57514 18912 57520 18964
rect 57572 18952 57578 18964
rect 57701 18955 57759 18961
rect 57701 18952 57713 18955
rect 57572 18924 57713 18952
rect 57572 18912 57578 18924
rect 57701 18921 57713 18924
rect 57747 18921 57759 18955
rect 57701 18915 57759 18921
rect 57333 18819 57391 18825
rect 57333 18816 57345 18819
rect 54527 18720 55996 18748
rect 56612 18788 57345 18816
rect 54527 18717 54539 18720
rect 54481 18711 54539 18717
rect 56612 18689 56640 18788
rect 57333 18785 57345 18788
rect 57379 18785 57391 18819
rect 57333 18779 57391 18785
rect 58250 18776 58256 18828
rect 58308 18776 58314 18828
rect 57149 18751 57207 18757
rect 57149 18717 57161 18751
rect 57195 18748 57207 18751
rect 57238 18748 57244 18760
rect 57195 18720 57244 18748
rect 57195 18717 57207 18720
rect 57149 18711 57207 18717
rect 57238 18708 57244 18720
rect 57296 18708 57302 18760
rect 56597 18683 56655 18689
rect 56597 18680 56609 18683
rect 53576 18652 56609 18680
rect 56597 18649 56609 18652
rect 56643 18649 56655 18683
rect 56597 18643 56655 18649
rect 47452 18584 49096 18612
rect 50157 18615 50215 18621
rect 47452 18572 47458 18584
rect 50157 18581 50169 18615
rect 50203 18581 50215 18615
rect 50157 18575 50215 18581
rect 53190 18572 53196 18624
rect 53248 18572 53254 18624
rect 53282 18572 53288 18624
rect 53340 18572 53346 18624
rect 53742 18572 53748 18624
rect 53800 18572 53806 18624
rect 54573 18615 54631 18621
rect 54573 18581 54585 18615
rect 54619 18612 54631 18615
rect 54662 18612 54668 18624
rect 54619 18584 54668 18612
rect 54619 18581 54631 18584
rect 54573 18575 54631 18581
rect 54662 18572 54668 18584
rect 54720 18612 54726 18624
rect 57241 18615 57299 18621
rect 57241 18612 57253 18615
rect 54720 18584 57253 18612
rect 54720 18572 54726 18584
rect 57241 18581 57253 18584
rect 57287 18612 57299 18615
rect 57606 18612 57612 18624
rect 57287 18584 57612 18612
rect 57287 18581 57299 18584
rect 57241 18575 57299 18581
rect 57606 18572 57612 18584
rect 57664 18572 57670 18624
rect 1104 18522 59040 18544
rect 1104 18470 15394 18522
rect 15446 18470 15458 18522
rect 15510 18470 15522 18522
rect 15574 18470 15586 18522
rect 15638 18470 15650 18522
rect 15702 18470 29838 18522
rect 29890 18470 29902 18522
rect 29954 18470 29966 18522
rect 30018 18470 30030 18522
rect 30082 18470 30094 18522
rect 30146 18470 44282 18522
rect 44334 18470 44346 18522
rect 44398 18470 44410 18522
rect 44462 18470 44474 18522
rect 44526 18470 44538 18522
rect 44590 18470 58726 18522
rect 58778 18470 58790 18522
rect 58842 18470 58854 18522
rect 58906 18470 58918 18522
rect 58970 18470 58982 18522
rect 59034 18470 59040 18522
rect 1104 18448 59040 18470
rect 4798 18368 4804 18420
rect 4856 18368 4862 18420
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 7524 18380 7849 18408
rect 7524 18368 7530 18380
rect 7837 18377 7849 18380
rect 7883 18377 7895 18411
rect 7837 18371 7895 18377
rect 10594 18368 10600 18420
rect 10652 18368 10658 18420
rect 10689 18411 10747 18417
rect 10689 18377 10701 18411
rect 10735 18408 10747 18411
rect 11054 18408 11060 18420
rect 10735 18380 11060 18408
rect 10735 18377 10747 18380
rect 10689 18371 10747 18377
rect 11054 18368 11060 18380
rect 11112 18368 11118 18420
rect 13817 18411 13875 18417
rect 13817 18377 13829 18411
rect 13863 18408 13875 18411
rect 13906 18408 13912 18420
rect 13863 18380 13912 18408
rect 13863 18377 13875 18380
rect 13817 18371 13875 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 19150 18368 19156 18420
rect 19208 18368 19214 18420
rect 20533 18411 20591 18417
rect 20533 18377 20545 18411
rect 20579 18408 20591 18411
rect 20806 18408 20812 18420
rect 20579 18380 20812 18408
rect 20579 18377 20591 18380
rect 20533 18371 20591 18377
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 21082 18368 21088 18420
rect 21140 18368 21146 18420
rect 21174 18368 21180 18420
rect 21232 18408 21238 18420
rect 27982 18408 27988 18420
rect 21232 18380 24992 18408
rect 21232 18368 21238 18380
rect 4816 18068 4844 18368
rect 6181 18343 6239 18349
rect 6181 18309 6193 18343
rect 6227 18340 6239 18343
rect 6227 18312 7788 18340
rect 6227 18309 6239 18312
rect 6181 18303 6239 18309
rect 7760 18284 7788 18312
rect 9232 18312 11008 18340
rect 6365 18275 6423 18281
rect 6365 18241 6377 18275
rect 6411 18272 6423 18275
rect 6454 18272 6460 18284
rect 6411 18244 6460 18272
rect 6411 18241 6423 18244
rect 6365 18235 6423 18241
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 6632 18275 6690 18281
rect 6632 18241 6644 18275
rect 6678 18272 6690 18275
rect 6914 18272 6920 18284
rect 6678 18244 6920 18272
rect 6678 18241 6690 18244
rect 6632 18235 6690 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7742 18232 7748 18284
rect 7800 18232 7806 18284
rect 9122 18232 9128 18284
rect 9180 18272 9186 18284
rect 9232 18281 9260 18312
rect 10980 18284 11008 18312
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 9180 18244 9229 18272
rect 9180 18232 9186 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9484 18275 9542 18281
rect 9484 18241 9496 18275
rect 9530 18272 9542 18275
rect 9766 18272 9772 18284
rect 9530 18244 9772 18272
rect 9530 18241 9542 18244
rect 9484 18235 9542 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 11882 18232 11888 18284
rect 11940 18232 11946 18284
rect 19168 18281 19196 18368
rect 20714 18300 20720 18352
rect 20772 18340 20778 18352
rect 20993 18343 21051 18349
rect 20993 18340 21005 18343
rect 20772 18312 21005 18340
rect 20772 18300 20778 18312
rect 20993 18309 21005 18312
rect 21039 18340 21051 18343
rect 22094 18340 22100 18352
rect 21039 18312 22100 18340
rect 21039 18309 21051 18312
rect 20993 18303 21051 18309
rect 22094 18300 22100 18312
rect 22152 18340 22158 18352
rect 22189 18343 22247 18349
rect 22189 18340 22201 18343
rect 22152 18312 22201 18340
rect 22152 18300 22158 18312
rect 22189 18309 22201 18312
rect 22235 18309 22247 18343
rect 22189 18303 22247 18309
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18272 13415 18275
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13403 18244 13737 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19420 18275 19478 18281
rect 19420 18241 19432 18275
rect 19466 18272 19478 18275
rect 19702 18272 19708 18284
rect 19466 18244 19708 18272
rect 19466 18241 19478 18244
rect 19420 18235 19478 18241
rect 19702 18232 19708 18244
rect 19760 18232 19766 18284
rect 21726 18232 21732 18284
rect 21784 18272 21790 18284
rect 22281 18275 22339 18281
rect 21784 18244 22241 18272
rect 21784 18232 21790 18244
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18173 8447 18207
rect 8389 18167 8447 18173
rect 7745 18139 7803 18145
rect 7745 18105 7757 18139
rect 7791 18136 7803 18139
rect 8404 18136 8432 18167
rect 11238 18164 11244 18216
rect 11296 18164 11302 18216
rect 11517 18207 11575 18213
rect 11517 18173 11529 18207
rect 11563 18204 11575 18207
rect 11900 18204 11928 18232
rect 11563 18176 11928 18204
rect 11563 18173 11575 18176
rect 11517 18167 11575 18173
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12124 18176 12449 18204
rect 12124 18164 12130 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12526 18164 12532 18216
rect 12584 18213 12590 18216
rect 12584 18207 12612 18213
rect 12600 18173 12612 18207
rect 12584 18167 12612 18173
rect 12584 18164 12590 18167
rect 12710 18164 12716 18216
rect 12768 18164 12774 18216
rect 13633 18207 13691 18213
rect 13633 18173 13645 18207
rect 13679 18204 13691 18207
rect 16390 18204 16396 18216
rect 13679 18176 16396 18204
rect 13679 18173 13691 18176
rect 13633 18167 13691 18173
rect 13740 18148 13768 18176
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 20990 18164 20996 18216
rect 21048 18204 21054 18216
rect 21177 18207 21235 18213
rect 21177 18204 21189 18207
rect 21048 18176 21189 18204
rect 21048 18164 21054 18176
rect 21177 18173 21189 18176
rect 21223 18204 21235 18207
rect 22002 18204 22008 18216
rect 21223 18176 22008 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 22002 18164 22008 18176
rect 22060 18164 22066 18216
rect 22213 18204 22241 18244
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 22649 18275 22707 18281
rect 22649 18272 22661 18275
rect 22327 18244 22661 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 22649 18241 22661 18244
rect 22695 18241 22707 18275
rect 24765 18275 24823 18281
rect 24765 18272 24777 18275
rect 22649 18235 22707 18241
rect 24044 18244 24777 18272
rect 22373 18207 22431 18213
rect 22373 18204 22385 18207
rect 22213 18176 22385 18204
rect 22373 18173 22385 18176
rect 22419 18173 22431 18207
rect 22373 18167 22431 18173
rect 22554 18164 22560 18216
rect 22612 18204 22618 18216
rect 23014 18204 23020 18216
rect 22612 18176 23020 18204
rect 22612 18164 22618 18176
rect 23014 18164 23020 18176
rect 23072 18164 23078 18216
rect 23201 18207 23259 18213
rect 23201 18173 23213 18207
rect 23247 18173 23259 18207
rect 23201 18167 23259 18173
rect 7791 18108 8432 18136
rect 8680 18108 9260 18136
rect 7791 18105 7803 18108
rect 7745 18099 7803 18105
rect 8680 18068 8708 18108
rect 4816 18040 8708 18068
rect 8754 18028 8760 18080
rect 8812 18028 8818 18080
rect 9232 18068 9260 18108
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 11112 18108 12173 18136
rect 11112 18096 11118 18108
rect 12161 18105 12173 18108
rect 12207 18136 12219 18139
rect 12250 18136 12256 18148
rect 12207 18108 12256 18136
rect 12207 18105 12219 18108
rect 12161 18099 12219 18105
rect 12250 18096 12256 18108
rect 12308 18096 12314 18148
rect 13722 18096 13728 18148
rect 13780 18096 13786 18148
rect 21910 18096 21916 18148
rect 21968 18136 21974 18148
rect 23216 18136 23244 18167
rect 21968 18108 23244 18136
rect 21968 18096 21974 18108
rect 9858 18068 9864 18080
rect 9232 18040 9864 18068
rect 9858 18028 9864 18040
rect 9916 18068 9922 18080
rect 14090 18068 14096 18080
rect 9916 18040 14096 18068
rect 9916 18028 9922 18040
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14182 18028 14188 18080
rect 14240 18028 14246 18080
rect 20625 18071 20683 18077
rect 20625 18037 20637 18071
rect 20671 18068 20683 18071
rect 20714 18068 20720 18080
rect 20671 18040 20720 18068
rect 20671 18037 20683 18040
rect 20625 18031 20683 18037
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 21818 18028 21824 18080
rect 21876 18028 21882 18080
rect 22462 18028 22468 18080
rect 22520 18068 22526 18080
rect 23382 18068 23388 18080
rect 22520 18040 23388 18068
rect 22520 18028 22526 18040
rect 23382 18028 23388 18040
rect 23440 18068 23446 18080
rect 24044 18077 24072 18244
rect 24765 18241 24777 18244
rect 24811 18272 24823 18275
rect 24854 18272 24860 18284
rect 24811 18244 24860 18272
rect 24811 18241 24823 18244
rect 24765 18235 24823 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 24964 18272 24992 18380
rect 26712 18380 27988 18408
rect 25038 18349 25044 18352
rect 25032 18303 25044 18349
rect 25096 18340 25102 18352
rect 26712 18349 26740 18380
rect 27982 18368 27988 18380
rect 28040 18408 28046 18420
rect 28166 18408 28172 18420
rect 28040 18380 28172 18408
rect 28040 18368 28046 18380
rect 28166 18368 28172 18380
rect 28224 18408 28230 18420
rect 28224 18380 29592 18408
rect 28224 18368 28230 18380
rect 26697 18343 26755 18349
rect 26697 18340 26709 18343
rect 25096 18312 25132 18340
rect 26160 18312 26709 18340
rect 25038 18300 25044 18303
rect 25096 18300 25102 18312
rect 26160 18272 26188 18312
rect 26697 18309 26709 18312
rect 26743 18309 26755 18343
rect 26697 18303 26755 18309
rect 28810 18300 28816 18352
rect 28868 18300 28874 18352
rect 29564 18340 29592 18380
rect 29638 18368 29644 18420
rect 29696 18408 29702 18420
rect 29696 18380 29960 18408
rect 29696 18368 29702 18380
rect 29822 18349 29828 18352
rect 29564 18312 29684 18340
rect 24964 18244 26188 18272
rect 26234 18232 26240 18284
rect 26292 18272 26298 18284
rect 27062 18272 27068 18284
rect 26292 18244 27068 18272
rect 26292 18232 26298 18244
rect 27062 18232 27068 18244
rect 27120 18272 27126 18284
rect 27120 18244 27292 18272
rect 27120 18232 27126 18244
rect 26878 18164 26884 18216
rect 26936 18204 26942 18216
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26936 18176 26985 18204
rect 26936 18164 26942 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 27154 18164 27160 18216
rect 27212 18164 27218 18216
rect 27264 18204 27292 18244
rect 28166 18232 28172 18284
rect 28224 18232 28230 18284
rect 29549 18275 29607 18281
rect 29549 18241 29561 18275
rect 29595 18241 29607 18275
rect 29656 18272 29684 18312
rect 29816 18303 29828 18349
rect 29822 18300 29828 18303
rect 29880 18300 29886 18352
rect 29932 18340 29960 18380
rect 30190 18368 30196 18420
rect 30248 18408 30254 18420
rect 31021 18411 31079 18417
rect 31021 18408 31033 18411
rect 30248 18380 31033 18408
rect 30248 18368 30254 18380
rect 31021 18377 31033 18380
rect 31067 18377 31079 18411
rect 31021 18371 31079 18377
rect 31389 18411 31447 18417
rect 31389 18377 31401 18411
rect 31435 18408 31447 18411
rect 31938 18408 31944 18420
rect 31435 18380 31944 18408
rect 31435 18377 31447 18380
rect 31389 18371 31447 18377
rect 31938 18368 31944 18380
rect 31996 18368 32002 18420
rect 32858 18368 32864 18420
rect 32916 18408 32922 18420
rect 34057 18411 34115 18417
rect 34057 18408 34069 18411
rect 32916 18380 34069 18408
rect 32916 18368 32922 18380
rect 34057 18377 34069 18380
rect 34103 18377 34115 18411
rect 34057 18371 34115 18377
rect 35986 18368 35992 18420
rect 36044 18368 36050 18420
rect 36078 18368 36084 18420
rect 36136 18368 36142 18420
rect 37918 18368 37924 18420
rect 37976 18368 37982 18420
rect 38470 18368 38476 18420
rect 38528 18368 38534 18420
rect 38930 18368 38936 18420
rect 38988 18368 38994 18420
rect 39022 18368 39028 18420
rect 39080 18408 39086 18420
rect 39301 18411 39359 18417
rect 39301 18408 39313 18411
rect 39080 18380 39313 18408
rect 39080 18368 39086 18380
rect 39301 18377 39313 18380
rect 39347 18377 39359 18411
rect 39301 18371 39359 18377
rect 39574 18368 39580 18420
rect 39632 18408 39638 18420
rect 40681 18411 40739 18417
rect 40681 18408 40693 18411
rect 39632 18380 40693 18408
rect 39632 18368 39638 18380
rect 40681 18377 40693 18380
rect 40727 18377 40739 18411
rect 40681 18371 40739 18377
rect 42245 18411 42303 18417
rect 42245 18377 42257 18411
rect 42291 18408 42303 18411
rect 42426 18408 42432 18420
rect 42291 18380 42432 18408
rect 42291 18377 42303 18380
rect 42245 18371 42303 18377
rect 29932 18312 31984 18340
rect 31956 18284 31984 18312
rect 32030 18300 32036 18352
rect 32088 18340 32094 18352
rect 34425 18343 34483 18349
rect 34425 18340 34437 18343
rect 32088 18312 33364 18340
rect 32088 18300 32094 18312
rect 29656 18244 31892 18272
rect 29549 18235 29607 18241
rect 27893 18207 27951 18213
rect 27893 18204 27905 18207
rect 27264 18176 27905 18204
rect 27893 18173 27905 18176
rect 27939 18173 27951 18207
rect 27893 18167 27951 18173
rect 27982 18164 27988 18216
rect 28040 18213 28046 18216
rect 28040 18207 28068 18213
rect 28056 18173 28068 18207
rect 28040 18167 28068 18173
rect 28040 18164 28046 18167
rect 28350 18164 28356 18216
rect 28408 18204 28414 18216
rect 29089 18207 29147 18213
rect 29089 18204 29101 18207
rect 28408 18176 29101 18204
rect 28408 18164 28414 18176
rect 29089 18173 29101 18176
rect 29135 18173 29147 18207
rect 29089 18167 29147 18173
rect 24029 18071 24087 18077
rect 24029 18068 24041 18071
rect 23440 18040 24041 18068
rect 23440 18028 23446 18040
rect 24029 18037 24041 18040
rect 24075 18037 24087 18071
rect 24029 18031 24087 18037
rect 26142 18028 26148 18080
rect 26200 18028 26206 18080
rect 27172 18068 27200 18164
rect 27614 18096 27620 18148
rect 27672 18096 27678 18148
rect 28994 18096 29000 18148
rect 29052 18136 29058 18148
rect 29564 18136 29592 18235
rect 31478 18164 31484 18216
rect 31536 18164 31542 18216
rect 31570 18164 31576 18216
rect 31628 18164 31634 18216
rect 29052 18108 29592 18136
rect 30929 18139 30987 18145
rect 29052 18096 29058 18108
rect 30929 18105 30941 18139
rect 30975 18136 30987 18139
rect 31386 18136 31392 18148
rect 30975 18108 31392 18136
rect 30975 18105 30987 18108
rect 30929 18099 30987 18105
rect 31386 18096 31392 18108
rect 31444 18096 31450 18148
rect 31496 18136 31524 18164
rect 31864 18136 31892 18244
rect 31938 18232 31944 18284
rect 31996 18232 32002 18284
rect 32122 18232 32128 18284
rect 32180 18232 32186 18284
rect 32392 18275 32450 18281
rect 32392 18241 32404 18275
rect 32438 18272 32450 18275
rect 33134 18272 33140 18284
rect 32438 18244 33140 18272
rect 32438 18241 32450 18244
rect 32392 18235 32450 18241
rect 33134 18232 33140 18244
rect 33192 18232 33198 18284
rect 33336 18204 33364 18312
rect 33428 18312 34437 18340
rect 33428 18284 33456 18312
rect 34425 18309 34437 18312
rect 34471 18309 34483 18343
rect 34425 18303 34483 18309
rect 33410 18232 33416 18284
rect 33468 18232 33474 18284
rect 33502 18232 33508 18284
rect 33560 18272 33566 18284
rect 33965 18275 34023 18281
rect 33965 18272 33977 18275
rect 33560 18244 33977 18272
rect 33560 18232 33566 18244
rect 33965 18241 33977 18244
rect 34011 18241 34023 18275
rect 36096 18272 36124 18368
rect 37274 18300 37280 18352
rect 37332 18340 37338 18352
rect 38948 18340 38976 18368
rect 37332 18312 38976 18340
rect 37332 18300 37338 18312
rect 36541 18275 36599 18281
rect 36541 18272 36553 18275
rect 33965 18235 34023 18241
rect 34072 18244 35112 18272
rect 36096 18244 36553 18272
rect 34072 18204 34100 18244
rect 33336 18176 34100 18204
rect 34241 18207 34299 18213
rect 34241 18173 34253 18207
rect 34287 18204 34299 18207
rect 34514 18204 34520 18216
rect 34287 18176 34520 18204
rect 34287 18173 34299 18176
rect 34241 18167 34299 18173
rect 34514 18164 34520 18176
rect 34572 18164 34578 18216
rect 34977 18207 35035 18213
rect 34977 18173 34989 18207
rect 35023 18173 35035 18207
rect 35084 18204 35112 18244
rect 36541 18241 36553 18244
rect 36587 18241 36599 18275
rect 36541 18235 36599 18241
rect 36722 18232 36728 18284
rect 36780 18272 36786 18284
rect 36909 18275 36967 18281
rect 36909 18272 36921 18275
rect 36780 18244 36921 18272
rect 36780 18232 36786 18244
rect 36909 18241 36921 18244
rect 36955 18241 36967 18275
rect 36909 18235 36967 18241
rect 37369 18275 37427 18281
rect 37369 18241 37381 18275
rect 37415 18272 37427 18275
rect 37550 18272 37556 18284
rect 37415 18244 37556 18272
rect 37415 18241 37427 18244
rect 37369 18235 37427 18241
rect 37550 18232 37556 18244
rect 37608 18232 37614 18284
rect 38838 18232 38844 18284
rect 38896 18272 38902 18284
rect 39025 18275 39083 18281
rect 39025 18272 39037 18275
rect 38896 18244 39037 18272
rect 38896 18232 38902 18244
rect 39025 18241 39037 18244
rect 39071 18241 39083 18275
rect 39025 18235 39083 18241
rect 39850 18232 39856 18284
rect 39908 18232 39914 18284
rect 40696 18272 40724 18371
rect 42426 18368 42432 18380
rect 42484 18368 42490 18420
rect 45002 18408 45008 18420
rect 43456 18380 45008 18408
rect 41132 18343 41190 18349
rect 41132 18309 41144 18343
rect 41178 18340 41190 18343
rect 41414 18340 41420 18352
rect 41178 18312 41420 18340
rect 41178 18309 41190 18312
rect 41132 18303 41190 18309
rect 41414 18300 41420 18312
rect 41472 18300 41478 18352
rect 42702 18300 42708 18352
rect 42760 18340 42766 18352
rect 42797 18343 42855 18349
rect 42797 18340 42809 18343
rect 42760 18312 42809 18340
rect 42760 18300 42766 18312
rect 42797 18309 42809 18312
rect 42843 18309 42855 18343
rect 42797 18303 42855 18309
rect 40862 18272 40868 18284
rect 40696 18244 40868 18272
rect 40862 18232 40868 18244
rect 40920 18232 40926 18284
rect 43456 18272 43484 18380
rect 45002 18368 45008 18380
rect 45060 18368 45066 18420
rect 45097 18411 45155 18417
rect 45097 18377 45109 18411
rect 45143 18408 45155 18411
rect 46290 18408 46296 18420
rect 45143 18380 46296 18408
rect 45143 18377 45155 18380
rect 45097 18371 45155 18377
rect 46290 18368 46296 18380
rect 46348 18368 46354 18420
rect 47762 18368 47768 18420
rect 47820 18368 47826 18420
rect 50062 18368 50068 18420
rect 50120 18408 50126 18420
rect 50157 18411 50215 18417
rect 50157 18408 50169 18411
rect 50120 18380 50169 18408
rect 50120 18368 50126 18380
rect 50157 18377 50169 18380
rect 50203 18377 50215 18411
rect 50157 18371 50215 18377
rect 51626 18368 51632 18420
rect 51684 18368 51690 18420
rect 52730 18368 52736 18420
rect 52788 18368 52794 18420
rect 53282 18368 53288 18420
rect 53340 18368 53346 18420
rect 53742 18368 53748 18420
rect 53800 18408 53806 18420
rect 54113 18411 54171 18417
rect 54113 18408 54125 18411
rect 53800 18380 54125 18408
rect 53800 18368 53806 18380
rect 54113 18377 54125 18380
rect 54159 18377 54171 18411
rect 54113 18371 54171 18377
rect 43530 18300 43536 18352
rect 43588 18340 43594 18352
rect 43962 18343 44020 18349
rect 43962 18340 43974 18343
rect 43588 18312 43974 18340
rect 43588 18300 43594 18312
rect 43962 18309 43974 18312
rect 44008 18309 44020 18343
rect 43962 18303 44020 18309
rect 45278 18300 45284 18352
rect 45336 18340 45342 18352
rect 45373 18343 45431 18349
rect 45373 18340 45385 18343
rect 45336 18312 45385 18340
rect 45336 18300 45342 18312
rect 45373 18309 45385 18312
rect 45419 18309 45431 18343
rect 45373 18303 45431 18309
rect 40972 18244 43484 18272
rect 40972 18204 41000 18244
rect 43622 18232 43628 18284
rect 43680 18272 43686 18284
rect 43717 18275 43775 18281
rect 43717 18272 43729 18275
rect 43680 18244 43729 18272
rect 43680 18232 43686 18244
rect 43717 18241 43729 18244
rect 43763 18241 43775 18275
rect 44818 18272 44824 18284
rect 43717 18235 43775 18241
rect 43824 18244 44824 18272
rect 35084 18176 41000 18204
rect 34977 18167 35035 18173
rect 32030 18136 32036 18148
rect 31496 18108 31754 18136
rect 31864 18108 32036 18136
rect 28166 18068 28172 18080
rect 27172 18040 28172 18068
rect 28166 18028 28172 18040
rect 28224 18028 28230 18080
rect 31726 18068 31754 18108
rect 32030 18096 32036 18108
rect 32088 18096 32094 18148
rect 33505 18139 33563 18145
rect 33505 18105 33517 18139
rect 33551 18136 33563 18139
rect 34992 18136 35020 18167
rect 42518 18164 42524 18216
rect 42576 18164 42582 18216
rect 42705 18207 42763 18213
rect 42705 18173 42717 18207
rect 42751 18204 42763 18207
rect 43824 18204 43852 18244
rect 44818 18232 44824 18244
rect 44876 18232 44882 18284
rect 53300 18281 53328 18368
rect 53285 18275 53343 18281
rect 53285 18241 53297 18275
rect 53331 18241 53343 18275
rect 53285 18235 53343 18241
rect 49881 18207 49939 18213
rect 49881 18204 49893 18207
rect 42751 18176 42840 18204
rect 42751 18173 42763 18176
rect 42705 18167 42763 18173
rect 42812 18148 42840 18176
rect 43088 18176 43852 18204
rect 49712 18176 49893 18204
rect 33551 18108 35020 18136
rect 33551 18105 33563 18108
rect 33505 18099 33563 18105
rect 35710 18096 35716 18148
rect 35768 18136 35774 18148
rect 39758 18136 39764 18148
rect 35768 18108 39764 18136
rect 35768 18096 35774 18108
rect 39758 18096 39764 18108
rect 39816 18096 39822 18148
rect 42794 18096 42800 18148
rect 42852 18096 42858 18148
rect 32766 18068 32772 18080
rect 31726 18040 32772 18068
rect 32766 18028 32772 18040
rect 32824 18028 32830 18080
rect 33594 18028 33600 18080
rect 33652 18028 33658 18080
rect 33686 18028 33692 18080
rect 33744 18068 33750 18080
rect 39942 18068 39948 18080
rect 33744 18040 39948 18068
rect 33744 18028 33750 18040
rect 39942 18028 39948 18040
rect 40000 18068 40006 18080
rect 40221 18071 40279 18077
rect 40221 18068 40233 18071
rect 40000 18040 40233 18068
rect 40000 18028 40006 18040
rect 40221 18037 40233 18040
rect 40267 18068 40279 18071
rect 43088 18068 43116 18176
rect 49712 18080 49740 18176
rect 49881 18173 49893 18176
rect 49927 18173 49939 18207
rect 49881 18167 49939 18173
rect 50065 18207 50123 18213
rect 50065 18173 50077 18207
rect 50111 18173 50123 18207
rect 50985 18207 51043 18213
rect 50985 18204 50997 18207
rect 50065 18167 50123 18173
rect 50540 18176 50997 18204
rect 40267 18040 43116 18068
rect 40267 18037 40279 18040
rect 40221 18031 40279 18037
rect 43162 18028 43168 18080
rect 43220 18028 43226 18080
rect 44082 18028 44088 18080
rect 44140 18068 44146 18080
rect 47302 18068 47308 18080
rect 44140 18040 47308 18068
rect 44140 18028 44146 18040
rect 47302 18028 47308 18040
rect 47360 18068 47366 18080
rect 47946 18068 47952 18080
rect 47360 18040 47952 18068
rect 47360 18028 47366 18040
rect 47946 18028 47952 18040
rect 48004 18068 48010 18080
rect 48133 18071 48191 18077
rect 48133 18068 48145 18071
rect 48004 18040 48145 18068
rect 48004 18028 48010 18040
rect 48133 18037 48145 18040
rect 48179 18068 48191 18071
rect 49602 18068 49608 18080
rect 48179 18040 49608 18068
rect 48179 18037 48191 18040
rect 48133 18031 48191 18037
rect 49602 18028 49608 18040
rect 49660 18028 49666 18080
rect 49694 18028 49700 18080
rect 49752 18028 49758 18080
rect 49878 18028 49884 18080
rect 49936 18068 49942 18080
rect 50080 18068 50108 18167
rect 50540 18145 50568 18176
rect 50985 18173 50997 18176
rect 51031 18173 51043 18207
rect 50985 18167 51043 18173
rect 52822 18164 52828 18216
rect 52880 18204 52886 18216
rect 53190 18204 53196 18216
rect 52880 18176 53196 18204
rect 52880 18164 52886 18176
rect 53190 18164 53196 18176
rect 53248 18204 53254 18216
rect 53469 18207 53527 18213
rect 53469 18204 53481 18207
rect 53248 18176 53481 18204
rect 53248 18164 53254 18176
rect 53469 18173 53481 18176
rect 53515 18173 53527 18207
rect 53469 18167 53527 18173
rect 58066 18164 58072 18216
rect 58124 18204 58130 18216
rect 58437 18207 58495 18213
rect 58437 18204 58449 18207
rect 58124 18176 58449 18204
rect 58124 18164 58130 18176
rect 58437 18173 58449 18176
rect 58483 18173 58495 18207
rect 58437 18167 58495 18173
rect 50525 18139 50583 18145
rect 50525 18105 50537 18139
rect 50571 18105 50583 18139
rect 50525 18099 50583 18105
rect 49936 18040 50108 18068
rect 52549 18071 52607 18077
rect 49936 18028 49942 18040
rect 52549 18037 52561 18071
rect 52595 18068 52607 18071
rect 52638 18068 52644 18080
rect 52595 18040 52644 18068
rect 52595 18037 52607 18040
rect 52549 18031 52607 18037
rect 52638 18028 52644 18040
rect 52696 18068 52702 18080
rect 53650 18068 53656 18080
rect 52696 18040 53656 18068
rect 52696 18028 52702 18040
rect 53650 18028 53656 18040
rect 53708 18028 53714 18080
rect 54478 18028 54484 18080
rect 54536 18028 54542 18080
rect 57882 18028 57888 18080
rect 57940 18028 57946 18080
rect 1104 17978 58880 18000
rect 1104 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 22616 17978
rect 22668 17926 22680 17978
rect 22732 17926 22744 17978
rect 22796 17926 22808 17978
rect 22860 17926 22872 17978
rect 22924 17926 37060 17978
rect 37112 17926 37124 17978
rect 37176 17926 37188 17978
rect 37240 17926 37252 17978
rect 37304 17926 37316 17978
rect 37368 17926 51504 17978
rect 51556 17926 51568 17978
rect 51620 17926 51632 17978
rect 51684 17926 51696 17978
rect 51748 17926 51760 17978
rect 51812 17926 58880 17978
rect 1104 17904 58880 17926
rect 6914 17824 6920 17876
rect 6972 17824 6978 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 11054 17864 11060 17876
rect 7975 17836 11060 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 7374 17796 7380 17808
rect 6880 17768 7380 17796
rect 6880 17756 6886 17768
rect 7374 17756 7380 17768
rect 7432 17796 7438 17808
rect 7944 17796 7972 17827
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11238 17824 11244 17876
rect 11296 17824 11302 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 13814 17864 13820 17876
rect 13495 17836 13820 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 16758 17824 16764 17876
rect 16816 17824 16822 17876
rect 19702 17824 19708 17876
rect 19760 17864 19766 17876
rect 20073 17867 20131 17873
rect 20073 17864 20085 17867
rect 19760 17836 20085 17864
rect 19760 17824 19766 17836
rect 20073 17833 20085 17836
rect 20119 17833 20131 17867
rect 20073 17827 20131 17833
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 22244 17836 22293 17864
rect 22244 17824 22250 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 22520 17836 22569 17864
rect 22520 17824 22526 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25314 17864 25320 17876
rect 24912 17836 25320 17864
rect 24912 17824 24918 17836
rect 25314 17824 25320 17836
rect 25372 17824 25378 17876
rect 25501 17867 25559 17873
rect 25501 17833 25513 17867
rect 25547 17864 25559 17867
rect 25590 17864 25596 17876
rect 25547 17836 25596 17864
rect 25547 17833 25559 17836
rect 25501 17827 25559 17833
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 27890 17864 27896 17876
rect 26988 17836 27896 17864
rect 7432 17768 7972 17796
rect 7432 17756 7438 17768
rect 10962 17756 10968 17808
rect 11020 17796 11026 17808
rect 16776 17796 16804 17824
rect 25332 17796 25360 17824
rect 26988 17796 27016 17836
rect 27890 17824 27896 17836
rect 27948 17864 27954 17876
rect 28074 17864 28080 17876
rect 27948 17836 28080 17864
rect 27948 17824 27954 17836
rect 28074 17824 28080 17836
rect 28132 17824 28138 17876
rect 28166 17824 28172 17876
rect 28224 17864 28230 17876
rect 28445 17867 28503 17873
rect 28445 17864 28457 17867
rect 28224 17836 28457 17864
rect 28224 17824 28230 17836
rect 28445 17833 28457 17836
rect 28491 17833 28503 17867
rect 28445 17827 28503 17833
rect 33134 17824 33140 17876
rect 33192 17864 33198 17876
rect 33321 17867 33379 17873
rect 33321 17864 33333 17867
rect 33192 17836 33333 17864
rect 33192 17824 33198 17836
rect 33321 17833 33333 17836
rect 33367 17833 33379 17867
rect 33321 17827 33379 17833
rect 33502 17824 33508 17876
rect 33560 17864 33566 17876
rect 33560 17836 34008 17864
rect 33560 17824 33566 17836
rect 11020 17768 12112 17796
rect 16776 17768 21588 17796
rect 25332 17768 27016 17796
rect 11020 17756 11026 17768
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17728 7619 17731
rect 7834 17728 7840 17740
rect 7607 17700 7840 17728
rect 7607 17697 7619 17700
rect 7561 17691 7619 17697
rect 7834 17688 7840 17700
rect 7892 17688 7898 17740
rect 9122 17688 9128 17740
rect 9180 17688 9186 17740
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17728 11207 17731
rect 11330 17728 11336 17740
rect 11195 17700 11336 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11330 17688 11336 17700
rect 11388 17728 11394 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11388 17700 11805 17728
rect 11388 17688 11394 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 11882 17688 11888 17740
rect 11940 17688 11946 17740
rect 12084 17737 12112 17768
rect 12069 17731 12127 17737
rect 12069 17697 12081 17731
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 13722 17688 13728 17740
rect 13780 17688 13786 17740
rect 20714 17688 20720 17740
rect 20772 17688 20778 17740
rect 3510 17620 3516 17672
rect 3568 17620 3574 17672
rect 3786 17620 3792 17672
rect 3844 17620 3850 17672
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 11900 17660 11928 17688
rect 11747 17632 11928 17660
rect 11992 17632 15240 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 9392 17595 9450 17601
rect 9392 17561 9404 17595
rect 9438 17592 9450 17595
rect 9582 17592 9588 17604
rect 9438 17564 9588 17592
rect 9438 17561 9450 17564
rect 9392 17555 9450 17561
rect 9582 17552 9588 17564
rect 9640 17552 9646 17604
rect 11992 17592 12020 17632
rect 9692 17564 12020 17592
rect 12336 17595 12394 17601
rect 2958 17484 2964 17536
rect 3016 17484 3022 17536
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 4304 17496 4445 17524
rect 4304 17484 4310 17496
rect 4433 17493 4445 17496
rect 4479 17493 4491 17527
rect 4433 17487 4491 17493
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 9692 17524 9720 17564
rect 12336 17561 12348 17595
rect 12382 17592 12394 17595
rect 12434 17592 12440 17604
rect 12382 17564 12440 17592
rect 12382 17561 12394 17564
rect 12336 17555 12394 17561
rect 12434 17552 12440 17564
rect 12492 17552 12498 17604
rect 15212 17592 15240 17632
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15344 17632 15669 17660
rect 15344 17620 15350 17632
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 15930 17620 15936 17672
rect 15988 17620 15994 17672
rect 16206 17620 16212 17672
rect 16264 17620 16270 17672
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 16224 17592 16252 17620
rect 15212 17564 16252 17592
rect 8444 17496 9720 17524
rect 8444 17484 8450 17496
rect 10502 17484 10508 17536
rect 10560 17484 10566 17536
rect 11609 17527 11667 17533
rect 11609 17493 11621 17527
rect 11655 17524 11667 17527
rect 12158 17524 12164 17536
rect 11655 17496 12164 17524
rect 11655 17493 11667 17496
rect 11609 17487 11667 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 15102 17484 15108 17536
rect 15160 17484 15166 17536
rect 16485 17527 16543 17533
rect 16485 17493 16497 17527
rect 16531 17524 16543 17527
rect 17218 17524 17224 17536
rect 16531 17496 17224 17524
rect 16531 17493 16543 17496
rect 16485 17487 16543 17493
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17589 17527 17647 17533
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 17770 17524 17776 17536
rect 17635 17496 17776 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 18046 17484 18052 17536
rect 18104 17524 18110 17536
rect 18141 17527 18199 17533
rect 18141 17524 18153 17527
rect 18104 17496 18153 17524
rect 18104 17484 18110 17496
rect 18141 17493 18153 17496
rect 18187 17493 18199 17527
rect 18141 17487 18199 17493
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 20990 17524 20996 17536
rect 20772 17496 20996 17524
rect 20772 17484 20778 17496
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21560 17533 21588 17768
rect 21729 17731 21787 17737
rect 21729 17697 21741 17731
rect 21775 17728 21787 17731
rect 21818 17728 21824 17740
rect 21775 17700 21824 17728
rect 21775 17697 21787 17700
rect 21729 17691 21787 17697
rect 21818 17688 21824 17700
rect 21876 17688 21882 17740
rect 26988 17737 27016 17768
rect 28353 17799 28411 17805
rect 28353 17765 28365 17799
rect 28399 17796 28411 17799
rect 33229 17799 33287 17805
rect 28399 17768 29040 17796
rect 28399 17765 28411 17768
rect 28353 17759 28411 17765
rect 29012 17737 29040 17768
rect 33229 17765 33241 17799
rect 33275 17796 33287 17799
rect 33980 17796 34008 17836
rect 34514 17824 34520 17876
rect 34572 17864 34578 17876
rect 35710 17864 35716 17876
rect 34572 17836 35716 17864
rect 34572 17824 34578 17836
rect 35710 17824 35716 17836
rect 35768 17824 35774 17876
rect 40862 17824 40868 17876
rect 40920 17864 40926 17876
rect 41141 17867 41199 17873
rect 41141 17864 41153 17867
rect 40920 17836 41153 17864
rect 40920 17824 40926 17836
rect 41141 17833 41153 17836
rect 41187 17833 41199 17867
rect 41141 17827 41199 17833
rect 33275 17768 33916 17796
rect 33980 17768 38148 17796
rect 33275 17765 33287 17768
rect 33229 17759 33287 17765
rect 26145 17731 26203 17737
rect 26145 17697 26157 17731
rect 26191 17697 26203 17731
rect 26145 17691 26203 17697
rect 26973 17731 27031 17737
rect 26973 17697 26985 17731
rect 27019 17697 27031 17731
rect 26973 17691 27031 17697
rect 28997 17731 29055 17737
rect 28997 17697 29009 17731
rect 29043 17697 29055 17731
rect 28997 17691 29055 17697
rect 24946 17620 24952 17672
rect 25004 17620 25010 17672
rect 26050 17620 26056 17672
rect 26108 17660 26114 17672
rect 26160 17660 26188 17691
rect 32674 17688 32680 17740
rect 32732 17688 32738 17740
rect 32769 17731 32827 17737
rect 32769 17697 32781 17731
rect 32815 17728 32827 17731
rect 33410 17728 33416 17740
rect 32815 17700 33416 17728
rect 32815 17697 32827 17700
rect 32769 17691 32827 17697
rect 33410 17688 33416 17700
rect 33468 17688 33474 17740
rect 33888 17737 33916 17768
rect 38120 17740 38148 17768
rect 33873 17731 33931 17737
rect 33873 17697 33885 17731
rect 33919 17697 33931 17731
rect 34238 17728 34244 17740
rect 33873 17691 33931 17697
rect 33980 17700 34244 17728
rect 26108 17632 26188 17660
rect 27240 17663 27298 17669
rect 26108 17620 26114 17632
rect 27240 17629 27252 17663
rect 27286 17660 27298 17663
rect 27522 17660 27528 17672
rect 27286 17632 27528 17660
rect 27286 17629 27298 17632
rect 27240 17623 27298 17629
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 31938 17620 31944 17672
rect 31996 17660 32002 17672
rect 33980 17660 34008 17700
rect 34238 17688 34244 17700
rect 34296 17728 34302 17740
rect 34296 17700 36492 17728
rect 34296 17688 34302 17700
rect 31996 17632 34008 17660
rect 31996 17620 32002 17632
rect 36078 17620 36084 17672
rect 36136 17660 36142 17672
rect 36357 17663 36415 17669
rect 36357 17660 36369 17663
rect 36136 17632 36369 17660
rect 36136 17620 36142 17632
rect 36357 17629 36369 17632
rect 36403 17629 36415 17663
rect 36464 17660 36492 17700
rect 38102 17688 38108 17740
rect 38160 17688 38166 17740
rect 41156 17728 41184 17827
rect 53650 17824 53656 17876
rect 53708 17864 53714 17876
rect 57054 17864 57060 17876
rect 53708 17836 57060 17864
rect 53708 17824 53714 17836
rect 57054 17824 57060 17836
rect 57112 17824 57118 17876
rect 42705 17799 42763 17805
rect 42705 17765 42717 17799
rect 42751 17796 42763 17799
rect 43806 17796 43812 17808
rect 42751 17768 43812 17796
rect 42751 17765 42763 17768
rect 42705 17759 42763 17765
rect 43806 17756 43812 17768
rect 43864 17756 43870 17808
rect 53466 17756 53472 17808
rect 53524 17796 53530 17808
rect 53837 17799 53895 17805
rect 53837 17796 53849 17799
rect 53524 17768 53849 17796
rect 53524 17756 53530 17768
rect 53837 17765 53849 17768
rect 53883 17765 53895 17799
rect 53837 17759 53895 17765
rect 41325 17731 41383 17737
rect 41325 17728 41337 17731
rect 41156 17700 41337 17728
rect 41325 17697 41337 17700
rect 41371 17697 41383 17731
rect 41325 17691 41383 17697
rect 43162 17688 43168 17740
rect 43220 17728 43226 17740
rect 43349 17731 43407 17737
rect 43349 17728 43361 17731
rect 43220 17700 43361 17728
rect 43220 17688 43226 17700
rect 43349 17697 43361 17700
rect 43395 17697 43407 17731
rect 43349 17691 43407 17697
rect 44174 17688 44180 17740
rect 44232 17728 44238 17740
rect 44453 17731 44511 17737
rect 44453 17728 44465 17731
rect 44232 17700 44465 17728
rect 44232 17688 44238 17700
rect 44453 17697 44465 17700
rect 44499 17697 44511 17731
rect 44453 17691 44511 17697
rect 44545 17731 44603 17737
rect 44545 17697 44557 17731
rect 44591 17697 44603 17731
rect 44545 17691 44603 17697
rect 43809 17663 43867 17669
rect 43809 17660 43821 17663
rect 36464 17632 43821 17660
rect 36357 17623 36415 17629
rect 43809 17629 43821 17632
rect 43855 17660 43867 17663
rect 44560 17660 44588 17691
rect 54570 17688 54576 17740
rect 54628 17728 54634 17740
rect 56873 17731 56931 17737
rect 56873 17728 56885 17731
rect 54628 17700 56885 17728
rect 54628 17688 54634 17700
rect 56873 17697 56885 17700
rect 56919 17697 56931 17731
rect 56873 17691 56931 17697
rect 43855 17632 44588 17660
rect 43855 17629 43867 17632
rect 43809 17623 43867 17629
rect 44726 17620 44732 17672
rect 44784 17620 44790 17672
rect 53006 17620 53012 17672
rect 53064 17620 53070 17672
rect 53098 17620 53104 17672
rect 53156 17620 53162 17672
rect 53834 17620 53840 17672
rect 53892 17660 53898 17672
rect 54389 17663 54447 17669
rect 54389 17660 54401 17663
rect 53892 17632 54401 17660
rect 53892 17620 53898 17632
rect 54389 17629 54401 17632
rect 54435 17629 54447 17663
rect 54389 17623 54447 17629
rect 55858 17620 55864 17672
rect 55916 17620 55922 17672
rect 56042 17620 56048 17672
rect 56100 17620 56106 17672
rect 26789 17595 26847 17601
rect 26789 17592 26801 17595
rect 24596 17564 26801 17592
rect 24596 17536 24624 17564
rect 26789 17561 26801 17564
rect 26835 17592 26847 17595
rect 27890 17592 27896 17604
rect 26835 17564 27896 17592
rect 26835 17561 26847 17564
rect 26789 17555 26847 17561
rect 27890 17552 27896 17564
rect 27948 17552 27954 17604
rect 30009 17595 30067 17601
rect 30009 17561 30021 17595
rect 30055 17561 30067 17595
rect 30009 17555 30067 17561
rect 31757 17595 31815 17601
rect 31757 17561 31769 17595
rect 31803 17592 31815 17595
rect 32033 17595 32091 17601
rect 32033 17592 32045 17595
rect 31803 17564 32045 17592
rect 31803 17561 31815 17564
rect 31757 17555 31815 17561
rect 32033 17561 32045 17564
rect 32079 17592 32091 17595
rect 37826 17592 37832 17604
rect 32079 17564 37832 17592
rect 32079 17561 32091 17564
rect 32033 17555 32091 17561
rect 21545 17527 21603 17533
rect 21545 17493 21557 17527
rect 21591 17524 21603 17527
rect 21726 17524 21732 17536
rect 21591 17496 21732 17524
rect 21591 17493 21603 17496
rect 21545 17487 21603 17493
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 24394 17484 24400 17536
rect 24452 17484 24458 17536
rect 24578 17484 24584 17536
rect 24636 17484 24642 17536
rect 25866 17484 25872 17536
rect 25924 17484 25930 17536
rect 25961 17527 26019 17533
rect 25961 17493 25973 17527
rect 26007 17524 26019 17527
rect 26418 17524 26424 17536
rect 26007 17496 26424 17524
rect 26007 17493 26019 17496
rect 25961 17487 26019 17493
rect 26418 17484 26424 17496
rect 26476 17484 26482 17536
rect 28994 17484 29000 17536
rect 29052 17524 29058 17536
rect 30024 17524 30052 17555
rect 37826 17552 37832 17564
rect 37884 17592 37890 17604
rect 41138 17592 41144 17604
rect 37884 17564 41144 17592
rect 37884 17552 37890 17564
rect 41138 17552 41144 17564
rect 41196 17552 41202 17604
rect 41592 17595 41650 17601
rect 41592 17561 41604 17595
rect 41638 17592 41650 17595
rect 42797 17595 42855 17601
rect 42797 17592 42809 17595
rect 41638 17564 42809 17592
rect 41638 17561 41650 17564
rect 41592 17555 41650 17561
rect 42797 17561 42809 17564
rect 42843 17561 42855 17595
rect 42797 17555 42855 17561
rect 44361 17595 44419 17601
rect 44361 17561 44373 17595
rect 44407 17592 44419 17595
rect 44744 17592 44772 17620
rect 44407 17564 44772 17592
rect 57140 17595 57198 17601
rect 44407 17561 44419 17564
rect 44361 17555 44419 17561
rect 57140 17561 57152 17595
rect 57186 17592 57198 17595
rect 57514 17592 57520 17604
rect 57186 17564 57520 17592
rect 57186 17561 57198 17564
rect 57140 17555 57198 17561
rect 57514 17552 57520 17564
rect 57572 17552 57578 17604
rect 30374 17524 30380 17536
rect 29052 17496 30380 17524
rect 29052 17484 29058 17496
rect 30374 17484 30380 17496
rect 30432 17484 30438 17536
rect 32766 17484 32772 17536
rect 32824 17524 32830 17536
rect 32861 17527 32919 17533
rect 32861 17524 32873 17527
rect 32824 17496 32873 17524
rect 32824 17484 32830 17496
rect 32861 17493 32873 17496
rect 32907 17493 32919 17527
rect 32861 17487 32919 17493
rect 35802 17484 35808 17536
rect 35860 17484 35866 17536
rect 37458 17484 37464 17536
rect 37516 17484 37522 17536
rect 43990 17484 43996 17536
rect 44048 17484 44054 17536
rect 52178 17484 52184 17536
rect 52236 17484 52242 17536
rect 52362 17484 52368 17536
rect 52420 17484 52426 17536
rect 53650 17484 53656 17536
rect 53708 17524 53714 17536
rect 53745 17527 53803 17533
rect 53745 17524 53757 17527
rect 53708 17496 53757 17524
rect 53708 17484 53714 17496
rect 53745 17493 53757 17496
rect 53791 17493 53803 17527
rect 53745 17487 53803 17493
rect 55306 17484 55312 17536
rect 55364 17484 55370 17536
rect 56594 17484 56600 17536
rect 56652 17524 56658 17536
rect 56689 17527 56747 17533
rect 56689 17524 56701 17527
rect 56652 17496 56701 17524
rect 56652 17484 56658 17496
rect 56689 17493 56701 17496
rect 56735 17493 56747 17527
rect 56689 17487 56747 17493
rect 58250 17484 58256 17536
rect 58308 17484 58314 17536
rect 1104 17434 59040 17456
rect 1104 17382 15394 17434
rect 15446 17382 15458 17434
rect 15510 17382 15522 17434
rect 15574 17382 15586 17434
rect 15638 17382 15650 17434
rect 15702 17382 29838 17434
rect 29890 17382 29902 17434
rect 29954 17382 29966 17434
rect 30018 17382 30030 17434
rect 30082 17382 30094 17434
rect 30146 17382 44282 17434
rect 44334 17382 44346 17434
rect 44398 17382 44410 17434
rect 44462 17382 44474 17434
rect 44526 17382 44538 17434
rect 44590 17382 58726 17434
rect 58778 17382 58790 17434
rect 58842 17382 58854 17434
rect 58906 17382 58918 17434
rect 58970 17382 58982 17434
rect 59034 17382 59040 17434
rect 1104 17360 59040 17382
rect 2958 17280 2964 17332
rect 3016 17280 3022 17332
rect 3786 17280 3792 17332
rect 3844 17280 3850 17332
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 9858 17320 9864 17332
rect 9732 17292 9864 17320
rect 9732 17280 9738 17292
rect 9858 17280 9864 17292
rect 9916 17320 9922 17332
rect 10318 17320 10324 17332
rect 9916 17292 10324 17320
rect 9916 17280 9922 17292
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 11790 17280 11796 17332
rect 11848 17280 11854 17332
rect 12434 17280 12440 17332
rect 12492 17280 12498 17332
rect 15286 17280 15292 17332
rect 15344 17280 15350 17332
rect 16669 17323 16727 17329
rect 16669 17289 16681 17323
rect 16715 17320 16727 17323
rect 16942 17320 16948 17332
rect 16715 17292 16948 17320
rect 16715 17289 16727 17292
rect 16669 17283 16727 17289
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 19392 17292 19809 17320
rect 19392 17280 19398 17292
rect 19797 17289 19809 17292
rect 19843 17320 19855 17323
rect 20530 17320 20536 17332
rect 19843 17292 20536 17320
rect 19843 17289 19855 17292
rect 19797 17283 19855 17289
rect 20530 17280 20536 17292
rect 20588 17280 20594 17332
rect 22370 17280 22376 17332
rect 22428 17320 22434 17332
rect 22741 17323 22799 17329
rect 22741 17320 22753 17323
rect 22428 17292 22753 17320
rect 22428 17280 22434 17292
rect 22741 17289 22753 17292
rect 22787 17289 22799 17323
rect 22741 17283 22799 17289
rect 24394 17280 24400 17332
rect 24452 17280 24458 17332
rect 25866 17280 25872 17332
rect 25924 17320 25930 17332
rect 26697 17323 26755 17329
rect 26697 17320 26709 17323
rect 25924 17292 26709 17320
rect 25924 17280 25930 17292
rect 26697 17289 26709 17292
rect 26743 17320 26755 17323
rect 27982 17320 27988 17332
rect 26743 17292 27988 17320
rect 26743 17289 26755 17292
rect 26697 17283 26755 17289
rect 27982 17280 27988 17292
rect 28040 17280 28046 17332
rect 30929 17323 30987 17329
rect 30929 17289 30941 17323
rect 30975 17320 30987 17323
rect 31570 17320 31576 17332
rect 30975 17292 31576 17320
rect 30975 17289 30987 17292
rect 30929 17283 30987 17289
rect 31570 17280 31576 17292
rect 31628 17280 31634 17332
rect 31754 17280 31760 17332
rect 31812 17320 31818 17332
rect 31849 17323 31907 17329
rect 31849 17320 31861 17323
rect 31812 17292 31861 17320
rect 31812 17280 31818 17292
rect 31849 17289 31861 17292
rect 31895 17289 31907 17323
rect 31849 17283 31907 17289
rect 32674 17280 32680 17332
rect 32732 17320 32738 17332
rect 33413 17323 33471 17329
rect 33413 17320 33425 17323
rect 32732 17292 33425 17320
rect 32732 17280 32738 17292
rect 33413 17289 33425 17292
rect 33459 17320 33471 17323
rect 33502 17320 33508 17332
rect 33459 17292 33508 17320
rect 33459 17289 33471 17292
rect 33413 17283 33471 17289
rect 33502 17280 33508 17292
rect 33560 17280 33566 17332
rect 35253 17323 35311 17329
rect 35253 17289 35265 17323
rect 35299 17320 35311 17323
rect 35802 17320 35808 17332
rect 35299 17292 35808 17320
rect 35299 17289 35311 17292
rect 35253 17283 35311 17289
rect 35802 17280 35808 17292
rect 35860 17280 35866 17332
rect 42794 17280 42800 17332
rect 42852 17280 42858 17332
rect 52362 17280 52368 17332
rect 52420 17280 52426 17332
rect 52549 17323 52607 17329
rect 52549 17289 52561 17323
rect 52595 17320 52607 17323
rect 53098 17320 53104 17332
rect 52595 17292 53104 17320
rect 52595 17289 52607 17292
rect 52549 17283 52607 17289
rect 53098 17280 53104 17292
rect 53156 17280 53162 17332
rect 53466 17280 53472 17332
rect 53524 17280 53530 17332
rect 55306 17280 55312 17332
rect 55364 17280 55370 17332
rect 55953 17323 56011 17329
rect 55953 17289 55965 17323
rect 55999 17320 56011 17323
rect 56042 17320 56048 17332
rect 55999 17292 56048 17320
rect 55999 17289 56011 17292
rect 55953 17283 56011 17289
rect 56042 17280 56048 17292
rect 56100 17280 56106 17332
rect 57422 17320 57428 17332
rect 56704 17292 57428 17320
rect 2676 17255 2734 17261
rect 2676 17221 2688 17255
rect 2722 17252 2734 17255
rect 2976 17252 3004 17280
rect 2722 17224 3004 17252
rect 2722 17221 2734 17224
rect 2676 17215 2734 17221
rect 8386 17212 8392 17264
rect 8444 17212 8450 17264
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 6914 17193 6920 17196
rect 6641 17187 6699 17193
rect 6641 17184 6653 17187
rect 6512 17156 6653 17184
rect 6512 17144 6518 17156
rect 6641 17153 6653 17156
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 6908 17147 6920 17193
rect 6914 17144 6920 17147
rect 6972 17144 6978 17196
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 8036 17156 8125 17184
rect 1578 17076 1584 17128
rect 1636 17116 1642 17128
rect 2406 17116 2412 17128
rect 1636 17088 2412 17116
rect 1636 17076 1642 17088
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 3878 17076 3884 17128
rect 3936 17076 3942 17128
rect 8036 17057 8064 17156
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10520 17184 10548 17280
rect 11241 17255 11299 17261
rect 11241 17221 11253 17255
rect 11287 17252 11299 17255
rect 12526 17252 12532 17264
rect 11287 17224 12532 17252
rect 11287 17221 11299 17224
rect 11241 17215 11299 17221
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10183 17156 10456 17184
rect 10520 17156 10609 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 10318 17076 10324 17128
rect 10376 17076 10382 17128
rect 10428 17116 10456 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 11256 17116 11284 17215
rect 12526 17212 12532 17224
rect 12584 17212 12590 17264
rect 15657 17255 15715 17261
rect 15657 17221 15669 17255
rect 15703 17252 15715 17255
rect 15838 17252 15844 17264
rect 15703 17224 15844 17252
rect 15703 17221 15715 17224
rect 15657 17215 15715 17221
rect 15838 17212 15844 17224
rect 15896 17212 15902 17264
rect 20548 17252 20576 17280
rect 23652 17255 23710 17261
rect 20548 17224 23612 17252
rect 12986 17144 12992 17196
rect 13044 17144 13050 17196
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 17218 17184 17224 17196
rect 15795 17156 17224 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 17793 17187 17851 17193
rect 17793 17153 17805 17187
rect 17839 17184 17851 17187
rect 19242 17184 19248 17196
rect 17839 17156 19248 17184
rect 17839 17153 17851 17156
rect 17793 17147 17851 17153
rect 19242 17144 19248 17156
rect 19300 17144 19306 17196
rect 23382 17144 23388 17196
rect 23440 17144 23446 17196
rect 23584 17184 23612 17224
rect 23652 17221 23664 17255
rect 23698 17252 23710 17255
rect 24412 17252 24440 17280
rect 23698 17224 24440 17252
rect 23698 17221 23710 17224
rect 23652 17215 23710 17221
rect 28074 17212 28080 17264
rect 28132 17252 28138 17264
rect 28994 17252 29000 17264
rect 28132 17224 29000 17252
rect 28132 17212 28138 17224
rect 28994 17212 29000 17224
rect 29052 17212 29058 17264
rect 39485 17255 39543 17261
rect 39485 17252 39497 17255
rect 31588 17224 39497 17252
rect 25777 17187 25835 17193
rect 25777 17184 25789 17187
rect 23584 17156 25789 17184
rect 25777 17153 25789 17156
rect 25823 17184 25835 17187
rect 26050 17184 26056 17196
rect 25823 17156 26056 17184
rect 25823 17153 25835 17156
rect 25777 17147 25835 17153
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 26142 17144 26148 17196
rect 26200 17144 26206 17196
rect 10428 17088 11284 17116
rect 15010 17076 15016 17128
rect 15068 17116 15074 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15068 17088 15853 17116
rect 15068 17076 15074 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 18046 17076 18052 17128
rect 18104 17076 18110 17128
rect 18874 17076 18880 17128
rect 18932 17076 18938 17128
rect 20898 17076 20904 17128
rect 20956 17076 20962 17128
rect 22370 17076 22376 17128
rect 22428 17076 22434 17128
rect 25409 17119 25467 17125
rect 25409 17116 25421 17119
rect 25056 17088 25421 17116
rect 8021 17051 8079 17057
rect 8021 17017 8033 17051
rect 8067 17017 8079 17051
rect 10244 17048 10272 17076
rect 12158 17048 12164 17060
rect 10244 17020 12164 17048
rect 8021 17011 8079 17017
rect 12158 17008 12164 17020
rect 12216 17008 12222 17060
rect 16298 17048 16304 17060
rect 12728 17020 16304 17048
rect 12728 16992 12756 17020
rect 16298 17008 16304 17020
rect 16356 17008 16362 17060
rect 21082 17048 21088 17060
rect 18248 17020 21088 17048
rect 4522 16940 4528 16992
rect 4580 16940 4586 16992
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 12710 16980 12716 16992
rect 11848 16952 12716 16980
rect 11848 16940 11854 16952
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 14829 16983 14887 16989
rect 14829 16949 14841 16983
rect 14875 16980 14887 16983
rect 15010 16980 15016 16992
rect 14875 16952 15016 16980
rect 14875 16949 14887 16952
rect 14829 16943 14887 16949
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15194 16940 15200 16992
rect 15252 16940 15258 16992
rect 16316 16980 16344 17008
rect 18248 16980 18276 17020
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 21637 17051 21695 17057
rect 21637 17017 21649 17051
rect 21683 17048 21695 17051
rect 21726 17048 21732 17060
rect 21683 17020 21732 17048
rect 21683 17017 21695 17020
rect 21637 17011 21695 17017
rect 21726 17008 21732 17020
rect 21784 17048 21790 17060
rect 24765 17051 24823 17057
rect 21784 17020 21956 17048
rect 21784 17008 21790 17020
rect 16316 16952 18276 16980
rect 18322 16940 18328 16992
rect 18380 16940 18386 16992
rect 20346 16940 20352 16992
rect 20404 16940 20410 16992
rect 21818 16940 21824 16992
rect 21876 16940 21882 16992
rect 21928 16980 21956 17020
rect 24765 17017 24777 17051
rect 24811 17048 24823 17051
rect 25056 17048 25084 17088
rect 25409 17085 25421 17088
rect 25455 17085 25467 17119
rect 25409 17079 25467 17085
rect 27614 17076 27620 17128
rect 27672 17116 27678 17128
rect 27801 17119 27859 17125
rect 27801 17116 27813 17119
rect 27672 17088 27813 17116
rect 27672 17076 27678 17088
rect 27801 17085 27813 17088
rect 27847 17085 27859 17119
rect 27801 17079 27859 17085
rect 28166 17076 28172 17128
rect 28224 17116 28230 17128
rect 28629 17119 28687 17125
rect 28629 17116 28641 17119
rect 28224 17088 28641 17116
rect 28224 17076 28230 17088
rect 28629 17085 28641 17088
rect 28675 17085 28687 17119
rect 28629 17079 28687 17085
rect 24811 17020 25084 17048
rect 24811 17017 24823 17020
rect 24765 17011 24823 17017
rect 25056 16992 25084 17020
rect 27890 17008 27896 17060
rect 27948 17048 27954 17060
rect 31588 17048 31616 17224
rect 39485 17221 39497 17224
rect 39531 17252 39543 17255
rect 39531 17224 39804 17252
rect 39531 17221 39543 17224
rect 39485 17215 39543 17221
rect 31662 17144 31668 17196
rect 31720 17184 31726 17196
rect 31720 17156 32435 17184
rect 31720 17144 31726 17156
rect 31938 17076 31944 17128
rect 31996 17116 32002 17128
rect 32309 17119 32367 17125
rect 32309 17116 32321 17119
rect 31996 17088 32321 17116
rect 31996 17076 32002 17088
rect 32309 17085 32321 17088
rect 32355 17085 32367 17119
rect 32407 17116 32435 17156
rect 33778 17144 33784 17196
rect 33836 17184 33842 17196
rect 34057 17187 34115 17193
rect 34057 17184 34069 17187
rect 33836 17156 34069 17184
rect 33836 17144 33842 17156
rect 34057 17153 34069 17156
rect 34103 17153 34115 17187
rect 34057 17147 34115 17153
rect 35250 17144 35256 17196
rect 35308 17184 35314 17196
rect 39776 17193 39804 17224
rect 44082 17212 44088 17264
rect 44140 17252 44146 17264
rect 51436 17255 51494 17261
rect 44140 17224 51396 17252
rect 44140 17212 44146 17224
rect 35345 17187 35403 17193
rect 35345 17184 35357 17187
rect 35308 17156 35357 17184
rect 35308 17144 35314 17156
rect 35345 17153 35357 17156
rect 35391 17153 35403 17187
rect 39761 17187 39819 17193
rect 35345 17147 35403 17153
rect 35636 17156 39712 17184
rect 34885 17119 34943 17125
rect 34885 17116 34897 17119
rect 32407 17088 34897 17116
rect 32309 17079 32367 17085
rect 34885 17085 34897 17088
rect 34931 17116 34943 17119
rect 35161 17119 35219 17125
rect 35161 17116 35173 17119
rect 34931 17088 35173 17116
rect 34931 17085 34943 17088
rect 34885 17079 34943 17085
rect 35161 17085 35173 17088
rect 35207 17116 35219 17119
rect 35636 17116 35664 17156
rect 36357 17119 36415 17125
rect 36357 17116 36369 17119
rect 35207 17088 35664 17116
rect 35728 17088 36369 17116
rect 35207 17085 35219 17088
rect 35161 17079 35219 17085
rect 35728 17057 35756 17088
rect 36357 17085 36369 17088
rect 36403 17085 36415 17119
rect 36357 17079 36415 17085
rect 37918 17076 37924 17128
rect 37976 17076 37982 17128
rect 38654 17076 38660 17128
rect 38712 17076 38718 17128
rect 27948 17020 31616 17048
rect 35713 17051 35771 17057
rect 27948 17008 27954 17020
rect 35713 17017 35725 17051
rect 35759 17017 35771 17051
rect 37458 17048 37464 17060
rect 35713 17011 35771 17017
rect 36740 17020 37464 17048
rect 22186 16980 22192 16992
rect 21928 16952 22192 16980
rect 22186 16940 22192 16952
rect 22244 16980 22250 16992
rect 24394 16980 24400 16992
rect 22244 16952 24400 16980
rect 22244 16940 22250 16952
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 24854 16940 24860 16992
rect 24912 16940 24918 16992
rect 25038 16940 25044 16992
rect 25096 16940 25102 16992
rect 27246 16940 27252 16992
rect 27304 16940 27310 16992
rect 27706 16940 27712 16992
rect 27764 16980 27770 16992
rect 28077 16983 28135 16989
rect 28077 16980 28089 16983
rect 27764 16952 28089 16980
rect 27764 16940 27770 16952
rect 28077 16949 28089 16952
rect 28123 16949 28135 16983
rect 28077 16943 28135 16949
rect 32950 16940 32956 16992
rect 33008 16940 33014 16992
rect 33778 16940 33784 16992
rect 33836 16980 33842 16992
rect 34514 16980 34520 16992
rect 33836 16952 34520 16980
rect 33836 16940 33842 16952
rect 34514 16940 34520 16952
rect 34572 16940 34578 16992
rect 35802 16940 35808 16992
rect 35860 16940 35866 16992
rect 36170 16940 36176 16992
rect 36228 16980 36234 16992
rect 36740 16989 36768 17020
rect 37458 17008 37464 17020
rect 37516 17008 37522 17060
rect 39684 17048 39712 17156
rect 39761 17153 39773 17187
rect 39807 17153 39819 17187
rect 39761 17147 39819 17153
rect 43441 17187 43499 17193
rect 43441 17153 43453 17187
rect 43487 17184 43499 17187
rect 43806 17184 43812 17196
rect 43487 17156 43812 17184
rect 43487 17153 43499 17156
rect 43441 17147 43499 17153
rect 43806 17144 43812 17156
rect 43864 17144 43870 17196
rect 48130 17144 48136 17196
rect 48188 17144 48194 17196
rect 48400 17187 48458 17193
rect 48400 17153 48412 17187
rect 48446 17184 48458 17187
rect 50341 17187 50399 17193
rect 50341 17184 50353 17187
rect 48446 17156 50353 17184
rect 48446 17153 48458 17156
rect 48400 17147 48458 17153
rect 50341 17153 50353 17156
rect 50387 17153 50399 17187
rect 50341 17147 50399 17153
rect 51166 17144 51172 17196
rect 51224 17144 51230 17196
rect 51368 17184 51396 17224
rect 51436 17221 51448 17255
rect 51482 17252 51494 17255
rect 52380 17252 52408 17280
rect 51482 17224 52408 17252
rect 51482 17221 51494 17224
rect 51436 17215 51494 17221
rect 52638 17212 52644 17264
rect 52696 17212 52702 17264
rect 52656 17184 52684 17212
rect 51368 17156 52684 17184
rect 53101 17187 53159 17193
rect 53101 17153 53113 17187
rect 53147 17184 53159 17187
rect 53484 17184 53512 17280
rect 54840 17255 54898 17261
rect 54840 17221 54852 17255
rect 54886 17252 54898 17255
rect 55324 17252 55352 17280
rect 54886 17224 55352 17252
rect 54886 17221 54898 17224
rect 54840 17215 54898 17221
rect 53147 17156 53512 17184
rect 53147 17153 53159 17156
rect 53101 17147 53159 17153
rect 54570 17144 54576 17196
rect 54628 17144 54634 17196
rect 40034 17076 40040 17128
rect 40092 17076 40098 17128
rect 40218 17076 40224 17128
rect 40276 17116 40282 17128
rect 41233 17119 41291 17125
rect 41233 17116 41245 17119
rect 40276 17088 41245 17116
rect 40276 17076 40282 17088
rect 41233 17085 41245 17088
rect 41279 17085 41291 17119
rect 41233 17079 41291 17085
rect 44174 17076 44180 17128
rect 44232 17076 44238 17128
rect 49605 17119 49663 17125
rect 49605 17116 49617 17119
rect 49528 17088 49617 17116
rect 40310 17048 40316 17060
rect 39684 17020 40316 17048
rect 40310 17008 40316 17020
rect 40368 17008 40374 17060
rect 49528 17057 49556 17088
rect 49605 17085 49617 17088
rect 49651 17085 49663 17119
rect 49605 17079 49663 17085
rect 50890 17076 50896 17128
rect 50948 17076 50954 17128
rect 52178 17076 52184 17128
rect 52236 17116 52242 17128
rect 52825 17119 52883 17125
rect 52825 17116 52837 17119
rect 52236 17088 52837 17116
rect 52236 17076 52242 17088
rect 52825 17085 52837 17088
rect 52871 17085 52883 17119
rect 52825 17079 52883 17085
rect 52914 17076 52920 17128
rect 52972 17116 52978 17128
rect 56704 17125 56732 17292
rect 57422 17280 57428 17292
rect 57480 17320 57486 17332
rect 57517 17323 57575 17329
rect 57517 17320 57529 17323
rect 57480 17292 57529 17320
rect 57480 17280 57486 17292
rect 57517 17289 57529 17292
rect 57563 17289 57575 17323
rect 57517 17283 57575 17289
rect 56781 17255 56839 17261
rect 56781 17221 56793 17255
rect 56827 17252 56839 17255
rect 57882 17252 57888 17264
rect 56827 17224 57888 17252
rect 56827 17221 56839 17224
rect 56781 17215 56839 17221
rect 57882 17212 57888 17224
rect 57940 17212 57946 17264
rect 56870 17144 56876 17196
rect 56928 17144 56934 17196
rect 53009 17119 53067 17125
rect 53009 17116 53021 17119
rect 52972 17088 53021 17116
rect 52972 17076 52978 17088
rect 53009 17085 53021 17088
rect 53055 17085 53067 17119
rect 54113 17119 54171 17125
rect 54113 17116 54125 17119
rect 53009 17079 53067 17085
rect 53484 17088 54125 17116
rect 53484 17057 53512 17088
rect 54113 17085 54125 17088
rect 54159 17085 54171 17119
rect 54113 17079 54171 17085
rect 56689 17119 56747 17125
rect 56689 17085 56701 17119
rect 56735 17085 56747 17119
rect 58437 17119 58495 17125
rect 58437 17116 58449 17119
rect 56689 17079 56747 17085
rect 57256 17088 58449 17116
rect 57256 17057 57284 17088
rect 58437 17085 58449 17088
rect 58483 17085 58495 17119
rect 58437 17079 58495 17085
rect 49513 17051 49571 17057
rect 49513 17017 49525 17051
rect 49559 17017 49571 17051
rect 49513 17011 49571 17017
rect 53469 17051 53527 17057
rect 53469 17017 53481 17051
rect 53515 17017 53527 17051
rect 53469 17011 53527 17017
rect 57241 17051 57299 17057
rect 57241 17017 57253 17051
rect 57287 17017 57299 17051
rect 57241 17011 57299 17017
rect 57330 17008 57336 17060
rect 57388 17048 57394 17060
rect 57885 17051 57943 17057
rect 57885 17048 57897 17051
rect 57388 17020 57897 17048
rect 57388 17008 57394 17020
rect 57885 17017 57897 17020
rect 57931 17017 57943 17051
rect 57885 17011 57943 17017
rect 36725 16983 36783 16989
rect 36725 16980 36737 16983
rect 36228 16952 36737 16980
rect 36228 16940 36234 16952
rect 36725 16949 36737 16952
rect 36771 16949 36783 16983
rect 36725 16943 36783 16949
rect 37277 16983 37335 16989
rect 37277 16949 37289 16983
rect 37323 16980 37335 16983
rect 37550 16980 37556 16992
rect 37323 16952 37556 16980
rect 37323 16949 37335 16952
rect 37277 16943 37335 16949
rect 37550 16940 37556 16952
rect 37608 16940 37614 16992
rect 38010 16940 38016 16992
rect 38068 16940 38074 16992
rect 40678 16940 40684 16992
rect 40736 16940 40742 16992
rect 43530 16940 43536 16992
rect 43588 16940 43594 16992
rect 50246 16940 50252 16992
rect 50304 16940 50310 16992
rect 53558 16940 53564 16992
rect 53616 16940 53622 16992
rect 56318 16940 56324 16992
rect 56376 16940 56382 16992
rect 56502 16940 56508 16992
rect 56560 16980 56566 16992
rect 56778 16980 56784 16992
rect 56560 16952 56784 16980
rect 56560 16940 56566 16952
rect 56778 16940 56784 16952
rect 56836 16940 56842 16992
rect 1104 16890 58880 16912
rect 1104 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 22616 16890
rect 22668 16838 22680 16890
rect 22732 16838 22744 16890
rect 22796 16838 22808 16890
rect 22860 16838 22872 16890
rect 22924 16838 37060 16890
rect 37112 16838 37124 16890
rect 37176 16838 37188 16890
rect 37240 16838 37252 16890
rect 37304 16838 37316 16890
rect 37368 16838 51504 16890
rect 51556 16838 51568 16890
rect 51620 16838 51632 16890
rect 51684 16838 51696 16890
rect 51748 16838 51760 16890
rect 51812 16838 58880 16890
rect 1104 16816 58880 16838
rect 6825 16779 6883 16785
rect 1596 16748 5304 16776
rect 1596 16652 1624 16748
rect 3878 16668 3884 16720
rect 3936 16668 3942 16720
rect 1578 16600 1584 16652
rect 1636 16600 1642 16652
rect 5276 16649 5304 16748
rect 6825 16745 6837 16779
rect 6871 16776 6883 16779
rect 6914 16776 6920 16788
rect 6871 16748 6920 16776
rect 6871 16745 6883 16748
rect 6825 16739 6883 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 8570 16736 8576 16788
rect 8628 16736 8634 16788
rect 9582 16736 9588 16788
rect 9640 16736 9646 16788
rect 11790 16736 11796 16788
rect 11848 16736 11854 16788
rect 15930 16736 15936 16788
rect 15988 16736 15994 16788
rect 16301 16779 16359 16785
rect 16301 16745 16313 16779
rect 16347 16776 16359 16779
rect 18138 16776 18144 16788
rect 16347 16748 18144 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18874 16776 18880 16788
rect 18279 16748 18880 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 19242 16736 19248 16788
rect 19300 16736 19306 16788
rect 21821 16779 21879 16785
rect 21821 16745 21833 16779
rect 21867 16776 21879 16779
rect 22370 16776 22376 16788
rect 21867 16748 22376 16776
rect 21867 16745 21879 16748
rect 21821 16739 21879 16745
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 22462 16736 22468 16788
rect 22520 16776 22526 16788
rect 22830 16776 22836 16788
rect 22520 16748 22836 16776
rect 22520 16736 22526 16748
rect 22830 16736 22836 16748
rect 22888 16736 22894 16788
rect 24854 16736 24860 16788
rect 24912 16736 24918 16788
rect 27249 16779 27307 16785
rect 27249 16745 27261 16779
rect 27295 16776 27307 16779
rect 27614 16776 27620 16788
rect 27295 16748 27620 16776
rect 27295 16745 27307 16748
rect 27249 16739 27307 16745
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 27706 16736 27712 16788
rect 27764 16736 27770 16788
rect 27890 16736 27896 16788
rect 27948 16736 27954 16788
rect 28074 16736 28080 16788
rect 28132 16776 28138 16788
rect 28445 16779 28503 16785
rect 28445 16776 28457 16779
rect 28132 16748 28457 16776
rect 28132 16736 28138 16748
rect 28445 16745 28457 16748
rect 28491 16745 28503 16779
rect 28445 16739 28503 16745
rect 30374 16736 30380 16788
rect 30432 16776 30438 16788
rect 30469 16779 30527 16785
rect 30469 16776 30481 16779
rect 30432 16748 30481 16776
rect 30432 16736 30438 16748
rect 30469 16745 30481 16748
rect 30515 16745 30527 16779
rect 35342 16776 35348 16788
rect 30469 16739 30527 16745
rect 34716 16748 35348 16776
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16640 6791 16643
rect 6779 16612 7328 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 3326 16572 3332 16584
rect 3283 16544 3332 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 7300 16581 7328 16612
rect 3513 16575 3571 16581
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 7009 16575 7067 16581
rect 7009 16572 7021 16575
rect 3559 16544 4660 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 1848 16507 1906 16513
rect 1848 16473 1860 16507
rect 1894 16504 1906 16507
rect 2498 16504 2504 16516
rect 1894 16476 2504 16504
rect 1894 16473 1906 16476
rect 1848 16467 1906 16473
rect 2498 16464 2504 16476
rect 2556 16464 2562 16516
rect 4632 16448 4660 16544
rect 5552 16544 7021 16572
rect 4890 16464 4896 16516
rect 4948 16504 4954 16516
rect 4994 16507 5052 16513
rect 4994 16504 5006 16507
rect 4948 16476 5006 16504
rect 4948 16464 4954 16476
rect 4994 16473 5006 16476
rect 5040 16473 5052 16507
rect 4994 16467 5052 16473
rect 5552 16448 5580 16544
rect 7009 16541 7021 16544
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16541 7251 16575
rect 7193 16535 7251 16541
rect 7285 16575 7343 16581
rect 7285 16541 7297 16575
rect 7331 16572 7343 16575
rect 7466 16572 7472 16584
rect 7331 16544 7472 16572
rect 7331 16541 7343 16544
rect 7285 16535 7343 16541
rect 2958 16396 2964 16448
rect 3016 16396 3022 16448
rect 3050 16396 3056 16448
rect 3108 16396 3114 16448
rect 3418 16396 3424 16448
rect 3476 16396 3482 16448
rect 4614 16396 4620 16448
rect 4672 16396 4678 16448
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 7208 16436 7236 16535
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 8297 16575 8355 16581
rect 8297 16541 8309 16575
rect 8343 16572 8355 16575
rect 8588 16572 8616 16736
rect 9217 16711 9275 16717
rect 9217 16708 9229 16711
rect 8343 16544 8616 16572
rect 8680 16680 9229 16708
rect 8343 16541 8355 16544
rect 8297 16535 8355 16541
rect 7561 16507 7619 16513
rect 7561 16473 7573 16507
rect 7607 16504 7619 16507
rect 8202 16504 8208 16516
rect 7607 16476 8208 16504
rect 7607 16473 7619 16476
rect 7561 16467 7619 16473
rect 8202 16464 8208 16476
rect 8260 16504 8266 16516
rect 8680 16504 8708 16680
rect 9217 16677 9229 16680
rect 9263 16708 9275 16711
rect 11808 16708 11836 16736
rect 9263 16680 11836 16708
rect 9263 16677 9275 16680
rect 9217 16671 9275 16677
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 17920 16680 19840 16708
rect 17920 16668 17926 16680
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9824 16612 10149 16640
rect 9824 16600 9830 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16356 16612 16957 16640
rect 16356 16600 16362 16612
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17218 16600 17224 16652
rect 17276 16600 17282 16652
rect 17497 16643 17555 16649
rect 17497 16609 17509 16643
rect 17543 16640 17555 16643
rect 17586 16640 17592 16652
rect 17543 16612 17592 16640
rect 17543 16609 17555 16612
rect 17497 16603 17555 16609
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 18141 16643 18199 16649
rect 18141 16640 18153 16643
rect 17788 16612 18153 16640
rect 17788 16584 17816 16612
rect 18141 16609 18153 16612
rect 18187 16609 18199 16643
rect 18141 16603 18199 16609
rect 18230 16600 18236 16652
rect 18288 16640 18294 16652
rect 19812 16649 19840 16680
rect 22204 16680 22508 16708
rect 22204 16652 22232 16680
rect 18693 16643 18751 16649
rect 18693 16640 18705 16643
rect 18288 16612 18705 16640
rect 18288 16600 18294 16612
rect 18693 16609 18705 16612
rect 18739 16609 18751 16643
rect 18693 16603 18751 16609
rect 18785 16643 18843 16649
rect 18785 16609 18797 16643
rect 18831 16609 18843 16643
rect 18785 16603 18843 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 14274 16532 14280 16584
rect 14332 16572 14338 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14332 16544 14565 16572
rect 14332 16532 14338 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 14820 16575 14878 16581
rect 14820 16541 14832 16575
rect 14866 16572 14878 16575
rect 15102 16572 15108 16584
rect 14866 16544 15108 16572
rect 14866 16541 14878 16544
rect 14820 16535 14878 16541
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 17034 16532 17040 16584
rect 17092 16581 17098 16584
rect 17092 16575 17141 16581
rect 17092 16541 17095 16575
rect 17129 16541 17141 16575
rect 17092 16535 17141 16541
rect 17092 16532 17098 16535
rect 17770 16532 17776 16584
rect 17828 16532 17834 16584
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16541 18015 16575
rect 17957 16535 18015 16541
rect 8260 16476 8708 16504
rect 17972 16504 18000 16535
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 18800 16572 18828 16603
rect 20530 16600 20536 16652
rect 20588 16600 20594 16652
rect 22186 16600 22192 16652
rect 22244 16600 22250 16652
rect 22480 16649 22508 16680
rect 22554 16668 22560 16720
rect 22612 16708 22618 16720
rect 23477 16711 23535 16717
rect 22612 16680 23060 16708
rect 22612 16668 22618 16680
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22830 16600 22836 16652
rect 22888 16600 22894 16652
rect 23032 16649 23060 16680
rect 23477 16677 23489 16711
rect 23523 16677 23535 16711
rect 23477 16671 23535 16677
rect 23017 16643 23075 16649
rect 23017 16609 23029 16643
rect 23063 16609 23075 16643
rect 23492 16640 23520 16671
rect 24872 16649 24900 16736
rect 24121 16643 24179 16649
rect 24121 16640 24133 16643
rect 23492 16612 24133 16640
rect 23017 16603 23075 16609
rect 24121 16609 24133 16612
rect 24167 16609 24179 16643
rect 24121 16603 24179 16609
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16609 25007 16643
rect 24949 16603 25007 16609
rect 18472 16544 18828 16572
rect 18472 16532 18478 16544
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20864 16544 21097 16572
rect 20864 16532 20870 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 22281 16575 22339 16581
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22922 16572 22928 16584
rect 22327 16544 22928 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 24486 16532 24492 16584
rect 24544 16572 24550 16584
rect 24765 16575 24823 16581
rect 24765 16572 24777 16575
rect 24544 16544 24777 16572
rect 24544 16532 24550 16544
rect 24765 16541 24777 16544
rect 24811 16541 24823 16575
rect 24964 16572 24992 16603
rect 25314 16600 25320 16652
rect 25372 16640 25378 16652
rect 27724 16649 27752 16736
rect 27908 16649 27936 16736
rect 25501 16643 25559 16649
rect 25501 16640 25513 16643
rect 25372 16612 25513 16640
rect 25372 16600 25378 16612
rect 25501 16609 25513 16612
rect 25547 16609 25559 16643
rect 25501 16603 25559 16609
rect 27709 16643 27767 16649
rect 27709 16609 27721 16643
rect 27755 16609 27767 16643
rect 27709 16603 27767 16609
rect 27893 16643 27951 16649
rect 27893 16609 27905 16643
rect 27939 16609 27951 16643
rect 27893 16603 27951 16609
rect 33134 16600 33140 16652
rect 33192 16640 33198 16652
rect 33321 16643 33379 16649
rect 33321 16640 33333 16643
rect 33192 16612 33333 16640
rect 33192 16600 33198 16612
rect 33321 16609 33333 16612
rect 33367 16640 33379 16643
rect 33686 16640 33692 16652
rect 33367 16612 33692 16640
rect 33367 16609 33379 16612
rect 33321 16603 33379 16609
rect 33686 16600 33692 16612
rect 33744 16600 33750 16652
rect 34514 16600 34520 16652
rect 34572 16640 34578 16652
rect 34716 16649 34744 16748
rect 35342 16736 35348 16748
rect 35400 16776 35406 16788
rect 36170 16776 36176 16788
rect 35400 16748 36176 16776
rect 35400 16736 35406 16748
rect 36170 16736 36176 16748
rect 36228 16736 36234 16788
rect 37458 16736 37464 16788
rect 37516 16776 37522 16788
rect 40678 16776 40684 16788
rect 37516 16748 39068 16776
rect 37516 16736 37522 16748
rect 36078 16668 36084 16720
rect 36136 16668 36142 16720
rect 36188 16649 36216 16736
rect 39040 16649 39068 16748
rect 40144 16748 40684 16776
rect 34701 16643 34759 16649
rect 34701 16640 34713 16643
rect 34572 16612 34713 16640
rect 34572 16600 34578 16612
rect 34701 16609 34713 16612
rect 34747 16609 34759 16643
rect 34701 16603 34759 16609
rect 36173 16643 36231 16649
rect 36173 16609 36185 16643
rect 36219 16609 36231 16643
rect 36173 16603 36231 16609
rect 39025 16643 39083 16649
rect 39025 16609 39037 16643
rect 39071 16609 39083 16643
rect 39025 16603 39083 16609
rect 40034 16600 40040 16652
rect 40092 16600 40098 16652
rect 40144 16649 40172 16748
rect 40678 16736 40684 16748
rect 40736 16736 40742 16788
rect 44545 16779 44603 16785
rect 44545 16776 44557 16779
rect 42904 16748 44557 16776
rect 40589 16711 40647 16717
rect 40589 16677 40601 16711
rect 40635 16677 40647 16711
rect 40589 16671 40647 16677
rect 40129 16643 40187 16649
rect 40129 16609 40141 16643
rect 40175 16609 40187 16643
rect 40604 16640 40632 16671
rect 41233 16643 41291 16649
rect 41233 16640 41245 16643
rect 40604 16612 41245 16640
rect 40129 16603 40187 16609
rect 41233 16609 41245 16612
rect 41279 16609 41291 16643
rect 41233 16603 41291 16609
rect 41414 16600 41420 16652
rect 41472 16600 41478 16652
rect 42904 16649 42932 16748
rect 44545 16745 44557 16748
rect 44591 16776 44603 16779
rect 45186 16776 45192 16788
rect 44591 16748 45192 16776
rect 44591 16745 44603 16748
rect 44545 16739 44603 16745
rect 45186 16736 45192 16748
rect 45244 16776 45250 16788
rect 45465 16779 45523 16785
rect 45465 16776 45477 16779
rect 45244 16748 45477 16776
rect 45244 16736 45250 16748
rect 45465 16745 45477 16748
rect 45511 16776 45523 16779
rect 48130 16776 48136 16788
rect 45511 16748 45692 16776
rect 45511 16745 45523 16748
rect 45465 16739 45523 16745
rect 45664 16649 45692 16748
rect 47872 16748 48136 16776
rect 47872 16649 47900 16748
rect 48130 16736 48136 16748
rect 48188 16736 48194 16788
rect 50157 16779 50215 16785
rect 50157 16745 50169 16779
rect 50203 16776 50215 16779
rect 50890 16776 50896 16788
rect 50203 16748 50896 16776
rect 50203 16745 50215 16748
rect 50157 16739 50215 16745
rect 50890 16736 50896 16748
rect 50948 16736 50954 16788
rect 53006 16736 53012 16788
rect 53064 16776 53070 16788
rect 53193 16779 53251 16785
rect 53193 16776 53205 16779
rect 53064 16748 53205 16776
rect 53064 16736 53070 16748
rect 53193 16745 53205 16748
rect 53239 16745 53251 16779
rect 53193 16739 53251 16745
rect 55125 16779 55183 16785
rect 55125 16745 55137 16779
rect 55171 16776 55183 16779
rect 55858 16776 55864 16788
rect 55171 16748 55864 16776
rect 55171 16745 55183 16748
rect 55125 16739 55183 16745
rect 55858 16736 55864 16748
rect 55916 16736 55922 16788
rect 56594 16776 56600 16788
rect 55968 16748 56600 16776
rect 54297 16711 54355 16717
rect 54297 16708 54309 16711
rect 53760 16680 54309 16708
rect 53760 16652 53788 16680
rect 54297 16677 54309 16680
rect 54343 16677 54355 16711
rect 55968 16708 55996 16748
rect 56594 16736 56600 16748
rect 56652 16736 56658 16788
rect 56778 16736 56784 16788
rect 56836 16736 56842 16788
rect 56870 16736 56876 16788
rect 56928 16776 56934 16788
rect 56928 16748 58112 16776
rect 56928 16736 56934 16748
rect 54297 16671 54355 16677
rect 54680 16680 55996 16708
rect 56796 16708 56824 16736
rect 56796 16680 56916 16708
rect 42889 16643 42947 16649
rect 42889 16640 42901 16643
rect 42812 16612 42901 16640
rect 24765 16535 24823 16541
rect 24872 16544 24992 16572
rect 18598 16504 18604 16516
rect 17972 16476 18604 16504
rect 8260 16464 8266 16476
rect 18598 16464 18604 16476
rect 18656 16464 18662 16516
rect 20349 16507 20407 16513
rect 20349 16473 20361 16507
rect 20395 16504 20407 16507
rect 21174 16504 21180 16516
rect 20395 16476 21180 16504
rect 20395 16473 20407 16476
rect 20349 16467 20407 16473
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 21729 16507 21787 16513
rect 21729 16473 21741 16507
rect 21775 16504 21787 16507
rect 21775 16476 22784 16504
rect 21775 16473 21787 16476
rect 21729 16467 21787 16473
rect 22756 16448 22784 16476
rect 24578 16464 24584 16516
rect 24636 16504 24642 16516
rect 24872 16504 24900 16544
rect 26050 16532 26056 16584
rect 26108 16572 26114 16584
rect 26108 16544 28672 16572
rect 26108 16532 26114 16544
rect 24636 16476 24900 16504
rect 24636 16464 24642 16476
rect 24946 16464 24952 16516
rect 25004 16464 25010 16516
rect 25768 16507 25826 16513
rect 25768 16473 25780 16507
rect 25814 16504 25826 16507
rect 25958 16504 25964 16516
rect 25814 16476 25964 16504
rect 25814 16473 25826 16476
rect 25768 16467 25826 16473
rect 25958 16464 25964 16476
rect 26016 16464 26022 16516
rect 27617 16507 27675 16513
rect 27617 16473 27629 16507
rect 27663 16504 27675 16507
rect 27798 16504 27804 16516
rect 27663 16476 27804 16504
rect 27663 16473 27675 16476
rect 27617 16467 27675 16473
rect 27798 16464 27804 16476
rect 27856 16464 27862 16516
rect 28644 16504 28672 16544
rect 28718 16532 28724 16584
rect 28776 16532 28782 16584
rect 30190 16532 30196 16584
rect 30248 16532 30254 16584
rect 31754 16532 31760 16584
rect 31812 16532 31818 16584
rect 32122 16532 32128 16584
rect 32180 16532 32186 16584
rect 32493 16575 32551 16581
rect 32493 16541 32505 16575
rect 32539 16541 32551 16575
rect 32493 16535 32551 16541
rect 29454 16504 29460 16516
rect 28644 16476 29460 16504
rect 29454 16464 29460 16476
rect 29512 16464 29518 16516
rect 29546 16464 29552 16516
rect 29604 16504 29610 16516
rect 31772 16504 31800 16532
rect 32508 16504 32536 16535
rect 29604 16476 31432 16504
rect 31772 16476 32536 16504
rect 33704 16504 33732 16600
rect 34146 16532 34152 16584
rect 34204 16532 34210 16584
rect 34968 16575 35026 16581
rect 34968 16541 34980 16575
rect 35014 16572 35026 16575
rect 35802 16572 35808 16584
rect 35014 16544 35808 16572
rect 35014 16541 35026 16544
rect 34968 16535 35026 16541
rect 35802 16532 35808 16544
rect 35860 16532 35866 16584
rect 36440 16575 36498 16581
rect 36440 16541 36452 16575
rect 36486 16572 36498 16575
rect 37550 16572 37556 16584
rect 36486 16544 37556 16572
rect 36486 16541 36498 16544
rect 36440 16535 36498 16541
rect 37550 16532 37556 16544
rect 37608 16532 37614 16584
rect 37458 16504 37464 16516
rect 33704 16476 37464 16504
rect 29604 16464 29610 16476
rect 6880 16408 7236 16436
rect 6880 16396 6886 16408
rect 19978 16396 19984 16448
rect 20036 16396 20042 16448
rect 20441 16439 20499 16445
rect 20441 16405 20453 16439
rect 20487 16436 20499 16439
rect 21266 16436 21272 16448
rect 20487 16408 21272 16436
rect 20487 16405 20499 16408
rect 20441 16399 20499 16405
rect 21266 16396 21272 16408
rect 21324 16436 21330 16448
rect 22186 16436 22192 16448
rect 21324 16408 22192 16436
rect 21324 16396 21330 16408
rect 22186 16396 22192 16408
rect 22244 16436 22250 16448
rect 22554 16436 22560 16448
rect 22244 16408 22560 16436
rect 22244 16396 22250 16408
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 22738 16396 22744 16448
rect 22796 16396 22802 16448
rect 23106 16396 23112 16448
rect 23164 16396 23170 16448
rect 23290 16396 23296 16448
rect 23348 16436 23354 16448
rect 23569 16439 23627 16445
rect 23569 16436 23581 16439
rect 23348 16408 23581 16436
rect 23348 16396 23354 16408
rect 23569 16405 23581 16408
rect 23615 16405 23627 16439
rect 23569 16399 23627 16405
rect 24397 16439 24455 16445
rect 24397 16405 24409 16439
rect 24443 16436 24455 16439
rect 24964 16436 24992 16464
rect 31404 16448 31432 16476
rect 37458 16464 37464 16476
rect 37516 16464 37522 16516
rect 38654 16504 38660 16516
rect 37568 16476 38660 16504
rect 24443 16408 24992 16436
rect 24443 16405 24455 16408
rect 24397 16399 24455 16405
rect 26878 16396 26884 16448
rect 26936 16396 26942 16448
rect 29362 16396 29368 16448
rect 29420 16396 29426 16448
rect 31294 16396 31300 16448
rect 31352 16396 31358 16448
rect 31386 16396 31392 16448
rect 31444 16396 31450 16448
rect 31478 16396 31484 16448
rect 31536 16396 31542 16448
rect 33594 16396 33600 16448
rect 33652 16396 33658 16448
rect 37568 16445 37596 16476
rect 38654 16464 38660 16476
rect 38712 16464 38718 16516
rect 38780 16507 38838 16513
rect 38780 16473 38792 16507
rect 38826 16504 38838 16507
rect 38930 16504 38936 16516
rect 38826 16476 38936 16504
rect 38826 16473 38838 16476
rect 38780 16467 38838 16473
rect 38930 16464 38936 16476
rect 38988 16464 38994 16516
rect 40052 16504 40080 16600
rect 40221 16575 40279 16581
rect 40221 16541 40233 16575
rect 40267 16572 40279 16575
rect 40586 16572 40592 16584
rect 40267 16544 40592 16572
rect 40267 16541 40279 16544
rect 40221 16535 40279 16541
rect 40586 16532 40592 16544
rect 40644 16532 40650 16584
rect 42150 16532 42156 16584
rect 42208 16572 42214 16584
rect 42812 16572 42840 16612
rect 42889 16609 42901 16612
rect 42935 16609 42947 16643
rect 42889 16603 42947 16609
rect 45649 16643 45707 16649
rect 45649 16609 45661 16643
rect 45695 16609 45707 16643
rect 45649 16603 45707 16609
rect 47857 16643 47915 16649
rect 47857 16609 47869 16643
rect 47903 16609 47915 16643
rect 47857 16603 47915 16609
rect 49050 16600 49056 16652
rect 49108 16640 49114 16652
rect 49881 16643 49939 16649
rect 49881 16640 49893 16643
rect 49108 16612 49893 16640
rect 49108 16600 49114 16612
rect 49881 16609 49893 16612
rect 49927 16609 49939 16643
rect 49881 16603 49939 16609
rect 50154 16600 50160 16652
rect 50212 16640 50218 16652
rect 50709 16643 50767 16649
rect 50709 16640 50721 16643
rect 50212 16612 50721 16640
rect 50212 16600 50218 16612
rect 50709 16609 50721 16612
rect 50755 16609 50767 16643
rect 50709 16603 50767 16609
rect 51166 16600 51172 16652
rect 51224 16640 51230 16652
rect 51718 16640 51724 16652
rect 51224 16612 51724 16640
rect 51224 16600 51230 16612
rect 51718 16600 51724 16612
rect 51776 16600 51782 16652
rect 53650 16600 53656 16652
rect 53708 16600 53714 16652
rect 53742 16600 53748 16652
rect 53800 16600 53806 16652
rect 53834 16600 53840 16652
rect 53892 16600 53898 16652
rect 54202 16600 54208 16652
rect 54260 16640 54266 16652
rect 54680 16649 54708 16680
rect 54481 16643 54539 16649
rect 54481 16640 54493 16643
rect 54260 16612 54493 16640
rect 54260 16600 54266 16612
rect 54481 16609 54493 16612
rect 54527 16640 54539 16643
rect 54665 16643 54723 16649
rect 54527 16612 54616 16640
rect 54527 16609 54539 16612
rect 54481 16603 54539 16609
rect 42208 16544 42840 16572
rect 43156 16575 43214 16581
rect 42208 16532 42214 16544
rect 43156 16541 43168 16575
rect 43202 16572 43214 16575
rect 43530 16572 43536 16584
rect 43202 16544 43536 16572
rect 43202 16541 43214 16544
rect 43156 16535 43214 16541
rect 43530 16532 43536 16544
rect 43588 16532 43594 16584
rect 47670 16532 47676 16584
rect 47728 16532 47734 16584
rect 48056 16544 49464 16572
rect 42061 16507 42119 16513
rect 40052 16476 40816 16504
rect 37553 16439 37611 16445
rect 37553 16405 37565 16439
rect 37599 16405 37611 16439
rect 37553 16399 37611 16405
rect 37642 16396 37648 16448
rect 37700 16396 37706 16448
rect 39022 16396 39028 16448
rect 39080 16436 39086 16448
rect 39577 16439 39635 16445
rect 39577 16436 39589 16439
rect 39080 16408 39589 16436
rect 39080 16396 39086 16408
rect 39577 16405 39589 16408
rect 39623 16405 39635 16439
rect 39577 16399 39635 16405
rect 40678 16396 40684 16448
rect 40736 16396 40742 16448
rect 40788 16436 40816 16476
rect 42061 16473 42073 16507
rect 42107 16504 42119 16507
rect 45916 16507 45974 16513
rect 42107 16476 43208 16504
rect 42107 16473 42119 16476
rect 42061 16467 42119 16473
rect 43180 16448 43208 16476
rect 45916 16473 45928 16507
rect 45962 16504 45974 16507
rect 47121 16507 47179 16513
rect 47121 16504 47133 16507
rect 45962 16476 47133 16504
rect 45962 16473 45974 16476
rect 45916 16467 45974 16473
rect 47121 16473 47133 16476
rect 47167 16473 47179 16507
rect 47121 16467 47179 16473
rect 42334 16436 42340 16448
rect 40788 16408 42340 16436
rect 42334 16396 42340 16408
rect 42392 16436 42398 16448
rect 42705 16439 42763 16445
rect 42705 16436 42717 16439
rect 42392 16408 42717 16436
rect 42392 16396 42398 16408
rect 42705 16405 42717 16408
rect 42751 16405 42763 16439
rect 42705 16399 42763 16405
rect 43162 16396 43168 16448
rect 43220 16396 43226 16448
rect 44269 16439 44327 16445
rect 44269 16405 44281 16439
rect 44315 16436 44327 16439
rect 45002 16436 45008 16448
rect 44315 16408 45008 16436
rect 44315 16405 44327 16408
rect 44269 16399 44327 16405
rect 45002 16396 45008 16408
rect 45060 16396 45066 16448
rect 47026 16396 47032 16448
rect 47084 16396 47090 16448
rect 48056 16436 48084 16544
rect 48124 16507 48182 16513
rect 48124 16473 48136 16507
rect 48170 16504 48182 16507
rect 49329 16507 49387 16513
rect 49329 16504 49341 16507
rect 48170 16476 49341 16504
rect 48170 16473 48182 16476
rect 48124 16467 48182 16473
rect 49329 16473 49341 16476
rect 49375 16473 49387 16507
rect 49436 16504 49464 16544
rect 50982 16532 50988 16584
rect 51040 16532 51046 16584
rect 51988 16575 52046 16581
rect 51988 16541 52000 16575
rect 52034 16572 52046 16575
rect 53558 16572 53564 16584
rect 52034 16544 53564 16572
rect 52034 16541 52046 16544
rect 51988 16535 52046 16541
rect 53558 16532 53564 16544
rect 53616 16532 53622 16584
rect 52362 16504 52368 16516
rect 49436 16476 52368 16504
rect 49329 16467 49387 16473
rect 52362 16464 52368 16476
rect 52420 16464 52426 16516
rect 53852 16504 53880 16600
rect 54588 16572 54616 16612
rect 54665 16609 54677 16643
rect 54711 16609 54723 16643
rect 55493 16643 55551 16649
rect 55493 16640 55505 16643
rect 54665 16603 54723 16609
rect 54772 16612 55505 16640
rect 54772 16572 54800 16612
rect 55493 16609 55505 16612
rect 55539 16609 55551 16643
rect 55493 16603 55551 16609
rect 55677 16643 55735 16649
rect 55677 16609 55689 16643
rect 55723 16640 55735 16643
rect 56778 16640 56784 16652
rect 55723 16612 56784 16640
rect 55723 16609 55735 16612
rect 55677 16603 55735 16609
rect 56778 16600 56784 16612
rect 56836 16600 56842 16652
rect 56888 16649 56916 16680
rect 56873 16643 56931 16649
rect 56873 16609 56885 16643
rect 56919 16609 56931 16643
rect 56873 16603 56931 16609
rect 57517 16643 57575 16649
rect 57517 16609 57529 16643
rect 57563 16640 57575 16643
rect 57882 16640 57888 16652
rect 57563 16612 57888 16640
rect 57563 16609 57575 16612
rect 57517 16603 57575 16609
rect 57882 16600 57888 16612
rect 57940 16600 57946 16652
rect 58084 16649 58112 16748
rect 58069 16643 58127 16649
rect 58069 16609 58081 16643
rect 58115 16609 58127 16643
rect 58069 16603 58127 16609
rect 58158 16600 58164 16652
rect 58216 16600 58222 16652
rect 54588 16544 54800 16572
rect 56318 16532 56324 16584
rect 56376 16532 56382 16584
rect 56410 16532 56416 16584
rect 56468 16581 56474 16584
rect 56468 16575 56517 16581
rect 56468 16541 56471 16575
rect 56505 16541 56517 16575
rect 56468 16535 56517 16541
rect 56468 16532 56474 16535
rect 56594 16532 56600 16584
rect 56652 16532 56658 16584
rect 57333 16575 57391 16581
rect 57333 16541 57345 16575
rect 57379 16541 57391 16575
rect 57333 16535 57391 16541
rect 53116 16476 53880 16504
rect 57348 16504 57376 16535
rect 57348 16476 57928 16504
rect 48222 16436 48228 16448
rect 48056 16408 48228 16436
rect 48222 16396 48228 16408
rect 48280 16396 48286 16448
rect 49234 16396 49240 16448
rect 49292 16396 49298 16448
rect 49418 16396 49424 16448
rect 49476 16436 49482 16448
rect 50246 16436 50252 16448
rect 49476 16408 50252 16436
rect 49476 16396 49482 16408
rect 50246 16396 50252 16408
rect 50304 16436 50310 16448
rect 50525 16439 50583 16445
rect 50525 16436 50537 16439
rect 50304 16408 50537 16436
rect 50304 16396 50310 16408
rect 50525 16405 50537 16408
rect 50571 16405 50583 16439
rect 50525 16399 50583 16405
rect 50614 16396 50620 16448
rect 50672 16396 50678 16448
rect 51629 16439 51687 16445
rect 51629 16405 51641 16439
rect 51675 16436 51687 16439
rect 52546 16436 52552 16448
rect 51675 16408 52552 16436
rect 51675 16405 51687 16408
rect 51629 16399 51687 16405
rect 52546 16396 52552 16408
rect 52604 16396 52610 16448
rect 53116 16445 53144 16476
rect 57900 16448 57928 16476
rect 53101 16439 53159 16445
rect 53101 16405 53113 16439
rect 53147 16405 53159 16439
rect 53101 16399 53159 16405
rect 53558 16396 53564 16448
rect 53616 16436 53622 16448
rect 54757 16439 54815 16445
rect 54757 16436 54769 16439
rect 53616 16408 54769 16436
rect 53616 16396 53622 16408
rect 54757 16405 54769 16408
rect 54803 16436 54815 16439
rect 55214 16436 55220 16448
rect 54803 16408 55220 16436
rect 54803 16405 54815 16408
rect 54757 16399 54815 16405
rect 55214 16396 55220 16408
rect 55272 16436 55278 16448
rect 56870 16436 56876 16448
rect 55272 16408 56876 16436
rect 55272 16396 55278 16408
rect 56870 16396 56876 16408
rect 56928 16396 56934 16448
rect 57606 16396 57612 16448
rect 57664 16396 57670 16448
rect 57882 16396 57888 16448
rect 57940 16436 57946 16448
rect 57977 16439 58035 16445
rect 57977 16436 57989 16439
rect 57940 16408 57989 16436
rect 57940 16396 57946 16408
rect 57977 16405 57989 16408
rect 58023 16405 58035 16439
rect 57977 16399 58035 16405
rect 1104 16346 59040 16368
rect 1104 16294 15394 16346
rect 15446 16294 15458 16346
rect 15510 16294 15522 16346
rect 15574 16294 15586 16346
rect 15638 16294 15650 16346
rect 15702 16294 29838 16346
rect 29890 16294 29902 16346
rect 29954 16294 29966 16346
rect 30018 16294 30030 16346
rect 30082 16294 30094 16346
rect 30146 16294 44282 16346
rect 44334 16294 44346 16346
rect 44398 16294 44410 16346
rect 44462 16294 44474 16346
rect 44526 16294 44538 16346
rect 44590 16294 58726 16346
rect 58778 16294 58790 16346
rect 58842 16294 58854 16346
rect 58906 16294 58918 16346
rect 58970 16294 58982 16346
rect 59034 16294 59040 16346
rect 1104 16272 59040 16294
rect 2498 16192 2504 16244
rect 2556 16192 2562 16244
rect 2958 16192 2964 16244
rect 3016 16192 3022 16244
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3476 16204 3893 16232
rect 3476 16192 3482 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 4890 16192 4896 16244
rect 4948 16192 4954 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16574 16232 16580 16244
rect 16163 16204 16580 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16574 16192 16580 16204
rect 16632 16232 16638 16244
rect 17034 16232 17040 16244
rect 16632 16204 17040 16232
rect 16632 16192 16638 16204
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 18598 16192 18604 16244
rect 18656 16192 18662 16244
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 20898 16192 20904 16244
rect 20956 16192 20962 16244
rect 21266 16192 21272 16244
rect 21324 16192 21330 16244
rect 21361 16235 21419 16241
rect 21361 16201 21373 16235
rect 21407 16232 21419 16235
rect 22738 16232 22744 16244
rect 21407 16204 22744 16232
rect 21407 16201 21419 16204
rect 21361 16195 21419 16201
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 24949 16235 25007 16241
rect 23164 16204 23520 16232
rect 23164 16192 23170 16204
rect 2976 16164 3004 16192
rect 2976 16136 3280 16164
rect 3050 16056 3056 16108
rect 3108 16056 3114 16108
rect 3252 16105 3280 16136
rect 4522 16124 4528 16176
rect 4580 16164 4586 16176
rect 5261 16167 5319 16173
rect 5261 16164 5273 16167
rect 4580 16136 5273 16164
rect 4580 16124 4586 16136
rect 5261 16133 5273 16136
rect 5307 16133 5319 16167
rect 8389 16167 8447 16173
rect 8389 16164 8401 16167
rect 5261 16127 5319 16133
rect 7116 16136 8401 16164
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16065 3295 16099
rect 3237 16059 3295 16065
rect 4614 16056 4620 16108
rect 4672 16096 4678 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4672 16068 5181 16096
rect 4672 16056 4678 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 5350 16056 5356 16108
rect 5408 16056 5414 16108
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5626 16096 5632 16108
rect 5583 16068 5632 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 5626 16056 5632 16068
rect 5684 16056 5690 16108
rect 7116 16105 7144 16136
rect 8389 16133 8401 16136
rect 8435 16133 8447 16167
rect 8389 16127 8447 16133
rect 17396 16167 17454 16173
rect 17396 16133 17408 16167
rect 17442 16164 17454 16167
rect 18322 16164 18328 16176
rect 17442 16136 18328 16164
rect 17442 16133 17454 16136
rect 17396 16127 17454 16133
rect 18322 16124 18328 16136
rect 18380 16124 18386 16176
rect 19696 16167 19754 16173
rect 19696 16133 19708 16167
rect 19742 16164 19754 16167
rect 20346 16164 20352 16176
rect 19742 16136 20352 16164
rect 19742 16133 19754 16136
rect 19696 16127 19754 16133
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 8202 16056 8208 16108
rect 8260 16056 8266 16108
rect 8754 16096 8760 16108
rect 8312 16068 8760 16096
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 15997 4399 16031
rect 4341 15991 4399 15997
rect 4356 15960 4384 15991
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 7282 16028 7288 16040
rect 6788 16000 7288 16028
rect 6788 15988 6794 16000
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 8312 16028 8340 16068
rect 8754 16056 8760 16068
rect 8812 16096 8818 16108
rect 14544 16099 14602 16105
rect 8812 16068 9536 16096
rect 8812 16056 8818 16068
rect 7524 16000 8340 16028
rect 9033 16031 9091 16037
rect 7524 15988 7530 16000
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9079 16000 9444 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 4985 15963 5043 15969
rect 4985 15960 4997 15963
rect 4356 15932 4997 15960
rect 4985 15929 4997 15932
rect 5031 15929 5043 15963
rect 4985 15923 5043 15929
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6181 15895 6239 15901
rect 6181 15892 6193 15895
rect 6052 15864 6193 15892
rect 6052 15852 6058 15864
rect 6181 15861 6193 15864
rect 6227 15892 6239 15895
rect 6546 15892 6552 15904
rect 6227 15864 6552 15892
rect 6227 15861 6239 15864
rect 6181 15855 6239 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 9416 15901 9444 16000
rect 9508 15972 9536 16068
rect 14544 16065 14556 16099
rect 14590 16096 14602 16099
rect 14826 16096 14832 16108
rect 14590 16068 14832 16096
rect 14590 16065 14602 16068
rect 14544 16059 14602 16065
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 16114 16096 16120 16108
rect 15580 16068 16120 16096
rect 15580 16040 15608 16068
rect 16114 16056 16120 16068
rect 16172 16096 16178 16108
rect 16172 16068 16344 16096
rect 16172 16056 16178 16068
rect 10870 15988 10876 16040
rect 10928 15988 10934 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12492 16000 13001 16028
rect 12492 15988 12498 16000
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 14274 15988 14280 16040
rect 14332 15988 14338 16040
rect 15562 15988 15568 16040
rect 15620 15988 15626 16040
rect 15838 15988 15844 16040
rect 15896 16028 15902 16040
rect 16316 16037 16344 16068
rect 20732 16068 21496 16096
rect 20732 16040 20760 16068
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15896 16000 16221 16028
rect 15896 15988 15902 16000
rect 16209 15997 16221 16000
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 16301 16031 16359 16037
rect 16301 15997 16313 16031
rect 16347 15997 16359 16031
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 16301 15991 16359 15997
rect 16868 16000 17141 16028
rect 9490 15920 9496 15972
rect 9548 15960 9554 15972
rect 9769 15963 9827 15969
rect 9769 15960 9781 15963
rect 9548 15932 9781 15960
rect 9548 15920 9554 15932
rect 9769 15929 9781 15932
rect 9815 15960 9827 15963
rect 15657 15963 15715 15969
rect 9815 15932 11652 15960
rect 9815 15929 9827 15932
rect 9769 15923 9827 15929
rect 11624 15904 11652 15932
rect 15657 15929 15669 15963
rect 15703 15960 15715 15963
rect 15930 15960 15936 15972
rect 15703 15932 15936 15960
rect 15703 15929 15715 15932
rect 15657 15923 15715 15929
rect 15930 15920 15936 15932
rect 15988 15920 15994 15972
rect 9401 15895 9459 15901
rect 9401 15861 9413 15895
rect 9447 15892 9459 15895
rect 9582 15892 9588 15904
rect 9447 15864 9588 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 10318 15852 10324 15904
rect 10376 15852 10382 15904
rect 11606 15852 11612 15904
rect 11664 15852 11670 15904
rect 11793 15895 11851 15901
rect 11793 15861 11805 15895
rect 11839 15892 11851 15895
rect 12066 15892 12072 15904
rect 11839 15864 12072 15892
rect 11839 15861 11851 15864
rect 11793 15855 11851 15861
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12437 15895 12495 15901
rect 12437 15892 12449 15895
rect 12400 15864 12449 15892
rect 12400 15852 12406 15864
rect 12437 15861 12449 15864
rect 12483 15861 12495 15895
rect 12437 15855 12495 15861
rect 13170 15852 13176 15904
rect 13228 15852 13234 15904
rect 15746 15852 15752 15904
rect 15804 15852 15810 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16868 15901 16896 16000
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 19153 16031 19211 16037
rect 19153 15997 19165 16031
rect 19199 15997 19211 16031
rect 19153 15991 19211 15997
rect 18509 15963 18567 15969
rect 18509 15929 18521 15963
rect 18555 15960 18567 15963
rect 19168 15960 19196 15991
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 19300 16000 19441 16028
rect 19300 15988 19306 16000
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 20714 15988 20720 16040
rect 20772 15988 20778 16040
rect 21174 15988 21180 16040
rect 21232 15988 21238 16040
rect 21468 16037 21496 16068
rect 22462 16056 22468 16108
rect 22520 16056 22526 16108
rect 22738 16056 22744 16108
rect 22796 16056 22802 16108
rect 23492 16105 23520 16204
rect 24949 16201 24961 16235
rect 24995 16232 25007 16235
rect 25314 16232 25320 16244
rect 24995 16204 25320 16232
rect 24995 16201 25007 16204
rect 24949 16195 25007 16201
rect 25314 16192 25320 16204
rect 25372 16232 25378 16244
rect 25869 16235 25927 16241
rect 25869 16232 25881 16235
rect 25372 16204 25881 16232
rect 25372 16192 25378 16204
rect 25869 16201 25881 16204
rect 25915 16201 25927 16235
rect 25869 16195 25927 16201
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23753 16099 23811 16105
rect 23753 16096 23765 16099
rect 23523 16068 23765 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23753 16065 23765 16068
rect 23799 16065 23811 16099
rect 25884 16096 25912 16195
rect 26418 16192 26424 16244
rect 26476 16232 26482 16244
rect 26476 16204 27108 16232
rect 26476 16192 26482 16204
rect 27080 16108 27108 16204
rect 29362 16192 29368 16244
rect 29420 16192 29426 16244
rect 29917 16235 29975 16241
rect 29917 16201 29929 16235
rect 29963 16232 29975 16235
rect 30190 16232 30196 16244
rect 29963 16204 30196 16232
rect 29963 16201 29975 16204
rect 29917 16195 29975 16201
rect 30190 16192 30196 16204
rect 30248 16192 30254 16244
rect 30374 16192 30380 16244
rect 30432 16192 30438 16244
rect 31478 16192 31484 16244
rect 31536 16192 31542 16244
rect 31938 16192 31944 16244
rect 31996 16192 32002 16244
rect 32122 16192 32128 16244
rect 32180 16192 32186 16244
rect 32490 16192 32496 16244
rect 32548 16232 32554 16244
rect 32585 16235 32643 16241
rect 32585 16232 32597 16235
rect 32548 16204 32597 16232
rect 32548 16192 32554 16204
rect 32585 16201 32597 16204
rect 32631 16232 32643 16235
rect 32950 16232 32956 16244
rect 32631 16204 32956 16232
rect 32631 16201 32643 16204
rect 32585 16195 32643 16201
rect 32950 16192 32956 16204
rect 33008 16192 33014 16244
rect 33689 16235 33747 16241
rect 33689 16201 33701 16235
rect 33735 16232 33747 16235
rect 34146 16232 34152 16244
rect 33735 16204 34152 16232
rect 33735 16201 33747 16204
rect 33689 16195 33747 16201
rect 34146 16192 34152 16204
rect 34204 16192 34210 16244
rect 37642 16192 37648 16244
rect 37700 16192 37706 16244
rect 37918 16192 37924 16244
rect 37976 16232 37982 16244
rect 38013 16235 38071 16241
rect 38013 16232 38025 16235
rect 37976 16204 38025 16232
rect 37976 16192 37982 16204
rect 38013 16201 38025 16204
rect 38059 16201 38071 16235
rect 38013 16195 38071 16201
rect 40678 16192 40684 16244
rect 40736 16192 40742 16244
rect 43809 16235 43867 16241
rect 43809 16201 43821 16235
rect 43855 16232 43867 16235
rect 43990 16232 43996 16244
rect 43855 16204 43996 16232
rect 43855 16201 43867 16204
rect 43809 16195 43867 16201
rect 43990 16192 43996 16204
rect 44048 16192 44054 16244
rect 45186 16192 45192 16244
rect 45244 16192 45250 16244
rect 47026 16192 47032 16244
rect 47084 16232 47090 16244
rect 50433 16235 50491 16241
rect 47084 16204 49556 16232
rect 47084 16192 47090 16204
rect 27246 16173 27252 16176
rect 27240 16164 27252 16173
rect 27207 16136 27252 16164
rect 27240 16127 27252 16136
rect 27246 16124 27252 16127
rect 27304 16124 27310 16176
rect 28804 16167 28862 16173
rect 28804 16133 28816 16167
rect 28850 16164 28862 16167
rect 29380 16164 29408 16192
rect 28850 16136 29408 16164
rect 28850 16133 28862 16136
rect 28804 16127 28862 16133
rect 26050 16096 26056 16108
rect 25884 16068 26056 16096
rect 23753 16059 23811 16065
rect 26050 16056 26056 16068
rect 26108 16096 26114 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26108 16068 26985 16096
rect 26108 16056 26114 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27062 16056 27068 16108
rect 27120 16056 27126 16108
rect 30392 16096 30420 16192
rect 30828 16167 30886 16173
rect 30828 16133 30840 16167
rect 30874 16164 30886 16167
rect 31496 16164 31524 16192
rect 30874 16136 31524 16164
rect 37660 16164 37688 16192
rect 39108 16167 39166 16173
rect 37660 16136 38700 16164
rect 30874 16133 30886 16136
rect 30828 16127 30886 16133
rect 30561 16099 30619 16105
rect 30561 16096 30573 16099
rect 28000 16068 29592 16096
rect 30392 16068 30573 16096
rect 21453 16031 21511 16037
rect 21453 15997 21465 16031
rect 21499 15997 21511 16031
rect 22603 16031 22661 16037
rect 22603 16028 22615 16031
rect 21453 15991 21511 15997
rect 22066 16000 22615 16028
rect 18555 15932 19196 15960
rect 21192 15960 21220 15988
rect 22066 15960 22094 16000
rect 22603 15997 22615 16000
rect 22649 15997 22661 16031
rect 22603 15991 22661 15997
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 23106 16028 23112 16040
rect 22980 16000 23112 16028
rect 22980 15988 22986 16000
rect 23106 15988 23112 16000
rect 23164 16028 23170 16040
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 23164 16000 23673 16028
rect 23164 15988 23170 16000
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 23661 15991 23719 15997
rect 24302 15988 24308 16040
rect 24360 15988 24366 16040
rect 24394 15988 24400 16040
rect 24452 16028 24458 16040
rect 26145 16031 26203 16037
rect 26145 16028 26157 16031
rect 24452 16000 26157 16028
rect 24452 15988 24458 16000
rect 21192 15932 22094 15960
rect 18555 15929 18567 15932
rect 18509 15923 18567 15929
rect 23014 15920 23020 15972
rect 23072 15920 23078 15972
rect 25516 15904 25544 16000
rect 26145 15997 26157 16000
rect 26191 15997 26203 16031
rect 26145 15991 26203 15997
rect 26160 15960 26188 15991
rect 26326 15988 26332 16040
rect 26384 15988 26390 16040
rect 26160 15932 27016 15960
rect 16853 15895 16911 15901
rect 16853 15892 16865 15895
rect 16448 15864 16865 15892
rect 16448 15852 16454 15864
rect 16853 15861 16865 15864
rect 16899 15861 16911 15895
rect 16853 15855 16911 15861
rect 21821 15895 21879 15901
rect 21821 15861 21833 15895
rect 21867 15892 21879 15895
rect 21910 15892 21916 15904
rect 21867 15864 21916 15892
rect 21867 15861 21879 15864
rect 21821 15855 21879 15861
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 23198 15892 23204 15904
rect 22520 15864 23204 15892
rect 22520 15852 22526 15864
rect 23198 15852 23204 15864
rect 23256 15852 23262 15904
rect 25498 15852 25504 15904
rect 25556 15852 25562 15904
rect 26786 15852 26792 15904
rect 26844 15852 26850 15904
rect 26988 15892 27016 15932
rect 28000 15892 28028 16068
rect 28074 15988 28080 16040
rect 28132 16028 28138 16040
rect 28534 16028 28540 16040
rect 28132 16000 28540 16028
rect 28132 15988 28138 16000
rect 28534 15988 28540 16000
rect 28592 15988 28598 16040
rect 29564 16028 29592 16068
rect 30561 16065 30573 16068
rect 30607 16065 30619 16099
rect 31294 16096 31300 16108
rect 30561 16059 30619 16065
rect 30668 16068 31300 16096
rect 30668 16028 30696 16068
rect 31294 16056 31300 16068
rect 31352 16096 31358 16108
rect 32493 16099 32551 16105
rect 31352 16068 31754 16096
rect 31352 16056 31358 16068
rect 29564 16000 30696 16028
rect 31726 16028 31754 16068
rect 32493 16065 32505 16099
rect 32539 16096 32551 16099
rect 33229 16099 33287 16105
rect 33229 16096 33241 16099
rect 32539 16068 33241 16096
rect 32539 16065 32551 16068
rect 32493 16059 32551 16065
rect 32968 16040 32996 16068
rect 33229 16065 33241 16068
rect 33275 16065 33287 16099
rect 33229 16059 33287 16065
rect 33321 16099 33379 16105
rect 33321 16065 33333 16099
rect 33367 16096 33379 16099
rect 33686 16096 33692 16108
rect 33367 16068 33692 16096
rect 33367 16065 33379 16068
rect 33321 16059 33379 16065
rect 33686 16056 33692 16068
rect 33744 16056 33750 16108
rect 34048 16099 34106 16105
rect 34048 16065 34060 16099
rect 34094 16096 34106 16099
rect 34422 16096 34428 16108
rect 34094 16068 34428 16096
rect 34094 16065 34106 16068
rect 34048 16059 34106 16065
rect 34422 16056 34428 16068
rect 34480 16056 34486 16108
rect 36170 16056 36176 16108
rect 36228 16056 36234 16108
rect 37093 16099 37151 16105
rect 36832 16068 37044 16096
rect 36832 16040 36860 16068
rect 32677 16031 32735 16037
rect 32677 16028 32689 16031
rect 31726 16000 32689 16028
rect 32677 15997 32689 16000
rect 32723 15997 32735 16031
rect 32677 15991 32735 15997
rect 32950 15988 32956 16040
rect 33008 15988 33014 16040
rect 33134 15988 33140 16040
rect 33192 15988 33198 16040
rect 33778 15988 33784 16040
rect 33836 15988 33842 16040
rect 35710 15988 35716 16040
rect 35768 16028 35774 16040
rect 35897 16031 35955 16037
rect 35897 16028 35909 16031
rect 35768 16000 35909 16028
rect 35768 15988 35774 16000
rect 35897 15997 35909 16000
rect 35943 15997 35955 16031
rect 35897 15991 35955 15997
rect 35986 15988 35992 16040
rect 36044 16037 36050 16040
rect 36044 16031 36093 16037
rect 36044 15997 36047 16031
rect 36081 15997 36093 16031
rect 36044 15991 36093 15997
rect 36044 15988 36050 15991
rect 36814 15988 36820 16040
rect 36872 15988 36878 16040
rect 36909 16031 36967 16037
rect 36909 15997 36921 16031
rect 36955 15997 36967 16031
rect 37016 16028 37044 16068
rect 37093 16065 37105 16099
rect 37139 16096 37151 16099
rect 37139 16068 37596 16096
rect 37139 16065 37151 16068
rect 37093 16059 37151 16065
rect 37568 16037 37596 16068
rect 37642 16056 37648 16108
rect 37700 16056 37706 16108
rect 38010 16056 38016 16108
rect 38068 16056 38074 16108
rect 38672 16105 38700 16136
rect 39108 16133 39120 16167
rect 39154 16164 39166 16167
rect 40696 16164 40724 16192
rect 39154 16136 40724 16164
rect 39154 16133 39166 16136
rect 39108 16127 39166 16133
rect 38657 16099 38715 16105
rect 38657 16065 38669 16099
rect 38703 16065 38715 16099
rect 38657 16059 38715 16065
rect 40773 16099 40831 16105
rect 40773 16065 40785 16099
rect 40819 16096 40831 16099
rect 43162 16096 43168 16108
rect 40819 16068 43168 16096
rect 40819 16065 40831 16068
rect 40773 16059 40831 16065
rect 43162 16056 43168 16068
rect 43220 16056 43226 16108
rect 43901 16099 43959 16105
rect 43901 16065 43913 16099
rect 43947 16096 43959 16099
rect 44269 16099 44327 16105
rect 44269 16096 44281 16099
rect 43947 16068 44281 16096
rect 43947 16065 43959 16068
rect 43901 16059 43959 16065
rect 44269 16065 44281 16068
rect 44315 16065 44327 16099
rect 45204 16096 45232 16192
rect 47302 16124 47308 16176
rect 47360 16124 47366 16176
rect 45462 16096 45468 16108
rect 45204 16068 45468 16096
rect 44269 16059 44327 16065
rect 45462 16056 45468 16068
rect 45520 16096 45526 16108
rect 45922 16105 45928 16108
rect 45649 16099 45707 16105
rect 45649 16096 45661 16099
rect 45520 16068 45661 16096
rect 45520 16056 45526 16068
rect 45649 16065 45661 16068
rect 45695 16065 45707 16099
rect 45649 16059 45707 16065
rect 45916 16059 45928 16105
rect 45922 16056 45928 16059
rect 45980 16056 45986 16108
rect 48222 16056 48228 16108
rect 48280 16056 48286 16108
rect 49528 16096 49556 16204
rect 50433 16201 50445 16235
rect 50479 16232 50491 16235
rect 50982 16232 50988 16244
rect 50479 16204 50988 16232
rect 50479 16201 50491 16204
rect 50433 16195 50491 16201
rect 50982 16192 50988 16204
rect 51040 16192 51046 16244
rect 52546 16192 52552 16244
rect 52604 16232 52610 16244
rect 53193 16235 53251 16241
rect 53193 16232 53205 16235
rect 52604 16204 53205 16232
rect 52604 16192 52610 16204
rect 53193 16201 53205 16204
rect 53239 16201 53251 16235
rect 53193 16195 53251 16201
rect 53558 16192 53564 16244
rect 53616 16192 53622 16244
rect 54570 16192 54576 16244
rect 54628 16192 54634 16244
rect 55306 16192 55312 16244
rect 55364 16232 55370 16244
rect 55861 16235 55919 16241
rect 55861 16232 55873 16235
rect 55364 16204 55873 16232
rect 55364 16192 55370 16204
rect 55861 16201 55873 16204
rect 55907 16232 55919 16235
rect 56502 16232 56508 16244
rect 55907 16204 56508 16232
rect 55907 16201 55919 16204
rect 55861 16195 55919 16201
rect 56502 16192 56508 16204
rect 56560 16192 56566 16244
rect 57514 16192 57520 16244
rect 57572 16192 57578 16244
rect 57606 16192 57612 16244
rect 57664 16232 57670 16244
rect 57664 16204 58480 16232
rect 57664 16192 57670 16204
rect 51568 16167 51626 16173
rect 51568 16133 51580 16167
rect 51614 16164 51626 16167
rect 51905 16167 51963 16173
rect 51905 16164 51917 16167
rect 51614 16136 51917 16164
rect 51614 16133 51626 16136
rect 51568 16127 51626 16133
rect 51905 16133 51917 16136
rect 51951 16133 51963 16167
rect 51905 16127 51963 16133
rect 53006 16124 53012 16176
rect 53064 16164 53070 16176
rect 53101 16167 53159 16173
rect 53101 16164 53113 16167
rect 53064 16136 53113 16164
rect 53064 16124 53070 16136
rect 53101 16133 53113 16136
rect 53147 16164 53159 16167
rect 53576 16164 53604 16192
rect 54588 16164 54616 16192
rect 56312 16167 56370 16173
rect 53147 16136 53604 16164
rect 54128 16136 56088 16164
rect 53147 16133 53159 16136
rect 53101 16127 53159 16133
rect 50065 16099 50123 16105
rect 50065 16096 50077 16099
rect 49528 16068 50077 16096
rect 50065 16065 50077 16068
rect 50111 16065 50123 16099
rect 50065 16059 50123 16065
rect 51718 16056 51724 16108
rect 51776 16096 51782 16108
rect 51813 16099 51871 16105
rect 51813 16096 51825 16099
rect 51776 16068 51825 16096
rect 51776 16056 51782 16068
rect 51813 16065 51825 16068
rect 51859 16065 51871 16099
rect 51813 16059 51871 16065
rect 52730 16056 52736 16108
rect 52788 16056 52794 16108
rect 54128 16105 54156 16136
rect 54386 16105 54392 16108
rect 54113 16099 54171 16105
rect 54113 16065 54125 16099
rect 54159 16065 54171 16099
rect 54113 16059 54171 16065
rect 54380 16059 54392 16105
rect 54386 16056 54392 16059
rect 54444 16056 54450 16108
rect 56060 16105 56088 16136
rect 56312 16133 56324 16167
rect 56358 16164 56370 16167
rect 57330 16164 57336 16176
rect 56358 16136 57336 16164
rect 56358 16133 56370 16136
rect 56312 16127 56370 16133
rect 57330 16124 57336 16136
rect 57388 16124 57394 16176
rect 57532 16164 57560 16192
rect 57885 16167 57943 16173
rect 57885 16164 57897 16167
rect 57532 16136 57897 16164
rect 57885 16133 57897 16136
rect 57931 16133 57943 16167
rect 57885 16127 57943 16133
rect 58452 16105 58480 16204
rect 56045 16099 56103 16105
rect 56045 16065 56057 16099
rect 56091 16065 56103 16099
rect 56045 16059 56103 16065
rect 58437 16099 58495 16105
rect 58437 16065 58449 16099
rect 58483 16065 58495 16099
rect 58437 16059 58495 16065
rect 37369 16031 37427 16037
rect 37369 16028 37381 16031
rect 37016 16000 37381 16028
rect 36909 15991 36967 15997
rect 37369 15997 37381 16000
rect 37415 15997 37427 16031
rect 37369 15991 37427 15997
rect 37553 16031 37611 16037
rect 37553 15997 37565 16031
rect 37599 16028 37611 16031
rect 38028 16028 38056 16056
rect 37599 16000 38056 16028
rect 38841 16031 38899 16037
rect 37599 15997 37611 16000
rect 37553 15991 37611 15997
rect 38841 15997 38853 16031
rect 38887 15997 38899 16031
rect 40497 16031 40555 16037
rect 40497 16028 40509 16031
rect 38841 15991 38899 15997
rect 39868 16000 40509 16028
rect 32582 15920 32588 15972
rect 32640 15960 32646 15972
rect 33796 15960 33824 15988
rect 35434 15960 35440 15972
rect 32640 15932 33824 15960
rect 35084 15932 35440 15960
rect 32640 15920 32646 15932
rect 26988 15864 28028 15892
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 28353 15895 28411 15901
rect 28353 15892 28365 15895
rect 28224 15864 28365 15892
rect 28224 15852 28230 15864
rect 28353 15861 28365 15864
rect 28399 15861 28411 15895
rect 28353 15855 28411 15861
rect 28902 15852 28908 15904
rect 28960 15892 28966 15904
rect 30466 15892 30472 15904
rect 28960 15864 30472 15892
rect 28960 15852 28966 15864
rect 30466 15852 30472 15864
rect 30524 15892 30530 15904
rect 31570 15892 31576 15904
rect 30524 15864 31576 15892
rect 30524 15852 30530 15864
rect 31570 15852 31576 15864
rect 31628 15892 31634 15904
rect 35084 15892 35112 15932
rect 35434 15920 35440 15932
rect 35492 15920 35498 15972
rect 36354 15920 36360 15972
rect 36412 15960 36418 15972
rect 36449 15963 36507 15969
rect 36449 15960 36461 15963
rect 36412 15932 36461 15960
rect 36412 15920 36418 15932
rect 36449 15929 36461 15932
rect 36495 15929 36507 15963
rect 36924 15960 36952 15991
rect 38105 15963 38163 15969
rect 38105 15960 38117 15963
rect 36924 15932 38117 15960
rect 36449 15923 36507 15929
rect 37568 15904 37596 15932
rect 38105 15929 38117 15932
rect 38151 15929 38163 15963
rect 38105 15923 38163 15929
rect 31628 15864 35112 15892
rect 31628 15852 31634 15864
rect 35158 15852 35164 15904
rect 35216 15852 35222 15904
rect 35253 15895 35311 15901
rect 35253 15861 35265 15895
rect 35299 15892 35311 15895
rect 36538 15892 36544 15904
rect 35299 15864 36544 15892
rect 35299 15861 35311 15864
rect 35253 15855 35311 15861
rect 36538 15852 36544 15864
rect 36596 15852 36602 15904
rect 37550 15852 37556 15904
rect 37608 15852 37614 15904
rect 38856 15892 38884 15991
rect 39022 15892 39028 15904
rect 38856 15864 39028 15892
rect 39022 15852 39028 15864
rect 39080 15852 39086 15904
rect 39574 15852 39580 15904
rect 39632 15892 39638 15904
rect 39868 15892 39896 16000
rect 40497 15997 40509 16000
rect 40543 15997 40555 16031
rect 40497 15991 40555 15997
rect 40681 16031 40739 16037
rect 40681 15997 40693 16031
rect 40727 16028 40739 16031
rect 41598 16028 41604 16040
rect 40727 16000 41604 16028
rect 40727 15997 40739 16000
rect 40681 15991 40739 15997
rect 41598 15988 41604 16000
rect 41656 15988 41662 16040
rect 41785 16031 41843 16037
rect 41785 15997 41797 16031
rect 41831 15997 41843 16031
rect 41785 15991 41843 15997
rect 41141 15963 41199 15969
rect 41141 15929 41153 15963
rect 41187 15960 41199 15963
rect 41800 15960 41828 15991
rect 41966 15988 41972 16040
rect 42024 16028 42030 16040
rect 42429 16031 42487 16037
rect 42429 16028 42441 16031
rect 42024 16000 42441 16028
rect 42024 15988 42030 16000
rect 42429 15997 42441 16000
rect 42475 15997 42487 16031
rect 42429 15991 42487 15997
rect 42794 15988 42800 16040
rect 42852 16028 42858 16040
rect 42981 16031 43039 16037
rect 42981 16028 42993 16031
rect 42852 16000 42993 16028
rect 42852 15988 42858 16000
rect 42981 15997 42993 16000
rect 43027 15997 43039 16031
rect 43993 16031 44051 16037
rect 43993 16028 44005 16031
rect 42981 15991 43039 15997
rect 43088 16000 44005 16028
rect 41187 15932 41828 15960
rect 41187 15929 41199 15932
rect 41141 15923 41199 15929
rect 42334 15920 42340 15972
rect 42392 15960 42398 15972
rect 43088 15960 43116 16000
rect 43993 15997 44005 16000
rect 44039 16028 44051 16031
rect 44082 16028 44088 16040
rect 44039 16000 44088 16028
rect 44039 15997 44051 16000
rect 43993 15991 44051 15997
rect 44082 15988 44088 16000
rect 44140 15988 44146 16040
rect 44174 15988 44180 16040
rect 44232 15988 44238 16040
rect 44913 16031 44971 16037
rect 44913 15997 44925 16031
rect 44959 16028 44971 16031
rect 45002 16028 45008 16040
rect 44959 16000 45008 16028
rect 44959 15997 44971 16000
rect 44913 15991 44971 15997
rect 45002 15988 45008 16000
rect 45060 15988 45066 16040
rect 48406 16037 48412 16040
rect 48384 16031 48412 16037
rect 48384 15997 48396 16031
rect 48384 15991 48412 15997
rect 48406 15988 48412 15991
rect 48464 15988 48470 16040
rect 48501 16031 48559 16037
rect 48501 15997 48513 16031
rect 48547 16028 48559 16031
rect 49237 16031 49295 16037
rect 48547 16000 48912 16028
rect 48547 15997 48559 16000
rect 48501 15991 48559 15997
rect 42392 15932 43116 15960
rect 43441 15963 43499 15969
rect 42392 15920 42398 15932
rect 43441 15929 43453 15963
rect 43487 15960 43499 15963
rect 44192 15960 44220 15988
rect 48884 15972 48912 16000
rect 49237 15997 49249 16031
rect 49283 16028 49295 16031
rect 49326 16028 49332 16040
rect 49283 16000 49332 16028
rect 49283 15997 49295 16000
rect 49237 15991 49295 15997
rect 49326 15988 49332 16000
rect 49384 15988 49390 16040
rect 49418 15988 49424 16040
rect 49476 15988 49482 16040
rect 52549 16031 52607 16037
rect 52549 15997 52561 16031
rect 52595 15997 52607 16031
rect 52748 16028 52776 16056
rect 53285 16031 53343 16037
rect 53285 16028 53297 16031
rect 52748 16000 53297 16028
rect 52549 15991 52607 15997
rect 53285 15997 53297 16000
rect 53331 16028 53343 16031
rect 53745 16031 53803 16037
rect 53745 16028 53757 16031
rect 53331 16000 53757 16028
rect 53331 15997 53343 16000
rect 53285 15991 53343 15997
rect 53745 15997 53757 16000
rect 53791 15997 53803 16031
rect 53745 15991 53803 15997
rect 43487 15932 44220 15960
rect 43487 15929 43499 15932
rect 43441 15923 43499 15929
rect 48682 15920 48688 15972
rect 48740 15960 48746 15972
rect 48777 15963 48835 15969
rect 48777 15960 48789 15963
rect 48740 15932 48789 15960
rect 48740 15920 48746 15932
rect 48777 15929 48789 15932
rect 48823 15929 48835 15963
rect 48777 15923 48835 15929
rect 48866 15920 48872 15972
rect 48924 15960 48930 15972
rect 49513 15963 49571 15969
rect 49513 15960 49525 15963
rect 48924 15932 49525 15960
rect 48924 15920 48930 15932
rect 49513 15929 49525 15932
rect 49559 15929 49571 15963
rect 52564 15960 52592 15991
rect 58066 15988 58072 16040
rect 58124 15988 58130 16040
rect 52733 15963 52791 15969
rect 52733 15960 52745 15963
rect 52564 15932 52745 15960
rect 49513 15923 49571 15929
rect 52733 15929 52745 15932
rect 52779 15929 52791 15963
rect 57425 15963 57483 15969
rect 52733 15923 52791 15929
rect 55048 15932 55904 15960
rect 39632 15864 39896 15892
rect 39632 15852 39638 15864
rect 40218 15852 40224 15904
rect 40276 15852 40282 15904
rect 41230 15852 41236 15904
rect 41288 15852 41294 15904
rect 42150 15852 42156 15904
rect 42208 15852 42214 15904
rect 47026 15852 47032 15904
rect 47084 15852 47090 15904
rect 47581 15895 47639 15901
rect 47581 15861 47593 15895
rect 47627 15892 47639 15895
rect 49786 15892 49792 15904
rect 47627 15864 49792 15892
rect 47627 15861 47639 15864
rect 47581 15855 47639 15861
rect 49786 15852 49792 15864
rect 49844 15852 49850 15904
rect 52362 15852 52368 15904
rect 52420 15892 52426 15904
rect 55048 15892 55076 15932
rect 52420 15864 55076 15892
rect 52420 15852 52426 15864
rect 55490 15852 55496 15904
rect 55548 15852 55554 15904
rect 55876 15892 55904 15932
rect 57425 15929 57437 15963
rect 57471 15960 57483 15963
rect 58084 15960 58112 15988
rect 57471 15932 58112 15960
rect 57471 15929 57483 15932
rect 57425 15923 57483 15929
rect 56318 15892 56324 15904
rect 55876 15864 56324 15892
rect 56318 15852 56324 15864
rect 56376 15852 56382 15904
rect 1104 15802 58880 15824
rect 1104 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 22616 15802
rect 22668 15750 22680 15802
rect 22732 15750 22744 15802
rect 22796 15750 22808 15802
rect 22860 15750 22872 15802
rect 22924 15750 37060 15802
rect 37112 15750 37124 15802
rect 37176 15750 37188 15802
rect 37240 15750 37252 15802
rect 37304 15750 37316 15802
rect 37368 15750 51504 15802
rect 51556 15750 51568 15802
rect 51620 15750 51632 15802
rect 51684 15750 51696 15802
rect 51748 15750 51760 15802
rect 51812 15750 58880 15802
rect 1104 15728 58880 15750
rect 3237 15691 3295 15697
rect 3237 15657 3249 15691
rect 3283 15688 3295 15691
rect 3510 15688 3516 15700
rect 3283 15660 3516 15688
rect 3283 15657 3295 15660
rect 3237 15651 3295 15657
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 3973 15691 4031 15697
rect 3973 15657 3985 15691
rect 4019 15688 4031 15691
rect 4801 15691 4859 15697
rect 4019 15660 4752 15688
rect 4019 15657 4031 15660
rect 3973 15651 4031 15657
rect 3418 15580 3424 15632
rect 3476 15620 3482 15632
rect 4249 15623 4307 15629
rect 4249 15620 4261 15623
rect 3476 15592 4261 15620
rect 3476 15580 3482 15592
rect 4249 15589 4261 15592
rect 4295 15589 4307 15623
rect 4249 15583 4307 15589
rect 4341 15623 4399 15629
rect 4341 15589 4353 15623
rect 4387 15620 4399 15623
rect 4522 15620 4528 15632
rect 4387 15592 4528 15620
rect 4387 15589 4399 15592
rect 4341 15583 4399 15589
rect 4522 15580 4528 15592
rect 4580 15580 4586 15632
rect 4724 15620 4752 15660
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5350 15688 5356 15700
rect 4847 15660 5356 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5534 15648 5540 15700
rect 5592 15648 5598 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 7466 15688 7472 15700
rect 6604 15660 7472 15688
rect 6604 15648 6610 15660
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10870 15688 10876 15700
rect 10459 15660 10876 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15688 13507 15691
rect 13722 15688 13728 15700
rect 13495 15660 13728 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15197 15691 15255 15697
rect 15197 15688 15209 15691
rect 14884 15660 15209 15688
rect 14884 15648 14890 15660
rect 15197 15657 15209 15660
rect 15243 15657 15255 15691
rect 15197 15651 15255 15657
rect 15746 15648 15752 15700
rect 15804 15648 15810 15700
rect 15930 15648 15936 15700
rect 15988 15648 15994 15700
rect 16574 15648 16580 15700
rect 16632 15648 16638 15700
rect 17497 15691 17555 15697
rect 17497 15657 17509 15691
rect 17543 15688 17555 15691
rect 17862 15688 17868 15700
rect 17543 15660 17868 15688
rect 17543 15657 17555 15660
rect 17497 15651 17555 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 21082 15648 21088 15700
rect 21140 15688 21146 15700
rect 21266 15688 21272 15700
rect 21140 15660 21272 15688
rect 21140 15648 21146 15660
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 24121 15691 24179 15697
rect 24121 15657 24133 15691
rect 24167 15688 24179 15691
rect 24302 15688 24308 15700
rect 24167 15660 24308 15688
rect 24167 15657 24179 15660
rect 24121 15651 24179 15657
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 25958 15648 25964 15700
rect 26016 15648 26022 15700
rect 26326 15648 26332 15700
rect 26384 15688 26390 15700
rect 26697 15691 26755 15697
rect 26697 15688 26709 15691
rect 26384 15660 26709 15688
rect 26384 15648 26390 15660
rect 26697 15657 26709 15660
rect 26743 15657 26755 15691
rect 26697 15651 26755 15657
rect 26786 15648 26792 15700
rect 26844 15648 26850 15700
rect 28537 15691 28595 15697
rect 28537 15657 28549 15691
rect 28583 15688 28595 15691
rect 28718 15688 28724 15700
rect 28583 15660 28724 15688
rect 28583 15657 28595 15660
rect 28537 15651 28595 15657
rect 28718 15648 28724 15660
rect 28776 15648 28782 15700
rect 28902 15648 28908 15700
rect 28960 15648 28966 15700
rect 29270 15688 29276 15700
rect 29196 15660 29276 15688
rect 6454 15620 6460 15632
rect 4724 15592 6132 15620
rect 5445 15555 5503 15561
rect 2976 15524 4200 15552
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 2685 15487 2743 15493
rect 2685 15484 2697 15487
rect 2648 15456 2697 15484
rect 2648 15444 2654 15456
rect 2685 15453 2697 15456
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 2866 15376 2872 15428
rect 2924 15376 2930 15428
rect 2976 15425 3004 15524
rect 4172 15493 4200 15524
rect 4356 15524 4936 15552
rect 4356 15496 4384 15524
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 4157 15487 4215 15493
rect 3099 15456 4108 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 2961 15419 3019 15425
rect 2961 15385 2973 15419
rect 3007 15385 3019 15419
rect 2961 15379 3019 15385
rect 4080 15348 4108 15456
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4246 15484 4252 15496
rect 4203 15456 4252 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 4338 15444 4344 15496
rect 4396 15444 4402 15496
rect 4430 15444 4436 15496
rect 4488 15444 4494 15496
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 4632 15416 4660 15447
rect 4706 15444 4712 15496
rect 4764 15444 4770 15496
rect 4908 15493 4936 15524
rect 5445 15521 5457 15555
rect 5491 15552 5503 15555
rect 5491 15524 6040 15552
rect 5491 15521 5503 15524
rect 5445 15515 5503 15521
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 5859 15456 5948 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 5166 15416 5172 15428
rect 4632 15388 5172 15416
rect 5166 15376 5172 15388
rect 5224 15376 5230 15428
rect 5534 15376 5540 15428
rect 5592 15376 5598 15428
rect 4614 15348 4620 15360
rect 4080 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5718 15308 5724 15360
rect 5776 15308 5782 15360
rect 5920 15357 5948 15456
rect 6012 15416 6040 15524
rect 6104 15496 6132 15592
rect 6288 15592 6460 15620
rect 6288 15561 6316 15592
rect 6454 15580 6460 15592
rect 6512 15620 6518 15632
rect 7374 15620 7380 15632
rect 6512 15592 7380 15620
rect 6512 15580 6518 15592
rect 7374 15580 7380 15592
rect 7432 15580 7438 15632
rect 9214 15580 9220 15632
rect 9272 15580 9278 15632
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 6822 15512 6828 15564
rect 6880 15552 6886 15564
rect 10321 15555 10379 15561
rect 6880 15524 8984 15552
rect 6880 15512 6886 15524
rect 6086 15444 6092 15496
rect 6144 15444 6150 15496
rect 6730 15484 6736 15496
rect 6380 15456 6736 15484
rect 6380 15425 6408 15456
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 6365 15419 6423 15425
rect 6365 15416 6377 15419
rect 6012 15388 6377 15416
rect 6365 15385 6377 15388
rect 6411 15385 6423 15419
rect 6365 15379 6423 15385
rect 6546 15376 6552 15428
rect 6604 15425 6610 15428
rect 6604 15419 6639 15425
rect 6627 15416 6639 15419
rect 6840 15416 6868 15512
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15484 6975 15487
rect 7006 15484 7012 15496
rect 6963 15456 7012 15484
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 8956 15493 8984 15524
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10410 15552 10416 15564
rect 10367 15524 10416 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10410 15512 10416 15524
rect 10468 15552 10474 15564
rect 15764 15561 15792 15648
rect 15948 15561 15976 15648
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 10468 15524 10977 15552
rect 10468 15512 10474 15524
rect 10965 15521 10977 15524
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 16758 15512 16764 15564
rect 16816 15552 16822 15564
rect 16853 15555 16911 15561
rect 16853 15552 16865 15555
rect 16816 15524 16865 15552
rect 16816 15512 16822 15524
rect 16853 15521 16865 15524
rect 16899 15521 16911 15555
rect 16853 15515 16911 15521
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15552 17095 15555
rect 17770 15552 17776 15564
rect 17083 15524 17776 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 26605 15555 26663 15561
rect 26605 15521 26617 15555
rect 26651 15552 26663 15555
rect 26804 15552 26832 15648
rect 28920 15620 28948 15648
rect 28000 15592 28948 15620
rect 26651 15524 26832 15552
rect 26651 15521 26663 15524
rect 26605 15515 26663 15521
rect 26878 15512 26884 15564
rect 26936 15552 26942 15564
rect 28000 15561 28028 15592
rect 29196 15561 29224 15660
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 30374 15648 30380 15700
rect 30432 15688 30438 15700
rect 30432 15660 32628 15688
rect 30432 15648 30438 15660
rect 29546 15620 29552 15632
rect 29288 15592 29552 15620
rect 27249 15555 27307 15561
rect 27249 15552 27261 15555
rect 26936 15524 27261 15552
rect 26936 15512 26942 15524
rect 27249 15521 27261 15524
rect 27295 15521 27307 15555
rect 27249 15515 27307 15521
rect 27985 15555 28043 15561
rect 27985 15521 27997 15555
rect 28031 15521 28043 15555
rect 29181 15555 29239 15561
rect 29181 15552 29193 15555
rect 27985 15515 28043 15521
rect 28092 15524 29193 15552
rect 7653 15487 7711 15493
rect 7653 15484 7665 15487
rect 7248 15456 7665 15484
rect 7248 15444 7254 15456
rect 7653 15453 7665 15456
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9033 15487 9091 15493
rect 9033 15453 9045 15487
rect 9079 15484 9091 15487
rect 9490 15484 9496 15496
rect 9079 15456 9496 15484
rect 9079 15453 9091 15456
rect 9033 15447 9091 15453
rect 9490 15444 9496 15456
rect 9548 15444 9554 15496
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11756 15456 11805 15484
rect 11756 15444 11762 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12066 15444 12072 15496
rect 12124 15444 12130 15496
rect 12342 15493 12348 15496
rect 12336 15447 12348 15493
rect 12342 15444 12348 15447
rect 12400 15444 12406 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 18104 15456 18613 15484
rect 18104 15444 18110 15456
rect 18601 15453 18613 15456
rect 18647 15484 18659 15487
rect 18969 15487 19027 15493
rect 18969 15484 18981 15487
rect 18647 15456 18981 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 18969 15453 18981 15456
rect 19015 15484 19027 15487
rect 19242 15484 19248 15496
rect 19015 15456 19248 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 21269 15487 21327 15493
rect 21269 15453 21281 15487
rect 21315 15484 21327 15487
rect 21358 15484 21364 15496
rect 21315 15456 21364 15484
rect 21315 15453 21327 15456
rect 21269 15447 21327 15453
rect 21358 15444 21364 15456
rect 21416 15484 21422 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 21416 15456 22753 15484
rect 21416 15444 21422 15456
rect 22741 15453 22753 15456
rect 22787 15484 22799 15487
rect 23474 15484 23480 15496
rect 22787 15456 23480 15484
rect 22787 15453 22799 15456
rect 22741 15447 22799 15453
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 27709 15487 27767 15493
rect 27709 15453 27721 15487
rect 27755 15484 27767 15487
rect 28092 15484 28120 15524
rect 29181 15521 29193 15524
rect 29227 15521 29239 15555
rect 29181 15515 29239 15521
rect 27755 15456 28120 15484
rect 28169 15487 28227 15493
rect 27755 15453 27767 15456
rect 27709 15447 27767 15453
rect 28169 15453 28181 15487
rect 28215 15484 28227 15487
rect 29288 15484 29316 15592
rect 29546 15580 29552 15592
rect 29604 15580 29610 15632
rect 31846 15512 31852 15564
rect 31904 15512 31910 15564
rect 32490 15512 32496 15564
rect 32548 15512 32554 15564
rect 32600 15496 32628 15660
rect 33594 15648 33600 15700
rect 33652 15648 33658 15700
rect 35158 15648 35164 15700
rect 35216 15648 35222 15700
rect 37550 15648 37556 15700
rect 37608 15648 37614 15700
rect 38930 15648 38936 15700
rect 38988 15688 38994 15700
rect 39025 15691 39083 15697
rect 39025 15688 39037 15691
rect 38988 15660 39037 15688
rect 38988 15648 38994 15660
rect 39025 15657 39037 15660
rect 39071 15657 39083 15691
rect 39025 15651 39083 15657
rect 42518 15648 42524 15700
rect 42576 15648 42582 15700
rect 45462 15648 45468 15700
rect 45520 15688 45526 15700
rect 45925 15691 45983 15697
rect 45925 15688 45937 15691
rect 45520 15660 45937 15688
rect 45520 15648 45526 15660
rect 45925 15657 45937 15660
rect 45971 15657 45983 15691
rect 45925 15651 45983 15657
rect 47029 15691 47087 15697
rect 47029 15657 47041 15691
rect 47075 15688 47087 15691
rect 47670 15688 47676 15700
rect 47075 15660 47676 15688
rect 47075 15657 47087 15660
rect 47029 15651 47087 15657
rect 47670 15648 47676 15660
rect 47728 15648 47734 15700
rect 48130 15648 48136 15700
rect 48188 15648 48194 15700
rect 48866 15648 48872 15700
rect 48924 15648 48930 15700
rect 49050 15648 49056 15700
rect 49108 15648 49114 15700
rect 49234 15648 49240 15700
rect 49292 15648 49298 15700
rect 51445 15691 51503 15697
rect 51445 15657 51457 15691
rect 51491 15688 51503 15691
rect 51491 15660 52960 15688
rect 51491 15657 51503 15660
rect 51445 15651 51503 15657
rect 28215 15456 29316 15484
rect 29549 15487 29607 15493
rect 28215 15453 28227 15456
rect 28169 15447 28227 15453
rect 29549 15453 29561 15487
rect 29595 15453 29607 15487
rect 29549 15447 29607 15453
rect 30377 15487 30435 15493
rect 30377 15453 30389 15487
rect 30423 15484 30435 15487
rect 30466 15484 30472 15496
rect 30423 15456 30472 15484
rect 30423 15453 30435 15456
rect 30377 15447 30435 15453
rect 6627 15388 6868 15416
rect 6627 15385 6639 15388
rect 6604 15379 6639 15385
rect 6604 15376 6610 15379
rect 7374 15376 7380 15428
rect 7432 15376 7438 15428
rect 8481 15419 8539 15425
rect 8481 15385 8493 15419
rect 8527 15416 8539 15419
rect 8662 15416 8668 15428
rect 8527 15388 8668 15416
rect 8527 15385 8539 15388
rect 8481 15379 8539 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 9122 15376 9128 15428
rect 9180 15416 9186 15428
rect 9217 15419 9275 15425
rect 9217 15416 9229 15419
rect 9180 15388 9229 15416
rect 9180 15376 9186 15388
rect 9217 15385 9229 15388
rect 9263 15385 9275 15419
rect 12084 15416 12112 15444
rect 13725 15419 13783 15425
rect 13725 15416 13737 15419
rect 12084 15388 13737 15416
rect 9217 15379 9275 15385
rect 13725 15385 13737 15388
rect 13771 15416 13783 15419
rect 14274 15416 14280 15428
rect 13771 15388 14280 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 18230 15416 18236 15428
rect 17972 15388 18236 15416
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 6564 15348 6592 15376
rect 17972 15360 18000 15388
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 19512 15419 19570 15425
rect 19512 15385 19524 15419
rect 19558 15416 19570 15419
rect 19794 15416 19800 15428
rect 19558 15388 19800 15416
rect 19558 15385 19570 15388
rect 19512 15379 19570 15385
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 21536 15419 21594 15425
rect 21536 15385 21548 15419
rect 21582 15416 21594 15419
rect 21818 15416 21824 15428
rect 21582 15388 21824 15416
rect 21582 15385 21594 15388
rect 21536 15379 21594 15385
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 23008 15419 23066 15425
rect 23008 15385 23020 15419
rect 23054 15416 23066 15419
rect 23290 15416 23296 15428
rect 23054 15388 23296 15416
rect 23054 15385 23066 15388
rect 23008 15379 23066 15385
rect 23290 15376 23296 15388
rect 23348 15376 23354 15428
rect 28077 15419 28135 15425
rect 28077 15385 28089 15419
rect 28123 15416 28135 15419
rect 28997 15419 29055 15425
rect 28997 15416 29009 15419
rect 28123 15388 29009 15416
rect 28123 15385 28135 15388
rect 28077 15379 28135 15385
rect 28997 15385 29009 15388
rect 29043 15416 29055 15419
rect 29043 15388 29316 15416
rect 29043 15385 29055 15388
rect 28997 15379 29055 15385
rect 29288 15360 29316 15388
rect 29454 15376 29460 15428
rect 29512 15416 29518 15428
rect 29564 15416 29592 15447
rect 30466 15444 30472 15456
rect 30524 15444 30530 15496
rect 31294 15444 31300 15496
rect 31352 15444 31358 15496
rect 31386 15444 31392 15496
rect 31444 15493 31450 15496
rect 31444 15487 31493 15493
rect 31444 15453 31447 15487
rect 31481 15453 31493 15487
rect 31444 15447 31493 15453
rect 31444 15444 31450 15447
rect 31570 15444 31576 15496
rect 31628 15444 31634 15496
rect 32309 15487 32367 15493
rect 32309 15453 32321 15487
rect 32355 15453 32367 15487
rect 32309 15447 32367 15453
rect 29512 15388 29592 15416
rect 32324 15416 32352 15447
rect 32582 15444 32588 15496
rect 32640 15444 32646 15496
rect 32852 15487 32910 15493
rect 32852 15453 32864 15487
rect 32898 15484 32910 15487
rect 33612 15484 33640 15648
rect 35066 15580 35072 15632
rect 35124 15580 35130 15632
rect 35176 15620 35204 15648
rect 35176 15592 35572 15620
rect 35084 15552 35112 15580
rect 35544 15561 35572 15592
rect 36078 15580 36084 15632
rect 36136 15620 36142 15632
rect 36814 15620 36820 15632
rect 36136 15592 36820 15620
rect 36136 15580 36142 15592
rect 36814 15580 36820 15592
rect 36872 15620 36878 15632
rect 37001 15623 37059 15629
rect 37001 15620 37013 15623
rect 36872 15592 37013 15620
rect 36872 15580 36878 15592
rect 37001 15589 37013 15592
rect 37047 15589 37059 15623
rect 37001 15583 37059 15589
rect 35253 15555 35311 15561
rect 35253 15552 35265 15555
rect 35084 15524 35265 15552
rect 35253 15521 35265 15524
rect 35299 15521 35311 15555
rect 35253 15515 35311 15521
rect 35529 15555 35587 15561
rect 35529 15521 35541 15555
rect 35575 15521 35587 15555
rect 35529 15515 35587 15521
rect 35802 15512 35808 15564
rect 35860 15552 35866 15564
rect 36354 15552 36360 15564
rect 35860 15524 36360 15552
rect 35860 15512 35866 15524
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 36630 15512 36636 15564
rect 36688 15552 36694 15564
rect 37277 15555 37335 15561
rect 37277 15552 37289 15555
rect 36688 15524 37289 15552
rect 36688 15512 36694 15524
rect 37277 15521 37289 15524
rect 37323 15521 37335 15555
rect 37277 15515 37335 15521
rect 32898 15456 33640 15484
rect 32898 15453 32910 15456
rect 32852 15447 32910 15453
rect 33686 15444 33692 15496
rect 33744 15444 33750 15496
rect 34330 15444 34336 15496
rect 34388 15444 34394 15496
rect 35069 15487 35127 15493
rect 35069 15453 35081 15487
rect 35115 15484 35127 15487
rect 35986 15484 35992 15496
rect 35115 15456 35992 15484
rect 35115 15453 35127 15456
rect 35069 15447 35127 15453
rect 35986 15444 35992 15456
rect 36044 15484 36050 15496
rect 37568 15493 37596 15648
rect 37921 15623 37979 15629
rect 37921 15589 37933 15623
rect 37967 15589 37979 15623
rect 42536 15620 42564 15648
rect 37921 15583 37979 15589
rect 41524 15592 42564 15620
rect 43993 15623 44051 15629
rect 37936 15552 37964 15583
rect 41524 15561 41552 15592
rect 43993 15589 44005 15623
rect 44039 15620 44051 15623
rect 48884 15620 48912 15648
rect 44039 15592 45600 15620
rect 44039 15589 44051 15592
rect 43993 15583 44051 15589
rect 38381 15555 38439 15561
rect 38381 15552 38393 15555
rect 37936 15524 38393 15552
rect 38381 15521 38393 15524
rect 38427 15521 38439 15555
rect 38381 15515 38439 15521
rect 41509 15555 41567 15561
rect 41509 15521 41521 15555
rect 41555 15521 41567 15555
rect 41509 15515 41567 15521
rect 41693 15555 41751 15561
rect 41693 15521 41705 15555
rect 41739 15552 41751 15555
rect 41966 15552 41972 15564
rect 41739 15524 41972 15552
rect 41739 15521 41751 15524
rect 41693 15515 41751 15521
rect 41966 15512 41972 15524
rect 42024 15512 42030 15564
rect 42150 15512 42156 15564
rect 42208 15552 42214 15564
rect 42613 15555 42671 15561
rect 42613 15552 42625 15555
rect 42208 15524 42625 15552
rect 42208 15512 42214 15524
rect 42613 15521 42625 15524
rect 42659 15521 42671 15555
rect 42613 15515 42671 15521
rect 44729 15555 44787 15561
rect 44729 15521 44741 15555
rect 44775 15552 44787 15555
rect 44910 15552 44916 15564
rect 44775 15524 44916 15552
rect 44775 15521 44787 15524
rect 44729 15515 44787 15521
rect 44910 15512 44916 15524
rect 44968 15512 44974 15564
rect 45572 15561 45600 15592
rect 47504 15592 48912 15620
rect 45557 15555 45615 15561
rect 45557 15521 45569 15555
rect 45603 15521 45615 15555
rect 45557 15515 45615 15521
rect 46842 15512 46848 15564
rect 46900 15512 46906 15564
rect 47504 15561 47532 15592
rect 47489 15555 47547 15561
rect 47489 15521 47501 15555
rect 47535 15521 47547 15555
rect 47489 15515 47547 15521
rect 47578 15512 47584 15564
rect 47636 15512 47642 15564
rect 48498 15512 48504 15564
rect 48556 15512 48562 15564
rect 49252 15561 49280 15648
rect 52932 15629 52960 15660
rect 55490 15648 55496 15700
rect 55548 15648 55554 15700
rect 55953 15691 56011 15697
rect 55953 15657 55965 15691
rect 55999 15688 56011 15691
rect 56410 15688 56416 15700
rect 55999 15660 56416 15688
rect 55999 15657 56011 15660
rect 55953 15651 56011 15657
rect 52917 15623 52975 15629
rect 52917 15589 52929 15623
rect 52963 15620 52975 15623
rect 55306 15620 55312 15632
rect 52963 15592 55312 15620
rect 52963 15589 52975 15592
rect 52917 15583 52975 15589
rect 55306 15580 55312 15592
rect 55364 15580 55370 15632
rect 49237 15555 49295 15561
rect 49237 15521 49249 15555
rect 49283 15521 49295 15555
rect 49237 15515 49295 15521
rect 52362 15512 52368 15564
rect 52420 15512 52426 15564
rect 52638 15512 52644 15564
rect 52696 15512 52702 15564
rect 53377 15555 53435 15561
rect 53377 15521 53389 15555
rect 53423 15552 53435 15555
rect 53466 15552 53472 15564
rect 53423 15524 53472 15552
rect 53423 15521 53435 15524
rect 53377 15515 53435 15521
rect 53466 15512 53472 15524
rect 53524 15512 53530 15564
rect 53561 15555 53619 15561
rect 53561 15521 53573 15555
rect 53607 15552 53619 15555
rect 53650 15552 53656 15564
rect 53607 15524 53656 15552
rect 53607 15521 53619 15524
rect 53561 15515 53619 15521
rect 53650 15512 53656 15524
rect 53708 15512 53714 15564
rect 54478 15552 54484 15564
rect 54220 15524 54484 15552
rect 36173 15487 36231 15493
rect 36173 15484 36185 15487
rect 36044 15456 36185 15484
rect 36044 15444 36050 15456
rect 36173 15453 36185 15456
rect 36219 15453 36231 15487
rect 36173 15447 36231 15453
rect 37553 15487 37611 15493
rect 37553 15453 37565 15487
rect 37599 15453 37611 15487
rect 37553 15447 37611 15453
rect 39850 15444 39856 15496
rect 39908 15484 39914 15496
rect 39945 15487 40003 15493
rect 39945 15484 39957 15487
rect 39908 15456 39957 15484
rect 39908 15444 39914 15456
rect 39945 15453 39957 15456
rect 39991 15453 40003 15487
rect 39945 15447 40003 15453
rect 41598 15444 41604 15496
rect 41656 15484 41662 15496
rect 41785 15487 41843 15493
rect 41785 15484 41797 15487
rect 41656 15456 41797 15484
rect 41656 15444 41662 15456
rect 41785 15453 41797 15456
rect 41831 15484 41843 15487
rect 42058 15484 42064 15496
rect 41831 15456 42064 15484
rect 41831 15453 41843 15456
rect 41785 15447 41843 15453
rect 42058 15444 42064 15456
rect 42116 15484 42122 15496
rect 43714 15484 43720 15496
rect 42116 15456 43720 15484
rect 42116 15444 42122 15456
rect 43714 15444 43720 15456
rect 43772 15484 43778 15496
rect 44453 15487 44511 15493
rect 44453 15484 44465 15487
rect 43772 15456 44465 15484
rect 43772 15444 43778 15456
rect 44453 15453 44465 15456
rect 44499 15453 44511 15487
rect 44453 15447 44511 15453
rect 46658 15444 46664 15496
rect 46716 15484 46722 15496
rect 47397 15487 47455 15493
rect 47397 15484 47409 15487
rect 46716 15456 47409 15484
rect 46716 15444 46722 15456
rect 47397 15453 47409 15456
rect 47443 15484 47455 15487
rect 48593 15487 48651 15493
rect 47443 15456 48544 15484
rect 47443 15453 47455 15456
rect 47397 15447 47455 15453
rect 33704 15416 33732 15444
rect 32324 15388 33732 15416
rect 34348 15416 34376 15444
rect 35161 15419 35219 15425
rect 34348 15388 35112 15416
rect 29512 15376 29518 15388
rect 5951 15320 6592 15348
rect 6733 15351 6791 15357
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 6733 15317 6745 15351
rect 6779 15348 6791 15351
rect 7834 15348 7840 15360
rect 6779 15320 7840 15348
rect 6779 15317 6791 15320
rect 6733 15311 6791 15317
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10744 15320 10793 15348
rect 10744 15308 10750 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10781 15311 10839 15317
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 11241 15351 11299 15357
rect 11241 15348 11253 15351
rect 10919 15320 11253 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 11241 15317 11253 15320
rect 11287 15317 11299 15351
rect 11241 15311 11299 15317
rect 14550 15308 14556 15360
rect 14608 15348 14614 15360
rect 15013 15351 15071 15357
rect 15013 15348 15025 15351
rect 14608 15320 15025 15348
rect 14608 15308 14614 15320
rect 15013 15317 15025 15320
rect 15059 15348 15071 15351
rect 15562 15348 15568 15360
rect 15059 15320 15568 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 15838 15308 15844 15360
rect 15896 15348 15902 15360
rect 17129 15351 17187 15357
rect 17129 15348 17141 15351
rect 15896 15320 17141 15348
rect 15896 15308 15902 15320
rect 17129 15317 17141 15320
rect 17175 15348 17187 15351
rect 17954 15348 17960 15360
rect 17175 15320 17960 15348
rect 17175 15317 17187 15320
rect 17129 15311 17187 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 18141 15351 18199 15357
rect 18141 15317 18153 15351
rect 18187 15348 18199 15351
rect 18322 15348 18328 15360
rect 18187 15320 18328 15348
rect 18187 15317 18199 15320
rect 18141 15311 18199 15317
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 21266 15308 21272 15360
rect 21324 15348 21330 15360
rect 21726 15348 21732 15360
rect 21324 15320 21732 15348
rect 21324 15308 21330 15320
rect 21726 15308 21732 15320
rect 21784 15348 21790 15360
rect 22462 15348 22468 15360
rect 21784 15320 22468 15348
rect 21784 15308 21790 15320
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 22646 15308 22652 15360
rect 22704 15308 22710 15360
rect 23750 15308 23756 15360
rect 23808 15348 23814 15360
rect 24578 15348 24584 15360
rect 23808 15320 24584 15348
rect 23808 15308 23814 15320
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 28258 15308 28264 15360
rect 28316 15348 28322 15360
rect 28629 15351 28687 15357
rect 28629 15348 28641 15351
rect 28316 15320 28641 15348
rect 28316 15308 28322 15320
rect 28629 15317 28641 15320
rect 28675 15317 28687 15351
rect 28629 15311 28687 15317
rect 29086 15308 29092 15360
rect 29144 15308 29150 15360
rect 29270 15308 29276 15360
rect 29328 15308 29334 15360
rect 30653 15351 30711 15357
rect 30653 15317 30665 15351
rect 30699 15348 30711 15351
rect 31754 15348 31760 15360
rect 30699 15320 31760 15348
rect 30699 15317 30711 15320
rect 30653 15311 30711 15317
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 33962 15308 33968 15360
rect 34020 15308 34026 15360
rect 34333 15351 34391 15357
rect 34333 15317 34345 15351
rect 34379 15348 34391 15351
rect 34606 15348 34612 15360
rect 34379 15320 34612 15348
rect 34379 15317 34391 15320
rect 34333 15311 34391 15317
rect 34606 15308 34612 15320
rect 34664 15308 34670 15360
rect 34698 15308 34704 15360
rect 34756 15308 34762 15360
rect 35084 15348 35112 15388
rect 35161 15385 35173 15419
rect 35207 15416 35219 15419
rect 35250 15416 35256 15428
rect 35207 15388 35256 15416
rect 35207 15385 35219 15388
rect 35161 15379 35219 15385
rect 35250 15376 35256 15388
rect 35308 15416 35314 15428
rect 37461 15419 37519 15425
rect 37461 15416 37473 15419
rect 35308 15388 37473 15416
rect 35308 15376 35314 15388
rect 37461 15385 37473 15388
rect 37507 15416 37519 15419
rect 37642 15416 37648 15428
rect 37507 15388 37648 15416
rect 37507 15385 37519 15388
rect 37461 15379 37519 15385
rect 37642 15376 37648 15388
rect 37700 15376 37706 15428
rect 40212 15419 40270 15425
rect 40212 15385 40224 15419
rect 40258 15416 40270 15419
rect 40770 15416 40776 15428
rect 40258 15388 40776 15416
rect 40258 15385 40270 15388
rect 40212 15379 40270 15385
rect 40770 15376 40776 15388
rect 40828 15376 40834 15428
rect 42880 15419 42938 15425
rect 41340 15388 42840 15416
rect 36630 15348 36636 15360
rect 35084 15320 36636 15348
rect 36630 15308 36636 15320
rect 36688 15308 36694 15360
rect 38470 15308 38476 15360
rect 38528 15348 38534 15360
rect 39574 15348 39580 15360
rect 38528 15320 39580 15348
rect 38528 15308 38534 15320
rect 39574 15308 39580 15320
rect 39632 15308 39638 15360
rect 41340 15357 41368 15388
rect 42812 15360 42840 15388
rect 42880 15385 42892 15419
rect 42926 15416 42938 15419
rect 44726 15416 44732 15428
rect 42926 15388 44732 15416
rect 42926 15385 42938 15388
rect 42880 15379 42938 15385
rect 44726 15376 44732 15388
rect 44784 15376 44790 15428
rect 46569 15419 46627 15425
rect 46569 15385 46581 15419
rect 46615 15416 46627 15419
rect 48222 15416 48228 15428
rect 46615 15388 48228 15416
rect 46615 15385 46627 15388
rect 46569 15379 46627 15385
rect 48222 15376 48228 15388
rect 48280 15376 48286 15428
rect 48516 15416 48544 15456
rect 48593 15453 48605 15487
rect 48639 15484 48651 15487
rect 49418 15484 49424 15496
rect 48639 15456 49424 15484
rect 48639 15453 48651 15456
rect 48593 15447 48651 15453
rect 49418 15444 49424 15456
rect 49476 15484 49482 15496
rect 49789 15487 49847 15493
rect 49789 15484 49801 15487
rect 49476 15456 49801 15484
rect 49476 15444 49482 15456
rect 49789 15453 49801 15456
rect 49835 15453 49847 15487
rect 49789 15447 49847 15453
rect 50614 15444 50620 15496
rect 50672 15444 50678 15496
rect 52546 15493 52552 15496
rect 52524 15487 52552 15493
rect 52524 15453 52536 15487
rect 52524 15447 52552 15453
rect 52546 15444 52552 15447
rect 52604 15444 52610 15496
rect 54220 15493 54248 15524
rect 54478 15512 54484 15524
rect 54536 15552 54542 15564
rect 54941 15555 54999 15561
rect 54941 15552 54953 15555
rect 54536 15524 54953 15552
rect 54536 15512 54542 15524
rect 54941 15521 54953 15524
rect 54987 15521 54999 15555
rect 54941 15515 54999 15521
rect 55401 15555 55459 15561
rect 55401 15521 55413 15555
rect 55447 15552 55459 15555
rect 55508 15552 55536 15648
rect 55447 15524 55536 15552
rect 55447 15521 55459 15524
rect 55401 15515 55459 15521
rect 54205 15487 54263 15493
rect 54205 15484 54217 15487
rect 53944 15456 54217 15484
rect 48685 15419 48743 15425
rect 48685 15416 48697 15419
rect 48516 15388 48697 15416
rect 48685 15385 48697 15388
rect 48731 15416 48743 15419
rect 49234 15416 49240 15428
rect 48731 15388 49240 15416
rect 48731 15385 48743 15388
rect 48685 15379 48743 15385
rect 49234 15376 49240 15388
rect 49292 15416 49298 15428
rect 50632 15416 50660 15444
rect 53944 15428 53972 15456
rect 54205 15453 54217 15456
rect 54251 15453 54263 15487
rect 54205 15447 54263 15453
rect 54757 15487 54815 15493
rect 54757 15453 54769 15487
rect 54803 15484 54815 15487
rect 55968 15484 55996 15651
rect 56410 15648 56416 15660
rect 56468 15648 56474 15700
rect 56778 15648 56784 15700
rect 56836 15688 56842 15700
rect 56836 15660 57100 15688
rect 56836 15648 56842 15660
rect 56778 15512 56784 15564
rect 56836 15552 56842 15564
rect 57072 15561 57100 15660
rect 57882 15648 57888 15700
rect 57940 15648 57946 15700
rect 56873 15555 56931 15561
rect 56873 15552 56885 15555
rect 56836 15524 56885 15552
rect 56836 15512 56842 15524
rect 56873 15521 56885 15524
rect 56919 15521 56931 15555
rect 56873 15515 56931 15521
rect 57057 15555 57115 15561
rect 57057 15521 57069 15555
rect 57103 15521 57115 15555
rect 57057 15515 57115 15521
rect 58250 15512 58256 15564
rect 58308 15552 58314 15564
rect 58437 15555 58495 15561
rect 58437 15552 58449 15555
rect 58308 15524 58449 15552
rect 58308 15512 58314 15524
rect 58437 15521 58449 15524
rect 58483 15521 58495 15555
rect 58437 15515 58495 15521
rect 54803 15456 55996 15484
rect 56060 15456 57192 15484
rect 54803 15453 54815 15456
rect 54757 15447 54815 15453
rect 49292 15388 50660 15416
rect 49292 15376 49298 15388
rect 53926 15376 53932 15428
rect 53984 15376 53990 15428
rect 56060 15416 56088 15456
rect 57164 15425 57192 15456
rect 54312 15388 56088 15416
rect 57149 15419 57207 15425
rect 41325 15351 41383 15357
rect 41325 15317 41337 15351
rect 41371 15317 41383 15351
rect 41325 15311 41383 15317
rect 41966 15308 41972 15360
rect 42024 15348 42030 15360
rect 42153 15351 42211 15357
rect 42153 15348 42165 15351
rect 42024 15320 42165 15348
rect 42024 15308 42030 15320
rect 42153 15317 42165 15320
rect 42199 15317 42211 15351
rect 42153 15311 42211 15317
rect 42794 15308 42800 15360
rect 42852 15348 42858 15360
rect 43346 15348 43352 15360
rect 42852 15320 43352 15348
rect 42852 15308 42858 15320
rect 43346 15308 43352 15320
rect 43404 15308 43410 15360
rect 44085 15351 44143 15357
rect 44085 15317 44097 15351
rect 44131 15348 44143 15351
rect 44174 15348 44180 15360
rect 44131 15320 44180 15348
rect 44131 15317 44143 15320
rect 44085 15311 44143 15317
rect 44174 15308 44180 15320
rect 44232 15308 44238 15360
rect 44545 15351 44603 15357
rect 44545 15317 44557 15351
rect 44591 15348 44603 15351
rect 44634 15348 44640 15360
rect 44591 15320 44640 15348
rect 44591 15317 44603 15320
rect 44545 15311 44603 15317
rect 44634 15308 44640 15320
rect 44692 15348 44698 15360
rect 45005 15351 45063 15357
rect 45005 15348 45017 15351
rect 44692 15320 45017 15348
rect 44692 15308 44698 15320
rect 45005 15317 45017 15320
rect 45051 15317 45063 15351
rect 45005 15311 45063 15317
rect 46198 15308 46204 15360
rect 46256 15308 46262 15360
rect 47302 15308 47308 15360
rect 47360 15348 47366 15360
rect 48590 15348 48596 15360
rect 47360 15320 48596 15348
rect 47360 15308 47366 15320
rect 48590 15308 48596 15320
rect 48648 15308 48654 15360
rect 50154 15308 50160 15360
rect 50212 15348 50218 15360
rect 50341 15351 50399 15357
rect 50341 15348 50353 15351
rect 50212 15320 50353 15348
rect 50212 15308 50218 15320
rect 50341 15317 50353 15320
rect 50387 15317 50399 15351
rect 50341 15311 50399 15317
rect 51721 15351 51779 15357
rect 51721 15317 51733 15351
rect 51767 15348 51779 15351
rect 54312 15348 54340 15388
rect 57149 15385 57161 15419
rect 57195 15385 57207 15419
rect 57149 15379 57207 15385
rect 51767 15320 54340 15348
rect 54389 15351 54447 15357
rect 51767 15317 51779 15320
rect 51721 15311 51779 15317
rect 54389 15317 54401 15351
rect 54435 15348 54447 15351
rect 54662 15348 54668 15360
rect 54435 15320 54668 15348
rect 54435 15317 54447 15320
rect 54389 15311 54447 15317
rect 54662 15308 54668 15320
rect 54720 15308 54726 15360
rect 54849 15351 54907 15357
rect 54849 15317 54861 15351
rect 54895 15348 54907 15351
rect 55214 15348 55220 15360
rect 54895 15320 55220 15348
rect 54895 15317 54907 15320
rect 54849 15311 54907 15317
rect 55214 15308 55220 15320
rect 55272 15348 55278 15360
rect 55766 15348 55772 15360
rect 55272 15320 55772 15348
rect 55272 15308 55278 15320
rect 55766 15308 55772 15320
rect 55824 15308 55830 15360
rect 56689 15351 56747 15357
rect 56689 15317 56701 15351
rect 56735 15348 56747 15351
rect 56778 15348 56784 15360
rect 56735 15320 56784 15348
rect 56735 15317 56747 15320
rect 56689 15311 56747 15317
rect 56778 15308 56784 15320
rect 56836 15308 56842 15360
rect 57514 15308 57520 15360
rect 57572 15308 57578 15360
rect 1104 15258 59040 15280
rect 1104 15206 15394 15258
rect 15446 15206 15458 15258
rect 15510 15206 15522 15258
rect 15574 15206 15586 15258
rect 15638 15206 15650 15258
rect 15702 15206 29838 15258
rect 29890 15206 29902 15258
rect 29954 15206 29966 15258
rect 30018 15206 30030 15258
rect 30082 15206 30094 15258
rect 30146 15206 44282 15258
rect 44334 15206 44346 15258
rect 44398 15206 44410 15258
rect 44462 15206 44474 15258
rect 44526 15206 44538 15258
rect 44590 15206 58726 15258
rect 58778 15206 58790 15258
rect 58842 15206 58854 15258
rect 58906 15206 58918 15258
rect 58970 15206 58982 15258
rect 59034 15206 59040 15258
rect 1104 15184 59040 15206
rect 2590 15104 2596 15156
rect 2648 15104 2654 15156
rect 2685 15147 2743 15153
rect 2685 15113 2697 15147
rect 2731 15113 2743 15147
rect 2685 15107 2743 15113
rect 2700 15076 2728 15107
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2924 15116 2973 15144
rect 2924 15104 2930 15116
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 2961 15107 3019 15113
rect 3050 15104 3056 15156
rect 3108 15104 3114 15156
rect 3510 15104 3516 15156
rect 3568 15144 3574 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3568 15116 3893 15144
rect 3568 15104 3574 15116
rect 3881 15113 3893 15116
rect 3927 15113 3939 15147
rect 4338 15144 4344 15156
rect 3881 15107 3939 15113
rect 3988 15116 4344 15144
rect 3068 15076 3096 15104
rect 2700 15048 3096 15076
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3142 15008 3148 15020
rect 2915 14980 3148 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 3234 14968 3240 15020
rect 3292 15008 3298 15020
rect 3789 15011 3847 15017
rect 3292 14980 3740 15008
rect 3292 14968 3298 14980
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14940 2559 14943
rect 3326 14940 3332 14952
rect 2547 14912 3332 14940
rect 2547 14909 2559 14912
rect 2501 14903 2559 14909
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 3712 14940 3740 14980
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 3988 15008 4016 15116
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4614 15104 4620 15156
rect 4672 15104 4678 15156
rect 4706 15104 4712 15156
rect 4764 15104 4770 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5776 15116 5825 15144
rect 5776 15104 5782 15116
rect 5813 15113 5825 15116
rect 5859 15144 5871 15147
rect 5994 15144 6000 15156
rect 5859 15116 6000 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 9214 15144 9220 15156
rect 6144 15116 6776 15144
rect 6144 15104 6150 15116
rect 4724 15076 4752 15104
rect 4080 15048 4752 15076
rect 4080 15017 4108 15048
rect 6748 15020 6776 15116
rect 7944 15116 9220 15144
rect 3835 14980 4016 15008
rect 4065 15011 4123 15017
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 4065 14977 4077 15011
rect 4111 14977 4123 15011
rect 4709 15011 4767 15017
rect 4709 15008 4721 15011
rect 4065 14971 4123 14977
rect 4264 14980 4721 15008
rect 3878 14940 3884 14952
rect 3712 14912 3884 14940
rect 3421 14903 3479 14909
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 3436 14872 3464 14903
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 4264 14940 4292 14980
rect 4709 14977 4721 14980
rect 4755 14977 4767 15011
rect 4709 14971 4767 14977
rect 5534 14968 5540 15020
rect 5592 15008 5598 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5592 14980 6377 15008
rect 5592 14968 5598 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 3988 14912 4292 14940
rect 4341 14943 4399 14949
rect 2832 14844 3464 14872
rect 2832 14832 2838 14844
rect 3988 14816 4016 14912
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 5552 14940 5580 14968
rect 4387 14912 5580 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 5626 14900 5632 14952
rect 5684 14900 5690 14952
rect 6380 14940 6408 14971
rect 6546 14968 6552 15020
rect 6604 14968 6610 15020
rect 6730 14968 6736 15020
rect 6788 14968 6794 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 6840 14980 7573 15008
rect 6840 14940 6868 14980
rect 7561 14977 7573 14980
rect 7607 15008 7619 15011
rect 7653 15011 7711 15017
rect 7653 15008 7665 15011
rect 7607 14980 7665 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 7653 14977 7665 14980
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 7834 14968 7840 15020
rect 7892 14968 7898 15020
rect 7944 15017 7972 15116
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9582 15104 9588 15156
rect 9640 15104 9646 15156
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 12618 15144 12624 15156
rect 11563 15116 12624 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 14274 15104 14280 15156
rect 14332 15144 14338 15156
rect 15749 15147 15807 15153
rect 15749 15144 15761 15147
rect 14332 15116 15761 15144
rect 14332 15104 14338 15116
rect 15749 15113 15761 15116
rect 15795 15144 15807 15147
rect 16390 15144 16396 15156
rect 15795 15116 16396 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16390 15104 16396 15116
rect 16448 15144 16454 15156
rect 17957 15147 18015 15153
rect 17957 15144 17969 15147
rect 16448 15116 17969 15144
rect 16448 15104 16454 15116
rect 17957 15113 17969 15116
rect 18003 15144 18015 15147
rect 18046 15144 18052 15156
rect 18003 15116 18052 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 18046 15104 18052 15116
rect 18104 15144 18110 15156
rect 18874 15144 18880 15156
rect 18104 15116 18880 15144
rect 18104 15104 18110 15116
rect 18874 15104 18880 15116
rect 18932 15144 18938 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 18932 15116 19073 15144
rect 18932 15104 18938 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 19794 15104 19800 15156
rect 19852 15104 19858 15156
rect 21174 15104 21180 15156
rect 21232 15104 21238 15156
rect 23106 15104 23112 15156
rect 23164 15104 23170 15156
rect 29086 15104 29092 15156
rect 29144 15144 29150 15156
rect 30193 15147 30251 15153
rect 30193 15144 30205 15147
rect 29144 15116 30205 15144
rect 29144 15104 29150 15116
rect 30193 15113 30205 15116
rect 30239 15113 30251 15147
rect 30193 15107 30251 15113
rect 31941 15147 31999 15153
rect 31941 15113 31953 15147
rect 31987 15144 31999 15147
rect 32030 15144 32036 15156
rect 31987 15116 32036 15144
rect 31987 15113 31999 15116
rect 31941 15107 31999 15113
rect 32030 15104 32036 15116
rect 32088 15104 32094 15156
rect 33686 15104 33692 15156
rect 33744 15104 33750 15156
rect 34422 15104 34428 15156
rect 34480 15104 34486 15156
rect 40770 15104 40776 15156
rect 40828 15144 40834 15156
rect 41325 15147 41383 15153
rect 41325 15144 41337 15147
rect 40828 15116 41337 15144
rect 40828 15104 40834 15116
rect 41325 15113 41337 15116
rect 41371 15113 41383 15147
rect 43254 15144 43260 15156
rect 41325 15107 41383 15113
rect 41524 15116 43260 15144
rect 10128 15079 10186 15085
rect 10128 15045 10140 15079
rect 10174 15076 10186 15079
rect 10318 15076 10324 15088
rect 10174 15048 10324 15076
rect 10174 15045 10186 15048
rect 10128 15039 10186 15045
rect 10318 15036 10324 15048
rect 10376 15036 10382 15088
rect 13170 15036 13176 15088
rect 13228 15036 13234 15088
rect 16669 15079 16727 15085
rect 16669 15045 16681 15079
rect 16715 15076 16727 15079
rect 17862 15076 17868 15088
rect 16715 15048 17868 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 17862 15036 17868 15048
rect 17920 15076 17926 15088
rect 18782 15076 18788 15088
rect 17920 15048 18788 15076
rect 17920 15036 17926 15048
rect 18782 15036 18788 15048
rect 18840 15036 18846 15088
rect 28629 15079 28687 15085
rect 28629 15045 28641 15079
rect 28675 15076 28687 15079
rect 28966 15079 29024 15085
rect 28966 15076 28978 15079
rect 28675 15048 28978 15076
rect 28675 15045 28687 15048
rect 28629 15039 28687 15045
rect 28966 15045 28978 15048
rect 29012 15045 29024 15079
rect 28966 15039 29024 15045
rect 29178 15036 29184 15088
rect 29236 15076 29242 15088
rect 29454 15076 29460 15088
rect 29236 15048 29460 15076
rect 29236 15036 29242 15048
rect 29454 15036 29460 15048
rect 29512 15076 29518 15088
rect 31113 15079 31171 15085
rect 31113 15076 31125 15079
rect 29512 15048 31125 15076
rect 29512 15036 29518 15048
rect 31113 15045 31125 15048
rect 31159 15045 31171 15079
rect 32048 15076 32076 15104
rect 32125 15079 32183 15085
rect 32125 15076 32137 15079
rect 32048 15048 32137 15076
rect 31113 15039 31171 15045
rect 32125 15045 32137 15048
rect 32171 15045 32183 15079
rect 32125 15039 32183 15045
rect 40120 15079 40178 15085
rect 40120 15045 40132 15079
rect 40166 15076 40178 15079
rect 41230 15076 41236 15088
rect 40166 15048 41236 15076
rect 40166 15045 40178 15048
rect 40120 15039 40178 15045
rect 41230 15036 41236 15048
rect 41288 15036 41294 15088
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 13188 15008 13216 15036
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 8067 14980 9674 15008
rect 13188 14980 13369 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 6380 14912 6868 14940
rect 7006 14900 7012 14952
rect 7064 14900 7070 14952
rect 7282 14900 7288 14952
rect 7340 14900 7346 14952
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 7944 14912 8309 14940
rect 4249 14875 4307 14881
rect 4249 14841 4261 14875
rect 4295 14872 4307 14875
rect 5644 14872 5672 14900
rect 4295 14844 5672 14872
rect 6181 14875 6239 14881
rect 4295 14841 4307 14844
rect 4249 14835 4307 14841
rect 6181 14841 6193 14875
rect 6227 14872 6239 14875
rect 7024 14872 7052 14900
rect 7944 14881 7972 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 9646 14940 9674 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 15008 13875 15011
rect 14277 15011 14335 15017
rect 14277 15008 14289 15011
rect 13863 14980 14289 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 14277 14977 14289 14980
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14752 14980 16068 15008
rect 9858 14940 9864 14952
rect 9646 14912 9864 14940
rect 8297 14903 8355 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11664 14912 12173 14940
rect 11664 14900 11670 14912
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 12250 14900 12256 14952
rect 12308 14949 12314 14952
rect 12308 14943 12357 14949
rect 12308 14909 12311 14943
rect 12345 14909 12357 14943
rect 12308 14903 12357 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 13173 14943 13231 14949
rect 12483 14912 12664 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 12308 14900 12314 14903
rect 6227 14844 7052 14872
rect 7929 14875 7987 14881
rect 6227 14841 6239 14844
rect 6181 14835 6239 14841
rect 7929 14841 7941 14875
rect 7975 14841 7987 14875
rect 7929 14835 7987 14841
rect 3970 14764 3976 14816
rect 4028 14764 4034 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4433 14807 4491 14813
rect 4433 14804 4445 14807
rect 4120 14776 4445 14804
rect 4120 14764 4126 14776
rect 4433 14773 4445 14776
rect 4479 14773 4491 14807
rect 4433 14767 4491 14773
rect 4522 14764 4528 14816
rect 4580 14764 4586 14816
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 11241 14807 11299 14813
rect 11241 14773 11253 14807
rect 11287 14804 11299 14807
rect 11698 14804 11704 14816
rect 11287 14776 11704 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11698 14764 11704 14776
rect 11756 14804 11762 14816
rect 12636 14804 12664 14912
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13832 14940 13860 14971
rect 13219 14912 13860 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13906 14900 13912 14952
rect 13964 14900 13970 14952
rect 14090 14900 14096 14952
rect 14148 14940 14154 14952
rect 14752 14940 14780 14980
rect 16040 14952 16068 14980
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20036 14980 20361 15008
rect 20036 14968 20042 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20622 14968 20628 15020
rect 20680 14968 20686 15020
rect 22557 15011 22615 15017
rect 22557 14977 22569 15011
rect 22603 15008 22615 15011
rect 22646 15008 22652 15020
rect 22603 14980 22652 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 28258 15008 28264 15020
rect 28123 14980 28264 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 28534 14968 28540 15020
rect 28592 15008 28598 15020
rect 28721 15011 28779 15017
rect 28721 15008 28733 15011
rect 28592 14980 28733 15008
rect 28592 14968 28598 14980
rect 28721 14977 28733 14980
rect 28767 14977 28779 15011
rect 28721 14971 28779 14977
rect 30837 15011 30895 15017
rect 30837 14977 30849 15011
rect 30883 15008 30895 15011
rect 31570 15008 31576 15020
rect 30883 14980 31576 15008
rect 30883 14977 30895 14980
rect 30837 14971 30895 14977
rect 14148 14912 14780 14940
rect 14148 14900 14154 14912
rect 14826 14900 14832 14952
rect 14884 14900 14890 14952
rect 15010 14900 15016 14952
rect 15068 14940 15074 14952
rect 15068 14912 15332 14940
rect 15068 14900 15074 14912
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 15194 14872 15200 14884
rect 12768 14844 15200 14872
rect 12768 14832 12774 14844
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15304 14872 15332 14912
rect 16022 14900 16028 14952
rect 16080 14900 16086 14952
rect 20070 14872 20076 14884
rect 15304 14844 20076 14872
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 30101 14875 30159 14881
rect 30101 14841 30113 14875
rect 30147 14872 30159 14875
rect 30852 14872 30880 14971
rect 31570 14968 31576 14980
rect 31628 14968 31634 15020
rect 33962 14968 33968 15020
rect 34020 15008 34026 15020
rect 34241 15011 34299 15017
rect 34241 15008 34253 15011
rect 34020 14980 34253 15008
rect 34020 14968 34026 14980
rect 34241 14977 34253 14980
rect 34287 14977 34299 15011
rect 34241 14971 34299 14977
rect 34698 14968 34704 15020
rect 34756 15008 34762 15020
rect 34977 15011 35035 15017
rect 34977 15008 34989 15011
rect 34756 14980 34989 15008
rect 34756 14968 34762 14980
rect 34977 14977 34989 14980
rect 35023 14977 35035 15011
rect 34977 14971 35035 14977
rect 41524 14952 41552 15116
rect 43254 15104 43260 15116
rect 43312 15104 43318 15156
rect 44361 15147 44419 15153
rect 44361 15113 44373 15147
rect 44407 15144 44419 15147
rect 44726 15144 44732 15156
rect 44407 15116 44732 15144
rect 44407 15113 44419 15116
rect 44361 15107 44419 15113
rect 44726 15104 44732 15116
rect 44784 15104 44790 15156
rect 45922 15104 45928 15156
rect 45980 15144 45986 15156
rect 46109 15147 46167 15153
rect 46109 15144 46121 15147
rect 45980 15116 46121 15144
rect 45980 15104 45986 15116
rect 46109 15113 46121 15116
rect 46155 15113 46167 15147
rect 46109 15107 46167 15113
rect 47121 15147 47179 15153
rect 47121 15113 47133 15147
rect 47167 15144 47179 15147
rect 47210 15144 47216 15156
rect 47167 15116 47216 15144
rect 47167 15113 47179 15116
rect 47121 15107 47179 15113
rect 47210 15104 47216 15116
rect 47268 15144 47274 15156
rect 47578 15144 47584 15156
rect 47268 15116 47584 15144
rect 47268 15104 47274 15116
rect 47578 15104 47584 15116
rect 47636 15104 47642 15156
rect 48222 15104 48228 15156
rect 48280 15104 48286 15156
rect 51629 15147 51687 15153
rect 51629 15113 51641 15147
rect 51675 15144 51687 15147
rect 52362 15144 52368 15156
rect 51675 15116 52368 15144
rect 51675 15113 51687 15116
rect 51629 15107 51687 15113
rect 52362 15104 52368 15116
rect 52420 15104 52426 15156
rect 54386 15104 54392 15156
rect 54444 15104 54450 15156
rect 41966 14968 41972 15020
rect 42024 14968 42030 15020
rect 43162 14968 43168 15020
rect 43220 15017 43226 15020
rect 43220 15011 43269 15017
rect 43220 14977 43223 15011
rect 43257 14977 43269 15011
rect 43220 14971 43269 14977
rect 43220 14968 43226 14971
rect 43346 14968 43352 15020
rect 43404 14968 43410 15020
rect 44174 14968 44180 15020
rect 44232 14968 44238 15020
rect 44269 15011 44327 15017
rect 44269 14977 44281 15011
rect 44315 15008 44327 15011
rect 44634 15008 44640 15020
rect 44315 14980 44640 15008
rect 44315 14977 44327 14980
rect 44269 14971 44327 14977
rect 44634 14968 44640 14980
rect 44692 14968 44698 15020
rect 46198 14968 46204 15020
rect 46256 15008 46262 15020
rect 46661 15011 46719 15017
rect 46661 15008 46673 15011
rect 46256 14980 46673 15008
rect 46256 14968 46262 14980
rect 46661 14977 46673 14980
rect 46707 14977 46719 15011
rect 46661 14971 46719 14977
rect 47026 14968 47032 15020
rect 47084 15008 47090 15020
rect 47581 15011 47639 15017
rect 47581 15008 47593 15011
rect 47084 14980 47593 15008
rect 47084 14968 47090 14980
rect 47581 14977 47593 14980
rect 47627 14977 47639 15011
rect 47581 14971 47639 14977
rect 48498 14968 48504 15020
rect 48556 15008 48562 15020
rect 48593 15011 48651 15017
rect 48593 15008 48605 15011
rect 48556 14980 48605 15008
rect 48556 14968 48562 14980
rect 48593 14977 48605 14980
rect 48639 15008 48651 15011
rect 54110 15008 54116 15020
rect 48639 14980 54116 15008
rect 48639 14977 48651 14980
rect 48593 14971 48651 14977
rect 54110 14968 54116 14980
rect 54168 14968 54174 15020
rect 54662 14968 54668 15020
rect 54720 15008 54726 15020
rect 54941 15011 54999 15017
rect 54941 15008 54953 15011
rect 54720 14980 54953 15008
rect 54720 14968 54726 14980
rect 54941 14977 54953 14980
rect 54987 14977 54999 15011
rect 54941 14971 54999 14977
rect 31294 14900 31300 14952
rect 31352 14940 31358 14952
rect 32306 14940 32312 14952
rect 31352 14912 32312 14940
rect 31352 14900 31358 14912
rect 32306 14900 32312 14912
rect 32364 14940 32370 14952
rect 32861 14943 32919 14949
rect 32861 14940 32873 14943
rect 32364 14912 32873 14940
rect 32364 14900 32370 14912
rect 32861 14909 32873 14912
rect 32907 14940 32919 14943
rect 33321 14943 33379 14949
rect 33321 14940 33333 14943
rect 32907 14912 33333 14940
rect 32907 14909 32919 14912
rect 32861 14903 32919 14909
rect 33321 14909 33333 14912
rect 33367 14940 33379 14943
rect 35710 14940 35716 14952
rect 33367 14912 35716 14940
rect 33367 14909 33379 14912
rect 33321 14903 33379 14909
rect 35710 14900 35716 14912
rect 35768 14900 35774 14952
rect 39022 14900 39028 14952
rect 39080 14940 39086 14952
rect 39850 14940 39856 14952
rect 39080 14912 39856 14940
rect 39080 14900 39086 14912
rect 39850 14900 39856 14912
rect 39908 14900 39914 14952
rect 41506 14900 41512 14952
rect 41564 14900 41570 14952
rect 41690 14900 41696 14952
rect 41748 14940 41754 14952
rect 43073 14943 43131 14949
rect 43073 14940 43085 14943
rect 41748 14912 43085 14940
rect 41748 14900 41754 14912
rect 43073 14909 43085 14912
rect 43119 14909 43131 14943
rect 44085 14943 44143 14949
rect 44085 14940 44097 14943
rect 43073 14903 43131 14909
rect 43824 14912 44097 14940
rect 30147 14844 30880 14872
rect 41233 14875 41291 14881
rect 30147 14841 30159 14844
rect 30101 14835 30159 14841
rect 41233 14841 41245 14875
rect 41279 14872 41291 14875
rect 41414 14872 41420 14884
rect 41279 14844 41420 14872
rect 41279 14841 41291 14844
rect 41233 14835 41291 14841
rect 41414 14832 41420 14844
rect 41472 14832 41478 14884
rect 42242 14832 42248 14884
rect 42300 14872 42306 14884
rect 43625 14875 43683 14881
rect 42300 14844 42564 14872
rect 42300 14832 42306 14844
rect 11756 14776 12664 14804
rect 11756 14764 11762 14776
rect 13446 14764 13452 14816
rect 13504 14764 13510 14816
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 16393 14807 16451 14813
rect 16393 14804 16405 14807
rect 13688 14776 16405 14804
rect 13688 14764 13694 14776
rect 16393 14773 16405 14776
rect 16439 14804 16451 14807
rect 16758 14804 16764 14816
rect 16439 14776 16764 14804
rect 16439 14773 16451 14776
rect 16393 14767 16451 14773
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 21266 14764 21272 14816
rect 21324 14804 21330 14816
rect 21453 14807 21511 14813
rect 21453 14804 21465 14807
rect 21324 14776 21465 14804
rect 21324 14764 21330 14776
rect 21453 14773 21465 14776
rect 21499 14773 21511 14807
rect 21453 14767 21511 14773
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 24210 14804 24216 14816
rect 23532 14776 24216 14804
rect 23532 14764 23538 14776
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 34606 14764 34612 14816
rect 34664 14804 34670 14816
rect 35345 14807 35403 14813
rect 35345 14804 35357 14807
rect 34664 14776 35357 14804
rect 34664 14764 34670 14776
rect 35345 14773 35357 14776
rect 35391 14804 35403 14807
rect 35802 14804 35808 14816
rect 35391 14776 35808 14804
rect 35391 14773 35403 14776
rect 35345 14767 35403 14773
rect 35802 14764 35808 14776
rect 35860 14764 35866 14816
rect 42426 14764 42432 14816
rect 42484 14764 42490 14816
rect 42536 14804 42564 14844
rect 43625 14841 43637 14875
rect 43671 14841 43683 14875
rect 43625 14835 43683 14841
rect 43640 14804 43668 14835
rect 43824 14816 43852 14912
rect 44085 14909 44097 14912
rect 44131 14909 44143 14943
rect 44192 14940 44220 14968
rect 44913 14943 44971 14949
rect 44913 14940 44925 14943
rect 44192 14912 44925 14940
rect 44085 14903 44143 14909
rect 44913 14909 44925 14912
rect 44959 14909 44971 14943
rect 44913 14903 44971 14909
rect 49602 14900 49608 14952
rect 49660 14900 49666 14952
rect 50246 14900 50252 14952
rect 50304 14900 50310 14952
rect 51902 14872 51908 14884
rect 51092 14844 51908 14872
rect 51092 14816 51120 14844
rect 51902 14832 51908 14844
rect 51960 14832 51966 14884
rect 42536 14776 43668 14804
rect 43806 14764 43812 14816
rect 43864 14764 43870 14816
rect 46017 14807 46075 14813
rect 46017 14773 46029 14807
rect 46063 14804 46075 14807
rect 46842 14804 46848 14816
rect 46063 14776 46848 14804
rect 46063 14773 46075 14776
rect 46017 14767 46075 14773
rect 46842 14764 46848 14776
rect 46900 14764 46906 14816
rect 48866 14764 48872 14816
rect 48924 14804 48930 14816
rect 48961 14807 49019 14813
rect 48961 14804 48973 14807
rect 48924 14776 48973 14804
rect 48924 14764 48930 14776
rect 48961 14773 48973 14776
rect 49007 14773 49019 14807
rect 48961 14767 49019 14773
rect 49326 14764 49332 14816
rect 49384 14804 49390 14816
rect 49697 14807 49755 14813
rect 49697 14804 49709 14807
rect 49384 14776 49709 14804
rect 49384 14764 49390 14776
rect 49697 14773 49709 14776
rect 49743 14773 49755 14807
rect 49697 14767 49755 14773
rect 51074 14764 51080 14816
rect 51132 14764 51138 14816
rect 57422 14764 57428 14816
rect 57480 14804 57486 14816
rect 58158 14804 58164 14816
rect 57480 14776 58164 14804
rect 57480 14764 57486 14776
rect 58158 14764 58164 14776
rect 58216 14764 58222 14816
rect 1104 14714 58880 14736
rect 1104 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 22616 14714
rect 22668 14662 22680 14714
rect 22732 14662 22744 14714
rect 22796 14662 22808 14714
rect 22860 14662 22872 14714
rect 22924 14662 37060 14714
rect 37112 14662 37124 14714
rect 37176 14662 37188 14714
rect 37240 14662 37252 14714
rect 37304 14662 37316 14714
rect 37368 14662 51504 14714
rect 51556 14662 51568 14714
rect 51620 14662 51632 14714
rect 51684 14662 51696 14714
rect 51748 14662 51760 14714
rect 51812 14662 58880 14714
rect 1104 14640 58880 14662
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 3200 14572 3249 14600
rect 3200 14560 3206 14572
rect 3237 14569 3249 14572
rect 3283 14569 3295 14603
rect 3237 14563 3295 14569
rect 3252 14532 3280 14563
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 4062 14600 4068 14612
rect 3384 14572 4068 14600
rect 3384 14560 3390 14572
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 4706 14600 4712 14612
rect 4571 14572 4712 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 6454 14560 6460 14612
rect 6512 14560 6518 14612
rect 6546 14560 6552 14612
rect 6604 14560 6610 14612
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 6788 14572 6929 14600
rect 6788 14560 6794 14572
rect 6917 14569 6929 14572
rect 6963 14569 6975 14603
rect 9858 14600 9864 14612
rect 6917 14563 6975 14569
rect 9692 14572 9864 14600
rect 3510 14532 3516 14544
rect 3252 14504 3516 14532
rect 3510 14492 3516 14504
rect 3568 14492 3574 14544
rect 4080 14532 4108 14560
rect 4080 14504 4384 14532
rect 3436 14436 4016 14464
rect 3436 14405 3464 14436
rect 3988 14408 4016 14436
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14396 3847 14399
rect 3878 14396 3884 14408
rect 3835 14368 3884 14396
rect 3835 14365 3847 14368
rect 3789 14359 3847 14365
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 3970 14356 3976 14408
rect 4028 14356 4034 14408
rect 4356 14405 4384 14504
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14365 4399 14399
rect 6472 14396 6500 14560
rect 6564 14464 6592 14560
rect 9692 14473 9720 14572
rect 9858 14560 9864 14572
rect 9916 14600 9922 14612
rect 11514 14600 11520 14612
rect 9916 14572 11520 14600
rect 9916 14560 9922 14572
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 14274 14560 14280 14612
rect 14332 14560 14338 14612
rect 14826 14560 14832 14612
rect 14884 14560 14890 14612
rect 18874 14560 18880 14612
rect 18932 14560 18938 14612
rect 21174 14560 21180 14612
rect 21232 14600 21238 14612
rect 21358 14600 21364 14612
rect 21232 14572 21364 14600
rect 21232 14560 21238 14572
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 27801 14603 27859 14609
rect 22066 14572 27752 14600
rect 11057 14535 11115 14541
rect 11057 14501 11069 14535
rect 11103 14501 11115 14535
rect 11057 14495 11115 14501
rect 9677 14467 9735 14473
rect 6564 14436 7144 14464
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6472 14368 6837 14396
rect 4341 14359 4399 14365
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 4080 14328 4108 14359
rect 3660 14300 4108 14328
rect 4172 14328 4200 14359
rect 7006 14356 7012 14408
rect 7064 14356 7070 14408
rect 7116 14405 7144 14436
rect 9677 14433 9689 14467
rect 9723 14433 9735 14467
rect 11072 14464 11100 14495
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 11072 14436 11161 14464
rect 9677 14427 9735 14433
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11532 14464 11560 14560
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 14844 14532 14872 14560
rect 13587 14504 14872 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 16114 14492 16120 14544
rect 16172 14532 16178 14544
rect 22066 14532 22094 14572
rect 16172 14504 22094 14532
rect 27724 14532 27752 14572
rect 27801 14569 27813 14603
rect 27847 14600 27859 14603
rect 28534 14600 28540 14612
rect 27847 14572 28540 14600
rect 27847 14569 27859 14572
rect 27801 14563 27859 14569
rect 28534 14560 28540 14572
rect 28592 14560 28598 14612
rect 28721 14603 28779 14609
rect 28721 14569 28733 14603
rect 28767 14600 28779 14603
rect 28902 14600 28908 14612
rect 28767 14572 28908 14600
rect 28767 14569 28779 14572
rect 28721 14563 28779 14569
rect 28902 14560 28908 14572
rect 28960 14560 28966 14612
rect 30653 14603 30711 14609
rect 30653 14569 30665 14603
rect 30699 14600 30711 14603
rect 32401 14603 32459 14609
rect 32401 14600 32413 14603
rect 30699 14572 32413 14600
rect 30699 14569 30711 14572
rect 30653 14563 30711 14569
rect 32401 14569 32413 14572
rect 32447 14600 32459 14603
rect 32582 14600 32588 14612
rect 32447 14572 32588 14600
rect 32447 14569 32459 14572
rect 32401 14563 32459 14569
rect 32582 14560 32588 14572
rect 32640 14560 32646 14612
rect 34977 14603 35035 14609
rect 34977 14569 34989 14603
rect 35023 14600 35035 14603
rect 35066 14600 35072 14612
rect 35023 14572 35072 14600
rect 35023 14569 35035 14572
rect 34977 14563 35035 14569
rect 35066 14560 35072 14572
rect 35124 14560 35130 14612
rect 35345 14603 35403 14609
rect 35345 14569 35357 14603
rect 35391 14600 35403 14603
rect 35434 14600 35440 14612
rect 35391 14572 35440 14600
rect 35391 14569 35403 14572
rect 35345 14563 35403 14569
rect 35434 14560 35440 14572
rect 35492 14560 35498 14612
rect 37458 14560 37464 14612
rect 37516 14600 37522 14612
rect 37737 14603 37795 14609
rect 37737 14600 37749 14603
rect 37516 14572 37749 14600
rect 37516 14560 37522 14572
rect 37737 14569 37749 14572
rect 37783 14600 37795 14603
rect 38194 14600 38200 14612
rect 37783 14572 38200 14600
rect 37783 14569 37795 14572
rect 37737 14563 37795 14569
rect 38194 14560 38200 14572
rect 38252 14560 38258 14612
rect 39850 14560 39856 14612
rect 39908 14600 39914 14612
rect 41417 14603 41475 14609
rect 41417 14600 41429 14603
rect 39908 14572 41429 14600
rect 39908 14560 39914 14572
rect 41417 14569 41429 14572
rect 41463 14600 41475 14603
rect 42150 14600 42156 14612
rect 41463 14572 42156 14600
rect 41463 14569 41475 14572
rect 41417 14563 41475 14569
rect 42150 14560 42156 14572
rect 42208 14560 42214 14612
rect 42426 14560 42432 14612
rect 42484 14560 42490 14612
rect 42610 14560 42616 14612
rect 42668 14600 42674 14612
rect 47210 14600 47216 14612
rect 42668 14572 47216 14600
rect 42668 14560 42674 14572
rect 47210 14560 47216 14572
rect 47268 14560 47274 14612
rect 48501 14603 48559 14609
rect 48501 14569 48513 14603
rect 48547 14600 48559 14603
rect 48590 14600 48596 14612
rect 48547 14572 48596 14600
rect 48547 14569 48559 14572
rect 48501 14563 48559 14569
rect 48590 14560 48596 14572
rect 48648 14600 48654 14612
rect 48648 14572 49280 14600
rect 48648 14560 48654 14572
rect 30929 14535 30987 14541
rect 30929 14532 30941 14535
rect 27724 14504 30941 14532
rect 16172 14492 16178 14504
rect 30929 14501 30941 14504
rect 30975 14501 30987 14535
rect 30929 14495 30987 14501
rect 12066 14464 12072 14476
rect 11532 14436 12072 14464
rect 11149 14427 11207 14433
rect 12066 14424 12072 14436
rect 12124 14464 12130 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 12124 14436 12173 14464
rect 12124 14424 12130 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 13909 14467 13967 14473
rect 13909 14433 13921 14467
rect 13955 14464 13967 14467
rect 14090 14464 14096 14476
rect 13955 14436 14096 14464
rect 13955 14433 13967 14436
rect 13909 14427 13967 14433
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 16132 14464 16160 14492
rect 15672 14436 16160 14464
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14396 8539 14399
rect 8662 14396 8668 14408
rect 8527 14368 8668 14396
rect 8527 14365 8539 14368
rect 8481 14359 8539 14365
rect 8662 14356 8668 14368
rect 8720 14396 8726 14408
rect 15672 14396 15700 14436
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 19058 14464 19064 14476
rect 16816 14436 19064 14464
rect 16816 14424 16822 14436
rect 19058 14424 19064 14436
rect 19116 14464 19122 14476
rect 21637 14467 21695 14473
rect 21637 14464 21649 14467
rect 19116 14436 21649 14464
rect 19116 14424 19122 14436
rect 21637 14433 21649 14436
rect 21683 14464 21695 14467
rect 22094 14464 22100 14476
rect 21683 14436 22100 14464
rect 21683 14433 21695 14436
rect 21637 14427 21695 14433
rect 22094 14424 22100 14436
rect 22152 14424 22158 14476
rect 26050 14424 26056 14476
rect 26108 14424 26114 14476
rect 30944 14464 30972 14495
rect 31018 14492 31024 14544
rect 31076 14532 31082 14544
rect 31076 14504 42380 14532
rect 31076 14492 31082 14504
rect 31110 14464 31116 14476
rect 30944 14436 31116 14464
rect 31110 14424 31116 14436
rect 31168 14464 31174 14476
rect 41506 14464 41512 14476
rect 31168 14436 41512 14464
rect 31168 14424 31174 14436
rect 41506 14424 41512 14436
rect 41564 14424 41570 14476
rect 42153 14467 42211 14473
rect 42153 14433 42165 14467
rect 42199 14464 42211 14467
rect 42242 14464 42248 14476
rect 42199 14436 42248 14464
rect 42199 14433 42211 14436
rect 42153 14427 42211 14433
rect 42242 14424 42248 14436
rect 42300 14424 42306 14476
rect 8720 14368 15700 14396
rect 15749 14399 15807 14405
rect 8720 14356 8726 14368
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 16022 14396 16028 14408
rect 15795 14368 16028 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16666 14396 16672 14408
rect 16623 14368 16672 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16666 14356 16672 14368
rect 16724 14396 16730 14408
rect 17310 14396 17316 14408
rect 16724 14368 17316 14396
rect 16724 14356 16730 14368
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17494 14356 17500 14408
rect 17552 14356 17558 14408
rect 17954 14356 17960 14408
rect 18012 14356 18018 14408
rect 22370 14356 22376 14408
rect 22428 14356 22434 14408
rect 24670 14356 24676 14408
rect 24728 14396 24734 14408
rect 24949 14399 25007 14405
rect 24949 14396 24961 14399
rect 24728 14368 24961 14396
rect 24728 14356 24734 14368
rect 24949 14365 24961 14368
rect 24995 14365 25007 14399
rect 24949 14359 25007 14365
rect 25314 14356 25320 14408
rect 25372 14356 25378 14408
rect 29730 14356 29736 14408
rect 29788 14356 29794 14408
rect 32398 14396 32404 14408
rect 29840 14368 32404 14396
rect 4522 14328 4528 14340
rect 4172 14300 4528 14328
rect 3660 14288 3666 14300
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 4172 14260 4200 14300
rect 4522 14288 4528 14300
rect 4580 14288 4586 14340
rect 7024 14328 7052 14356
rect 9950 14337 9956 14340
rect 7653 14331 7711 14337
rect 7653 14328 7665 14331
rect 7024 14300 7665 14328
rect 7653 14297 7665 14300
rect 7699 14328 7711 14331
rect 7699 14300 9904 14328
rect 7699 14297 7711 14300
rect 7653 14291 7711 14297
rect 3384 14232 4200 14260
rect 3384 14220 3390 14232
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 9122 14220 9128 14272
rect 9180 14220 9186 14272
rect 9876 14260 9904 14300
rect 9944 14291 9956 14337
rect 9950 14288 9956 14291
rect 10008 14288 10014 14340
rect 10870 14328 10876 14340
rect 10520 14300 10876 14328
rect 10520 14260 10548 14300
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 12428 14331 12486 14337
rect 12428 14297 12440 14331
rect 12474 14328 12486 14331
rect 13262 14328 13268 14340
rect 12474 14300 13268 14328
rect 12474 14297 12486 14300
rect 12428 14291 12486 14297
rect 13262 14288 13268 14300
rect 13320 14288 13326 14340
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 20714 14328 20720 14340
rect 15344 14300 20720 14328
rect 15344 14288 15350 14300
rect 20714 14288 20720 14300
rect 20772 14328 20778 14340
rect 21542 14328 21548 14340
rect 20772 14300 21548 14328
rect 20772 14288 20778 14300
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 26142 14288 26148 14340
rect 26200 14328 26206 14340
rect 26298 14331 26356 14337
rect 26298 14328 26310 14331
rect 26200 14300 26310 14328
rect 26200 14288 26206 14300
rect 26298 14297 26310 14300
rect 26344 14297 26356 14331
rect 26298 14291 26356 14297
rect 27246 14288 27252 14340
rect 27304 14328 27310 14340
rect 29840 14328 29868 14368
rect 32398 14356 32404 14368
rect 32456 14396 32462 14408
rect 32769 14399 32827 14405
rect 32769 14396 32781 14399
rect 32456 14368 32781 14396
rect 32456 14356 32462 14368
rect 32769 14365 32781 14368
rect 32815 14365 32827 14399
rect 32769 14359 32827 14365
rect 36078 14356 36084 14408
rect 36136 14356 36142 14408
rect 36170 14356 36176 14408
rect 36228 14396 36234 14408
rect 37093 14399 37151 14405
rect 37093 14396 37105 14399
rect 36228 14368 37105 14396
rect 36228 14356 36234 14368
rect 37093 14365 37105 14368
rect 37139 14396 37151 14399
rect 37826 14396 37832 14408
rect 37139 14368 37832 14396
rect 37139 14365 37151 14368
rect 37093 14359 37151 14365
rect 37826 14356 37832 14368
rect 37884 14356 37890 14408
rect 38565 14399 38623 14405
rect 38565 14365 38577 14399
rect 38611 14396 38623 14399
rect 38654 14396 38660 14408
rect 38611 14368 38660 14396
rect 38611 14365 38623 14368
rect 38565 14359 38623 14365
rect 38654 14356 38660 14368
rect 38712 14356 38718 14408
rect 42352 14396 42380 14504
rect 42444 14464 42472 14560
rect 42518 14492 42524 14544
rect 42576 14532 42582 14544
rect 49142 14532 49148 14544
rect 42576 14504 42932 14532
rect 42576 14492 42582 14504
rect 42904 14473 42932 14504
rect 42996 14504 49148 14532
rect 42797 14467 42855 14473
rect 42797 14464 42809 14467
rect 42444 14436 42809 14464
rect 42797 14433 42809 14436
rect 42843 14433 42855 14467
rect 42797 14427 42855 14433
rect 42889 14467 42947 14473
rect 42889 14433 42901 14467
rect 42935 14433 42947 14467
rect 42889 14427 42947 14433
rect 42996 14396 43024 14504
rect 49142 14492 49148 14504
rect 49200 14492 49206 14544
rect 49252 14532 49280 14572
rect 49602 14560 49608 14612
rect 49660 14600 49666 14612
rect 49697 14603 49755 14609
rect 49697 14600 49709 14603
rect 49660 14572 49709 14600
rect 49660 14560 49666 14572
rect 49697 14569 49709 14572
rect 49743 14569 49755 14603
rect 49697 14563 49755 14569
rect 54110 14560 54116 14612
rect 54168 14560 54174 14612
rect 56594 14560 56600 14612
rect 56652 14600 56658 14612
rect 56781 14603 56839 14609
rect 56781 14600 56793 14603
rect 56652 14572 56793 14600
rect 56652 14560 56658 14572
rect 56781 14569 56793 14572
rect 56827 14569 56839 14603
rect 56781 14563 56839 14569
rect 51997 14535 52055 14541
rect 49252 14504 50660 14532
rect 43625 14467 43683 14473
rect 43625 14433 43637 14467
rect 43671 14433 43683 14467
rect 43625 14427 43683 14433
rect 42352 14368 43024 14396
rect 43640 14396 43668 14427
rect 43714 14424 43720 14476
rect 43772 14424 43778 14476
rect 44818 14424 44824 14476
rect 44876 14464 44882 14476
rect 45189 14467 45247 14473
rect 45189 14464 45201 14467
rect 44876 14436 45201 14464
rect 44876 14424 44882 14436
rect 45189 14433 45201 14436
rect 45235 14464 45247 14467
rect 48777 14467 48835 14473
rect 48777 14464 48789 14467
rect 45235 14436 48789 14464
rect 45235 14433 45247 14436
rect 45189 14427 45247 14433
rect 48777 14433 48789 14436
rect 48823 14464 48835 14467
rect 49053 14467 49111 14473
rect 49053 14464 49065 14467
rect 48823 14436 49065 14464
rect 48823 14433 48835 14436
rect 48777 14427 48835 14433
rect 44836 14396 44864 14424
rect 43640 14368 44864 14396
rect 44910 14356 44916 14408
rect 44968 14356 44974 14408
rect 46658 14356 46664 14408
rect 46716 14356 46722 14408
rect 27304 14300 29868 14328
rect 30285 14331 30343 14337
rect 27304 14288 27310 14300
rect 30285 14297 30297 14331
rect 30331 14328 30343 14331
rect 30374 14328 30380 14340
rect 30331 14300 30380 14328
rect 30331 14297 30343 14300
rect 30285 14291 30343 14297
rect 30374 14288 30380 14300
rect 30432 14328 30438 14340
rect 33689 14331 33747 14337
rect 30432 14300 31616 14328
rect 30432 14288 30438 14300
rect 31588 14272 31616 14300
rect 33689 14297 33701 14331
rect 33735 14328 33747 14331
rect 34422 14328 34428 14340
rect 33735 14300 34428 14328
rect 33735 14297 33747 14300
rect 33689 14291 33747 14297
rect 34422 14288 34428 14300
rect 34480 14328 34486 14340
rect 35989 14331 36047 14337
rect 35989 14328 36001 14331
rect 34480 14300 36001 14328
rect 34480 14288 34486 14300
rect 35989 14297 36001 14300
rect 36035 14328 36047 14331
rect 38378 14328 38384 14340
rect 36035 14300 36952 14328
rect 36035 14297 36047 14300
rect 35989 14291 36047 14297
rect 36924 14272 36952 14300
rect 37016 14300 38384 14328
rect 37016 14272 37044 14300
rect 38378 14288 38384 14300
rect 38436 14328 38442 14340
rect 41690 14328 41696 14340
rect 38436 14300 41696 14328
rect 38436 14288 38442 14300
rect 41690 14288 41696 14300
rect 41748 14288 41754 14340
rect 41782 14288 41788 14340
rect 41840 14328 41846 14340
rect 44545 14331 44603 14337
rect 41840 14300 42748 14328
rect 41840 14288 41846 14300
rect 9876 14232 10548 14260
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 11793 14263 11851 14269
rect 11793 14260 11805 14263
rect 10652 14232 11805 14260
rect 10652 14220 10658 14232
rect 11793 14229 11805 14232
rect 11839 14260 11851 14263
rect 12250 14260 12256 14272
rect 11839 14232 12256 14260
rect 11839 14229 11851 14232
rect 11793 14223 11851 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14976 14232 15117 14260
rect 14976 14220 14982 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 15930 14220 15936 14272
rect 15988 14220 15994 14272
rect 16942 14220 16948 14272
rect 17000 14220 17006 14272
rect 18598 14220 18604 14272
rect 18656 14220 18662 14272
rect 21818 14220 21824 14272
rect 21876 14220 21882 14272
rect 24029 14263 24087 14269
rect 24029 14229 24041 14263
rect 24075 14260 24087 14263
rect 24210 14260 24216 14272
rect 24075 14232 24216 14260
rect 24075 14229 24087 14232
rect 24029 14223 24087 14229
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 25869 14263 25927 14269
rect 25869 14229 25881 14263
rect 25915 14260 25927 14263
rect 26050 14260 26056 14272
rect 25915 14232 26056 14260
rect 25915 14229 25927 14232
rect 25869 14223 25927 14229
rect 26050 14220 26056 14232
rect 26108 14220 26114 14272
rect 27430 14220 27436 14272
rect 27488 14220 27494 14272
rect 29365 14263 29423 14269
rect 29365 14229 29377 14263
rect 29411 14260 29423 14263
rect 29638 14260 29644 14272
rect 29411 14232 29644 14260
rect 29411 14229 29423 14232
rect 29365 14223 29423 14229
rect 29638 14220 29644 14232
rect 29696 14260 29702 14272
rect 31018 14260 31024 14272
rect 29696 14232 31024 14260
rect 29696 14220 29702 14232
rect 31018 14220 31024 14232
rect 31076 14220 31082 14272
rect 31570 14220 31576 14272
rect 31628 14220 31634 14272
rect 36725 14263 36783 14269
rect 36725 14229 36737 14263
rect 36771 14260 36783 14263
rect 36814 14260 36820 14272
rect 36771 14232 36820 14260
rect 36771 14229 36783 14232
rect 36725 14223 36783 14229
rect 36814 14220 36820 14232
rect 36872 14220 36878 14272
rect 36906 14220 36912 14272
rect 36964 14220 36970 14272
rect 36998 14220 37004 14272
rect 37056 14220 37062 14272
rect 37918 14220 37924 14272
rect 37976 14220 37982 14272
rect 42334 14220 42340 14272
rect 42392 14220 42398 14272
rect 42720 14269 42748 14300
rect 44545 14297 44557 14331
rect 44591 14328 44603 14331
rect 44928 14328 44956 14356
rect 44591 14300 44956 14328
rect 44591 14297 44603 14300
rect 44545 14291 44603 14297
rect 42705 14263 42763 14269
rect 42705 14229 42717 14263
rect 42751 14229 42763 14263
rect 42705 14223 42763 14229
rect 43806 14220 43812 14272
rect 43864 14220 43870 14272
rect 44174 14220 44180 14272
rect 44232 14220 44238 14272
rect 45922 14220 45928 14272
rect 45980 14260 45986 14272
rect 46109 14263 46167 14269
rect 46109 14260 46121 14263
rect 45980 14232 46121 14260
rect 45980 14220 45986 14232
rect 46109 14229 46121 14232
rect 46155 14229 46167 14263
rect 46109 14223 46167 14229
rect 46198 14220 46204 14272
rect 46256 14260 46262 14272
rect 48590 14260 48596 14272
rect 46256 14232 48596 14260
rect 46256 14220 46262 14232
rect 48590 14220 48596 14232
rect 48648 14220 48654 14272
rect 48976 14260 49004 14436
rect 49053 14433 49065 14436
rect 49099 14433 49111 14467
rect 49053 14427 49111 14433
rect 49234 14356 49240 14408
rect 49292 14356 49298 14408
rect 49326 14356 49332 14408
rect 49384 14356 49390 14408
rect 50632 14405 50660 14504
rect 51997 14501 52009 14535
rect 52043 14532 52055 14535
rect 52546 14532 52552 14544
rect 52043 14504 52552 14532
rect 52043 14501 52055 14504
rect 51997 14495 52055 14501
rect 52546 14492 52552 14504
rect 52604 14532 52610 14544
rect 52604 14504 53512 14532
rect 52604 14492 52610 14504
rect 51902 14424 51908 14476
rect 51960 14464 51966 14476
rect 53484 14473 53512 14504
rect 52641 14467 52699 14473
rect 52641 14464 52653 14467
rect 51960 14436 52653 14464
rect 51960 14424 51966 14436
rect 52641 14433 52653 14436
rect 52687 14433 52699 14467
rect 52641 14427 52699 14433
rect 53469 14467 53527 14473
rect 53469 14433 53481 14467
rect 53515 14433 53527 14467
rect 53469 14427 53527 14433
rect 50617 14399 50675 14405
rect 50617 14365 50629 14399
rect 50663 14365 50675 14399
rect 50617 14359 50675 14365
rect 49694 14260 49700 14272
rect 48976 14232 49700 14260
rect 49694 14220 49700 14232
rect 49752 14220 49758 14272
rect 50525 14263 50583 14269
rect 50525 14229 50537 14263
rect 50571 14260 50583 14263
rect 50632 14260 50660 14359
rect 54846 14356 54852 14408
rect 54904 14356 54910 14408
rect 58434 14356 58440 14408
rect 58492 14356 58498 14408
rect 50884 14331 50942 14337
rect 50884 14297 50896 14331
rect 50930 14328 50942 14331
rect 51534 14328 51540 14340
rect 50930 14300 51540 14328
rect 50930 14297 50942 14300
rect 50884 14291 50942 14297
rect 51534 14288 51540 14300
rect 51592 14288 51598 14340
rect 52457 14331 52515 14337
rect 52457 14297 52469 14331
rect 52503 14328 52515 14331
rect 52917 14331 52975 14337
rect 52917 14328 52929 14331
rect 52503 14300 52929 14328
rect 52503 14297 52515 14300
rect 52457 14291 52515 14297
rect 52917 14297 52929 14300
rect 52963 14297 52975 14331
rect 52917 14291 52975 14297
rect 53006 14288 53012 14340
rect 53064 14288 53070 14340
rect 51902 14260 51908 14272
rect 50571 14232 51908 14260
rect 50571 14229 50583 14232
rect 50525 14223 50583 14229
rect 51902 14220 51908 14232
rect 51960 14220 51966 14272
rect 52086 14220 52092 14272
rect 52144 14220 52150 14272
rect 52549 14263 52607 14269
rect 52549 14229 52561 14263
rect 52595 14260 52607 14263
rect 53024 14260 53052 14288
rect 52595 14232 53052 14260
rect 52595 14229 52607 14232
rect 52549 14223 52607 14229
rect 54294 14220 54300 14272
rect 54352 14220 54358 14272
rect 56870 14220 56876 14272
rect 56928 14260 56934 14272
rect 57149 14263 57207 14269
rect 57149 14260 57161 14263
rect 56928 14232 57161 14260
rect 56928 14220 56934 14232
rect 57149 14229 57161 14232
rect 57195 14229 57207 14263
rect 57149 14223 57207 14229
rect 57238 14220 57244 14272
rect 57296 14260 57302 14272
rect 57885 14263 57943 14269
rect 57885 14260 57897 14263
rect 57296 14232 57897 14260
rect 57296 14220 57302 14232
rect 57885 14229 57897 14232
rect 57931 14229 57943 14263
rect 57885 14223 57943 14229
rect 1104 14170 59040 14192
rect 1104 14118 15394 14170
rect 15446 14118 15458 14170
rect 15510 14118 15522 14170
rect 15574 14118 15586 14170
rect 15638 14118 15650 14170
rect 15702 14118 29838 14170
rect 29890 14118 29902 14170
rect 29954 14118 29966 14170
rect 30018 14118 30030 14170
rect 30082 14118 30094 14170
rect 30146 14118 44282 14170
rect 44334 14118 44346 14170
rect 44398 14118 44410 14170
rect 44462 14118 44474 14170
rect 44526 14118 44538 14170
rect 44590 14118 58726 14170
rect 58778 14118 58790 14170
rect 58842 14118 58854 14170
rect 58906 14118 58918 14170
rect 58970 14118 58982 14170
rect 59034 14118 59040 14170
rect 1104 14096 59040 14118
rect 3326 14016 3332 14068
rect 3384 14016 3390 14068
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 4338 14056 4344 14068
rect 3835 14028 4344 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7190 14056 7196 14068
rect 6871 14028 7196 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 8662 14016 8668 14068
rect 8720 14016 8726 14068
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9858 14056 9864 14068
rect 9079 14028 9864 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 3970 13988 3976 14000
rect 3804 13960 3976 13988
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 2746 13892 3249 13920
rect 2746 13784 2774 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 3602 13880 3608 13932
rect 3660 13880 3666 13932
rect 3804 13929 3832 13960
rect 3970 13948 3976 13960
rect 4028 13988 4034 14000
rect 5261 13991 5319 13997
rect 5261 13988 5273 13991
rect 4028 13960 5273 13988
rect 4028 13948 4034 13960
rect 5261 13957 5273 13960
rect 5307 13957 5319 13991
rect 7300 13988 7328 14016
rect 7938 13991 7996 13997
rect 7938 13988 7950 13991
rect 7300 13960 7950 13988
rect 5261 13951 5319 13957
rect 7938 13957 7950 13960
rect 7984 13957 7996 13991
rect 7938 13951 7996 13957
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 3936 13892 5181 13920
rect 3936 13880 3942 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 6362 13920 6368 13932
rect 5399 13892 6368 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 3620 13852 3648 13880
rect 4062 13852 4068 13864
rect 3620 13824 4068 13852
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 5184 13852 5212 13883
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 8205 13923 8263 13929
rect 8205 13889 8217 13923
rect 8251 13920 8263 13923
rect 9048 13920 9076 14019
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 9950 14016 9956 14068
rect 10008 14016 10014 14068
rect 10229 14059 10287 14065
rect 10229 14025 10241 14059
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 9493 13991 9551 13997
rect 9493 13957 9505 13991
rect 9539 13988 9551 13991
rect 9968 13988 9996 14016
rect 9539 13960 9996 13988
rect 9539 13957 9551 13960
rect 9493 13951 9551 13957
rect 8251 13892 9076 13920
rect 9401 13923 9459 13929
rect 8251 13889 8263 13892
rect 8205 13883 8263 13889
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9674 13920 9680 13932
rect 9447 13892 9680 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 10244 13920 10272 14019
rect 10594 14016 10600 14068
rect 10652 14016 10658 14068
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 10928 14028 11253 14056
rect 10928 14016 10934 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 11241 14019 11299 14025
rect 10183 13892 10272 13920
rect 10704 13920 10732 14016
rect 11256 13988 11284 14019
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 12250 14056 12256 14068
rect 11388 14028 12256 14056
rect 11388 14016 11394 14028
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12434 14016 12440 14068
rect 12492 14016 12498 14068
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 12897 14059 12955 14065
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 13170 14056 13176 14068
rect 12943 14028 13176 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13262 14016 13268 14068
rect 13320 14016 13326 14068
rect 13446 14016 13452 14068
rect 13504 14016 13510 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 15930 14056 15936 14068
rect 15611 14028 15936 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16022 14016 16028 14068
rect 16080 14016 16086 14068
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 16264 14028 16405 14056
rect 16264 14016 16270 14028
rect 16393 14025 16405 14028
rect 16439 14025 16451 14059
rect 16393 14019 16451 14025
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 18509 14059 18567 14065
rect 18509 14025 18521 14059
rect 18555 14056 18567 14059
rect 18598 14056 18604 14068
rect 18555 14028 18604 14056
rect 18555 14025 18567 14028
rect 18509 14019 18567 14025
rect 12728 13988 12756 14016
rect 11256 13960 12756 13988
rect 12805 13923 12863 13929
rect 12805 13920 12817 13923
rect 10704 13892 12817 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 12805 13889 12817 13892
rect 12851 13920 12863 13923
rect 13464 13920 13492 14016
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 16574 13988 16580 14000
rect 15252 13960 16580 13988
rect 15252 13948 15258 13960
rect 16574 13948 16580 13960
rect 16632 13948 16638 14000
rect 16942 13997 16948 14000
rect 16925 13991 16948 13997
rect 16925 13957 16937 13991
rect 16925 13951 16948 13957
rect 16942 13948 16948 13951
rect 17000 13948 17006 14000
rect 18064 13988 18092 14019
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 18877 14059 18935 14065
rect 18877 14025 18889 14059
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 22557 14059 22615 14065
rect 22557 14025 22569 14059
rect 22603 14025 22615 14059
rect 22557 14019 22615 14025
rect 18064 13960 18828 13988
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 12851 13892 13308 13920
rect 13464 13892 13829 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 5902 13852 5908 13864
rect 5184 13824 5908 13852
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 9122 13852 9128 13864
rect 8312 13824 9128 13852
rect 8312 13784 8340 13824
rect 9122 13812 9128 13824
rect 9180 13852 9186 13864
rect 10502 13852 10508 13864
rect 9180 13824 10508 13852
rect 9180 13812 9186 13824
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10612 13824 10793 13852
rect 2608 13756 2774 13784
rect 8220 13756 8340 13784
rect 2608 13728 2636 13756
rect 2590 13676 2596 13728
rect 2648 13676 2654 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 8220 13716 8248 13756
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 10612 13784 10640 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13821 13139 13855
rect 13280 13852 13308 13892
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 15746 13920 15752 13932
rect 15703 13892 15752 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18417 13923 18475 13929
rect 18417 13920 18429 13923
rect 18104 13892 18429 13920
rect 18104 13880 18110 13892
rect 18417 13889 18429 13892
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 13924 13852 13952 13880
rect 13280 13824 13952 13852
rect 13081 13815 13139 13821
rect 9732 13756 10640 13784
rect 9732 13744 9738 13756
rect 12250 13744 12256 13796
rect 12308 13784 12314 13796
rect 13096 13784 13124 13815
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14424 13824 14749 13852
rect 14424 13812 14430 13824
rect 14737 13821 14749 13824
rect 14783 13852 14795 13855
rect 15286 13852 15292 13864
rect 14783 13824 15292 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 15286 13812 15292 13824
rect 15344 13852 15350 13864
rect 15381 13855 15439 13861
rect 15381 13852 15393 13855
rect 15344 13824 15393 13852
rect 15344 13812 15350 13824
rect 15381 13821 15393 13824
rect 15427 13821 15439 13855
rect 15381 13815 15439 13821
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 16390 13812 16396 13864
rect 16448 13852 16454 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16448 13824 16681 13852
rect 16448 13812 16454 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 18233 13855 18291 13861
rect 18233 13852 18245 13855
rect 16669 13815 16727 13821
rect 17972 13824 18245 13852
rect 12308 13756 15332 13784
rect 12308 13744 12314 13756
rect 15304 13728 15332 13756
rect 6880 13688 8248 13716
rect 6880 13676 6886 13688
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 11606 13716 11612 13728
rect 11388 13688 11612 13716
rect 11388 13676 11394 13688
rect 11606 13676 11612 13688
rect 11664 13716 11670 13728
rect 11701 13719 11759 13725
rect 11701 13716 11713 13719
rect 11664 13688 11713 13716
rect 11664 13676 11670 13688
rect 11701 13685 11713 13688
rect 11747 13685 11759 13719
rect 11701 13679 11759 13685
rect 15286 13676 15292 13728
rect 15344 13676 15350 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16224 13716 16252 13812
rect 17972 13716 18000 13824
rect 18233 13821 18245 13824
rect 18279 13821 18291 13855
rect 18800 13852 18828 13960
rect 18892 13920 18920 14019
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 18892 13892 19533 13920
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 21818 13920 21824 13932
rect 20956 13892 21824 13920
rect 20956 13880 20962 13892
rect 21818 13880 21824 13892
rect 21876 13920 21882 13932
rect 22097 13923 22155 13929
rect 22097 13920 22109 13923
rect 21876 13892 22109 13920
rect 21876 13880 21882 13892
rect 22097 13889 22109 13892
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22572 13920 22600 14019
rect 25314 14016 25320 14068
rect 25372 14056 25378 14068
rect 25501 14059 25559 14065
rect 25501 14056 25513 14059
rect 25372 14028 25513 14056
rect 25372 14016 25378 14028
rect 25501 14025 25513 14028
rect 25547 14025 25559 14059
rect 25501 14019 25559 14025
rect 26142 14016 26148 14068
rect 26200 14016 26206 14068
rect 27246 14016 27252 14068
rect 27304 14016 27310 14068
rect 27430 14016 27436 14068
rect 27488 14016 27494 14068
rect 28813 14059 28871 14065
rect 28813 14025 28825 14059
rect 28859 14025 28871 14059
rect 28813 14019 28871 14025
rect 29273 14059 29331 14065
rect 29273 14025 29285 14059
rect 29319 14056 29331 14059
rect 30374 14056 30380 14068
rect 29319 14028 30380 14056
rect 29319 14025 29331 14028
rect 29273 14019 29331 14025
rect 24210 13948 24216 14000
rect 24268 13988 24274 14000
rect 24268 13960 26740 13988
rect 24268 13948 24274 13960
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 22572 13892 23213 13920
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 19794 13852 19800 13864
rect 18800 13824 19800 13852
rect 18233 13815 18291 13821
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 19978 13812 19984 13864
rect 20036 13852 20042 13864
rect 20165 13855 20223 13861
rect 20165 13852 20177 13855
rect 20036 13824 20177 13852
rect 20036 13812 20042 13824
rect 20165 13821 20177 13824
rect 20211 13821 20223 13855
rect 20165 13815 20223 13821
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 20404 13824 20729 13852
rect 20404 13812 20410 13824
rect 20717 13821 20729 13824
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 20990 13812 20996 13864
rect 21048 13812 21054 13864
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13852 22063 13855
rect 22051 13824 23428 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22112 13796 22140 13824
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18322 13784 18328 13796
rect 18104 13756 18328 13784
rect 18104 13744 18110 13756
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 21266 13744 21272 13796
rect 21324 13784 21330 13796
rect 21324 13756 22057 13784
rect 21324 13744 21330 13756
rect 16080 13688 18000 13716
rect 16080 13676 16086 13688
rect 18966 13676 18972 13728
rect 19024 13676 19030 13728
rect 20070 13676 20076 13728
rect 20128 13716 20134 13728
rect 20714 13716 20720 13728
rect 20128 13688 20720 13716
rect 20128 13676 20134 13688
rect 20714 13676 20720 13688
rect 20772 13676 20778 13728
rect 20806 13676 20812 13728
rect 20864 13716 20870 13728
rect 21637 13719 21695 13725
rect 21637 13716 21649 13719
rect 20864 13688 21649 13716
rect 20864 13676 20870 13688
rect 21637 13685 21649 13688
rect 21683 13685 21695 13719
rect 22029 13716 22057 13756
rect 22094 13744 22100 13796
rect 22152 13744 22158 13796
rect 22462 13744 22468 13796
rect 22520 13784 22526 13796
rect 22649 13787 22707 13793
rect 22649 13784 22661 13787
rect 22520 13756 22661 13784
rect 22520 13744 22526 13756
rect 22649 13753 22661 13756
rect 22695 13753 22707 13787
rect 23400 13784 23428 13824
rect 23474 13812 23480 13864
rect 23532 13812 23538 13864
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24228 13852 24256 13948
rect 24394 13929 24400 13932
rect 24388 13920 24400 13929
rect 24355 13892 24400 13920
rect 24388 13883 24400 13892
rect 24394 13880 24400 13883
rect 24452 13880 24458 13932
rect 26712 13864 26740 13960
rect 27448 13929 27476 14016
rect 27433 13923 27491 13929
rect 27433 13889 27445 13923
rect 27479 13889 27491 13923
rect 27433 13883 27491 13889
rect 28169 13923 28227 13929
rect 28169 13889 28181 13923
rect 28215 13920 28227 13923
rect 28828 13920 28856 14019
rect 30374 14016 30380 14028
rect 30432 14016 30438 14068
rect 32398 14016 32404 14068
rect 32456 14016 32462 14068
rect 35805 14059 35863 14065
rect 35805 14025 35817 14059
rect 35851 14056 35863 14059
rect 36078 14056 36084 14068
rect 35851 14028 36084 14056
rect 35851 14025 35863 14028
rect 35805 14019 35863 14025
rect 36078 14016 36084 14028
rect 36136 14016 36142 14068
rect 36538 14016 36544 14068
rect 36596 14016 36602 14068
rect 37277 14059 37335 14065
rect 37277 14025 37289 14059
rect 37323 14056 37335 14059
rect 38378 14056 38384 14068
rect 37323 14028 38384 14056
rect 37323 14025 37335 14028
rect 37277 14019 37335 14025
rect 38378 14016 38384 14028
rect 38436 14016 38442 14068
rect 38841 14059 38899 14065
rect 38841 14025 38853 14059
rect 38887 14025 38899 14059
rect 38841 14019 38899 14025
rect 30469 13991 30527 13997
rect 30469 13988 30481 13991
rect 29472 13960 30481 13988
rect 28215 13892 28856 13920
rect 29181 13923 29239 13929
rect 28215 13889 28227 13892
rect 28169 13883 28227 13889
rect 29181 13889 29193 13923
rect 29227 13920 29239 13923
rect 29270 13920 29276 13932
rect 29227 13892 29276 13920
rect 29227 13889 29239 13892
rect 29181 13883 29239 13889
rect 29270 13880 29276 13892
rect 29328 13880 29334 13932
rect 29472 13864 29500 13960
rect 30469 13957 30481 13960
rect 30515 13988 30527 13991
rect 30926 13988 30932 14000
rect 30515 13960 30932 13988
rect 30515 13957 30527 13960
rect 30469 13951 30527 13957
rect 30926 13948 30932 13960
rect 30984 13988 30990 14000
rect 31662 13988 31668 14000
rect 30984 13960 31668 13988
rect 30984 13948 30990 13960
rect 31662 13948 31668 13960
rect 31720 13948 31726 14000
rect 29638 13880 29644 13932
rect 29696 13880 29702 13932
rect 31110 13880 31116 13932
rect 31168 13880 31174 13932
rect 32416 13929 32444 14016
rect 33229 13991 33287 13997
rect 33229 13957 33241 13991
rect 33275 13988 33287 13991
rect 34054 13988 34060 14000
rect 33275 13960 34060 13988
rect 33275 13957 33287 13960
rect 33229 13951 33287 13957
rect 34054 13948 34060 13960
rect 34112 13988 34118 14000
rect 34330 13988 34336 14000
rect 34112 13960 34336 13988
rect 34112 13948 34118 13960
rect 34330 13948 34336 13960
rect 34388 13948 34394 14000
rect 36556 13988 36584 14016
rect 37645 13991 37703 13997
rect 37645 13988 37657 13991
rect 36556 13960 37657 13988
rect 37645 13957 37657 13960
rect 37691 13957 37703 13991
rect 37645 13951 37703 13957
rect 37844 13960 38654 13988
rect 32401 13923 32459 13929
rect 32401 13889 32413 13923
rect 32447 13889 32459 13923
rect 32401 13883 32459 13889
rect 34422 13880 34428 13932
rect 34480 13880 34486 13932
rect 34692 13923 34750 13929
rect 34692 13889 34704 13923
rect 34738 13920 34750 13923
rect 35897 13923 35955 13929
rect 35897 13920 35909 13923
rect 34738 13892 35909 13920
rect 34738 13889 34750 13892
rect 34692 13883 34750 13889
rect 35897 13889 35909 13892
rect 35943 13889 35955 13923
rect 35897 13883 35955 13889
rect 24167 13824 24256 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 25866 13812 25872 13864
rect 25924 13812 25930 13864
rect 26694 13812 26700 13864
rect 26752 13812 26758 13864
rect 26786 13812 26792 13864
rect 26844 13812 26850 13864
rect 27522 13812 27528 13864
rect 27580 13852 27586 13864
rect 27985 13855 28043 13861
rect 27985 13852 27997 13855
rect 27580 13824 27997 13852
rect 27580 13812 27586 13824
rect 27985 13821 27997 13824
rect 28031 13821 28043 13855
rect 27985 13815 28043 13821
rect 29454 13812 29460 13864
rect 29512 13812 29518 13864
rect 23400 13756 24164 13784
rect 22649 13747 22707 13753
rect 23014 13716 23020 13728
rect 22029 13688 23020 13716
rect 21637 13679 21695 13685
rect 23014 13676 23020 13688
rect 23072 13716 23078 13728
rect 23290 13716 23296 13728
rect 23072 13688 23296 13716
rect 23072 13676 23078 13688
rect 23290 13676 23296 13688
rect 23348 13676 23354 13728
rect 24026 13676 24032 13728
rect 24084 13676 24090 13728
rect 24136 13716 24164 13756
rect 25130 13744 25136 13796
rect 25188 13784 25194 13796
rect 29656 13784 29684 13880
rect 37844 13864 37872 13960
rect 37918 13880 37924 13932
rect 37976 13920 37982 13932
rect 38473 13923 38531 13929
rect 38473 13920 38485 13923
rect 37976 13892 38485 13920
rect 37976 13880 37982 13892
rect 38473 13889 38485 13892
rect 38519 13889 38531 13923
rect 38473 13883 38531 13889
rect 31665 13855 31723 13861
rect 31665 13821 31677 13855
rect 31711 13852 31723 13855
rect 31846 13852 31852 13864
rect 31711 13824 31852 13852
rect 31711 13821 31723 13824
rect 31665 13815 31723 13821
rect 31846 13812 31852 13824
rect 31904 13852 31910 13864
rect 32858 13852 32864 13864
rect 31904 13824 32864 13852
rect 31904 13812 31910 13824
rect 32858 13812 32864 13824
rect 32916 13812 32922 13864
rect 33502 13812 33508 13864
rect 33560 13812 33566 13864
rect 34146 13812 34152 13864
rect 34204 13812 34210 13864
rect 36078 13812 36084 13864
rect 36136 13852 36142 13864
rect 36449 13855 36507 13861
rect 36449 13852 36461 13855
rect 36136 13824 36461 13852
rect 36136 13812 36142 13824
rect 36449 13821 36461 13824
rect 36495 13821 36507 13855
rect 36449 13815 36507 13821
rect 36630 13812 36636 13864
rect 36688 13852 36694 13864
rect 37737 13855 37795 13861
rect 37737 13852 37749 13855
rect 36688 13824 37749 13852
rect 36688 13812 36694 13824
rect 37737 13821 37749 13824
rect 37783 13821 37795 13855
rect 37737 13815 37795 13821
rect 37826 13812 37832 13864
rect 37884 13812 37890 13864
rect 38010 13812 38016 13864
rect 38068 13852 38074 13864
rect 38194 13852 38200 13864
rect 38068 13824 38200 13852
rect 38068 13812 38074 13824
rect 38194 13812 38200 13824
rect 38252 13812 38258 13864
rect 38381 13855 38439 13861
rect 38381 13821 38393 13855
rect 38427 13821 38439 13855
rect 38626 13852 38654 13960
rect 38856 13920 38884 14019
rect 39758 14016 39764 14068
rect 39816 14016 39822 14068
rect 40310 14016 40316 14068
rect 40368 14056 40374 14068
rect 40773 14059 40831 14065
rect 40773 14056 40785 14059
rect 40368 14028 40785 14056
rect 40368 14016 40374 14028
rect 40773 14025 40785 14028
rect 40819 14056 40831 14059
rect 42150 14056 42156 14068
rect 40819 14028 42156 14056
rect 40819 14025 40831 14028
rect 40773 14019 40831 14025
rect 42150 14016 42156 14028
rect 42208 14016 42214 14068
rect 42245 14059 42303 14065
rect 42245 14025 42257 14059
rect 42291 14056 42303 14059
rect 42518 14056 42524 14068
rect 42291 14028 42524 14056
rect 42291 14025 42303 14028
rect 42245 14019 42303 14025
rect 39485 13923 39543 13929
rect 39485 13920 39497 13923
rect 38856 13892 39497 13920
rect 39485 13889 39497 13892
rect 39531 13889 39543 13923
rect 39485 13883 39543 13889
rect 39776 13920 39804 14016
rect 42260 13920 42288 14019
rect 42518 14016 42524 14028
rect 42576 14016 42582 14068
rect 43806 14016 43812 14068
rect 43864 14056 43870 14068
rect 45005 14059 45063 14065
rect 45005 14056 45017 14059
rect 43864 14028 45017 14056
rect 43864 14016 43870 14028
rect 45005 14025 45017 14028
rect 45051 14025 45063 14059
rect 45005 14019 45063 14025
rect 46017 14059 46075 14065
rect 46017 14025 46029 14059
rect 46063 14056 46075 14059
rect 46198 14056 46204 14068
rect 46063 14028 46204 14056
rect 46063 14025 46075 14028
rect 46017 14019 46075 14025
rect 46198 14016 46204 14028
rect 46256 14016 46262 14068
rect 46293 14059 46351 14065
rect 46293 14025 46305 14059
rect 46339 14056 46351 14059
rect 46658 14056 46664 14068
rect 46339 14028 46664 14056
rect 46339 14025 46351 14028
rect 46293 14019 46351 14025
rect 46658 14016 46664 14028
rect 46716 14016 46722 14068
rect 46750 14016 46756 14068
rect 46808 14016 46814 14068
rect 49973 14059 50031 14065
rect 49973 14025 49985 14059
rect 50019 14056 50031 14059
rect 50246 14056 50252 14068
rect 50019 14028 50252 14056
rect 50019 14025 50031 14028
rect 49973 14019 50031 14025
rect 50246 14016 50252 14028
rect 50304 14016 50310 14068
rect 51534 14016 51540 14068
rect 51592 14016 51598 14068
rect 54481 14059 54539 14065
rect 54481 14025 54493 14059
rect 54527 14056 54539 14059
rect 54846 14056 54852 14068
rect 54527 14028 54852 14056
rect 54527 14025 54539 14028
rect 54481 14019 54539 14025
rect 54846 14016 54852 14028
rect 54904 14016 54910 14068
rect 56594 14016 56600 14068
rect 56652 14016 56658 14068
rect 57238 14016 57244 14068
rect 57296 14016 57302 14068
rect 57333 14059 57391 14065
rect 57333 14025 57345 14059
rect 57379 14056 57391 14059
rect 57514 14056 57520 14068
rect 57379 14028 57520 14056
rect 57379 14025 57391 14028
rect 57333 14019 57391 14025
rect 57514 14016 57520 14028
rect 57572 14016 57578 14068
rect 57701 14059 57759 14065
rect 57701 14025 57713 14059
rect 57747 14056 57759 14059
rect 57747 14028 58480 14056
rect 57747 14025 57759 14028
rect 57701 14019 57759 14025
rect 42429 13991 42487 13997
rect 42429 13957 42441 13991
rect 42475 13988 42487 13991
rect 42702 13988 42708 14000
rect 42475 13960 42708 13988
rect 42475 13957 42487 13960
rect 42429 13951 42487 13957
rect 42702 13948 42708 13960
rect 42760 13988 42766 14000
rect 52454 13988 52460 14000
rect 42760 13960 52460 13988
rect 42760 13948 42766 13960
rect 52454 13948 52460 13960
rect 52512 13948 52518 14000
rect 55122 13988 55128 14000
rect 54864 13960 55128 13988
rect 39776 13892 41276 13920
rect 39776 13852 39804 13892
rect 38626 13824 39804 13852
rect 38381 13815 38439 13821
rect 25188 13756 29684 13784
rect 25188 13744 25194 13756
rect 33962 13744 33968 13796
rect 34020 13784 34026 13796
rect 34330 13784 34336 13796
rect 34020 13756 34336 13784
rect 34020 13744 34026 13756
rect 34330 13744 34336 13756
rect 34388 13744 34394 13796
rect 36817 13787 36875 13793
rect 36817 13784 36829 13787
rect 35728 13756 36829 13784
rect 35728 13728 35756 13756
rect 36817 13753 36829 13756
rect 36863 13784 36875 13787
rect 36998 13784 37004 13796
rect 36863 13756 37004 13784
rect 36863 13753 36875 13756
rect 36817 13747 36875 13753
rect 36998 13744 37004 13756
rect 37056 13744 37062 13796
rect 37642 13744 37648 13796
rect 37700 13784 37706 13796
rect 38396 13784 38424 13815
rect 41046 13812 41052 13864
rect 41104 13812 41110 13864
rect 41248 13852 41276 13892
rect 41524 13892 42288 13920
rect 41524 13852 41552 13892
rect 44082 13880 44088 13932
rect 44140 13880 44146 13932
rect 44174 13880 44180 13932
rect 44232 13920 44238 13932
rect 44821 13923 44879 13929
rect 44821 13920 44833 13923
rect 44232 13892 44833 13920
rect 44232 13880 44238 13892
rect 44821 13889 44833 13892
rect 44867 13889 44879 13923
rect 44821 13883 44879 13889
rect 46661 13923 46719 13929
rect 46661 13889 46673 13923
rect 46707 13920 46719 13923
rect 48225 13923 48283 13929
rect 48225 13920 48237 13923
rect 46707 13892 48237 13920
rect 46707 13889 46719 13892
rect 46661 13883 46719 13889
rect 48225 13889 48237 13892
rect 48271 13920 48283 13923
rect 48314 13920 48320 13932
rect 48271 13892 48320 13920
rect 48271 13889 48283 13892
rect 48225 13883 48283 13889
rect 48314 13880 48320 13892
rect 48372 13880 48378 13932
rect 48590 13880 48596 13932
rect 48648 13880 48654 13932
rect 48866 13929 48872 13932
rect 48860 13920 48872 13929
rect 48827 13892 48872 13920
rect 48860 13883 48872 13892
rect 48866 13880 48872 13883
rect 48924 13880 48930 13932
rect 49142 13880 49148 13932
rect 49200 13920 49206 13932
rect 49200 13892 51304 13920
rect 49200 13880 49206 13892
rect 41248 13824 41552 13852
rect 41598 13812 41604 13864
rect 41656 13812 41662 13864
rect 42242 13812 42248 13864
rect 42300 13852 42306 13864
rect 42518 13852 42524 13864
rect 42300 13824 42524 13852
rect 42300 13812 42306 13824
rect 42518 13812 42524 13824
rect 42576 13812 42582 13864
rect 45554 13812 45560 13864
rect 45612 13812 45618 13864
rect 46845 13855 46903 13861
rect 46845 13821 46857 13855
rect 46891 13852 46903 13855
rect 47397 13855 47455 13861
rect 47397 13852 47409 13855
rect 46891 13824 47409 13852
rect 46891 13821 46903 13824
rect 46845 13815 46903 13821
rect 37700 13756 38424 13784
rect 37700 13744 37706 13756
rect 26418 13716 26424 13728
rect 24136 13688 26424 13716
rect 26418 13676 26424 13688
rect 26476 13676 26482 13728
rect 28721 13719 28779 13725
rect 28721 13685 28733 13719
rect 28767 13716 28779 13719
rect 28810 13716 28816 13728
rect 28767 13688 28816 13716
rect 28767 13685 28779 13688
rect 28721 13679 28779 13685
rect 28810 13676 28816 13688
rect 28868 13676 28874 13728
rect 35710 13676 35716 13728
rect 35768 13676 35774 13728
rect 35802 13676 35808 13728
rect 35860 13716 35866 13728
rect 36722 13716 36728 13728
rect 35860 13688 36728 13716
rect 35860 13676 35866 13688
rect 36722 13676 36728 13688
rect 36780 13676 36786 13728
rect 38746 13676 38752 13728
rect 38804 13716 38810 13728
rect 38933 13719 38991 13725
rect 38933 13716 38945 13719
rect 38804 13688 38945 13716
rect 38804 13676 38810 13688
rect 38933 13685 38945 13688
rect 38979 13685 38991 13719
rect 38933 13679 38991 13685
rect 44266 13676 44272 13728
rect 44324 13676 44330 13728
rect 46474 13676 46480 13728
rect 46532 13716 46538 13728
rect 47044 13716 47072 13824
rect 47397 13821 47409 13824
rect 47443 13821 47455 13855
rect 47397 13815 47455 13821
rect 47412 13784 47440 13815
rect 47578 13812 47584 13864
rect 47636 13812 47642 13864
rect 47762 13812 47768 13864
rect 47820 13812 47826 13864
rect 50062 13812 50068 13864
rect 50120 13812 50126 13864
rect 47780 13784 47808 13812
rect 47412 13756 47808 13784
rect 51276 13784 51304 13892
rect 52086 13880 52092 13932
rect 52144 13880 52150 13932
rect 54864 13929 54892 13960
rect 55122 13948 55128 13960
rect 55180 13948 55186 14000
rect 54849 13923 54907 13929
rect 54849 13889 54861 13923
rect 54895 13889 54907 13923
rect 54849 13883 54907 13889
rect 54941 13923 54999 13929
rect 54941 13889 54953 13923
rect 54987 13920 54999 13923
rect 55858 13920 55864 13932
rect 54987 13892 55864 13920
rect 54987 13889 54999 13892
rect 54941 13883 54999 13889
rect 55858 13880 55864 13892
rect 55916 13920 55922 13932
rect 55953 13923 56011 13929
rect 55953 13920 55965 13923
rect 55916 13892 55965 13920
rect 55916 13880 55922 13892
rect 55953 13889 55965 13892
rect 55999 13889 56011 13923
rect 56612 13920 56640 14016
rect 58452 13929 58480 14028
rect 58437 13923 58495 13929
rect 56612 13892 57100 13920
rect 55953 13883 56011 13889
rect 52362 13812 52368 13864
rect 52420 13852 52426 13864
rect 52733 13855 52791 13861
rect 52733 13852 52745 13855
rect 52420 13824 52745 13852
rect 52420 13812 52426 13824
rect 52733 13821 52745 13824
rect 52779 13821 52791 13855
rect 52733 13815 52791 13821
rect 53282 13812 53288 13864
rect 53340 13812 53346 13864
rect 53466 13812 53472 13864
rect 53524 13812 53530 13864
rect 54110 13812 54116 13864
rect 54168 13852 54174 13864
rect 55033 13855 55091 13861
rect 55033 13852 55045 13855
rect 54168 13824 55045 13852
rect 54168 13812 54174 13824
rect 55033 13821 55045 13824
rect 55079 13821 55091 13855
rect 55033 13815 55091 13821
rect 55306 13812 55312 13864
rect 55364 13812 55370 13864
rect 56594 13812 56600 13864
rect 56652 13812 56658 13864
rect 57072 13861 57100 13892
rect 58437 13889 58449 13923
rect 58483 13889 58495 13923
rect 58437 13883 58495 13889
rect 57057 13855 57115 13861
rect 57057 13821 57069 13855
rect 57103 13821 57115 13855
rect 57057 13815 57115 13821
rect 52457 13787 52515 13793
rect 52457 13784 52469 13787
rect 51276 13756 52469 13784
rect 52457 13753 52469 13756
rect 52503 13784 52515 13787
rect 53098 13784 53104 13796
rect 52503 13756 53104 13784
rect 52503 13753 52515 13756
rect 52457 13747 52515 13753
rect 53098 13744 53104 13756
rect 53156 13744 53162 13796
rect 46532 13688 47072 13716
rect 46532 13676 46538 13688
rect 50706 13676 50712 13728
rect 50764 13676 50770 13728
rect 54018 13676 54024 13728
rect 54076 13716 54082 13728
rect 54113 13719 54171 13725
rect 54113 13716 54125 13719
rect 54076 13688 54125 13716
rect 54076 13676 54082 13688
rect 54113 13685 54125 13688
rect 54159 13685 54171 13719
rect 54113 13679 54171 13685
rect 56042 13676 56048 13728
rect 56100 13676 56106 13728
rect 57882 13676 57888 13728
rect 57940 13676 57946 13728
rect 1104 13626 58880 13648
rect 1104 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 22616 13626
rect 22668 13574 22680 13626
rect 22732 13574 22744 13626
rect 22796 13574 22808 13626
rect 22860 13574 22872 13626
rect 22924 13574 37060 13626
rect 37112 13574 37124 13626
rect 37176 13574 37188 13626
rect 37240 13574 37252 13626
rect 37304 13574 37316 13626
rect 37368 13574 51504 13626
rect 51556 13574 51568 13626
rect 51620 13574 51632 13626
rect 51684 13574 51696 13626
rect 51748 13574 51760 13626
rect 51812 13574 58880 13626
rect 1104 13552 58880 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2832 13484 2881 13512
rect 2832 13472 2838 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 3418 13472 3424 13524
rect 3476 13472 3482 13524
rect 4062 13472 4068 13524
rect 4120 13472 4126 13524
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4488 13484 4629 13512
rect 4488 13472 4494 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 4617 13475 4675 13481
rect 6362 13472 6368 13524
rect 6420 13512 6426 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 6420 13484 6561 13512
rect 6420 13472 6426 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 6549 13475 6607 13481
rect 6822 13472 6828 13524
rect 6880 13512 6886 13524
rect 7009 13515 7067 13521
rect 7009 13512 7021 13515
rect 6880 13484 7021 13512
rect 6880 13472 6886 13484
rect 7009 13481 7021 13484
rect 7055 13481 7067 13515
rect 7009 13475 7067 13481
rect 7374 13472 7380 13524
rect 7432 13472 7438 13524
rect 10686 13512 10692 13524
rect 10152 13484 10692 13512
rect 2746 13416 3832 13444
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 2746 13376 2774 13416
rect 2648 13348 2774 13376
rect 2648 13336 2654 13348
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2958 13308 2964 13320
rect 2547 13280 2964 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2958 13268 2964 13280
rect 3016 13308 3022 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 3016 13280 3249 13308
rect 3016 13268 3022 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 3252 13240 3280 13271
rect 3510 13268 3516 13320
rect 3568 13268 3574 13320
rect 3804 13317 3832 13416
rect 5902 13404 5908 13456
rect 5960 13404 5966 13456
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 6840 13376 6868 13472
rect 9769 13447 9827 13453
rect 9769 13444 9781 13447
rect 9692 13416 9781 13444
rect 9692 13385 9720 13416
rect 9769 13413 9781 13416
rect 9815 13413 9827 13447
rect 9769 13407 9827 13413
rect 5859 13348 6316 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4706 13268 4712 13320
rect 4764 13268 4770 13320
rect 6288 13317 6316 13348
rect 6656 13348 6868 13376
rect 9677 13379 9735 13385
rect 6656 13317 6684 13348
rect 9677 13345 9689 13379
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 10152 13317 10180 13484
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11514 13472 11520 13524
rect 11572 13472 11578 13524
rect 12158 13472 12164 13524
rect 12216 13472 12222 13524
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 15010 13512 15016 13524
rect 13412 13484 15016 13512
rect 13412 13472 13418 13484
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16632 13484 17540 13512
rect 16632 13472 16638 13484
rect 16025 13447 16083 13453
rect 10244 13416 11284 13444
rect 10244 13385 10272 13416
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 10459 13348 11100 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 6180 13311 6238 13317
rect 6180 13277 6192 13311
rect 6226 13277 6238 13311
rect 6180 13271 6238 13277
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 6640 13311 6698 13317
rect 6640 13308 6652 13311
rect 6319 13280 6652 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6640 13277 6652 13280
rect 6686 13277 6698 13311
rect 6640 13271 6698 13277
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13277 6791 13311
rect 6733 13271 6791 13277
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 3881 13243 3939 13249
rect 3881 13240 3893 13243
rect 3252 13212 3893 13240
rect 3881 13209 3893 13212
rect 3927 13209 3939 13243
rect 3881 13203 3939 13209
rect 4062 13200 4068 13252
rect 4120 13200 4126 13252
rect 6196 13240 6224 13271
rect 6748 13240 6776 13271
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 6196 13212 6776 13240
rect 6656 13184 6684 13212
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 8812 13212 10456 13240
rect 8812 13200 8818 13212
rect 10428 13184 10456 13212
rect 11072 13184 11100 13348
rect 6638 13132 6644 13184
rect 6696 13132 6702 13184
rect 9030 13132 9036 13184
rect 9088 13132 9094 13184
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 11054 13132 11060 13184
rect 11112 13132 11118 13184
rect 11256 13181 11284 13416
rect 16025 13413 16037 13447
rect 16071 13413 16083 13447
rect 16025 13407 16083 13413
rect 12621 13379 12679 13385
rect 12621 13345 12633 13379
rect 12667 13376 12679 13379
rect 12894 13376 12900 13388
rect 12667 13348 12900 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 12894 13336 12900 13348
rect 12952 13376 12958 13388
rect 13722 13376 13728 13388
rect 12952 13348 13728 13376
rect 12952 13336 12958 13348
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 14332 13348 14657 13376
rect 14332 13336 14338 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 16040 13376 16068 13407
rect 16298 13404 16304 13456
rect 16356 13444 16362 13456
rect 17512 13444 17540 13484
rect 18322 13472 18328 13524
rect 18380 13472 18386 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 18932 13484 20269 13512
rect 18932 13472 18938 13484
rect 20257 13481 20269 13484
rect 20303 13512 20315 13515
rect 21174 13512 21180 13524
rect 20303 13484 21180 13512
rect 20303 13481 20315 13484
rect 20257 13475 20315 13481
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 21361 13515 21419 13521
rect 21361 13481 21373 13515
rect 21407 13512 21419 13515
rect 22370 13512 22376 13524
rect 21407 13484 22376 13512
rect 21407 13481 21419 13484
rect 21361 13475 21419 13481
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 23290 13472 23296 13524
rect 23348 13472 23354 13524
rect 23474 13472 23480 13524
rect 23532 13472 23538 13524
rect 24397 13515 24455 13521
rect 24397 13481 24409 13515
rect 24443 13512 24455 13515
rect 24670 13512 24676 13524
rect 24443 13484 24676 13512
rect 24443 13481 24455 13484
rect 24397 13475 24455 13481
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 26050 13512 26056 13524
rect 24872 13484 26056 13512
rect 17586 13444 17592 13456
rect 16356 13416 16620 13444
rect 17512 13416 17592 13444
rect 16356 13404 16362 13416
rect 16482 13376 16488 13388
rect 16040 13348 16488 13376
rect 14645 13339 14703 13345
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 16592 13376 16620 13416
rect 17586 13404 17592 13416
rect 17644 13444 17650 13456
rect 17644 13416 19380 13444
rect 17644 13404 17650 13416
rect 16592 13348 17080 13376
rect 14918 13317 14924 13320
rect 14912 13308 14924 13317
rect 11532 13280 12434 13308
rect 14879 13280 14924 13308
rect 11532 13252 11560 13280
rect 11514 13200 11520 13252
rect 11572 13200 11578 13252
rect 12066 13200 12072 13252
rect 12124 13200 12130 13252
rect 12406 13240 12434 13280
rect 14912 13271 14924 13280
rect 14918 13268 14924 13271
rect 14976 13268 14982 13320
rect 17052 13317 17080 13348
rect 17310 13336 17316 13388
rect 17368 13336 17374 13388
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 18598 13376 18604 13388
rect 18095 13348 18604 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 18874 13336 18880 13388
rect 18932 13336 18938 13388
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 17126 13268 17132 13320
rect 17184 13317 17190 13320
rect 17184 13311 17233 13317
rect 17184 13277 17187 13311
rect 17221 13277 17233 13311
rect 17184 13271 17233 13277
rect 17184 13268 17190 13271
rect 18230 13268 18236 13320
rect 18288 13308 18294 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18288 13280 19257 13308
rect 18288 13268 18294 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 12986 13240 12992 13252
rect 12406 13212 12992 13240
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 18785 13243 18843 13249
rect 18785 13240 18797 13243
rect 18064 13212 18797 13240
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11606 13172 11612 13184
rect 11287 13144 11612 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 16393 13175 16451 13181
rect 16393 13141 16405 13175
rect 16439 13172 16451 13175
rect 18064 13172 18092 13212
rect 18785 13209 18797 13212
rect 18831 13209 18843 13243
rect 19352 13240 19380 13416
rect 20346 13404 20352 13456
rect 20404 13404 20410 13456
rect 20714 13404 20720 13456
rect 20772 13444 20778 13456
rect 20772 13416 21036 13444
rect 20772 13404 20778 13416
rect 19794 13336 19800 13388
rect 19852 13336 19858 13388
rect 20806 13336 20812 13388
rect 20864 13336 20870 13388
rect 21008 13385 21036 13416
rect 22756 13416 24256 13444
rect 22756 13385 22784 13416
rect 24228 13388 24256 13416
rect 20993 13379 21051 13385
rect 20993 13345 21005 13379
rect 21039 13376 21051 13379
rect 22741 13379 22799 13385
rect 21039 13348 21772 13376
rect 21039 13345 21051 13348
rect 20993 13339 21051 13345
rect 20824 13308 20852 13336
rect 21634 13308 21640 13320
rect 20824 13280 21640 13308
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 21744 13308 21772 13348
rect 22741 13345 22753 13379
rect 22787 13345 22799 13379
rect 24029 13379 24087 13385
rect 24029 13376 24041 13379
rect 22741 13339 22799 13345
rect 23768 13348 24041 13376
rect 21744 13280 22324 13308
rect 19794 13240 19800 13252
rect 19352 13212 19800 13240
rect 18785 13203 18843 13209
rect 19794 13200 19800 13212
rect 19852 13200 19858 13252
rect 16439 13144 18092 13172
rect 16439 13141 16451 13144
rect 16393 13135 16451 13141
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 18196 13144 18705 13172
rect 18196 13132 18202 13144
rect 18693 13141 18705 13144
rect 18739 13141 18751 13175
rect 18693 13135 18751 13141
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 22186 13172 22192 13184
rect 20772 13144 22192 13172
rect 20772 13132 20778 13144
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 22296 13172 22324 13280
rect 22462 13268 22468 13320
rect 22520 13317 22526 13320
rect 22520 13308 22532 13317
rect 23768 13308 23796 13348
rect 24029 13345 24041 13348
rect 24075 13345 24087 13379
rect 24029 13339 24087 13345
rect 24210 13336 24216 13388
rect 24268 13336 24274 13388
rect 24872 13385 24900 13484
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 26786 13472 26792 13524
rect 26844 13512 26850 13524
rect 27157 13515 27215 13521
rect 27157 13512 27169 13515
rect 26844 13484 27169 13512
rect 26844 13472 26850 13484
rect 27157 13481 27169 13484
rect 27203 13481 27215 13515
rect 27157 13475 27215 13481
rect 29365 13515 29423 13521
rect 29365 13481 29377 13515
rect 29411 13512 29423 13515
rect 29454 13512 29460 13524
rect 29411 13484 29460 13512
rect 29411 13481 29423 13484
rect 29365 13475 29423 13481
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 34238 13472 34244 13524
rect 34296 13512 34302 13524
rect 34333 13515 34391 13521
rect 34333 13512 34345 13515
rect 34296 13484 34345 13512
rect 34296 13472 34302 13484
rect 34333 13481 34345 13484
rect 34379 13481 34391 13515
rect 34333 13475 34391 13481
rect 35805 13515 35863 13521
rect 35805 13481 35817 13515
rect 35851 13512 35863 13515
rect 36630 13512 36636 13524
rect 35851 13484 36636 13512
rect 35851 13481 35863 13484
rect 35805 13475 35863 13481
rect 36630 13472 36636 13484
rect 36688 13472 36694 13524
rect 37734 13512 37740 13524
rect 37016 13484 37740 13512
rect 25130 13444 25136 13456
rect 24964 13416 25136 13444
rect 24964 13388 24992 13416
rect 25130 13404 25136 13416
rect 25188 13404 25194 13456
rect 26326 13404 26332 13456
rect 26384 13444 26390 13456
rect 26421 13447 26479 13453
rect 26421 13444 26433 13447
rect 26384 13416 26433 13444
rect 26384 13404 26390 13416
rect 26421 13413 26433 13416
rect 26467 13413 26479 13447
rect 33042 13444 33048 13456
rect 26421 13407 26479 13413
rect 32232 13416 33048 13444
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 24946 13336 24952 13388
rect 25004 13336 25010 13388
rect 26007 13379 26065 13385
rect 26007 13376 26019 13379
rect 25056 13348 26019 13376
rect 22520 13280 22565 13308
rect 23308 13280 23796 13308
rect 23845 13311 23903 13317
rect 22520 13271 22532 13280
rect 22520 13268 22526 13271
rect 23308 13252 23336 13280
rect 23845 13277 23857 13311
rect 23891 13308 23903 13311
rect 24486 13308 24492 13320
rect 23891 13280 24492 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 24486 13268 24492 13280
rect 24544 13308 24550 13320
rect 25056 13308 25084 13348
rect 26007 13345 26019 13348
rect 26053 13345 26065 13379
rect 26007 13339 26065 13345
rect 26142 13336 26148 13388
rect 26200 13336 26206 13388
rect 27246 13336 27252 13388
rect 27304 13376 27310 13388
rect 27709 13379 27767 13385
rect 27709 13376 27721 13379
rect 27304 13348 27721 13376
rect 27304 13336 27310 13348
rect 27709 13345 27721 13348
rect 27755 13345 27767 13379
rect 27709 13339 27767 13345
rect 24544 13280 25084 13308
rect 24544 13268 24550 13280
rect 25866 13268 25872 13320
rect 25924 13268 25930 13320
rect 26881 13311 26939 13317
rect 26881 13277 26893 13311
rect 26927 13277 26939 13311
rect 26881 13271 26939 13277
rect 27065 13311 27123 13317
rect 27065 13277 27077 13311
rect 27111 13308 27123 13311
rect 27430 13308 27436 13320
rect 27111 13280 27436 13308
rect 27111 13277 27123 13280
rect 27065 13271 27123 13277
rect 23290 13200 23296 13252
rect 23348 13200 23354 13252
rect 26896 13240 26924 13271
rect 27430 13268 27436 13280
rect 27488 13308 27494 13320
rect 27985 13311 28043 13317
rect 27985 13308 27997 13311
rect 27488 13280 27997 13308
rect 27488 13268 27494 13280
rect 27985 13277 27997 13280
rect 28031 13277 28043 13311
rect 27985 13271 28043 13277
rect 28534 13268 28540 13320
rect 28592 13268 28598 13320
rect 28626 13268 28632 13320
rect 28684 13308 28690 13320
rect 31849 13311 31907 13317
rect 31849 13308 31861 13311
rect 28684 13280 31861 13308
rect 28684 13268 28690 13280
rect 31849 13277 31861 13280
rect 31895 13308 31907 13311
rect 32125 13311 32183 13317
rect 32125 13308 32137 13311
rect 31895 13280 32137 13308
rect 31895 13277 31907 13280
rect 31849 13271 31907 13277
rect 32125 13277 32137 13280
rect 32171 13308 32183 13311
rect 32232 13308 32260 13416
rect 33042 13404 33048 13416
rect 33100 13404 33106 13456
rect 32582 13336 32588 13388
rect 32640 13336 32646 13388
rect 33413 13379 33471 13385
rect 33413 13376 33425 13379
rect 33152 13348 33425 13376
rect 32171 13280 32260 13308
rect 32171 13277 32183 13280
rect 32125 13271 32183 13277
rect 33152 13252 33180 13348
rect 33413 13345 33425 13348
rect 33459 13345 33471 13379
rect 33413 13339 33471 13345
rect 33229 13311 33287 13317
rect 33229 13277 33241 13311
rect 33275 13308 33287 13311
rect 34256 13308 34284 13472
rect 37016 13456 37044 13484
rect 37734 13472 37740 13484
rect 37792 13512 37798 13524
rect 39114 13512 39120 13524
rect 37792 13484 39120 13512
rect 37792 13472 37798 13484
rect 39114 13472 39120 13484
rect 39172 13472 39178 13524
rect 41138 13472 41144 13524
rect 41196 13472 41202 13524
rect 41690 13472 41696 13524
rect 41748 13512 41754 13524
rect 42058 13512 42064 13524
rect 41748 13484 42064 13512
rect 41748 13472 41754 13484
rect 42058 13472 42064 13484
rect 42116 13472 42122 13524
rect 44637 13515 44695 13521
rect 44637 13481 44649 13515
rect 44683 13512 44695 13515
rect 45554 13512 45560 13524
rect 44683 13484 45560 13512
rect 44683 13481 44695 13484
rect 44637 13475 44695 13481
rect 45554 13472 45560 13484
rect 45612 13472 45618 13524
rect 47029 13515 47087 13521
rect 47029 13481 47041 13515
rect 47075 13512 47087 13515
rect 47578 13512 47584 13524
rect 47075 13484 47584 13512
rect 47075 13481 47087 13484
rect 47029 13475 47087 13481
rect 47578 13472 47584 13484
rect 47636 13472 47642 13524
rect 51902 13472 51908 13524
rect 51960 13512 51966 13524
rect 53561 13515 53619 13521
rect 53561 13512 53573 13515
rect 51960 13484 53573 13512
rect 51960 13472 51966 13484
rect 53561 13481 53573 13484
rect 53607 13481 53619 13515
rect 53561 13475 53619 13481
rect 55125 13515 55183 13521
rect 55125 13481 55137 13515
rect 55171 13512 55183 13515
rect 55306 13512 55312 13524
rect 55171 13484 55312 13512
rect 55171 13481 55183 13484
rect 55125 13475 55183 13481
rect 35986 13444 35992 13456
rect 34348 13416 35992 13444
rect 34348 13388 34376 13416
rect 35986 13404 35992 13416
rect 36044 13404 36050 13456
rect 36998 13404 37004 13456
rect 37056 13404 37062 13456
rect 47394 13404 47400 13456
rect 47452 13404 47458 13456
rect 48777 13447 48835 13453
rect 48777 13413 48789 13447
rect 48823 13444 48835 13447
rect 48958 13444 48964 13456
rect 48823 13416 48964 13444
rect 48823 13413 48835 13416
rect 48777 13407 48835 13413
rect 48958 13404 48964 13416
rect 49016 13444 49022 13456
rect 49697 13447 49755 13453
rect 49697 13444 49709 13447
rect 49016 13416 49709 13444
rect 49016 13404 49022 13416
rect 49697 13413 49709 13416
rect 49743 13413 49755 13447
rect 51350 13444 51356 13456
rect 49697 13407 49755 13413
rect 50356 13416 51356 13444
rect 34330 13336 34336 13388
rect 34388 13336 34394 13388
rect 35250 13336 35256 13388
rect 35308 13336 35314 13388
rect 35434 13336 35440 13388
rect 35492 13336 35498 13388
rect 35710 13336 35716 13388
rect 35768 13376 35774 13388
rect 36449 13379 36507 13385
rect 36449 13376 36461 13379
rect 35768 13348 36461 13376
rect 35768 13336 35774 13348
rect 36449 13345 36461 13348
rect 36495 13345 36507 13379
rect 36449 13339 36507 13345
rect 36722 13336 36728 13388
rect 36780 13336 36786 13388
rect 37461 13379 37519 13385
rect 37461 13345 37473 13379
rect 37507 13376 37519 13379
rect 37918 13376 37924 13388
rect 37507 13348 37924 13376
rect 37507 13345 37519 13348
rect 37461 13339 37519 13345
rect 37918 13336 37924 13348
rect 37976 13336 37982 13388
rect 42150 13336 42156 13388
rect 42208 13376 42214 13388
rect 42337 13379 42395 13385
rect 42337 13376 42349 13379
rect 42208 13348 42349 13376
rect 42208 13336 42214 13348
rect 42337 13345 42349 13348
rect 42383 13376 42395 13379
rect 42610 13376 42616 13388
rect 42383 13348 42616 13376
rect 42383 13345 42395 13348
rect 42337 13339 42395 13345
rect 42610 13336 42616 13348
rect 42668 13336 42674 13388
rect 47412 13376 47440 13404
rect 48222 13376 48228 13388
rect 47412 13348 48228 13376
rect 48222 13336 48228 13348
rect 48280 13336 48286 13388
rect 48314 13336 48320 13388
rect 48372 13385 48378 13388
rect 48372 13379 48421 13385
rect 48372 13345 48375 13379
rect 48409 13345 48421 13379
rect 48372 13339 48421 13345
rect 49237 13379 49295 13385
rect 49237 13345 49249 13379
rect 49283 13376 49295 13379
rect 49326 13376 49332 13388
rect 49283 13348 49332 13376
rect 49283 13345 49295 13348
rect 49237 13339 49295 13345
rect 48372 13336 48378 13339
rect 49326 13336 49332 13348
rect 49384 13336 49390 13388
rect 50356 13385 50384 13416
rect 51350 13404 51356 13416
rect 51408 13404 51414 13456
rect 52549 13447 52607 13453
rect 52549 13413 52561 13447
rect 52595 13444 52607 13447
rect 53282 13444 53288 13456
rect 52595 13416 53288 13444
rect 52595 13413 52607 13416
rect 52549 13407 52607 13413
rect 53282 13404 53288 13416
rect 53340 13404 53346 13456
rect 50341 13379 50399 13385
rect 50341 13345 50353 13379
rect 50387 13345 50399 13379
rect 50341 13339 50399 13345
rect 50433 13379 50491 13385
rect 50433 13345 50445 13379
rect 50479 13376 50491 13379
rect 50706 13376 50712 13388
rect 50479 13348 50712 13376
rect 50479 13345 50491 13348
rect 50433 13339 50491 13345
rect 36630 13317 36636 13320
rect 33275 13280 34284 13308
rect 36608 13311 36636 13317
rect 33275 13277 33287 13280
rect 33229 13271 33287 13277
rect 36608 13277 36620 13311
rect 36608 13271 36636 13277
rect 36630 13268 36636 13271
rect 36688 13268 36694 13320
rect 37642 13268 37648 13320
rect 37700 13268 37706 13320
rect 39022 13268 39028 13320
rect 39080 13308 39086 13320
rect 39117 13311 39175 13317
rect 39117 13308 39129 13311
rect 39080 13280 39129 13308
rect 39080 13268 39086 13280
rect 39117 13277 39129 13280
rect 39163 13308 39175 13311
rect 39393 13311 39451 13317
rect 39393 13308 39405 13311
rect 39163 13280 39405 13308
rect 39163 13277 39175 13280
rect 39117 13271 39175 13277
rect 39393 13277 39405 13280
rect 39439 13277 39451 13311
rect 43073 13311 43131 13317
rect 43073 13308 43085 13311
rect 39393 13271 39451 13277
rect 41386 13280 43085 13308
rect 41386 13252 41414 13280
rect 43073 13277 43085 13280
rect 43119 13277 43131 13311
rect 43073 13271 43131 13277
rect 43254 13268 43260 13320
rect 43312 13308 43318 13320
rect 44082 13308 44088 13320
rect 43312 13280 44088 13308
rect 43312 13268 43318 13280
rect 44082 13268 44088 13280
rect 44140 13308 44146 13320
rect 45281 13311 45339 13317
rect 45281 13308 45293 13311
rect 44140 13280 45293 13308
rect 44140 13268 44146 13280
rect 45281 13277 45293 13280
rect 45327 13308 45339 13311
rect 45554 13308 45560 13320
rect 45327 13280 45560 13308
rect 45327 13277 45339 13280
rect 45281 13271 45339 13277
rect 45554 13268 45560 13280
rect 45612 13308 45618 13320
rect 45922 13317 45928 13320
rect 45649 13311 45707 13317
rect 45649 13308 45661 13311
rect 45612 13280 45661 13308
rect 45612 13268 45618 13280
rect 45649 13277 45661 13280
rect 45695 13277 45707 13311
rect 45916 13308 45928 13317
rect 45883 13280 45928 13308
rect 45649 13271 45707 13277
rect 45916 13271 45928 13280
rect 27522 13240 27528 13252
rect 26896 13212 27528 13240
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 29546 13200 29552 13252
rect 29604 13200 29610 13252
rect 31726 13212 32720 13240
rect 22922 13172 22928 13184
rect 22296 13144 22928 13172
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 23937 13175 23995 13181
rect 23937 13141 23949 13175
rect 23983 13172 23995 13175
rect 24765 13175 24823 13181
rect 24765 13172 24777 13175
rect 23983 13144 24777 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 24765 13141 24777 13144
rect 24811 13172 24823 13175
rect 25130 13172 25136 13184
rect 24811 13144 25136 13172
rect 24811 13141 24823 13144
rect 24765 13135 24823 13141
rect 25130 13132 25136 13144
rect 25188 13132 25194 13184
rect 25225 13175 25283 13181
rect 25225 13141 25237 13175
rect 25271 13172 25283 13175
rect 26602 13172 26608 13184
rect 25271 13144 26608 13172
rect 25271 13141 25283 13144
rect 25225 13135 25283 13141
rect 26602 13132 26608 13144
rect 26660 13132 26666 13184
rect 27338 13132 27344 13184
rect 27396 13172 27402 13184
rect 27617 13175 27675 13181
rect 27617 13172 27629 13175
rect 27396 13144 27629 13172
rect 27396 13132 27402 13144
rect 27617 13141 27629 13144
rect 27663 13141 27675 13175
rect 27617 13135 27675 13141
rect 30742 13132 30748 13184
rect 30800 13172 30806 13184
rect 30837 13175 30895 13181
rect 30837 13172 30849 13175
rect 30800 13144 30849 13172
rect 30800 13132 30806 13144
rect 30837 13141 30849 13144
rect 30883 13172 30895 13175
rect 31726 13172 31754 13212
rect 30883 13144 31754 13172
rect 32692 13172 32720 13212
rect 33134 13200 33140 13252
rect 33192 13200 33198 13252
rect 34256 13212 36032 13240
rect 34256 13172 34284 13212
rect 32692 13144 34284 13172
rect 30883 13141 30895 13144
rect 30837 13135 30895 13141
rect 34790 13132 34796 13184
rect 34848 13132 34854 13184
rect 35158 13132 35164 13184
rect 35216 13132 35222 13184
rect 36004 13172 36032 13212
rect 37476 13212 38792 13240
rect 37476 13172 37504 13212
rect 36004 13144 37504 13172
rect 37737 13175 37795 13181
rect 37737 13141 37749 13175
rect 37783 13172 37795 13175
rect 38562 13172 38568 13184
rect 37783 13144 38568 13172
rect 37783 13141 37795 13144
rect 37737 13135 37795 13141
rect 38562 13132 38568 13144
rect 38620 13132 38626 13184
rect 38764 13172 38792 13212
rect 38838 13200 38844 13252
rect 38896 13249 38902 13252
rect 38896 13203 38908 13249
rect 39666 13240 39672 13252
rect 38948 13212 39672 13240
rect 38896 13200 38902 13203
rect 38948 13172 38976 13212
rect 39666 13200 39672 13212
rect 39724 13240 39730 13252
rect 39853 13243 39911 13249
rect 39853 13240 39865 13243
rect 39724 13212 39865 13240
rect 39724 13200 39730 13212
rect 39853 13209 39865 13212
rect 39899 13209 39911 13243
rect 39853 13203 39911 13209
rect 41322 13200 41328 13252
rect 41380 13212 41414 13252
rect 41380 13200 41386 13212
rect 41966 13200 41972 13252
rect 42024 13240 42030 13252
rect 42061 13243 42119 13249
rect 42061 13240 42073 13243
rect 42024 13212 42073 13240
rect 42024 13200 42030 13212
rect 42061 13209 42073 13212
rect 42107 13240 42119 13243
rect 42610 13240 42616 13252
rect 42107 13212 42616 13240
rect 42107 13209 42119 13212
rect 42061 13203 42119 13209
rect 42610 13200 42616 13212
rect 42668 13200 42674 13252
rect 43524 13243 43582 13249
rect 43524 13209 43536 13243
rect 43570 13240 43582 13243
rect 44266 13240 44272 13252
rect 43570 13212 44272 13240
rect 43570 13209 43582 13212
rect 43524 13203 43582 13209
rect 44266 13200 44272 13212
rect 44324 13200 44330 13252
rect 45664 13240 45692 13271
rect 45922 13268 45928 13271
rect 45980 13268 45986 13320
rect 46198 13268 46204 13320
rect 46256 13268 46262 13320
rect 48498 13268 48504 13320
rect 48556 13268 48562 13320
rect 49421 13311 49479 13317
rect 49421 13277 49433 13311
rect 49467 13308 49479 13311
rect 50448 13308 50476 13339
rect 50706 13336 50712 13348
rect 50764 13336 50770 13388
rect 53098 13336 53104 13388
rect 53156 13336 53162 13388
rect 53576 13376 53604 13475
rect 55306 13472 55312 13484
rect 55364 13472 55370 13524
rect 58253 13515 58311 13521
rect 58253 13481 58265 13515
rect 58299 13512 58311 13515
rect 58434 13512 58440 13524
rect 58299 13484 58440 13512
rect 58299 13481 58311 13484
rect 58253 13475 58311 13481
rect 58434 13472 58440 13484
rect 58492 13472 58498 13524
rect 53745 13379 53803 13385
rect 53745 13376 53757 13379
rect 53576 13348 53757 13376
rect 53745 13345 53757 13348
rect 53791 13345 53803 13379
rect 53745 13339 53803 13345
rect 51537 13311 51595 13317
rect 51537 13308 51549 13311
rect 49467 13280 50476 13308
rect 50908 13280 51549 13308
rect 49467 13277 49479 13280
rect 49421 13271 49479 13277
rect 46216 13240 46244 13268
rect 45664 13212 46244 13240
rect 49234 13200 49240 13252
rect 49292 13240 49298 13252
rect 50525 13243 50583 13249
rect 50525 13240 50537 13243
rect 49292 13212 50537 13240
rect 49292 13200 49298 13212
rect 50525 13209 50537 13212
rect 50571 13209 50583 13243
rect 50525 13203 50583 13209
rect 38764 13144 38976 13172
rect 41690 13132 41696 13184
rect 41748 13132 41754 13184
rect 42153 13175 42211 13181
rect 42153 13141 42165 13175
rect 42199 13172 42211 13175
rect 42334 13172 42340 13184
rect 42199 13144 42340 13172
rect 42199 13141 42211 13144
rect 42153 13135 42211 13141
rect 42334 13132 42340 13144
rect 42392 13172 42398 13184
rect 42521 13175 42579 13181
rect 42521 13172 42533 13175
rect 42392 13144 42533 13172
rect 42392 13132 42398 13144
rect 42521 13141 42533 13144
rect 42567 13141 42579 13175
rect 42521 13135 42579 13141
rect 47578 13132 47584 13184
rect 47636 13132 47642 13184
rect 48406 13132 48412 13184
rect 48464 13172 48470 13184
rect 49252 13172 49280 13200
rect 50908 13181 50936 13280
rect 51537 13277 51549 13280
rect 51583 13277 51595 13311
rect 51537 13271 51595 13277
rect 52454 13268 52460 13320
rect 52512 13268 52518 13320
rect 53760 13308 53788 13339
rect 55306 13308 55312 13320
rect 53760 13280 55312 13308
rect 55306 13268 55312 13280
rect 55364 13308 55370 13320
rect 56870 13308 56876 13320
rect 55364 13280 56876 13308
rect 55364 13268 55370 13280
rect 56870 13268 56876 13280
rect 56928 13268 56934 13320
rect 57140 13311 57198 13317
rect 57140 13277 57152 13311
rect 57186 13308 57198 13311
rect 57882 13308 57888 13320
rect 57186 13280 57888 13308
rect 57186 13277 57198 13280
rect 57140 13271 57198 13277
rect 57882 13268 57888 13280
rect 57940 13268 57946 13320
rect 52917 13243 52975 13249
rect 52917 13209 52929 13243
rect 52963 13240 52975 13243
rect 53190 13240 53196 13252
rect 52963 13212 53196 13240
rect 52963 13209 52975 13212
rect 52917 13203 52975 13209
rect 53190 13200 53196 13212
rect 53248 13240 53254 13252
rect 54012 13243 54070 13249
rect 53248 13212 53880 13240
rect 53248 13200 53254 13212
rect 48464 13144 49280 13172
rect 50893 13175 50951 13181
rect 48464 13132 48470 13144
rect 50893 13141 50905 13175
rect 50939 13141 50951 13175
rect 50893 13135 50951 13141
rect 50982 13132 50988 13184
rect 51040 13132 51046 13184
rect 51810 13132 51816 13184
rect 51868 13132 51874 13184
rect 53009 13175 53067 13181
rect 53009 13141 53021 13175
rect 53055 13172 53067 13175
rect 53742 13172 53748 13184
rect 53055 13144 53748 13172
rect 53055 13141 53067 13144
rect 53009 13135 53067 13141
rect 53742 13132 53748 13144
rect 53800 13132 53806 13184
rect 53852 13172 53880 13212
rect 54012 13209 54024 13243
rect 54058 13240 54070 13243
rect 54294 13240 54300 13252
rect 54058 13212 54300 13240
rect 54058 13209 54070 13212
rect 54012 13203 54070 13209
rect 54294 13200 54300 13212
rect 54352 13200 54358 13252
rect 55576 13243 55634 13249
rect 55576 13209 55588 13243
rect 55622 13240 55634 13243
rect 56042 13240 56048 13252
rect 55622 13212 56048 13240
rect 55622 13209 55634 13212
rect 55576 13203 55634 13209
rect 56042 13200 56048 13212
rect 56100 13200 56106 13252
rect 55122 13172 55128 13184
rect 53852 13144 55128 13172
rect 55122 13132 55128 13144
rect 55180 13132 55186 13184
rect 56686 13132 56692 13184
rect 56744 13132 56750 13184
rect 1104 13082 59040 13104
rect 1104 13030 15394 13082
rect 15446 13030 15458 13082
rect 15510 13030 15522 13082
rect 15574 13030 15586 13082
rect 15638 13030 15650 13082
rect 15702 13030 29838 13082
rect 29890 13030 29902 13082
rect 29954 13030 29966 13082
rect 30018 13030 30030 13082
rect 30082 13030 30094 13082
rect 30146 13030 44282 13082
rect 44334 13030 44346 13082
rect 44398 13030 44410 13082
rect 44462 13030 44474 13082
rect 44526 13030 44538 13082
rect 44590 13030 58726 13082
rect 58778 13030 58790 13082
rect 58842 13030 58854 13082
rect 58906 13030 58918 13082
rect 58970 13030 58982 13082
rect 59034 13030 59040 13082
rect 1104 13008 59040 13030
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12968 3571 12971
rect 4062 12968 4068 12980
rect 3559 12940 4068 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 7285 12971 7343 12977
rect 7285 12968 7297 12971
rect 6840 12940 7297 12968
rect 6454 12860 6460 12912
rect 6512 12900 6518 12912
rect 6742 12903 6800 12909
rect 6742 12900 6754 12903
rect 6512 12872 6754 12900
rect 6512 12860 6518 12872
rect 6742 12869 6754 12872
rect 6788 12900 6800 12903
rect 6840 12900 6868 12940
rect 7285 12937 7297 12940
rect 7331 12937 7343 12971
rect 7285 12931 7343 12937
rect 7469 12971 7527 12977
rect 7469 12937 7481 12971
rect 7515 12937 7527 12971
rect 7469 12931 7527 12937
rect 7101 12903 7159 12909
rect 7101 12900 7113 12903
rect 6788 12872 6868 12900
rect 6932 12872 7113 12900
rect 6788 12869 6800 12872
rect 6742 12863 6800 12869
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 6638 12832 6644 12844
rect 6411 12804 6644 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6638 12792 6644 12804
rect 6696 12832 6702 12844
rect 6932 12832 6960 12872
rect 7101 12869 7113 12872
rect 7147 12869 7159 12903
rect 7484 12900 7512 12931
rect 16298 12928 16304 12980
rect 16356 12928 16362 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 16853 12971 16911 12977
rect 16853 12968 16865 12971
rect 16448 12940 16865 12968
rect 16448 12928 16454 12940
rect 16853 12937 16865 12940
rect 16899 12937 16911 12971
rect 16853 12931 16911 12937
rect 17313 12971 17371 12977
rect 17313 12937 17325 12971
rect 17359 12968 17371 12971
rect 17954 12968 17960 12980
rect 17359 12940 17960 12968
rect 17359 12937 17371 12940
rect 17313 12931 17371 12937
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 21048 12940 21097 12968
rect 21048 12928 21054 12940
rect 21085 12937 21097 12940
rect 21131 12937 21143 12971
rect 21085 12931 21143 12937
rect 21910 12928 21916 12980
rect 21968 12968 21974 12980
rect 22557 12971 22615 12977
rect 22557 12968 22569 12971
rect 21968 12940 22569 12968
rect 21968 12928 21974 12940
rect 22557 12937 22569 12940
rect 22603 12937 22615 12971
rect 22557 12931 22615 12937
rect 22922 12928 22928 12980
rect 22980 12968 22986 12980
rect 23661 12971 23719 12977
rect 23661 12968 23673 12971
rect 22980 12940 23673 12968
rect 22980 12928 22986 12940
rect 23661 12937 23673 12940
rect 23707 12968 23719 12971
rect 24946 12968 24952 12980
rect 23707 12940 24952 12968
rect 23707 12937 23719 12940
rect 23661 12931 23719 12937
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 25130 12928 25136 12980
rect 25188 12968 25194 12980
rect 26789 12971 26847 12977
rect 25188 12940 26280 12968
rect 25188 12928 25194 12940
rect 9214 12900 9220 12912
rect 7484 12872 9220 12900
rect 7101 12863 7159 12869
rect 9214 12860 9220 12872
rect 9272 12860 9278 12912
rect 10134 12900 10140 12912
rect 9692 12872 10140 12900
rect 6696 12804 6960 12832
rect 7009 12835 7067 12841
rect 6696 12792 6702 12804
rect 7009 12801 7021 12835
rect 7055 12832 7067 12835
rect 9692 12832 9720 12872
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 13354 12900 13360 12912
rect 11112 12872 13360 12900
rect 11112 12860 11118 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 18448 12903 18506 12909
rect 18448 12869 18460 12903
rect 18494 12900 18506 12903
rect 18966 12900 18972 12912
rect 18494 12872 18972 12900
rect 18494 12869 18506 12872
rect 18448 12863 18506 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 19720 12872 23612 12900
rect 19720 12844 19748 12872
rect 7055 12804 9720 12832
rect 7055 12801 7067 12804
rect 7009 12795 7067 12801
rect 9766 12792 9772 12844
rect 9824 12841 9830 12844
rect 9824 12795 9836 12841
rect 9824 12792 9830 12795
rect 10410 12792 10416 12844
rect 10468 12792 10474 12844
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 12894 12792 12900 12844
rect 12952 12792 12958 12844
rect 13630 12832 13636 12844
rect 13464 12804 13636 12832
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3786 12764 3792 12776
rect 3099 12736 3792 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 10962 12764 10968 12776
rect 10091 12736 10968 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 3418 12656 3424 12708
rect 3476 12656 3482 12708
rect 8036 12696 8064 12727
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 12216 12736 12357 12764
rect 12216 12724 12222 12736
rect 12345 12733 12357 12736
rect 12391 12764 12403 12767
rect 13464 12764 13492 12804
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 14728 12835 14786 12841
rect 14728 12801 14740 12835
rect 14774 12832 14786 12835
rect 15010 12832 15016 12844
rect 14774 12804 15016 12832
rect 14774 12801 14786 12804
rect 14728 12795 14786 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 18693 12835 18751 12841
rect 15160 12804 18644 12832
rect 15160 12792 15166 12804
rect 12391 12736 13492 12764
rect 13541 12767 13599 12773
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 13541 12733 13553 12767
rect 13587 12764 13599 12767
rect 13814 12764 13820 12776
rect 13587 12736 13820 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14458 12724 14464 12776
rect 14516 12724 14522 12776
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 17126 12764 17132 12776
rect 15620 12736 17132 12764
rect 15620 12724 15626 12736
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 18616 12764 18644 12804
rect 18693 12801 18705 12835
rect 18739 12832 18751 12835
rect 19702 12832 19708 12844
rect 18739 12804 19708 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 19702 12792 19708 12804
rect 19760 12792 19766 12844
rect 19978 12841 19984 12844
rect 19972 12832 19984 12841
rect 19939 12804 19984 12832
rect 19972 12795 19984 12804
rect 19978 12792 19984 12795
rect 20036 12792 20042 12844
rect 22462 12792 22468 12844
rect 22520 12792 22526 12844
rect 23584 12832 23612 12872
rect 23768 12872 25452 12900
rect 23768 12841 23796 12872
rect 24026 12841 24032 12844
rect 23753 12835 23811 12841
rect 23753 12832 23765 12835
rect 23584 12804 23765 12832
rect 23753 12801 23765 12804
rect 23799 12801 23811 12835
rect 24020 12832 24032 12841
rect 23987 12804 24032 12832
rect 23753 12795 23811 12801
rect 24020 12795 24032 12804
rect 24026 12792 24032 12795
rect 24084 12792 24090 12844
rect 25424 12841 25452 12872
rect 25409 12835 25467 12841
rect 25409 12801 25421 12835
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 25676 12835 25734 12841
rect 25676 12801 25688 12835
rect 25722 12832 25734 12835
rect 26142 12832 26148 12844
rect 25722 12804 26148 12832
rect 25722 12801 25734 12804
rect 25676 12795 25734 12801
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 26252 12832 26280 12940
rect 26789 12937 26801 12971
rect 26835 12968 26847 12971
rect 28534 12968 28540 12980
rect 26835 12940 28540 12968
rect 26835 12937 26847 12940
rect 26789 12931 26847 12937
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 28626 12928 28632 12980
rect 28684 12928 28690 12980
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 29917 12971 29975 12977
rect 29917 12968 29929 12971
rect 29788 12940 29929 12968
rect 29788 12928 29794 12940
rect 29917 12937 29929 12940
rect 29963 12937 29975 12971
rect 29917 12931 29975 12937
rect 33502 12928 33508 12980
rect 33560 12928 33566 12980
rect 35250 12928 35256 12980
rect 35308 12928 35314 12980
rect 35805 12971 35863 12977
rect 35805 12937 35817 12971
rect 35851 12968 35863 12971
rect 36078 12968 36084 12980
rect 35851 12940 36084 12968
rect 35851 12937 35863 12940
rect 35805 12931 35863 12937
rect 36078 12928 36084 12940
rect 36136 12928 36142 12980
rect 36265 12971 36323 12977
rect 36265 12937 36277 12971
rect 36311 12968 36323 12971
rect 36722 12968 36728 12980
rect 36311 12940 36728 12968
rect 36311 12937 36323 12940
rect 36265 12931 36323 12937
rect 36722 12928 36728 12940
rect 36780 12928 36786 12980
rect 36814 12928 36820 12980
rect 36872 12968 36878 12980
rect 36909 12971 36967 12977
rect 36909 12968 36921 12971
rect 36872 12940 36921 12968
rect 36872 12928 36878 12940
rect 36909 12937 36921 12940
rect 36955 12968 36967 12971
rect 36998 12968 37004 12980
rect 36955 12940 37004 12968
rect 36955 12937 36967 12940
rect 36909 12931 36967 12937
rect 36998 12928 37004 12940
rect 37056 12928 37062 12980
rect 38654 12928 38660 12980
rect 38712 12928 38718 12980
rect 38749 12971 38807 12977
rect 38749 12937 38761 12971
rect 38795 12968 38807 12971
rect 38838 12968 38844 12980
rect 38795 12940 38844 12968
rect 38795 12937 38807 12940
rect 38749 12931 38807 12937
rect 38838 12928 38844 12940
rect 38896 12928 38902 12980
rect 39666 12928 39672 12980
rect 39724 12928 39730 12980
rect 41046 12928 41052 12980
rect 41104 12968 41110 12980
rect 41233 12971 41291 12977
rect 41233 12968 41245 12971
rect 41104 12940 41245 12968
rect 41104 12928 41110 12940
rect 41233 12937 41245 12940
rect 41279 12937 41291 12971
rect 41233 12931 41291 12937
rect 42702 12928 42708 12980
rect 42760 12928 42766 12980
rect 43254 12928 43260 12980
rect 43312 12928 43318 12980
rect 45554 12928 45560 12980
rect 45612 12928 45618 12980
rect 47578 12928 47584 12980
rect 47636 12968 47642 12980
rect 49605 12971 49663 12977
rect 47636 12940 48912 12968
rect 47636 12928 47642 12940
rect 26694 12860 26700 12912
rect 26752 12900 26758 12912
rect 26752 12872 28488 12900
rect 26752 12860 26758 12872
rect 27338 12832 27344 12844
rect 26252 12804 27344 12832
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 27430 12792 27436 12844
rect 27488 12792 27494 12844
rect 28460 12841 28488 12872
rect 28445 12835 28503 12841
rect 28445 12801 28457 12835
rect 28491 12832 28503 12835
rect 28537 12835 28595 12841
rect 28537 12832 28549 12835
rect 28491 12804 28549 12832
rect 28491 12801 28503 12804
rect 28445 12795 28503 12801
rect 28537 12801 28549 12804
rect 28583 12801 28595 12835
rect 28537 12795 28595 12801
rect 18874 12764 18880 12776
rect 18616 12736 18880 12764
rect 18874 12724 18880 12736
rect 18932 12764 18938 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 18932 12736 18981 12764
rect 18932 12724 18938 12736
rect 18969 12733 18981 12736
rect 19015 12764 19027 12767
rect 22649 12767 22707 12773
rect 19015 12736 19334 12764
rect 19015 12733 19027 12736
rect 18969 12727 19027 12733
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 6748 12668 7328 12696
rect 8036 12668 8677 12696
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 6748 12637 6776 12668
rect 7300 12637 7328 12668
rect 8665 12665 8677 12668
rect 8711 12665 8723 12699
rect 8665 12659 8723 12665
rect 6733 12631 6791 12637
rect 6733 12628 6745 12631
rect 5776 12600 6745 12628
rect 5776 12588 5782 12600
rect 6733 12597 6745 12600
rect 6779 12597 6791 12631
rect 6733 12591 6791 12597
rect 7285 12631 7343 12637
rect 7285 12597 7297 12631
rect 7331 12597 7343 12631
rect 7285 12591 7343 12597
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12628 8631 12631
rect 8938 12628 8944 12640
rect 8619 12600 8944 12628
rect 8619 12597 8631 12600
rect 8573 12591 8631 12597
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 10502 12588 10508 12640
rect 10560 12628 10566 12640
rect 11698 12628 11704 12640
rect 10560 12600 11704 12628
rect 10560 12588 10566 12600
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 15841 12631 15899 12637
rect 15841 12597 15853 12631
rect 15887 12628 15899 12631
rect 16206 12628 16212 12640
rect 15887 12600 16212 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 19306 12628 19334 12736
rect 22649 12733 22661 12767
rect 22695 12733 22707 12767
rect 22649 12727 22707 12733
rect 21637 12699 21695 12705
rect 21637 12665 21649 12699
rect 21683 12696 21695 12699
rect 22664 12696 22692 12727
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 25130 12764 25136 12776
rect 24912 12736 25136 12764
rect 24912 12724 24918 12736
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 26418 12724 26424 12776
rect 26476 12764 26482 12776
rect 27522 12764 27528 12776
rect 26476 12736 27528 12764
rect 26476 12724 26482 12736
rect 27522 12724 27528 12736
rect 27580 12764 27586 12776
rect 28644 12764 28672 12928
rect 28810 12909 28816 12912
rect 28804 12863 28816 12909
rect 28868 12900 28874 12912
rect 35268 12900 35296 12928
rect 36173 12903 36231 12909
rect 36173 12900 36185 12903
rect 28868 12872 28904 12900
rect 30576 12872 34376 12900
rect 35268 12872 36185 12900
rect 28810 12860 28816 12863
rect 28868 12860 28874 12872
rect 30576 12841 30604 12872
rect 30469 12835 30527 12841
rect 30469 12801 30481 12835
rect 30515 12832 30527 12835
rect 30561 12835 30619 12841
rect 30561 12832 30573 12835
rect 30515 12804 30573 12832
rect 30515 12801 30527 12804
rect 30469 12795 30527 12801
rect 30561 12801 30573 12804
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 30828 12835 30886 12841
rect 30828 12801 30840 12835
rect 30874 12832 30886 12835
rect 31846 12832 31852 12844
rect 30874 12804 31852 12832
rect 30874 12801 30886 12804
rect 30828 12795 30886 12801
rect 31846 12792 31852 12804
rect 31904 12792 31910 12844
rect 32140 12841 32168 12872
rect 32125 12835 32183 12841
rect 32125 12801 32137 12835
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 32392 12835 32450 12841
rect 32392 12801 32404 12835
rect 32438 12832 32450 12835
rect 33226 12832 33232 12844
rect 32438 12804 33232 12832
rect 32438 12801 32450 12804
rect 32392 12795 32450 12801
rect 33226 12792 33232 12804
rect 33284 12792 33290 12844
rect 34348 12841 34376 12872
rect 36173 12869 36185 12872
rect 36219 12900 36231 12903
rect 36538 12900 36544 12912
rect 36219 12872 36544 12900
rect 36219 12869 36231 12872
rect 36173 12863 36231 12869
rect 36538 12860 36544 12872
rect 36596 12860 36602 12912
rect 40120 12903 40178 12909
rect 40120 12869 40132 12903
rect 40166 12900 40178 12903
rect 41325 12903 41383 12909
rect 41325 12900 41337 12903
rect 40166 12872 41337 12900
rect 40166 12869 40178 12872
rect 40120 12863 40178 12869
rect 41325 12869 41337 12872
rect 41371 12869 41383 12903
rect 41325 12863 41383 12869
rect 34333 12835 34391 12841
rect 34333 12801 34345 12835
rect 34379 12832 34391 12835
rect 34422 12832 34428 12844
rect 34379 12804 34428 12832
rect 34379 12801 34391 12804
rect 34333 12795 34391 12801
rect 34422 12792 34428 12804
rect 34480 12792 34486 12844
rect 34606 12841 34612 12844
rect 34600 12795 34612 12841
rect 34606 12792 34612 12795
rect 34664 12792 34670 12844
rect 37544 12835 37602 12841
rect 37544 12801 37556 12835
rect 37590 12832 37602 12835
rect 38746 12832 38752 12844
rect 37590 12804 38752 12832
rect 37590 12801 37602 12804
rect 37544 12795 37602 12801
rect 38746 12792 38752 12804
rect 38804 12792 38810 12844
rect 38930 12792 38936 12844
rect 38988 12832 38994 12844
rect 39853 12835 39911 12841
rect 39853 12832 39865 12835
rect 38988 12804 39865 12832
rect 38988 12792 38994 12804
rect 39853 12801 39865 12804
rect 39899 12801 39911 12835
rect 39853 12795 39911 12801
rect 40678 12792 40684 12844
rect 40736 12832 40742 12844
rect 41138 12832 41144 12844
rect 40736 12804 41144 12832
rect 40736 12792 40742 12804
rect 41138 12792 41144 12804
rect 41196 12832 41202 12844
rect 42720 12832 42748 12928
rect 41196 12804 42748 12832
rect 41196 12792 41202 12804
rect 42886 12792 42892 12844
rect 42944 12832 42950 12844
rect 43073 12835 43131 12841
rect 43073 12832 43085 12835
rect 42944 12804 43085 12832
rect 42944 12792 42950 12804
rect 43073 12801 43085 12804
rect 43119 12832 43131 12835
rect 43272 12832 43300 12928
rect 47765 12903 47823 12909
rect 47765 12900 47777 12903
rect 45756 12872 47777 12900
rect 43119 12804 43300 12832
rect 43340 12835 43398 12841
rect 43119 12801 43131 12804
rect 43073 12795 43131 12801
rect 43340 12801 43352 12835
rect 43386 12832 43398 12835
rect 44545 12835 44603 12841
rect 44545 12832 44557 12835
rect 43386 12804 44557 12832
rect 43386 12801 43398 12804
rect 43340 12795 43398 12801
rect 44545 12801 44557 12804
rect 44591 12801 44603 12835
rect 44545 12795 44603 12801
rect 45756 12776 45784 12872
rect 47765 12869 47777 12872
rect 47811 12900 47823 12903
rect 47811 12872 48268 12900
rect 47811 12869 47823 12872
rect 47765 12863 47823 12869
rect 46014 12841 46020 12844
rect 46008 12795 46020 12841
rect 46014 12792 46020 12795
rect 46072 12792 46078 12844
rect 48240 12841 48268 12872
rect 48314 12860 48320 12912
rect 48372 12860 48378 12912
rect 48884 12900 48912 12940
rect 49605 12937 49617 12971
rect 49651 12968 49663 12971
rect 50062 12968 50068 12980
rect 49651 12940 50068 12968
rect 49651 12937 49663 12940
rect 49605 12931 49663 12937
rect 50062 12928 50068 12940
rect 50120 12928 50126 12980
rect 50982 12928 50988 12980
rect 51040 12928 51046 12980
rect 51810 12928 51816 12980
rect 51868 12928 51874 12980
rect 52454 12928 52460 12980
rect 52512 12968 52518 12980
rect 52733 12971 52791 12977
rect 52733 12968 52745 12971
rect 52512 12940 52745 12968
rect 52512 12928 52518 12940
rect 52733 12937 52745 12940
rect 52779 12937 52791 12971
rect 52733 12931 52791 12937
rect 53101 12971 53159 12977
rect 53101 12937 53113 12971
rect 53147 12968 53159 12971
rect 54018 12968 54024 12980
rect 53147 12940 54024 12968
rect 53147 12937 53159 12940
rect 53101 12931 53159 12937
rect 54018 12928 54024 12940
rect 54076 12968 54082 12980
rect 54754 12968 54760 12980
rect 54076 12940 54760 12968
rect 54076 12928 54082 12940
rect 54754 12928 54760 12940
rect 54812 12928 54818 12980
rect 55953 12971 56011 12977
rect 55953 12937 55965 12971
rect 55999 12968 56011 12971
rect 56594 12968 56600 12980
rect 55999 12940 56600 12968
rect 55999 12937 56011 12940
rect 55953 12931 56011 12937
rect 56594 12928 56600 12940
rect 56652 12928 56658 12980
rect 56686 12928 56692 12980
rect 56744 12928 56750 12980
rect 50157 12903 50215 12909
rect 50157 12900 50169 12903
rect 48884 12872 50169 12900
rect 50157 12869 50169 12872
rect 50203 12869 50215 12903
rect 50157 12863 50215 12869
rect 48225 12835 48283 12841
rect 48225 12801 48237 12835
rect 48271 12801 48283 12835
rect 48225 12795 48283 12801
rect 34149 12767 34207 12773
rect 34149 12764 34161 12767
rect 27580 12736 28672 12764
rect 33152 12736 34161 12764
rect 27580 12724 27586 12736
rect 27798 12696 27804 12708
rect 21683 12668 22692 12696
rect 24688 12668 25268 12696
rect 21683 12665 21695 12668
rect 21637 12659 21695 12665
rect 21450 12628 21456 12640
rect 19306 12600 21456 12628
rect 21450 12588 21456 12600
rect 21508 12628 21514 12640
rect 21652 12628 21680 12659
rect 21508 12600 21680 12628
rect 21508 12588 21514 12600
rect 22094 12588 22100 12640
rect 22152 12588 22158 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 24688 12628 24716 12668
rect 23348 12600 24716 12628
rect 23348 12588 23354 12600
rect 25130 12588 25136 12640
rect 25188 12588 25194 12640
rect 25240 12628 25268 12668
rect 26344 12668 27804 12696
rect 26344 12628 26372 12668
rect 27798 12656 27804 12668
rect 27856 12656 27862 12708
rect 25240 12600 26372 12628
rect 26970 12588 26976 12640
rect 27028 12588 27034 12640
rect 31941 12631 31999 12637
rect 31941 12597 31953 12631
rect 31987 12628 31999 12631
rect 33152 12628 33180 12736
rect 34149 12733 34161 12736
rect 34195 12733 34207 12767
rect 34149 12727 34207 12733
rect 35802 12724 35808 12776
rect 35860 12764 35866 12776
rect 36446 12764 36452 12776
rect 35860 12736 36452 12764
rect 35860 12724 35866 12736
rect 36446 12724 36452 12736
rect 36504 12724 36510 12776
rect 36906 12724 36912 12776
rect 36964 12764 36970 12776
rect 37277 12767 37335 12773
rect 37277 12764 37289 12767
rect 36964 12736 37289 12764
rect 36964 12724 36970 12736
rect 37277 12733 37289 12736
rect 37323 12733 37335 12767
rect 37277 12727 37335 12733
rect 39298 12724 39304 12776
rect 39356 12724 39362 12776
rect 41414 12724 41420 12776
rect 41472 12764 41478 12776
rect 41877 12767 41935 12773
rect 41877 12764 41889 12767
rect 41472 12736 41889 12764
rect 41472 12724 41478 12736
rect 41877 12733 41889 12736
rect 41923 12733 41935 12767
rect 41877 12727 41935 12733
rect 45094 12724 45100 12776
rect 45152 12724 45158 12776
rect 45738 12724 45744 12776
rect 45796 12724 45802 12776
rect 47486 12764 47492 12776
rect 47136 12736 47492 12764
rect 47136 12705 47164 12736
rect 47486 12724 47492 12736
rect 47544 12764 47550 12776
rect 48332 12764 48360 12860
rect 48492 12835 48550 12841
rect 48492 12801 48504 12835
rect 48538 12832 48550 12835
rect 48538 12804 49740 12832
rect 48538 12801 48550 12804
rect 48492 12795 48550 12801
rect 47544 12736 48360 12764
rect 49712 12764 49740 12804
rect 49786 12792 49792 12844
rect 49844 12832 49850 12844
rect 50065 12835 50123 12841
rect 50065 12832 50077 12835
rect 49844 12804 50077 12832
rect 49844 12792 49850 12804
rect 50065 12801 50077 12804
rect 50111 12801 50123 12835
rect 51000 12832 51028 12928
rect 51436 12903 51494 12909
rect 51436 12869 51448 12903
rect 51482 12900 51494 12903
rect 51828 12900 51856 12928
rect 51482 12872 51856 12900
rect 53024 12872 53328 12900
rect 51482 12869 51494 12872
rect 51436 12863 51494 12869
rect 53024 12832 53052 12872
rect 50065 12795 50123 12801
rect 50172 12804 51028 12832
rect 51092 12804 53052 12832
rect 50172 12764 50200 12804
rect 49712 12736 50200 12764
rect 47544 12724 47550 12736
rect 50338 12724 50344 12776
rect 50396 12724 50402 12776
rect 51092 12764 51120 12804
rect 53190 12792 53196 12844
rect 53248 12792 53254 12844
rect 51046 12736 51120 12764
rect 47121 12699 47179 12705
rect 47121 12665 47133 12699
rect 47167 12665 47179 12699
rect 51046 12696 51074 12736
rect 51166 12724 51172 12776
rect 51224 12724 51230 12776
rect 53300 12773 53328 12872
rect 53742 12860 53748 12912
rect 53800 12900 53806 12912
rect 53926 12900 53932 12912
rect 53800 12872 53932 12900
rect 53800 12860 53806 12872
rect 53926 12860 53932 12872
rect 53984 12860 53990 12912
rect 54754 12792 54760 12844
rect 54812 12841 54818 12844
rect 54812 12835 54861 12841
rect 54812 12801 54815 12835
rect 54849 12801 54861 12835
rect 54812 12795 54861 12801
rect 55677 12835 55735 12841
rect 55677 12801 55689 12835
rect 55723 12832 55735 12835
rect 56321 12835 56379 12841
rect 56321 12832 56333 12835
rect 55723 12804 56333 12832
rect 55723 12801 55735 12804
rect 55677 12795 55735 12801
rect 56321 12801 56333 12804
rect 56367 12832 56379 12835
rect 56704 12832 56732 12928
rect 57333 12835 57391 12841
rect 57333 12832 57345 12835
rect 56367 12804 56640 12832
rect 56704 12804 57345 12832
rect 56367 12801 56379 12804
rect 56321 12795 56379 12801
rect 54812 12792 54818 12795
rect 53285 12767 53343 12773
rect 53285 12733 53297 12767
rect 53331 12764 53343 12767
rect 53745 12767 53803 12773
rect 53745 12764 53757 12767
rect 53331 12736 53757 12764
rect 53331 12733 53343 12736
rect 53285 12727 53343 12733
rect 53745 12733 53757 12736
rect 53791 12733 53803 12767
rect 53745 12727 53803 12733
rect 54662 12724 54668 12776
rect 54720 12724 54726 12776
rect 54938 12724 54944 12776
rect 54996 12724 55002 12776
rect 55122 12724 55128 12776
rect 55180 12764 55186 12776
rect 55180 12736 55352 12764
rect 55180 12724 55186 12736
rect 47121 12659 47179 12665
rect 49160 12668 51074 12696
rect 31987 12600 33180 12628
rect 31987 12597 31999 12600
rect 31941 12591 31999 12597
rect 33594 12588 33600 12640
rect 33652 12588 33658 12640
rect 35710 12588 35716 12640
rect 35768 12588 35774 12640
rect 42426 12588 42432 12640
rect 42484 12628 42490 12640
rect 42702 12628 42708 12640
rect 42484 12600 42708 12628
rect 42484 12588 42490 12600
rect 42702 12588 42708 12600
rect 42760 12588 42766 12640
rect 44450 12588 44456 12640
rect 44508 12588 44514 12640
rect 46750 12588 46756 12640
rect 46808 12628 46814 12640
rect 49160 12628 49188 12668
rect 53466 12656 53472 12708
rect 53524 12656 53530 12708
rect 55214 12656 55220 12708
rect 55272 12656 55278 12708
rect 55324 12696 55352 12736
rect 55858 12724 55864 12776
rect 55916 12724 55922 12776
rect 56413 12767 56471 12773
rect 56413 12733 56425 12767
rect 56459 12733 56471 12767
rect 56413 12727 56471 12733
rect 56428 12696 56456 12727
rect 56502 12724 56508 12776
rect 56560 12724 56566 12776
rect 56612 12764 56640 12804
rect 57333 12801 57345 12804
rect 57379 12801 57391 12835
rect 57333 12795 57391 12801
rect 56781 12767 56839 12773
rect 56781 12764 56793 12767
rect 56612 12736 56793 12764
rect 56781 12733 56793 12736
rect 56827 12733 56839 12767
rect 56781 12727 56839 12733
rect 57146 12724 57152 12776
rect 57204 12724 57210 12776
rect 57164 12696 57192 12724
rect 55324 12668 57192 12696
rect 46808 12600 49188 12628
rect 46808 12588 46814 12600
rect 49694 12588 49700 12640
rect 49752 12588 49758 12640
rect 50801 12631 50859 12637
rect 50801 12597 50813 12631
rect 50847 12628 50859 12631
rect 51350 12628 51356 12640
rect 50847 12600 51356 12628
rect 50847 12597 50859 12600
rect 50801 12591 50859 12597
rect 51350 12588 51356 12600
rect 51408 12588 51414 12640
rect 52549 12631 52607 12637
rect 52549 12597 52561 12631
rect 52595 12628 52607 12631
rect 53484 12628 53512 12656
rect 52595 12600 53512 12628
rect 54021 12631 54079 12637
rect 52595 12597 52607 12600
rect 52549 12591 52607 12597
rect 54021 12597 54033 12631
rect 54067 12628 54079 12631
rect 56134 12628 56140 12640
rect 54067 12600 56140 12628
rect 54067 12597 54079 12600
rect 54021 12591 54079 12597
rect 56134 12588 56140 12600
rect 56192 12588 56198 12640
rect 1104 12538 58880 12560
rect 1104 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 22616 12538
rect 22668 12486 22680 12538
rect 22732 12486 22744 12538
rect 22796 12486 22808 12538
rect 22860 12486 22872 12538
rect 22924 12486 37060 12538
rect 37112 12486 37124 12538
rect 37176 12486 37188 12538
rect 37240 12486 37252 12538
rect 37304 12486 37316 12538
rect 37368 12486 51504 12538
rect 51556 12486 51568 12538
rect 51620 12486 51632 12538
rect 51684 12486 51696 12538
rect 51748 12486 51760 12538
rect 51812 12486 58880 12538
rect 1104 12464 58880 12486
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 5166 12424 5172 12436
rect 4304 12396 5172 12424
rect 4304 12384 4310 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 8757 12427 8815 12433
rect 8757 12393 8769 12427
rect 8803 12424 8815 12427
rect 9766 12424 9772 12436
rect 8803 12396 9772 12424
rect 8803 12393 8815 12396
rect 8757 12387 8815 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 10413 12427 10471 12433
rect 10413 12393 10425 12427
rect 10459 12424 10471 12427
rect 10594 12424 10600 12436
rect 10459 12396 10600 12424
rect 10459 12393 10471 12396
rect 10413 12387 10471 12393
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 11790 12384 11796 12436
rect 11848 12384 11854 12436
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 14550 12424 14556 12436
rect 12308 12396 14556 12424
rect 12308 12384 12314 12396
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 16945 12427 17003 12433
rect 16945 12393 16957 12427
rect 16991 12424 17003 12427
rect 17494 12424 17500 12436
rect 16991 12396 17500 12424
rect 16991 12393 17003 12396
rect 16945 12387 17003 12393
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 19702 12424 19708 12436
rect 19444 12396 19708 12424
rect 3510 12316 3516 12368
rect 3568 12356 3574 12368
rect 3789 12359 3847 12365
rect 3789 12356 3801 12359
rect 3568 12328 3801 12356
rect 3568 12316 3574 12328
rect 3789 12325 3801 12328
rect 3835 12325 3847 12359
rect 3789 12319 3847 12325
rect 5077 12359 5135 12365
rect 5077 12325 5089 12359
rect 5123 12325 5135 12359
rect 5077 12319 5135 12325
rect 2590 12248 2596 12300
rect 2648 12248 2654 12300
rect 5092 12288 5120 12319
rect 3344 12260 3832 12288
rect 3344 12229 3372 12260
rect 3804 12232 3832 12260
rect 4080 12260 5120 12288
rect 5184 12288 5212 12384
rect 6454 12316 6460 12368
rect 6512 12316 6518 12368
rect 11808 12356 11836 12384
rect 15102 12356 15108 12368
rect 11808 12328 15108 12356
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 5184 12260 5549 12288
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3510 12180 3516 12232
rect 3568 12180 3574 12232
rect 3786 12180 3792 12232
rect 3844 12180 3850 12232
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 4080 12229 4108 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 6472 12288 6500 12316
rect 5537 12251 5595 12257
rect 6288 12260 6500 12288
rect 4064 12223 4122 12229
rect 4064 12220 4076 12223
rect 3936 12192 4076 12220
rect 3936 12180 3942 12192
rect 4064 12189 4076 12192
rect 4110 12189 4122 12223
rect 4064 12183 4122 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4172 12096 4200 12183
rect 5718 12180 5724 12232
rect 5776 12180 5782 12232
rect 6288 12229 6316 12260
rect 7558 12248 7564 12300
rect 7616 12248 7622 12300
rect 10962 12288 10968 12300
rect 10796 12260 10968 12288
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12220 5871 12223
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5859 12192 6285 12220
rect 5859 12189 5871 12192
rect 5813 12183 5871 12189
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 5077 12155 5135 12161
rect 5077 12121 5089 12155
rect 5123 12152 5135 12155
rect 5166 12152 5172 12164
rect 5123 12124 5172 12152
rect 5123 12121 5135 12124
rect 5077 12115 5135 12121
rect 5166 12112 5172 12124
rect 5224 12112 5230 12164
rect 5736 12152 5764 12180
rect 6822 12152 6828 12164
rect 5736 12124 6828 12152
rect 6822 12112 6828 12124
rect 6880 12152 6886 12164
rect 6932 12152 6960 12183
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9033 12223 9091 12229
rect 9033 12220 9045 12223
rect 8996 12192 9045 12220
rect 8996 12180 9002 12192
rect 9033 12189 9045 12192
rect 9079 12220 9091 12223
rect 10796 12220 10824 12260
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11146 12248 11152 12300
rect 11204 12288 11210 12300
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11204 12260 11345 12288
rect 11204 12248 11210 12260
rect 11333 12257 11345 12260
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 11606 12248 11612 12300
rect 11664 12248 11670 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11848 12260 11897 12288
rect 11848 12248 11854 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 11885 12251 11943 12257
rect 12176 12260 12541 12288
rect 12176 12232 12204 12260
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 13188 12297 13216 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 16669 12359 16727 12365
rect 16669 12325 16681 12359
rect 16715 12356 16727 12359
rect 17126 12356 17132 12368
rect 16715 12328 17132 12356
rect 16715 12325 16727 12328
rect 16669 12319 16727 12325
rect 17126 12316 17132 12328
rect 17184 12316 17190 12368
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 12676 12260 13093 12288
rect 12676 12248 12682 12260
rect 13081 12257 13093 12260
rect 13127 12257 13139 12291
rect 13081 12251 13139 12257
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12257 13231 12291
rect 13173 12251 13231 12257
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 15838 12297 15844 12300
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 13964 12260 14565 12288
rect 13964 12248 13970 12260
rect 14553 12257 14565 12260
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 14645 12291 14703 12297
rect 14645 12257 14657 12291
rect 14691 12257 14703 12291
rect 14645 12251 14703 12257
rect 15795 12291 15844 12297
rect 15795 12257 15807 12291
rect 15841 12257 15844 12291
rect 15795 12251 15844 12257
rect 9079 12192 10824 12220
rect 9079 12189 9091 12192
rect 9033 12183 9091 12189
rect 11422 12180 11428 12232
rect 11480 12229 11486 12232
rect 11480 12223 11529 12229
rect 11480 12189 11483 12223
rect 11517 12189 11529 12223
rect 11480 12183 11529 12189
rect 11480 12180 11486 12183
rect 12158 12180 12164 12232
rect 12216 12180 12222 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 12391 12192 14473 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 13924 12164 13952 12192
rect 14461 12189 14473 12192
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 6880 12124 6960 12152
rect 6880 12112 6886 12124
rect 9122 12112 9128 12164
rect 9180 12152 9186 12164
rect 9278 12155 9336 12161
rect 9278 12152 9290 12155
rect 9180 12124 9290 12152
rect 9180 12112 9186 12124
rect 9278 12121 9290 12124
rect 9324 12121 9336 12155
rect 9278 12115 9336 12121
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12121 10747 12155
rect 12989 12155 13047 12161
rect 12989 12152 13001 12155
rect 10689 12115 10747 12121
rect 12406 12124 13001 12152
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 4212 12056 4445 12084
rect 4212 12044 4218 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 5629 12087 5687 12093
rect 5629 12084 5641 12087
rect 4672 12056 5641 12084
rect 4672 12044 4678 12056
rect 5629 12053 5641 12056
rect 5675 12053 5687 12087
rect 10704 12084 10732 12115
rect 12406 12084 12434 12124
rect 12989 12121 13001 12124
rect 13035 12121 13047 12155
rect 12989 12115 13047 12121
rect 13906 12112 13912 12164
rect 13964 12112 13970 12164
rect 14660 12152 14688 12251
rect 15838 12248 15844 12251
rect 15896 12248 15902 12300
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12288 16175 12291
rect 16206 12288 16212 12300
rect 16163 12260 16212 12288
rect 16163 12257 16175 12260
rect 16117 12251 16175 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 16482 12248 16488 12300
rect 16540 12288 16546 12300
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 16540 12260 17509 12288
rect 16540 12248 16546 12260
rect 17497 12257 17509 12260
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 18230 12248 18236 12300
rect 18288 12248 18294 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19444 12297 19472 12396
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 22741 12427 22799 12433
rect 22741 12424 22753 12427
rect 22520 12396 22753 12424
rect 22520 12384 22526 12396
rect 22741 12393 22753 12396
rect 22787 12393 22799 12427
rect 22741 12387 22799 12393
rect 24486 12384 24492 12436
rect 24544 12384 24550 12436
rect 26234 12384 26240 12436
rect 26292 12424 26298 12436
rect 26329 12427 26387 12433
rect 26329 12424 26341 12427
rect 26292 12396 26341 12424
rect 26292 12384 26298 12396
rect 26329 12393 26341 12396
rect 26375 12393 26387 12427
rect 26329 12387 26387 12393
rect 27341 12427 27399 12433
rect 27341 12393 27353 12427
rect 27387 12424 27399 12427
rect 27522 12424 27528 12436
rect 27387 12396 27528 12424
rect 27387 12393 27399 12396
rect 27341 12387 27399 12393
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 29730 12384 29736 12436
rect 29788 12424 29794 12436
rect 44085 12427 44143 12433
rect 29788 12396 44036 12424
rect 29788 12384 29794 12396
rect 28629 12359 28687 12365
rect 28629 12356 28641 12359
rect 28000 12328 28641 12356
rect 19429 12291 19487 12297
rect 19429 12288 19441 12291
rect 19392 12260 19441 12288
rect 19392 12248 19398 12260
rect 19429 12257 19441 12260
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 20898 12248 20904 12300
rect 20956 12248 20962 12300
rect 21266 12288 21272 12300
rect 21008 12260 21272 12288
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 18248 12220 18276 12248
rect 17451 12192 18276 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 14016 12124 14688 12152
rect 19696 12155 19754 12161
rect 14016 12096 14044 12124
rect 19696 12121 19708 12155
rect 19742 12152 19754 12155
rect 19886 12152 19892 12164
rect 19742 12124 19892 12152
rect 19742 12121 19754 12124
rect 19696 12115 19754 12121
rect 19886 12112 19892 12124
rect 19944 12112 19950 12164
rect 21008 12152 21036 12260
rect 21266 12248 21272 12260
rect 21324 12288 21330 12300
rect 21545 12291 21603 12297
rect 21545 12288 21557 12291
rect 21324 12260 21557 12288
rect 21324 12248 21330 12260
rect 21545 12257 21557 12260
rect 21591 12257 21603 12291
rect 21545 12251 21603 12257
rect 21634 12248 21640 12300
rect 21692 12288 21698 12300
rect 21821 12291 21879 12297
rect 21821 12288 21833 12291
rect 21692 12260 21833 12288
rect 21692 12248 21698 12260
rect 21821 12257 21833 12260
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 25130 12248 25136 12300
rect 25188 12248 25194 12300
rect 26970 12248 26976 12300
rect 27028 12248 27034 12300
rect 28000 12297 28028 12328
rect 28629 12325 28641 12328
rect 28675 12325 28687 12359
rect 30374 12356 30380 12368
rect 28629 12319 28687 12325
rect 29288 12328 30380 12356
rect 29288 12297 29316 12328
rect 30374 12316 30380 12328
rect 30432 12316 30438 12368
rect 32674 12316 32680 12368
rect 32732 12356 32738 12368
rect 34330 12356 34336 12368
rect 32732 12328 34336 12356
rect 32732 12316 32738 12328
rect 27985 12291 28043 12297
rect 27985 12257 27997 12291
rect 28031 12257 28043 12291
rect 27985 12251 28043 12257
rect 29273 12291 29331 12297
rect 29273 12257 29285 12291
rect 29319 12257 29331 12291
rect 31435 12291 31493 12297
rect 31435 12288 31447 12291
rect 29273 12251 29331 12257
rect 30300 12260 31447 12288
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21910 12180 21916 12232
rect 21968 12229 21974 12232
rect 21968 12223 21996 12229
rect 21984 12189 21996 12223
rect 21968 12183 21996 12189
rect 21968 12180 21974 12183
rect 22094 12180 22100 12232
rect 22152 12180 22158 12232
rect 27798 12180 27804 12232
rect 27856 12220 27862 12232
rect 29730 12220 29736 12232
rect 27856 12192 29736 12220
rect 27856 12180 27862 12192
rect 29730 12180 29736 12192
rect 29788 12180 29794 12232
rect 30300 12152 30328 12260
rect 31435 12257 31447 12260
rect 31481 12257 31493 12291
rect 31435 12251 31493 12257
rect 31570 12248 31576 12300
rect 31628 12248 31634 12300
rect 31849 12291 31907 12297
rect 31849 12257 31861 12291
rect 31895 12288 31907 12291
rect 31938 12288 31944 12300
rect 31895 12260 31944 12288
rect 31895 12257 31907 12260
rect 31849 12251 31907 12257
rect 31938 12248 31944 12260
rect 31996 12248 32002 12300
rect 32784 12297 32812 12328
rect 34330 12316 34336 12328
rect 34388 12316 34394 12368
rect 34606 12316 34612 12368
rect 34664 12356 34670 12368
rect 34701 12359 34759 12365
rect 34701 12356 34713 12359
rect 34664 12328 34713 12356
rect 34664 12316 34670 12328
rect 34701 12325 34713 12328
rect 34747 12325 34759 12359
rect 34701 12319 34759 12325
rect 35158 12316 35164 12368
rect 35216 12356 35222 12368
rect 36173 12359 36231 12365
rect 36173 12356 36185 12359
rect 35216 12328 36185 12356
rect 35216 12316 35222 12328
rect 36173 12325 36185 12328
rect 36219 12356 36231 12359
rect 36630 12356 36636 12368
rect 36219 12328 36636 12356
rect 36219 12325 36231 12328
rect 36173 12319 36231 12325
rect 36630 12316 36636 12328
rect 36688 12316 36694 12368
rect 37921 12359 37979 12365
rect 37921 12325 37933 12359
rect 37967 12356 37979 12359
rect 39298 12356 39304 12368
rect 37967 12328 39304 12356
rect 37967 12325 37979 12328
rect 37921 12319 37979 12325
rect 39298 12316 39304 12328
rect 39356 12316 39362 12368
rect 41322 12316 41328 12368
rect 41380 12316 41386 12368
rect 41417 12359 41475 12365
rect 41417 12325 41429 12359
rect 41463 12356 41475 12359
rect 41598 12356 41604 12368
rect 41463 12328 41604 12356
rect 41463 12325 41475 12328
rect 41417 12319 41475 12325
rect 41598 12316 41604 12328
rect 41656 12316 41662 12368
rect 42613 12359 42671 12365
rect 42613 12325 42625 12359
rect 42659 12356 42671 12359
rect 42702 12356 42708 12368
rect 42659 12328 42708 12356
rect 42659 12325 42671 12328
rect 42613 12319 42671 12325
rect 42702 12316 42708 12328
rect 42760 12316 42766 12368
rect 44008 12356 44036 12396
rect 44085 12393 44097 12427
rect 44131 12424 44143 12427
rect 45094 12424 45100 12436
rect 44131 12396 45100 12424
rect 44131 12393 44143 12396
rect 44085 12387 44143 12393
rect 45094 12384 45100 12396
rect 45152 12384 45158 12436
rect 47026 12384 47032 12436
rect 47084 12384 47090 12436
rect 47302 12384 47308 12436
rect 47360 12424 47366 12436
rect 48041 12427 48099 12433
rect 48041 12424 48053 12427
rect 47360 12396 48053 12424
rect 47360 12384 47366 12396
rect 48041 12393 48053 12396
rect 48087 12393 48099 12427
rect 48041 12387 48099 12393
rect 49605 12427 49663 12433
rect 49605 12393 49617 12427
rect 49651 12424 49663 12427
rect 50338 12424 50344 12436
rect 49651 12396 50344 12424
rect 49651 12393 49663 12396
rect 49605 12387 49663 12393
rect 44008 12328 47256 12356
rect 32769 12291 32827 12297
rect 32769 12257 32781 12291
rect 32815 12257 32827 12291
rect 32769 12251 32827 12257
rect 32861 12291 32919 12297
rect 32861 12257 32873 12291
rect 32907 12288 32919 12291
rect 33594 12288 33600 12300
rect 32907 12260 33600 12288
rect 32907 12257 32919 12260
rect 32861 12251 32919 12257
rect 30374 12180 30380 12232
rect 30432 12180 30438 12232
rect 31294 12180 31300 12232
rect 31352 12180 31358 12232
rect 32309 12223 32367 12229
rect 32309 12189 32321 12223
rect 32355 12189 32367 12223
rect 32309 12183 32367 12189
rect 32493 12223 32551 12229
rect 32493 12189 32505 12223
rect 32539 12220 32551 12223
rect 32876 12220 32904 12251
rect 33594 12248 33600 12260
rect 33652 12248 33658 12300
rect 34054 12248 34060 12300
rect 34112 12248 34118 12300
rect 34790 12248 34796 12300
rect 34848 12288 34854 12300
rect 35253 12291 35311 12297
rect 35253 12288 35265 12291
rect 34848 12260 35265 12288
rect 34848 12248 34854 12260
rect 35253 12257 35265 12260
rect 35299 12257 35311 12291
rect 35253 12251 35311 12257
rect 35621 12291 35679 12297
rect 35621 12257 35633 12291
rect 35667 12288 35679 12291
rect 35710 12288 35716 12300
rect 35667 12260 35716 12288
rect 35667 12257 35679 12260
rect 35621 12251 35679 12257
rect 35710 12248 35716 12260
rect 35768 12248 35774 12300
rect 35894 12248 35900 12300
rect 35952 12288 35958 12300
rect 36722 12288 36728 12300
rect 35952 12260 36728 12288
rect 35952 12248 35958 12260
rect 36722 12248 36728 12260
rect 36780 12248 36786 12300
rect 36814 12248 36820 12300
rect 36872 12288 36878 12300
rect 37093 12291 37151 12297
rect 37093 12288 37105 12291
rect 36872 12260 37105 12288
rect 36872 12248 36878 12260
rect 37093 12257 37105 12260
rect 37139 12288 37151 12291
rect 37369 12291 37427 12297
rect 37369 12288 37381 12291
rect 37139 12260 37381 12288
rect 37139 12257 37151 12260
rect 37093 12251 37151 12257
rect 37369 12257 37381 12260
rect 37415 12288 37427 12291
rect 38102 12288 38108 12300
rect 37415 12260 38108 12288
rect 37415 12257 37427 12260
rect 37369 12251 37427 12257
rect 38102 12248 38108 12260
rect 38160 12248 38166 12300
rect 38654 12248 38660 12300
rect 38712 12248 38718 12300
rect 41506 12248 41512 12300
rect 41564 12288 41570 12300
rect 42199 12291 42257 12297
rect 42199 12288 42211 12291
rect 41564 12260 42211 12288
rect 41564 12248 41570 12260
rect 42199 12257 42211 12260
rect 42245 12257 42257 12291
rect 42199 12251 42257 12257
rect 42334 12248 42340 12300
rect 42392 12248 42398 12300
rect 43441 12291 43499 12297
rect 43441 12257 43453 12291
rect 43487 12257 43499 12291
rect 43441 12251 43499 12257
rect 32539 12192 32904 12220
rect 32539 12189 32551 12192
rect 32493 12183 32551 12189
rect 32324 12152 32352 12183
rect 32950 12180 32956 12232
rect 33008 12220 33014 12232
rect 33873 12223 33931 12229
rect 33873 12220 33885 12223
rect 33008 12192 33885 12220
rect 33008 12180 33014 12192
rect 33873 12189 33885 12192
rect 33919 12189 33931 12223
rect 33873 12183 33931 12189
rect 37461 12223 37519 12229
rect 37461 12189 37473 12223
rect 37507 12220 37519 12223
rect 37642 12220 37648 12232
rect 37507 12192 37648 12220
rect 37507 12189 37519 12192
rect 37461 12183 37519 12189
rect 37642 12180 37648 12192
rect 37700 12220 37706 12232
rect 38013 12223 38071 12229
rect 38013 12220 38025 12223
rect 37700 12192 38025 12220
rect 37700 12180 37706 12192
rect 38013 12189 38025 12192
rect 38059 12189 38071 12223
rect 39942 12220 39948 12232
rect 38013 12183 38071 12189
rect 38948 12192 39948 12220
rect 33781 12155 33839 12161
rect 33781 12152 33793 12155
rect 20732 12124 21036 12152
rect 29012 12124 30328 12152
rect 30392 12124 30880 12152
rect 32324 12124 33793 12152
rect 10704 12056 12434 12084
rect 12621 12087 12679 12093
rect 5629 12047 5687 12053
rect 12621 12053 12633 12087
rect 12667 12084 12679 12087
rect 12710 12084 12716 12096
rect 12667 12056 12716 12084
rect 12667 12053 12679 12056
rect 12621 12047 12679 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 13998 12084 14004 12096
rect 13872 12056 14004 12084
rect 13872 12044 13878 12056
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 14090 12044 14096 12096
rect 14148 12044 14154 12096
rect 15194 12044 15200 12096
rect 15252 12044 15258 12096
rect 15657 12087 15715 12093
rect 15657 12053 15669 12087
rect 15703 12084 15715 12087
rect 15746 12084 15752 12096
rect 15703 12056 15752 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 15746 12044 15752 12056
rect 15804 12084 15810 12096
rect 17310 12084 17316 12096
rect 15804 12056 17316 12084
rect 15804 12044 15810 12056
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 20732 12084 20760 12124
rect 29012 12096 29040 12124
rect 19852 12056 20760 12084
rect 19852 12044 19858 12056
rect 20806 12044 20812 12096
rect 20864 12044 20870 12096
rect 28534 12044 28540 12096
rect 28592 12044 28598 12096
rect 28994 12044 29000 12096
rect 29052 12044 29058 12096
rect 29089 12087 29147 12093
rect 29089 12053 29101 12087
rect 29135 12084 29147 12087
rect 29270 12084 29276 12096
rect 29135 12056 29276 12084
rect 29135 12053 29147 12056
rect 29089 12047 29147 12053
rect 29270 12044 29276 12056
rect 29328 12084 29334 12096
rect 30392 12084 30420 12124
rect 30852 12096 30880 12124
rect 33781 12121 33793 12124
rect 33827 12152 33839 12155
rect 34146 12152 34152 12164
rect 33827 12124 34152 12152
rect 33827 12121 33839 12124
rect 33781 12115 33839 12121
rect 34146 12112 34152 12124
rect 34204 12112 34210 12164
rect 37553 12155 37611 12161
rect 37553 12152 37565 12155
rect 36556 12124 37565 12152
rect 36556 12096 36584 12124
rect 37553 12121 37565 12124
rect 37599 12121 37611 12155
rect 37553 12115 37611 12121
rect 38948 12096 38976 12192
rect 39942 12180 39948 12192
rect 40000 12180 40006 12232
rect 42058 12180 42064 12232
rect 42116 12180 42122 12232
rect 43073 12223 43131 12229
rect 43073 12189 43085 12223
rect 43119 12189 43131 12223
rect 43073 12183 43131 12189
rect 40212 12155 40270 12161
rect 40212 12121 40224 12155
rect 40258 12152 40270 12155
rect 40954 12152 40960 12164
rect 40258 12124 40960 12152
rect 40258 12121 40270 12124
rect 40212 12115 40270 12121
rect 40954 12112 40960 12124
rect 41012 12112 41018 12164
rect 43088 12152 43116 12183
rect 43162 12180 43168 12232
rect 43220 12220 43226 12232
rect 43257 12223 43315 12229
rect 43257 12220 43269 12223
rect 43220 12192 43269 12220
rect 43220 12180 43226 12192
rect 43257 12189 43269 12192
rect 43303 12189 43315 12223
rect 43456 12220 43484 12251
rect 44450 12248 44456 12300
rect 44508 12288 44514 12300
rect 44729 12291 44787 12297
rect 44729 12288 44741 12291
rect 44508 12260 44741 12288
rect 44508 12248 44514 12260
rect 44729 12257 44741 12260
rect 44775 12257 44787 12291
rect 46385 12291 46443 12297
rect 46385 12288 46397 12291
rect 44729 12251 44787 12257
rect 46124 12260 46397 12288
rect 43530 12220 43536 12232
rect 43456 12192 43536 12220
rect 43257 12183 43315 12189
rect 43530 12180 43536 12192
rect 43588 12180 43594 12232
rect 43717 12155 43775 12161
rect 43717 12152 43729 12155
rect 43088 12124 43729 12152
rect 43717 12121 43729 12124
rect 43763 12152 43775 12155
rect 44177 12155 44235 12161
rect 44177 12152 44189 12155
rect 43763 12124 44189 12152
rect 43763 12121 43775 12124
rect 43717 12115 43775 12121
rect 44177 12121 44189 12124
rect 44223 12121 44235 12155
rect 44177 12115 44235 12121
rect 29328 12056 30420 12084
rect 29328 12044 29334 12056
rect 30650 12044 30656 12096
rect 30708 12044 30714 12096
rect 30834 12044 30840 12096
rect 30892 12084 30898 12096
rect 32950 12084 32956 12096
rect 30892 12056 32956 12084
rect 30892 12044 30898 12056
rect 32950 12044 32956 12056
rect 33008 12044 33014 12096
rect 33318 12044 33324 12096
rect 33376 12044 33382 12096
rect 33410 12044 33416 12096
rect 33468 12044 33474 12096
rect 34517 12087 34575 12093
rect 34517 12053 34529 12087
rect 34563 12084 34575 12087
rect 35894 12084 35900 12096
rect 34563 12056 35900 12084
rect 34563 12053 34575 12056
rect 34517 12047 34575 12053
rect 35894 12044 35900 12056
rect 35952 12044 35958 12096
rect 36446 12044 36452 12096
rect 36504 12044 36510 12096
rect 36538 12044 36544 12096
rect 36596 12044 36602 12096
rect 38930 12044 38936 12096
rect 38988 12044 38994 12096
rect 39114 12044 39120 12096
rect 39172 12084 39178 12096
rect 39669 12087 39727 12093
rect 39669 12084 39681 12087
rect 39172 12056 39681 12084
rect 39172 12044 39178 12056
rect 39669 12053 39681 12056
rect 39715 12084 39727 12087
rect 42426 12084 42432 12096
rect 39715 12056 42432 12084
rect 39715 12053 39727 12056
rect 39669 12047 39727 12053
rect 42426 12044 42432 12056
rect 42484 12044 42490 12096
rect 42518 12044 42524 12096
rect 42576 12084 42582 12096
rect 43625 12087 43683 12093
rect 43625 12084 43637 12087
rect 42576 12056 43637 12084
rect 42576 12044 42582 12056
rect 43625 12053 43637 12056
rect 43671 12053 43683 12087
rect 43625 12047 43683 12053
rect 45554 12044 45560 12096
rect 45612 12084 45618 12096
rect 46124 12093 46152 12260
rect 46385 12257 46397 12260
rect 46431 12288 46443 12291
rect 46750 12288 46756 12300
rect 46431 12260 46756 12288
rect 46431 12257 46443 12260
rect 46385 12251 46443 12257
rect 46750 12248 46756 12260
rect 46808 12248 46814 12300
rect 46569 12155 46627 12161
rect 46569 12121 46581 12155
rect 46615 12152 46627 12155
rect 47121 12155 47179 12161
rect 47121 12152 47133 12155
rect 46615 12124 47133 12152
rect 46615 12121 46627 12124
rect 46569 12115 46627 12121
rect 47121 12121 47133 12124
rect 47167 12121 47179 12155
rect 47228 12152 47256 12328
rect 47670 12248 47676 12300
rect 47728 12248 47734 12300
rect 48056 12220 48084 12387
rect 50338 12384 50344 12396
rect 50396 12384 50402 12436
rect 53926 12384 53932 12436
rect 53984 12424 53990 12436
rect 54938 12424 54944 12436
rect 53984 12396 54944 12424
rect 53984 12384 53990 12396
rect 54938 12384 54944 12396
rect 54996 12384 55002 12436
rect 55490 12384 55496 12436
rect 55548 12384 55554 12436
rect 53193 12359 53251 12365
rect 53193 12325 53205 12359
rect 53239 12356 53251 12359
rect 53239 12328 53328 12356
rect 53239 12325 53251 12328
rect 53193 12319 53251 12325
rect 48498 12248 48504 12300
rect 48556 12288 48562 12300
rect 48593 12291 48651 12297
rect 48593 12288 48605 12291
rect 48556 12260 48605 12288
rect 48556 12248 48562 12260
rect 48593 12257 48605 12260
rect 48639 12288 48651 12291
rect 48958 12288 48964 12300
rect 48639 12260 48964 12288
rect 48639 12257 48651 12260
rect 48593 12251 48651 12257
rect 48958 12248 48964 12260
rect 49016 12248 49022 12300
rect 53300 12297 53328 12328
rect 53285 12291 53343 12297
rect 53285 12257 53297 12291
rect 53331 12257 53343 12291
rect 53285 12251 53343 12257
rect 48225 12223 48283 12229
rect 48225 12220 48237 12223
rect 48056 12192 48237 12220
rect 48225 12189 48237 12192
rect 48271 12189 48283 12223
rect 51074 12220 51080 12232
rect 48225 12183 48283 12189
rect 48332 12192 51080 12220
rect 48332 12152 48360 12192
rect 51074 12180 51080 12192
rect 51132 12180 51138 12232
rect 51813 12223 51871 12229
rect 51813 12220 51825 12223
rect 51644 12192 51825 12220
rect 47228 12124 48360 12152
rect 47121 12115 47179 12121
rect 46109 12087 46167 12093
rect 46109 12084 46121 12087
rect 45612 12056 46121 12084
rect 45612 12044 45618 12056
rect 46109 12053 46121 12056
rect 46155 12053 46167 12087
rect 46109 12047 46167 12053
rect 46661 12087 46719 12093
rect 46661 12053 46673 12087
rect 46707 12084 46719 12087
rect 48406 12084 48412 12096
rect 46707 12056 48412 12084
rect 46707 12053 46719 12056
rect 46661 12047 46719 12053
rect 48406 12044 48412 12056
rect 48464 12044 48470 12096
rect 49878 12044 49884 12096
rect 49936 12084 49942 12096
rect 50890 12084 50896 12096
rect 49936 12056 50896 12084
rect 49936 12044 49942 12056
rect 50890 12044 50896 12056
rect 50948 12084 50954 12096
rect 50985 12087 51043 12093
rect 50985 12084 50997 12087
rect 50948 12056 50997 12084
rect 50948 12044 50954 12056
rect 50985 12053 50997 12056
rect 51031 12084 51043 12087
rect 51258 12084 51264 12096
rect 51031 12056 51264 12084
rect 51031 12053 51043 12056
rect 50985 12047 51043 12053
rect 51258 12044 51264 12056
rect 51316 12084 51322 12096
rect 51644 12093 51672 12192
rect 51813 12189 51825 12192
rect 51859 12189 51871 12223
rect 51813 12183 51871 12189
rect 52080 12223 52138 12229
rect 52080 12189 52092 12223
rect 52126 12220 52138 12223
rect 52362 12220 52368 12232
rect 52126 12192 52368 12220
rect 52126 12189 52138 12192
rect 52080 12183 52138 12189
rect 52362 12180 52368 12192
rect 52420 12180 52426 12232
rect 56042 12180 56048 12232
rect 56100 12180 56106 12232
rect 56686 12180 56692 12232
rect 56744 12180 56750 12232
rect 55214 12152 55220 12164
rect 54404 12124 55220 12152
rect 54404 12096 54432 12124
rect 55214 12112 55220 12124
rect 55272 12112 55278 12164
rect 56597 12155 56655 12161
rect 56597 12121 56609 12155
rect 56643 12152 56655 12155
rect 56934 12155 56992 12161
rect 56934 12152 56946 12155
rect 56643 12124 56946 12152
rect 56643 12121 56655 12124
rect 56597 12115 56655 12121
rect 56934 12121 56946 12124
rect 56980 12121 56992 12155
rect 56934 12115 56992 12121
rect 51629 12087 51687 12093
rect 51629 12084 51641 12087
rect 51316 12056 51641 12084
rect 51316 12044 51322 12056
rect 51629 12053 51641 12056
rect 51675 12053 51687 12087
rect 51629 12047 51687 12053
rect 54297 12087 54355 12093
rect 54297 12053 54309 12087
rect 54343 12084 54355 12087
rect 54386 12084 54392 12096
rect 54343 12056 54392 12084
rect 54343 12053 54355 12056
rect 54297 12047 54355 12053
rect 54386 12044 54392 12056
rect 54444 12044 54450 12096
rect 54662 12044 54668 12096
rect 54720 12084 54726 12096
rect 56226 12084 56232 12096
rect 54720 12056 56232 12084
rect 54720 12044 54726 12056
rect 56226 12044 56232 12056
rect 56284 12044 56290 12096
rect 57514 12044 57520 12096
rect 57572 12084 57578 12096
rect 58069 12087 58127 12093
rect 58069 12084 58081 12087
rect 57572 12056 58081 12084
rect 57572 12044 57578 12056
rect 58069 12053 58081 12056
rect 58115 12053 58127 12087
rect 58069 12047 58127 12053
rect 1104 11994 59040 12016
rect 1104 11942 15394 11994
rect 15446 11942 15458 11994
rect 15510 11942 15522 11994
rect 15574 11942 15586 11994
rect 15638 11942 15650 11994
rect 15702 11942 29838 11994
rect 29890 11942 29902 11994
rect 29954 11942 29966 11994
rect 30018 11942 30030 11994
rect 30082 11942 30094 11994
rect 30146 11942 44282 11994
rect 44334 11942 44346 11994
rect 44398 11942 44410 11994
rect 44462 11942 44474 11994
rect 44526 11942 44538 11994
rect 44590 11942 58726 11994
rect 58778 11942 58790 11994
rect 58842 11942 58854 11994
rect 58906 11942 58918 11994
rect 58970 11942 58982 11994
rect 59034 11942 59040 11994
rect 1104 11920 59040 11942
rect 2958 11840 2964 11892
rect 3016 11840 3022 11892
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 5534 11880 5540 11892
rect 3844 11852 5540 11880
rect 3844 11840 3850 11852
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 5810 11880 5816 11892
rect 5767 11852 5816 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8260 11852 8861 11880
rect 8260 11840 8266 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 9180 11852 9229 11880
rect 9180 11840 9186 11852
rect 9217 11849 9229 11852
rect 9263 11880 9275 11883
rect 11422 11880 11428 11892
rect 9263 11852 11428 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11756 11852 11805 11880
rect 11756 11840 11762 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 12250 11880 12256 11892
rect 11793 11843 11851 11849
rect 11900 11852 12256 11880
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6549 11815 6607 11821
rect 6549 11812 6561 11815
rect 6512 11784 6561 11812
rect 6512 11772 6518 11784
rect 6549 11781 6561 11784
rect 6595 11781 6607 11815
rect 6549 11775 6607 11781
rect 6638 11772 6644 11824
rect 6696 11772 6702 11824
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 7101 11815 7159 11821
rect 7101 11812 7113 11815
rect 6880 11784 7113 11812
rect 6880 11772 6886 11784
rect 7101 11781 7113 11784
rect 7147 11781 7159 11815
rect 7101 11775 7159 11781
rect 9309 11815 9367 11821
rect 9309 11781 9321 11815
rect 9355 11812 9367 11815
rect 10686 11812 10692 11824
rect 9355 11784 10692 11812
rect 9355 11781 9367 11784
rect 9309 11775 9367 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 10778 11772 10784 11824
rect 10836 11812 10842 11824
rect 11900 11812 11928 11852
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 15010 11840 15016 11892
rect 15068 11840 15074 11892
rect 15194 11840 15200 11892
rect 15252 11840 15258 11892
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 21545 11883 21603 11889
rect 21545 11880 21557 11883
rect 20487 11852 21557 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 21545 11849 21557 11852
rect 21591 11880 21603 11883
rect 21910 11880 21916 11892
rect 21591 11852 21916 11880
rect 21591 11849 21603 11852
rect 21545 11843 21603 11849
rect 21910 11840 21916 11852
rect 21968 11840 21974 11892
rect 28534 11840 28540 11892
rect 28592 11840 28598 11892
rect 28994 11840 29000 11892
rect 29052 11840 29058 11892
rect 30650 11840 30656 11892
rect 30708 11880 30714 11892
rect 32493 11883 32551 11889
rect 32493 11880 32505 11883
rect 30708 11852 32505 11880
rect 30708 11840 30714 11852
rect 32493 11849 32505 11852
rect 32539 11849 32551 11883
rect 32493 11843 32551 11849
rect 33318 11840 33324 11892
rect 33376 11840 33382 11892
rect 33410 11840 33416 11892
rect 33468 11840 33474 11892
rect 35897 11883 35955 11889
rect 35897 11849 35909 11883
rect 35943 11880 35955 11883
rect 36906 11880 36912 11892
rect 35943 11852 36912 11880
rect 35943 11849 35955 11852
rect 35897 11843 35955 11849
rect 36906 11840 36912 11852
rect 36964 11840 36970 11892
rect 38102 11840 38108 11892
rect 38160 11880 38166 11892
rect 39114 11880 39120 11892
rect 38160 11852 39120 11880
rect 38160 11840 38166 11852
rect 39114 11840 39120 11852
rect 39172 11840 39178 11892
rect 39942 11840 39948 11892
rect 40000 11880 40006 11892
rect 41969 11883 42027 11889
rect 41969 11880 41981 11883
rect 40000 11852 41981 11880
rect 40000 11840 40006 11852
rect 41969 11849 41981 11852
rect 42015 11880 42027 11883
rect 42242 11880 42248 11892
rect 42015 11852 42248 11880
rect 42015 11849 42027 11852
rect 41969 11843 42027 11849
rect 42242 11840 42248 11852
rect 42300 11880 42306 11892
rect 42886 11880 42892 11892
rect 42300 11852 42892 11880
rect 42300 11840 42306 11852
rect 42886 11840 42892 11852
rect 42944 11840 42950 11892
rect 46014 11840 46020 11892
rect 46072 11880 46078 11892
rect 46201 11883 46259 11889
rect 46201 11880 46213 11883
rect 46072 11852 46213 11880
rect 46072 11840 46078 11852
rect 46201 11849 46213 11852
rect 46247 11849 46259 11883
rect 46201 11843 46259 11849
rect 47026 11840 47032 11892
rect 47084 11840 47090 11892
rect 49513 11883 49571 11889
rect 49513 11849 49525 11883
rect 49559 11880 49571 11883
rect 49786 11880 49792 11892
rect 49559 11852 49792 11880
rect 49559 11849 49571 11852
rect 49513 11843 49571 11849
rect 49786 11840 49792 11852
rect 49844 11840 49850 11892
rect 50154 11840 50160 11892
rect 50212 11840 50218 11892
rect 50890 11840 50896 11892
rect 50948 11840 50954 11892
rect 52917 11883 52975 11889
rect 52917 11849 52929 11883
rect 52963 11880 52975 11883
rect 54570 11880 54576 11892
rect 52963 11852 54576 11880
rect 52963 11849 52975 11852
rect 52917 11843 52975 11849
rect 54570 11840 54576 11852
rect 54628 11840 54634 11892
rect 56042 11840 56048 11892
rect 56100 11840 56106 11892
rect 56597 11883 56655 11889
rect 56597 11849 56609 11883
rect 56643 11880 56655 11883
rect 56686 11880 56692 11892
rect 56643 11852 56692 11880
rect 56643 11849 56655 11852
rect 56597 11843 56655 11849
rect 56686 11840 56692 11852
rect 56744 11840 56750 11892
rect 56781 11883 56839 11889
rect 56781 11849 56793 11883
rect 56827 11849 56839 11883
rect 56781 11843 56839 11849
rect 14458 11812 14464 11824
rect 10836 11784 11928 11812
rect 11992 11784 14464 11812
rect 10836 11772 10842 11784
rect 6643 11769 6701 11772
rect 3236 11747 3294 11753
rect 3236 11713 3248 11747
rect 3282 11713 3294 11747
rect 3236 11707 3294 11713
rect 3252 11676 3280 11707
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3878 11744 3884 11756
rect 3384 11716 3884 11744
rect 3384 11704 3390 11716
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 5626 11704 5632 11756
rect 5684 11704 5690 11756
rect 6643 11735 6655 11769
rect 6689 11735 6701 11769
rect 6643 11729 6701 11735
rect 7006 11704 7012 11756
rect 7064 11704 7070 11756
rect 9944 11747 10002 11753
rect 9944 11713 9956 11747
rect 9990 11744 10002 11747
rect 10502 11744 10508 11756
rect 9990 11716 10508 11744
rect 9990 11713 10002 11716
rect 9944 11707 10002 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 11992 11753 12020 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11020 11716 11989 11744
rect 11020 11704 11026 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12244 11747 12302 11753
rect 12244 11713 12256 11747
rect 12290 11744 12302 11747
rect 13633 11747 13691 11753
rect 13633 11744 13645 11747
rect 12290 11716 13645 11744
rect 12290 11713 12302 11716
rect 12244 11707 12302 11713
rect 13633 11713 13645 11716
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 14148 11716 14197 11744
rect 14148 11704 14154 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 15212 11744 15240 11840
rect 20806 11772 20812 11824
rect 20864 11772 20870 11824
rect 28552 11812 28580 11840
rect 28782 11815 28840 11821
rect 28782 11812 28794 11815
rect 28552 11784 28794 11812
rect 28782 11781 28794 11784
rect 28828 11781 28840 11815
rect 28782 11775 28840 11781
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15212 11716 15577 11744
rect 14185 11707 14243 11713
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 20824 11744 20852 11772
rect 20901 11747 20959 11753
rect 20901 11744 20913 11747
rect 15565 11707 15623 11713
rect 19536 11716 20668 11744
rect 20824 11716 20913 11744
rect 9493 11679 9551 11685
rect 3252 11648 4200 11676
rect 4172 11552 4200 11648
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9582 11676 9588 11688
rect 9539 11648 9588 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9692 11608 9720 11639
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 19536 11685 19564 11716
rect 20640 11685 20668 11716
rect 20901 11713 20913 11716
rect 20947 11713 20959 11747
rect 29012 11744 29040 11840
rect 31754 11772 31760 11824
rect 31812 11812 31818 11824
rect 32585 11815 32643 11821
rect 32585 11812 32597 11815
rect 31812 11784 32597 11812
rect 31812 11772 31818 11784
rect 32585 11781 32597 11784
rect 32631 11781 32643 11815
rect 32585 11775 32643 11781
rect 30653 11747 30711 11753
rect 30653 11744 30665 11747
rect 29012 11716 30665 11744
rect 20901 11707 20959 11713
rect 30653 11713 30665 11716
rect 30699 11713 30711 11747
rect 30653 11707 30711 11713
rect 31846 11704 31852 11756
rect 31904 11744 31910 11756
rect 32953 11747 33011 11753
rect 32953 11744 32965 11747
rect 31904 11716 32965 11744
rect 31904 11704 31910 11716
rect 32953 11713 32965 11716
rect 32999 11713 33011 11747
rect 33336 11744 33364 11840
rect 33428 11812 33456 11840
rect 33428 11784 34284 11812
rect 34256 11753 34284 11784
rect 40954 11772 40960 11824
rect 41012 11772 41018 11824
rect 42058 11772 42064 11824
rect 42116 11812 42122 11824
rect 42613 11815 42671 11821
rect 42613 11812 42625 11815
rect 42116 11784 42625 11812
rect 42116 11772 42122 11784
rect 42613 11781 42625 11784
rect 42659 11781 42671 11815
rect 42613 11775 42671 11781
rect 33505 11747 33563 11753
rect 33505 11744 33517 11747
rect 33336 11716 33517 11744
rect 32953 11707 33011 11713
rect 33505 11713 33517 11716
rect 33551 11713 33563 11747
rect 33505 11707 33563 11713
rect 34241 11747 34299 11753
rect 34241 11713 34253 11747
rect 34287 11713 34299 11747
rect 34241 11707 34299 11713
rect 34330 11704 34336 11756
rect 34388 11744 34394 11756
rect 35069 11747 35127 11753
rect 35069 11744 35081 11747
rect 34388 11716 35081 11744
rect 34388 11704 34394 11716
rect 35069 11713 35081 11716
rect 35115 11744 35127 11747
rect 36170 11744 36176 11756
rect 35115 11716 36176 11744
rect 35115 11713 35127 11716
rect 35069 11707 35127 11713
rect 36170 11704 36176 11716
rect 36228 11704 36234 11756
rect 40497 11747 40555 11753
rect 40497 11713 40509 11747
rect 40543 11744 40555 11747
rect 41506 11744 41512 11756
rect 40543 11716 41512 11744
rect 40543 11713 40555 11716
rect 40497 11707 40555 11713
rect 41506 11704 41512 11716
rect 41564 11704 41570 11756
rect 41601 11747 41659 11753
rect 41601 11713 41613 11747
rect 41647 11744 41659 11747
rect 41690 11744 41696 11756
rect 41647 11716 41696 11744
rect 41647 11713 41659 11716
rect 41601 11707 41659 11713
rect 41690 11704 41696 11716
rect 41748 11704 41754 11756
rect 46845 11747 46903 11753
rect 46845 11713 46857 11747
rect 46891 11744 46903 11747
rect 47044 11744 47072 11840
rect 50172 11812 50200 11840
rect 55769 11815 55827 11821
rect 55769 11812 55781 11815
rect 50172 11784 55781 11812
rect 46891 11716 47072 11744
rect 46891 11713 46903 11716
rect 46845 11707 46903 11713
rect 49234 11704 49240 11756
rect 49292 11744 49298 11756
rect 49421 11747 49479 11753
rect 49421 11744 49433 11747
rect 49292 11716 49433 11744
rect 49292 11704 49298 11716
rect 49421 11713 49433 11716
rect 49467 11713 49479 11747
rect 49421 11707 49479 11713
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 14608 11648 19533 11676
rect 14608 11636 14614 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11676 20683 11679
rect 23290 11676 23296 11688
rect 20671 11648 23296 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 11790 11608 11796 11620
rect 8996 11580 9720 11608
rect 10612 11580 11796 11608
rect 8996 11568 9002 11580
rect 10612 11552 10640 11580
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 15838 11608 15844 11620
rect 14844 11580 15844 11608
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 6362 11540 6368 11552
rect 4212 11512 6368 11540
rect 4212 11500 4218 11512
rect 6362 11500 6368 11512
rect 6420 11540 6426 11552
rect 7374 11540 7380 11552
rect 6420 11512 7380 11540
rect 6420 11500 6426 11512
rect 7374 11500 7380 11512
rect 7432 11540 7438 11552
rect 10594 11540 10600 11552
rect 7432 11512 10600 11540
rect 7432 11500 7438 11512
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11330 11540 11336 11552
rect 11103 11512 11336 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 13354 11500 13360 11552
rect 13412 11500 13418 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 14844 11549 14872 11580
rect 15838 11568 15844 11580
rect 15896 11608 15902 11620
rect 16390 11608 16396 11620
rect 15896 11580 16396 11608
rect 15896 11568 15902 11580
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 20548 11608 20576 11639
rect 23290 11636 23296 11648
rect 23348 11636 23354 11688
rect 23566 11636 23572 11688
rect 23624 11636 23630 11688
rect 25406 11636 25412 11688
rect 25464 11636 25470 11688
rect 28537 11679 28595 11685
rect 28537 11676 28549 11679
rect 28368 11648 28549 11676
rect 20714 11608 20720 11620
rect 20548 11580 20720 11608
rect 20714 11568 20720 11580
rect 20772 11608 20778 11620
rect 22094 11608 22100 11620
rect 20772 11580 22100 11608
rect 20772 11568 20778 11580
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 25225 11611 25283 11617
rect 25225 11577 25237 11611
rect 25271 11608 25283 11611
rect 25498 11608 25504 11620
rect 25271 11580 25504 11608
rect 25271 11577 25283 11580
rect 25225 11571 25283 11577
rect 25498 11568 25504 11580
rect 25556 11608 25562 11620
rect 25556 11580 26188 11608
rect 25556 11568 25562 11580
rect 26160 11552 26188 11580
rect 14829 11543 14887 11549
rect 14829 11540 14841 11543
rect 13596 11512 14841 11540
rect 13596 11500 13602 11512
rect 14829 11509 14841 11512
rect 14875 11509 14887 11543
rect 14829 11503 14887 11509
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16482 11540 16488 11552
rect 16080 11512 16488 11540
rect 16080 11500 16086 11512
rect 16482 11500 16488 11512
rect 16540 11540 16546 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16540 11512 16865 11540
rect 16540 11500 16546 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 16853 11503 16911 11509
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 19852 11512 19901 11540
rect 19852 11500 19858 11512
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 19889 11503 19947 11509
rect 20070 11500 20076 11552
rect 20128 11500 20134 11552
rect 23014 11500 23020 11552
rect 23072 11500 23078 11552
rect 25961 11543 26019 11549
rect 25961 11509 25973 11543
rect 26007 11540 26019 11543
rect 26050 11540 26056 11552
rect 26007 11512 26056 11540
rect 26007 11509 26019 11512
rect 25961 11503 26019 11509
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 26142 11500 26148 11552
rect 26200 11500 26206 11552
rect 28166 11500 28172 11552
rect 28224 11540 28230 11552
rect 28368 11549 28396 11648
rect 28537 11645 28549 11648
rect 28583 11645 28595 11679
rect 28537 11639 28595 11645
rect 30009 11679 30067 11685
rect 30009 11645 30021 11679
rect 30055 11645 30067 11679
rect 30009 11639 30067 11645
rect 29917 11611 29975 11617
rect 29917 11577 29929 11611
rect 29963 11608 29975 11611
rect 30024 11608 30052 11639
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 32677 11679 32735 11685
rect 32677 11676 32689 11679
rect 32640 11648 32689 11676
rect 32640 11636 32646 11648
rect 32677 11645 32689 11648
rect 32723 11676 32735 11679
rect 33134 11676 33140 11688
rect 32723 11648 33140 11676
rect 32723 11645 32735 11648
rect 32677 11639 32735 11645
rect 33134 11636 33140 11648
rect 33192 11636 33198 11688
rect 33226 11636 33232 11688
rect 33284 11676 33290 11688
rect 33689 11679 33747 11685
rect 33689 11676 33701 11679
rect 33284 11648 33701 11676
rect 33284 11636 33290 11648
rect 33689 11645 33701 11648
rect 33735 11645 33747 11679
rect 36262 11676 36268 11688
rect 33689 11639 33747 11645
rect 33980 11648 36268 11676
rect 29963 11580 30052 11608
rect 29963 11577 29975 11580
rect 29917 11571 29975 11577
rect 31846 11568 31852 11620
rect 31904 11608 31910 11620
rect 32858 11608 32864 11620
rect 31904 11580 32864 11608
rect 31904 11568 31910 11580
rect 32858 11568 32864 11580
rect 32916 11568 32922 11620
rect 33152 11608 33180 11636
rect 33980 11608 34008 11648
rect 36262 11636 36268 11648
rect 36320 11636 36326 11688
rect 40221 11679 40279 11685
rect 40221 11676 40233 11679
rect 40052 11648 40233 11676
rect 33152 11580 34008 11608
rect 34054 11568 34060 11620
rect 34112 11608 34118 11620
rect 34701 11611 34759 11617
rect 34701 11608 34713 11611
rect 34112 11580 34713 11608
rect 34112 11568 34118 11580
rect 34701 11577 34713 11580
rect 34747 11608 34759 11611
rect 34747 11580 35756 11608
rect 34747 11577 34759 11580
rect 34701 11571 34759 11577
rect 35728 11552 35756 11580
rect 38930 11568 38936 11620
rect 38988 11568 38994 11620
rect 40052 11552 40080 11648
rect 40221 11645 40233 11648
rect 40267 11645 40279 11679
rect 40221 11639 40279 11645
rect 40405 11679 40463 11685
rect 40405 11645 40417 11679
rect 40451 11676 40463 11679
rect 42518 11676 42524 11688
rect 40451 11648 42524 11676
rect 40451 11645 40463 11648
rect 40405 11639 40463 11645
rect 42518 11636 42524 11648
rect 42576 11636 42582 11688
rect 43257 11679 43315 11685
rect 43257 11645 43269 11679
rect 43303 11676 43315 11679
rect 43530 11676 43536 11688
rect 43303 11648 43536 11676
rect 43303 11645 43315 11648
rect 43257 11639 43315 11645
rect 43530 11636 43536 11648
rect 43588 11676 43594 11688
rect 50172 11676 50200 11784
rect 55769 11781 55781 11784
rect 55815 11781 55827 11815
rect 56060 11812 56088 11840
rect 56796 11812 56824 11843
rect 56060 11784 56824 11812
rect 55769 11775 55827 11781
rect 52825 11747 52883 11753
rect 52825 11713 52837 11747
rect 52871 11744 52883 11747
rect 53098 11744 53104 11756
rect 52871 11716 53104 11744
rect 52871 11713 52883 11716
rect 52825 11707 52883 11713
rect 53098 11704 53104 11716
rect 53156 11704 53162 11756
rect 55784 11744 55812 11775
rect 56502 11744 56508 11756
rect 55784 11716 56508 11744
rect 56502 11704 56508 11716
rect 56560 11704 56566 11756
rect 56962 11704 56968 11756
rect 57020 11744 57026 11756
rect 57146 11744 57152 11756
rect 57020 11716 57152 11744
rect 57020 11704 57026 11716
rect 57146 11704 57152 11716
rect 57204 11704 57210 11756
rect 57241 11747 57299 11753
rect 57241 11713 57253 11747
rect 57287 11744 57299 11747
rect 57885 11747 57943 11753
rect 57885 11744 57897 11747
rect 57287 11716 57897 11744
rect 57287 11713 57299 11716
rect 57241 11707 57299 11713
rect 57885 11713 57897 11716
rect 57931 11713 57943 11747
rect 57885 11707 57943 11713
rect 43588 11648 50200 11676
rect 43588 11636 43594 11648
rect 51442 11636 51448 11688
rect 51500 11676 51506 11688
rect 52362 11676 52368 11688
rect 51500 11648 52368 11676
rect 51500 11636 51506 11648
rect 52362 11636 52368 11648
rect 52420 11676 52426 11688
rect 56229 11679 56287 11685
rect 56229 11676 56241 11679
rect 52420 11648 56241 11676
rect 52420 11636 52426 11648
rect 56229 11645 56241 11648
rect 56275 11676 56287 11679
rect 57422 11676 57428 11688
rect 56275 11648 57428 11676
rect 56275 11645 56287 11648
rect 56229 11639 56287 11645
rect 57422 11636 57428 11648
rect 57480 11636 57486 11688
rect 57514 11636 57520 11688
rect 57572 11676 57578 11688
rect 58437 11679 58495 11685
rect 58437 11676 58449 11679
rect 57572 11648 58449 11676
rect 57572 11636 57578 11648
rect 58437 11645 58449 11648
rect 58483 11645 58495 11679
rect 58437 11639 58495 11645
rect 40865 11611 40923 11617
rect 40865 11577 40877 11611
rect 40911 11608 40923 11611
rect 41414 11608 41420 11620
rect 40911 11580 41420 11608
rect 40911 11577 40923 11580
rect 40865 11571 40923 11577
rect 41414 11568 41420 11580
rect 41472 11568 41478 11620
rect 46842 11568 46848 11620
rect 46900 11608 46906 11620
rect 50525 11611 50583 11617
rect 50525 11608 50537 11611
rect 46900 11580 50537 11608
rect 46900 11568 46906 11580
rect 50525 11577 50537 11580
rect 50571 11608 50583 11611
rect 50571 11580 51074 11608
rect 50571 11577 50583 11580
rect 50525 11571 50583 11577
rect 28353 11543 28411 11549
rect 28353 11540 28365 11543
rect 28224 11512 28365 11540
rect 28224 11500 28230 11512
rect 28353 11509 28365 11512
rect 28399 11509 28411 11543
rect 28353 11503 28411 11509
rect 31294 11500 31300 11552
rect 31352 11540 31358 11552
rect 31941 11543 31999 11549
rect 31941 11540 31953 11543
rect 31352 11512 31953 11540
rect 31352 11500 31358 11512
rect 31941 11509 31953 11512
rect 31987 11540 31999 11543
rect 32030 11540 32036 11552
rect 31987 11512 32036 11540
rect 31987 11509 31999 11512
rect 31941 11503 31999 11509
rect 32030 11500 32036 11512
rect 32088 11500 32094 11552
rect 32125 11543 32183 11549
rect 32125 11509 32137 11543
rect 32171 11540 32183 11543
rect 32490 11540 32496 11552
rect 32171 11512 32496 11540
rect 32171 11509 32183 11512
rect 32125 11503 32183 11509
rect 32490 11500 32496 11512
rect 32548 11500 32554 11552
rect 35342 11500 35348 11552
rect 35400 11500 35406 11552
rect 35710 11500 35716 11552
rect 35768 11500 35774 11552
rect 40034 11500 40040 11552
rect 40092 11500 40098 11552
rect 45646 11500 45652 11552
rect 45704 11500 45710 11552
rect 51046 11540 51074 11580
rect 51350 11540 51356 11552
rect 51046 11512 51356 11540
rect 51350 11500 51356 11512
rect 51408 11500 51414 11552
rect 1104 11450 58880 11472
rect 1104 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 22616 11450
rect 22668 11398 22680 11450
rect 22732 11398 22744 11450
rect 22796 11398 22808 11450
rect 22860 11398 22872 11450
rect 22924 11398 37060 11450
rect 37112 11398 37124 11450
rect 37176 11398 37188 11450
rect 37240 11398 37252 11450
rect 37304 11398 37316 11450
rect 37368 11398 51504 11450
rect 51556 11398 51568 11450
rect 51620 11398 51632 11450
rect 51684 11398 51696 11450
rect 51748 11398 51760 11450
rect 51812 11398 58880 11450
rect 1104 11376 58880 11398
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11336 4031 11339
rect 4614 11336 4620 11348
rect 4019 11308 4620 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 5077 11339 5135 11345
rect 5077 11305 5089 11339
rect 5123 11336 5135 11339
rect 9861 11339 9919 11345
rect 5123 11308 7236 11336
rect 5123 11305 5135 11308
rect 5077 11299 5135 11305
rect 4154 11228 4160 11280
rect 4212 11228 4218 11280
rect 6454 11228 6460 11280
rect 6512 11268 6518 11280
rect 6549 11271 6607 11277
rect 6549 11268 6561 11271
rect 6512 11240 6561 11268
rect 6512 11228 6518 11240
rect 6549 11237 6561 11240
rect 6595 11237 6607 11271
rect 6549 11231 6607 11237
rect 6641 11271 6699 11277
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 6687 11240 6868 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 4172 11132 4200 11228
rect 6840 11212 6868 11240
rect 4706 11200 4712 11212
rect 4356 11172 4712 11200
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 4172 11104 4261 11132
rect 4249 11101 4261 11104
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 3786 11024 3792 11076
rect 3844 11024 3850 11076
rect 4356 11073 4384 11172
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 5776 11172 6745 11200
rect 5776 11160 5782 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 6822 11160 6828 11212
rect 6880 11160 6886 11212
rect 7208 11209 7236 11308
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 11146 11336 11152 11348
rect 9907 11308 11152 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 13354 11296 13360 11348
rect 13412 11296 13418 11348
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 16022 11336 16028 11348
rect 15344 11308 16028 11336
rect 15344 11296 15350 11308
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 19886 11296 19892 11348
rect 19944 11296 19950 11348
rect 20070 11296 20076 11348
rect 20128 11296 20134 11348
rect 22278 11296 22284 11348
rect 22336 11336 22342 11348
rect 23293 11339 23351 11345
rect 23293 11336 23305 11339
rect 22336 11308 23305 11336
rect 22336 11296 22342 11308
rect 23293 11305 23305 11308
rect 23339 11305 23351 11339
rect 23293 11299 23351 11305
rect 25406 11296 25412 11348
rect 25464 11296 25470 11348
rect 29825 11339 29883 11345
rect 29825 11305 29837 11339
rect 29871 11336 29883 11339
rect 30374 11336 30380 11348
rect 29871 11308 30380 11336
rect 29871 11305 29883 11308
rect 29825 11299 29883 11305
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 32582 11296 32588 11348
rect 32640 11296 32646 11348
rect 32766 11296 32772 11348
rect 32824 11296 32830 11348
rect 35728 11308 36952 11336
rect 12066 11268 12072 11280
rect 11716 11240 12072 11268
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10778 11200 10784 11212
rect 10367 11172 10784 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4341 11067 4399 11073
rect 4341 11064 4353 11067
rect 3896 11036 4353 11064
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 3896 10996 3924 11036
rect 4341 11033 4353 11036
rect 4387 11033 4399 11067
rect 4341 11027 4399 11033
rect 4448 11008 4476 11095
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6135 11104 6193 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6181 11101 6193 11104
rect 6227 11132 6239 11135
rect 6638 11132 6644 11144
rect 6227 11104 6644 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 5077 11067 5135 11073
rect 5077 11033 5089 11067
rect 5123 11033 5135 11067
rect 5077 11027 5135 11033
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5810 11064 5816 11076
rect 5307 11036 5816 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 2648 10968 3924 10996
rect 3999 10999 4057 11005
rect 2648 10956 2654 10968
rect 3999 10965 4011 10999
rect 4045 10996 4057 10999
rect 4246 10996 4252 11008
rect 4045 10968 4252 10996
rect 4045 10965 4057 10968
rect 3999 10959 4057 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 4430 10956 4436 11008
rect 4488 10956 4494 11008
rect 5092 10996 5120 11027
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7098 11024 7104 11076
rect 7156 11024 7162 11076
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 9582 11064 9588 11076
rect 9539 11036 9588 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 9582 11024 9588 11036
rect 9640 11064 9646 11076
rect 10336 11064 10364 11163
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11716 11209 11744 11240
rect 12066 11228 12072 11240
rect 12124 11268 12130 11280
rect 12124 11240 12296 11268
rect 12124 11228 12130 11240
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 12158 11160 12164 11212
rect 12216 11160 12222 11212
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11132 11575 11135
rect 12176 11132 12204 11160
rect 11563 11104 12204 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 12268 11076 12296 11240
rect 13372 11209 13400 11296
rect 14182 11228 14188 11280
rect 14240 11268 14246 11280
rect 14366 11268 14372 11280
rect 14240 11240 14372 11268
rect 14240 11228 14246 11240
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11169 13415 11203
rect 20088 11200 20116 11296
rect 35728 11280 35756 11308
rect 21910 11228 21916 11280
rect 21968 11268 21974 11280
rect 27246 11268 27252 11280
rect 21968 11240 27252 11268
rect 21968 11228 21974 11240
rect 27246 11228 27252 11240
rect 27304 11228 27310 11280
rect 35710 11228 35716 11280
rect 35768 11228 35774 11280
rect 36924 11268 36952 11308
rect 40126 11296 40132 11348
rect 40184 11336 40190 11348
rect 40313 11339 40371 11345
rect 40313 11336 40325 11339
rect 40184 11308 40325 11336
rect 40184 11296 40190 11308
rect 40313 11305 40325 11308
rect 40359 11305 40371 11339
rect 40313 11299 40371 11305
rect 42242 11296 42248 11348
rect 42300 11296 42306 11348
rect 42610 11296 42616 11348
rect 42668 11296 42674 11348
rect 43530 11296 43536 11348
rect 43588 11296 43594 11348
rect 57054 11296 57060 11348
rect 57112 11336 57118 11348
rect 57609 11339 57667 11345
rect 57609 11336 57621 11339
rect 57112 11308 57621 11336
rect 57112 11296 57118 11308
rect 57609 11305 57621 11308
rect 57655 11336 57667 11339
rect 57977 11339 58035 11345
rect 57977 11336 57989 11339
rect 57655 11308 57989 11336
rect 57655 11305 57667 11308
rect 57609 11299 57667 11305
rect 57977 11305 57989 11308
rect 58023 11305 58035 11339
rect 57977 11299 58035 11305
rect 43548 11268 43576 11296
rect 36924 11240 43576 11268
rect 45646 11228 45652 11280
rect 45704 11268 45710 11280
rect 47489 11271 47547 11277
rect 47489 11268 47501 11271
rect 45704 11240 47501 11268
rect 45704 11228 45710 11240
rect 47489 11237 47501 11240
rect 47535 11237 47547 11271
rect 47489 11231 47547 11237
rect 50356 11240 51074 11268
rect 20441 11203 20499 11209
rect 20441 11200 20453 11203
rect 20088 11172 20453 11200
rect 13357 11163 13415 11169
rect 20441 11169 20453 11172
rect 20487 11169 20499 11203
rect 22002 11200 22008 11212
rect 20441 11163 20499 11169
rect 20824 11172 22008 11200
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 14366 11092 14372 11144
rect 14424 11092 14430 11144
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15381 11135 15439 11141
rect 15381 11132 15393 11135
rect 15252 11104 15393 11132
rect 15252 11092 15258 11104
rect 15381 11101 15393 11104
rect 15427 11132 15439 11135
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 15427 11104 17417 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 17405 11101 17417 11104
rect 17451 11132 17463 11135
rect 17862 11132 17868 11144
rect 17451 11104 17868 11132
rect 17451 11101 17463 11104
rect 17405 11095 17463 11101
rect 17862 11092 17868 11104
rect 17920 11132 17926 11144
rect 18230 11132 18236 11144
rect 17920 11104 18236 11132
rect 17920 11092 17926 11104
rect 18230 11092 18236 11104
rect 18288 11092 18294 11144
rect 20824 11076 20852 11172
rect 22002 11160 22008 11172
rect 22060 11200 22066 11212
rect 24118 11200 24124 11212
rect 22060 11172 24124 11200
rect 22060 11160 22066 11172
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 26053 11203 26111 11209
rect 26053 11169 26065 11203
rect 26099 11200 26111 11203
rect 26142 11200 26148 11212
rect 26099 11172 26148 11200
rect 26099 11169 26111 11172
rect 26053 11163 26111 11169
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 36078 11160 36084 11212
rect 36136 11200 36142 11212
rect 36173 11203 36231 11209
rect 36173 11200 36185 11203
rect 36136 11172 36185 11200
rect 36136 11160 36142 11172
rect 36173 11169 36185 11172
rect 36219 11200 36231 11203
rect 36814 11200 36820 11212
rect 36219 11172 36820 11200
rect 36219 11169 36231 11172
rect 36173 11163 36231 11169
rect 36814 11160 36820 11172
rect 36872 11160 36878 11212
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 21910 11132 21916 11144
rect 21775 11104 21916 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22554 11092 22560 11144
rect 22612 11092 22618 11144
rect 24210 11092 24216 11144
rect 24268 11132 24274 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 24268 11104 24409 11132
rect 24268 11092 24274 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24854 11092 24860 11144
rect 24912 11132 24918 11144
rect 25590 11132 25596 11144
rect 24912 11104 25596 11132
rect 24912 11092 24918 11104
rect 25590 11092 25596 11104
rect 25648 11132 25654 11144
rect 25777 11135 25835 11141
rect 25777 11132 25789 11135
rect 25648 11104 25789 11132
rect 25648 11092 25654 11104
rect 25777 11101 25789 11104
rect 25823 11101 25835 11135
rect 25777 11095 25835 11101
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11132 25927 11135
rect 26237 11135 26295 11141
rect 26237 11132 26249 11135
rect 25915 11104 26249 11132
rect 25915 11101 25927 11104
rect 25869 11095 25927 11101
rect 26237 11101 26249 11104
rect 26283 11101 26295 11135
rect 26237 11095 26295 11101
rect 26418 11092 26424 11144
rect 26476 11132 26482 11144
rect 26789 11135 26847 11141
rect 26789 11132 26801 11135
rect 26476 11104 26801 11132
rect 26476 11092 26482 11104
rect 26789 11101 26801 11104
rect 26835 11101 26847 11135
rect 26789 11095 26847 11101
rect 29086 11092 29092 11144
rect 29144 11092 29150 11144
rect 33594 11092 33600 11144
rect 33652 11092 33658 11144
rect 34330 11092 34336 11144
rect 34388 11092 34394 11144
rect 35342 11092 35348 11144
rect 35400 11092 35406 11144
rect 36446 11092 36452 11144
rect 36504 11092 36510 11144
rect 36722 11092 36728 11144
rect 36780 11132 36786 11144
rect 37001 11135 37059 11141
rect 37001 11132 37013 11135
rect 36780 11104 37013 11132
rect 36780 11092 36786 11104
rect 37001 11101 37013 11104
rect 37047 11101 37059 11135
rect 37001 11095 37059 11101
rect 37274 11092 37280 11144
rect 37332 11132 37338 11144
rect 37737 11135 37795 11141
rect 37737 11132 37749 11135
rect 37332 11104 37749 11132
rect 37332 11092 37338 11104
rect 37737 11101 37749 11104
rect 37783 11101 37795 11135
rect 37737 11095 37795 11101
rect 38746 11092 38752 11144
rect 38804 11092 38810 11144
rect 39574 11092 39580 11144
rect 39632 11092 39638 11144
rect 40126 11092 40132 11144
rect 40184 11132 40190 11144
rect 40589 11135 40647 11141
rect 40589 11132 40601 11135
rect 40184 11104 40601 11132
rect 40184 11092 40190 11104
rect 40589 11101 40601 11104
rect 40635 11101 40647 11135
rect 40589 11095 40647 11101
rect 41230 11092 41236 11144
rect 41288 11132 41294 11144
rect 41877 11135 41935 11141
rect 41877 11132 41889 11135
rect 41288 11104 41889 11132
rect 41288 11092 41294 11104
rect 41877 11101 41889 11104
rect 41923 11101 41935 11135
rect 41877 11095 41935 11101
rect 43806 11092 43812 11144
rect 43864 11092 43870 11144
rect 44174 11092 44180 11144
rect 44232 11132 44238 11144
rect 44453 11135 44511 11141
rect 44453 11132 44465 11135
rect 44232 11104 44465 11132
rect 44232 11092 44238 11104
rect 44453 11101 44465 11104
rect 44499 11101 44511 11135
rect 44453 11095 44511 11101
rect 44818 11092 44824 11144
rect 44876 11132 44882 11144
rect 45557 11135 45615 11141
rect 45557 11132 45569 11135
rect 44876 11104 45569 11132
rect 44876 11092 44882 11104
rect 45557 11101 45569 11104
rect 45603 11101 45615 11135
rect 45557 11095 45615 11101
rect 45830 11092 45836 11144
rect 45888 11092 45894 11144
rect 47026 11092 47032 11144
rect 47084 11092 47090 11144
rect 9640 11036 10364 11064
rect 9640 11024 9646 11036
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 11425 11067 11483 11073
rect 11425 11064 11437 11067
rect 10928 11036 11437 11064
rect 10928 11024 10934 11036
rect 11425 11033 11437 11036
rect 11471 11064 11483 11067
rect 11606 11064 11612 11076
rect 11471 11036 11612 11064
rect 11471 11033 11483 11036
rect 11425 11027 11483 11033
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 12161 11067 12219 11073
rect 12161 11033 12173 11067
rect 12207 11064 12219 11067
rect 12250 11064 12256 11076
rect 12207 11036 12256 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 13170 11024 13176 11076
rect 13228 11024 13234 11076
rect 13998 11024 14004 11076
rect 14056 11064 14062 11076
rect 16482 11064 16488 11076
rect 14056 11036 16488 11064
rect 14056 11024 14062 11036
rect 16482 11024 16488 11036
rect 16540 11064 16546 11076
rect 18046 11064 18052 11076
rect 16540 11036 18052 11064
rect 16540 11024 16546 11036
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 20806 11024 20812 11076
rect 20864 11024 20870 11076
rect 23106 11024 23112 11076
rect 23164 11064 23170 11076
rect 23201 11067 23259 11073
rect 23201 11064 23213 11067
rect 23164 11036 23213 11064
rect 23164 11024 23170 11036
rect 23201 11033 23213 11036
rect 23247 11033 23259 11067
rect 23201 11027 23259 11033
rect 24029 11067 24087 11073
rect 24029 11033 24041 11067
rect 24075 11064 24087 11067
rect 24075 11036 26188 11064
rect 24075 11033 24087 11036
rect 24029 11027 24087 11033
rect 5166 10996 5172 11008
rect 5092 10968 5172 10996
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5442 10956 5448 11008
rect 5500 10956 5506 11008
rect 7834 10956 7840 11008
rect 7892 10956 7898 11008
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 14921 10999 14979 11005
rect 14921 10965 14933 10999
rect 14967 10996 14979 10999
rect 15010 10996 15016 11008
rect 14967 10968 15016 10996
rect 14967 10965 14979 10968
rect 14921 10959 14979 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 16853 10999 16911 11005
rect 16853 10965 16865 10999
rect 16899 10996 16911 10999
rect 17678 10996 17684 11008
rect 16899 10968 17684 10996
rect 16899 10965 16911 10968
rect 16853 10959 16911 10965
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 22002 10956 22008 11008
rect 22060 10956 22066 11008
rect 25041 10999 25099 11005
rect 25041 10965 25053 10999
rect 25087 10996 25099 10999
rect 25498 10996 25504 11008
rect 25087 10968 25504 10996
rect 25087 10965 25099 10968
rect 25041 10959 25099 10965
rect 25498 10956 25504 10968
rect 25556 10956 25562 11008
rect 26160 10996 26188 11036
rect 28534 11024 28540 11076
rect 28592 11024 28598 11076
rect 32861 11067 32919 11073
rect 32861 11033 32873 11067
rect 32907 11064 32919 11067
rect 33318 11064 33324 11076
rect 32907 11036 33324 11064
rect 32907 11033 32919 11036
rect 32861 11027 32919 11033
rect 33318 11024 33324 11036
rect 33376 11024 33382 11076
rect 36464 11064 36492 11092
rect 36814 11064 36820 11076
rect 33704 11036 33916 11064
rect 26326 10996 26332 11008
rect 26160 10968 26332 10996
rect 26326 10956 26332 10968
rect 26384 10956 26390 11008
rect 32674 10956 32680 11008
rect 32732 10996 32738 11008
rect 33045 10999 33103 11005
rect 33045 10996 33057 10999
rect 32732 10968 33057 10996
rect 32732 10956 32738 10968
rect 33045 10965 33057 10968
rect 33091 10965 33103 10999
rect 33045 10959 33103 10965
rect 33226 10956 33232 11008
rect 33284 10996 33290 11008
rect 33704 10996 33732 11036
rect 33284 10968 33732 10996
rect 33284 10956 33290 10968
rect 33778 10956 33784 11008
rect 33836 10956 33842 11008
rect 33888 10996 33916 11036
rect 34808 11036 35020 11064
rect 36464 11036 36820 11064
rect 34808 10996 34836 11036
rect 33888 10968 34836 10996
rect 34882 10956 34888 11008
rect 34940 10956 34946 11008
rect 34992 10996 35020 11036
rect 36814 11024 36820 11036
rect 36872 11024 36878 11076
rect 40402 11024 40408 11076
rect 40460 11024 40466 11076
rect 42058 11024 42064 11076
rect 42116 11064 42122 11076
rect 42521 11067 42579 11073
rect 42521 11064 42533 11067
rect 42116 11036 42533 11064
rect 42116 11024 42122 11036
rect 42521 11033 42533 11036
rect 42567 11033 42579 11067
rect 46385 11067 46443 11073
rect 46385 11064 46397 11067
rect 42521 11027 42579 11033
rect 46216 11036 46397 11064
rect 46216 11008 46244 11036
rect 46385 11033 46397 11036
rect 46431 11033 46443 11067
rect 46385 11027 46443 11033
rect 35434 10996 35440 11008
rect 34992 10968 35440 10996
rect 35434 10956 35440 10968
rect 35492 10996 35498 11008
rect 35802 10996 35808 11008
rect 35492 10968 35808 10996
rect 35492 10956 35498 10968
rect 35802 10956 35808 10968
rect 35860 10956 35866 11008
rect 36446 10956 36452 11008
rect 36504 10956 36510 11008
rect 36630 10956 36636 11008
rect 36688 10996 36694 11008
rect 37185 10999 37243 11005
rect 37185 10996 37197 10999
rect 36688 10968 37197 10996
rect 36688 10956 36694 10968
rect 37185 10965 37197 10968
rect 37231 10965 37243 10999
rect 37185 10959 37243 10965
rect 38194 10956 38200 11008
rect 38252 10956 38258 11008
rect 38933 10999 38991 11005
rect 38933 10965 38945 10999
rect 38979 10996 38991 10999
rect 39022 10996 39028 11008
rect 38979 10968 39028 10996
rect 38979 10965 38991 10968
rect 38933 10959 38991 10965
rect 39022 10956 39028 10968
rect 39080 10956 39086 11008
rect 41138 10956 41144 11008
rect 41196 10996 41202 11008
rect 41233 10999 41291 11005
rect 41233 10996 41245 10999
rect 41196 10968 41245 10996
rect 41196 10956 41202 10968
rect 41233 10965 41245 10968
rect 41279 10965 41291 10999
rect 41233 10959 41291 10965
rect 41322 10956 41328 11008
rect 41380 10956 41386 11008
rect 43162 10956 43168 11008
rect 43220 10956 43226 11008
rect 43898 10956 43904 11008
rect 43956 10956 43962 11008
rect 44634 10956 44640 11008
rect 44692 10996 44698 11008
rect 45005 10999 45063 11005
rect 45005 10996 45017 10999
rect 44692 10968 45017 10996
rect 44692 10956 44698 10968
rect 45005 10965 45017 10968
rect 45051 10965 45063 10999
rect 45005 10959 45063 10965
rect 46198 10956 46204 11008
rect 46256 10956 46262 11008
rect 46474 10956 46480 11008
rect 46532 10956 46538 11008
rect 47504 10996 47532 11231
rect 50356 11212 50384 11240
rect 50338 11160 50344 11212
rect 50396 11160 50402 11212
rect 50614 11160 50620 11212
rect 50672 11200 50678 11212
rect 50893 11203 50951 11209
rect 50893 11200 50905 11203
rect 50672 11172 50905 11200
rect 50672 11160 50678 11172
rect 50893 11169 50905 11172
rect 50939 11169 50951 11203
rect 51046 11200 51074 11240
rect 52086 11200 52092 11212
rect 51046 11172 52092 11200
rect 50893 11163 50951 11169
rect 52086 11160 52092 11172
rect 52144 11200 52150 11212
rect 56505 11203 56563 11209
rect 56505 11200 56517 11203
rect 52144 11172 56517 11200
rect 52144 11160 52150 11172
rect 56505 11169 56517 11172
rect 56551 11200 56563 11203
rect 56778 11200 56784 11212
rect 56551 11172 56784 11200
rect 56551 11169 56563 11172
rect 56505 11163 56563 11169
rect 56778 11160 56784 11172
rect 56836 11160 56842 11212
rect 50706 11092 50712 11144
rect 50764 11092 50770 11144
rect 52178 11092 52184 11144
rect 52236 11092 52242 11144
rect 56134 11092 56140 11144
rect 56192 11132 56198 11144
rect 56965 11135 57023 11141
rect 56965 11132 56977 11135
rect 56192 11104 56977 11132
rect 56192 11092 56198 11104
rect 56965 11101 56977 11104
rect 57011 11101 57023 11135
rect 56965 11095 57023 11101
rect 49602 11064 49608 11076
rect 48516 11036 49608 11064
rect 48516 11008 48544 11036
rect 49602 11024 49608 11036
rect 49660 11064 49666 11076
rect 49881 11067 49939 11073
rect 49881 11064 49893 11067
rect 49660 11036 49893 11064
rect 49660 11024 49666 11036
rect 49881 11033 49893 11036
rect 49927 11033 49939 11067
rect 49881 11027 49939 11033
rect 51074 11024 51080 11076
rect 51132 11064 51138 11076
rect 51629 11067 51687 11073
rect 51629 11064 51641 11067
rect 51132 11036 51641 11064
rect 51132 11024 51138 11036
rect 51629 11033 51641 11036
rect 51675 11033 51687 11067
rect 51629 11027 51687 11033
rect 54386 11024 54392 11076
rect 54444 11064 54450 11076
rect 55493 11067 55551 11073
rect 55493 11064 55505 11067
rect 54444 11036 55505 11064
rect 54444 11024 54450 11036
rect 55493 11033 55505 11036
rect 55539 11064 55551 11067
rect 56778 11064 56784 11076
rect 55539 11036 56784 11064
rect 55539 11033 55551 11036
rect 55493 11027 55551 11033
rect 56778 11024 56784 11036
rect 56836 11024 56842 11076
rect 48314 10996 48320 11008
rect 47504 10968 48320 10996
rect 48314 10956 48320 10968
rect 48372 10956 48378 11008
rect 48498 10956 48504 11008
rect 48556 10956 48562 11008
rect 50154 10956 50160 11008
rect 50212 10956 50218 11008
rect 51166 10956 51172 11008
rect 51224 10996 51230 11008
rect 51537 10999 51595 11005
rect 51537 10996 51549 10999
rect 51224 10968 51549 10996
rect 51224 10956 51230 10968
rect 51537 10965 51549 10968
rect 51583 10965 51595 10999
rect 51537 10959 51595 10965
rect 55953 10999 56011 11005
rect 55953 10965 55965 10999
rect 55999 10996 56011 10999
rect 56226 10996 56232 11008
rect 55999 10968 56232 10996
rect 55999 10965 56011 10968
rect 55953 10959 56011 10965
rect 56226 10956 56232 10968
rect 56284 10956 56290 11008
rect 56870 10956 56876 11008
rect 56928 10956 56934 11008
rect 57330 10956 57336 11008
rect 57388 10956 57394 11008
rect 1104 10906 59040 10928
rect 1104 10854 15394 10906
rect 15446 10854 15458 10906
rect 15510 10854 15522 10906
rect 15574 10854 15586 10906
rect 15638 10854 15650 10906
rect 15702 10854 29838 10906
rect 29890 10854 29902 10906
rect 29954 10854 29966 10906
rect 30018 10854 30030 10906
rect 30082 10854 30094 10906
rect 30146 10854 44282 10906
rect 44334 10854 44346 10906
rect 44398 10854 44410 10906
rect 44462 10854 44474 10906
rect 44526 10854 44538 10906
rect 44590 10854 58726 10906
rect 58778 10854 58790 10906
rect 58842 10854 58854 10906
rect 58906 10854 58918 10906
rect 58970 10854 58982 10906
rect 59034 10854 59040 10906
rect 1104 10832 59040 10854
rect 5350 10752 5356 10804
rect 5408 10752 5414 10804
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 6638 10792 6644 10804
rect 6503 10764 6644 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 2593 10727 2651 10733
rect 2593 10693 2605 10727
rect 2639 10724 2651 10727
rect 5166 10724 5172 10736
rect 2639 10696 5172 10724
rect 2639 10693 2651 10696
rect 2593 10687 2651 10693
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3528 10628 3801 10656
rect 3528 10600 3556 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3510 10548 3516 10600
rect 3568 10548 3574 10600
rect 3694 10548 3700 10600
rect 3752 10548 3758 10600
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 2682 10520 2688 10532
rect 1636 10492 2688 10520
rect 1636 10480 1642 10492
rect 2682 10480 2688 10492
rect 2740 10520 2746 10532
rect 2961 10523 3019 10529
rect 2961 10520 2973 10523
rect 2740 10492 2973 10520
rect 2740 10480 2746 10492
rect 2961 10489 2973 10492
rect 3007 10489 3019 10523
rect 3804 10520 3832 10619
rect 4890 10616 4896 10668
rect 4948 10656 4954 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 4948 10628 5457 10656
rect 4948 10616 4954 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10588 5871 10591
rect 5994 10588 6000 10600
rect 5859 10560 6000 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 5994 10548 6000 10560
rect 6052 10588 6058 10600
rect 6472 10588 6500 10755
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7834 10752 7840 10804
rect 7892 10752 7898 10804
rect 9861 10795 9919 10801
rect 9861 10761 9873 10795
rect 9907 10792 9919 10795
rect 10134 10792 10140 10804
rect 9907 10764 10140 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10502 10752 10508 10804
rect 10560 10752 10566 10804
rect 12618 10752 12624 10804
rect 12676 10792 12682 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 12676 10764 13645 10792
rect 12676 10752 12682 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 14093 10795 14151 10801
rect 14093 10761 14105 10795
rect 14139 10792 14151 10795
rect 15010 10792 15016 10804
rect 14139 10764 15016 10792
rect 14139 10761 14151 10764
rect 14093 10755 14151 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 17034 10792 17040 10804
rect 16899 10764 17040 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 18230 10752 18236 10804
rect 18288 10792 18294 10804
rect 18509 10795 18567 10801
rect 18509 10792 18521 10795
rect 18288 10764 18521 10792
rect 18288 10752 18294 10764
rect 18509 10761 18521 10764
rect 18555 10761 18567 10795
rect 39209 10795 39267 10801
rect 18509 10755 18567 10761
rect 18616 10764 38332 10792
rect 7592 10727 7650 10733
rect 7592 10693 7604 10727
rect 7638 10724 7650 10727
rect 7852 10724 7880 10752
rect 7638 10696 7880 10724
rect 7638 10693 7650 10696
rect 7592 10687 7650 10693
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 18616 10724 18644 10764
rect 9088 10696 18644 10724
rect 19981 10727 20039 10733
rect 9088 10684 9094 10696
rect 19981 10693 19993 10727
rect 20027 10724 20039 10727
rect 20530 10724 20536 10736
rect 20027 10696 20536 10724
rect 20027 10693 20039 10696
rect 19981 10687 20039 10693
rect 20530 10684 20536 10696
rect 20588 10724 20594 10736
rect 30742 10724 30748 10736
rect 20588 10696 30748 10724
rect 20588 10684 20594 10696
rect 30742 10684 30748 10696
rect 30800 10684 30806 10736
rect 33045 10727 33103 10733
rect 33045 10693 33057 10727
rect 33091 10724 33103 10727
rect 33778 10724 33784 10736
rect 33091 10696 33784 10724
rect 33091 10693 33103 10696
rect 33045 10687 33103 10693
rect 33778 10684 33784 10696
rect 33836 10684 33842 10736
rect 34238 10684 34244 10736
rect 34296 10724 34302 10736
rect 34333 10727 34391 10733
rect 34333 10724 34345 10727
rect 34296 10696 34345 10724
rect 34296 10684 34302 10696
rect 34333 10693 34345 10696
rect 34379 10724 34391 10727
rect 35060 10727 35118 10733
rect 34379 10696 35011 10724
rect 34379 10693 34391 10696
rect 34333 10687 34391 10693
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 8938 10656 8944 10668
rect 7883 10628 8944 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 11054 10616 11060 10668
rect 11112 10616 11118 10668
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 13173 10659 13231 10665
rect 13173 10656 13185 10659
rect 12759 10628 13185 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 13173 10625 13185 10628
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13311 10628 14013 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 14001 10625 14013 10628
rect 14047 10656 14059 10659
rect 14550 10656 14556 10668
rect 14047 10628 14556 10656
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 6052 10560 6500 10588
rect 10413 10591 10471 10597
rect 6052 10548 6058 10560
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10594 10588 10600 10600
rect 10459 10560 10600 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13188 10588 13216 10619
rect 14550 10616 14556 10628
rect 14608 10656 14614 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 14608 10628 15853 10656
rect 14608 10616 14614 10628
rect 15841 10625 15853 10628
rect 15887 10656 15899 10659
rect 15887 10628 16528 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 13449 10591 13507 10597
rect 12676 10560 12848 10588
rect 13188 10560 13308 10588
rect 12676 10548 12682 10560
rect 5718 10520 5724 10532
rect 3804 10492 5724 10520
rect 2961 10483 3019 10489
rect 5718 10480 5724 10492
rect 5776 10480 5782 10532
rect 11532 10520 11560 10548
rect 12820 10529 12848 10560
rect 8680 10492 11560 10520
rect 12805 10523 12863 10529
rect 2406 10412 2412 10464
rect 2464 10412 2470 10464
rect 2590 10412 2596 10464
rect 2648 10412 2654 10464
rect 3050 10412 3056 10464
rect 3108 10412 3114 10464
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4982 10452 4988 10464
rect 4488 10424 4988 10452
rect 4488 10412 4494 10424
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 5583 10455 5641 10461
rect 5583 10452 5595 10455
rect 5316 10424 5595 10452
rect 5316 10412 5322 10424
rect 5583 10421 5595 10424
rect 5629 10452 5641 10455
rect 5902 10452 5908 10464
rect 5629 10424 5908 10452
rect 5629 10421 5641 10424
rect 5583 10415 5641 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10452 6147 10455
rect 8680 10452 8708 10492
rect 12805 10489 12817 10523
rect 12851 10489 12863 10523
rect 13280 10520 13308 10560
rect 13449 10557 13461 10591
rect 13495 10588 13507 10591
rect 13538 10588 13544 10600
rect 13495 10560 13544 10588
rect 13495 10557 13507 10560
rect 13449 10551 13507 10557
rect 13538 10548 13544 10560
rect 13596 10548 13602 10600
rect 14182 10548 14188 10600
rect 14240 10548 14246 10600
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10588 15439 10591
rect 15427 10560 15516 10588
rect 15427 10557 15439 10560
rect 15381 10551 15439 10557
rect 15488 10529 15516 10560
rect 15930 10548 15936 10600
rect 15988 10548 15994 10600
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16500 10588 16528 10628
rect 16758 10616 16764 10668
rect 16816 10616 16822 10668
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 21683 10628 22201 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 23474 10616 23480 10668
rect 23532 10656 23538 10668
rect 23569 10659 23627 10665
rect 23569 10656 23581 10659
rect 23532 10628 23581 10656
rect 23532 10616 23538 10628
rect 23569 10625 23581 10628
rect 23615 10625 23627 10659
rect 23569 10619 23627 10625
rect 23661 10659 23719 10665
rect 23661 10625 23673 10659
rect 23707 10656 23719 10659
rect 24670 10656 24676 10668
rect 23707 10628 24676 10656
rect 23707 10625 23719 10628
rect 23661 10619 23719 10625
rect 24670 10616 24676 10628
rect 24728 10616 24734 10668
rect 25682 10656 25688 10668
rect 25332 10628 25688 10656
rect 16850 10588 16856 10600
rect 16500 10560 16856 10588
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20036 10560 20729 10588
rect 20036 10548 20042 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 21910 10548 21916 10600
rect 21968 10548 21974 10600
rect 22094 10548 22100 10600
rect 22152 10548 22158 10600
rect 23753 10591 23811 10597
rect 23753 10588 23765 10591
rect 23308 10560 23765 10588
rect 15473 10523 15531 10529
rect 13280 10492 15424 10520
rect 12805 10483 12863 10489
rect 15396 10464 15424 10492
rect 15473 10489 15485 10523
rect 15519 10489 15531 10523
rect 16040 10520 16068 10548
rect 23308 10532 23336 10560
rect 23753 10557 23765 10560
rect 23799 10557 23811 10591
rect 23753 10551 23811 10557
rect 24026 10548 24032 10600
rect 24084 10548 24090 10600
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 25332 10588 25360 10628
rect 25682 10616 25688 10628
rect 25740 10616 25746 10668
rect 26050 10616 26056 10668
rect 26108 10665 26114 10668
rect 26108 10656 26120 10665
rect 29089 10659 29147 10665
rect 26108 10628 26153 10656
rect 26108 10619 26120 10628
rect 29089 10625 29101 10659
rect 29135 10656 29147 10659
rect 30193 10659 30251 10665
rect 30193 10656 30205 10659
rect 29135 10628 30205 10656
rect 29135 10625 29147 10628
rect 29089 10619 29147 10625
rect 30193 10625 30205 10628
rect 30239 10656 30251 10659
rect 30558 10656 30564 10668
rect 30239 10628 30564 10656
rect 30239 10625 30251 10628
rect 30193 10619 30251 10625
rect 26108 10616 26114 10619
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 30837 10659 30895 10665
rect 30837 10625 30849 10659
rect 30883 10656 30895 10659
rect 31202 10656 31208 10668
rect 30883 10628 31208 10656
rect 30883 10625 30895 10628
rect 30837 10619 30895 10625
rect 31202 10616 31208 10628
rect 31260 10616 31266 10668
rect 33505 10659 33563 10665
rect 33505 10656 33517 10659
rect 31864 10628 33517 10656
rect 24176 10560 25360 10588
rect 24176 10548 24182 10560
rect 26326 10548 26332 10600
rect 26384 10588 26390 10600
rect 26384 10560 26740 10588
rect 26384 10548 26390 10560
rect 19610 10520 19616 10532
rect 16040 10492 19616 10520
rect 15473 10483 15531 10489
rect 19610 10480 19616 10492
rect 19668 10480 19674 10532
rect 21818 10480 21824 10532
rect 21876 10520 21882 10532
rect 23109 10523 23167 10529
rect 23109 10520 23121 10523
rect 21876 10492 23121 10520
rect 21876 10480 21882 10492
rect 23109 10489 23121 10492
rect 23155 10520 23167 10523
rect 23290 10520 23296 10532
rect 23155 10492 23296 10520
rect 23155 10489 23167 10492
rect 23109 10483 23167 10489
rect 23290 10480 23296 10492
rect 23348 10480 23354 10532
rect 23566 10480 23572 10532
rect 23624 10480 23630 10532
rect 26418 10480 26424 10532
rect 26476 10480 26482 10532
rect 6135 10424 8708 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 10560 10424 11897 10452
rect 10560 10412 10566 10424
rect 11885 10421 11897 10424
rect 11931 10452 11943 10455
rect 14182 10452 14188 10464
rect 11931 10424 14188 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14737 10455 14795 10461
rect 14737 10421 14749 10455
rect 14783 10452 14795 10455
rect 15286 10452 15292 10464
rect 14783 10424 15292 10452
rect 14783 10421 14795 10424
rect 14737 10415 14795 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 15838 10412 15844 10464
rect 15896 10452 15902 10464
rect 16022 10452 16028 10464
rect 15896 10424 16028 10452
rect 15896 10412 15902 10424
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 19484 10424 20085 10452
rect 19484 10412 19490 10424
rect 20073 10421 20085 10424
rect 20119 10421 20131 10455
rect 20073 10415 20131 10421
rect 22554 10412 22560 10464
rect 22612 10412 22618 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 23584 10452 23612 10480
rect 23247 10424 23612 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 24578 10412 24584 10464
rect 24636 10452 24642 10464
rect 24949 10455 25007 10461
rect 24949 10452 24961 10455
rect 24636 10424 24961 10452
rect 24636 10412 24642 10424
rect 24949 10421 24961 10424
rect 24995 10452 25007 10455
rect 26436 10452 26464 10480
rect 26712 10464 26740 10560
rect 28994 10548 29000 10600
rect 29052 10588 29058 10600
rect 29181 10591 29239 10597
rect 29181 10588 29193 10591
rect 29052 10560 29193 10588
rect 29052 10548 29058 10560
rect 29181 10557 29193 10560
rect 29227 10557 29239 10591
rect 29181 10551 29239 10557
rect 29270 10548 29276 10600
rect 29328 10548 29334 10600
rect 29454 10548 29460 10600
rect 29512 10588 29518 10600
rect 29549 10591 29607 10597
rect 29549 10588 29561 10591
rect 29512 10560 29561 10588
rect 29512 10548 29518 10560
rect 29549 10557 29561 10560
rect 29595 10557 29607 10591
rect 29549 10551 29607 10557
rect 28629 10523 28687 10529
rect 28629 10489 28641 10523
rect 28675 10520 28687 10523
rect 29288 10520 29316 10548
rect 28675 10492 29316 10520
rect 28675 10489 28687 10492
rect 28629 10483 28687 10489
rect 31864 10464 31892 10628
rect 33505 10625 33517 10628
rect 33551 10625 33563 10659
rect 33505 10619 33563 10625
rect 34793 10659 34851 10665
rect 34793 10625 34805 10659
rect 34839 10656 34851 10659
rect 34882 10656 34888 10668
rect 34839 10628 34888 10656
rect 34839 10625 34851 10628
rect 34793 10619 34851 10625
rect 34882 10616 34888 10628
rect 34940 10616 34946 10668
rect 34983 10656 35011 10696
rect 35060 10693 35072 10727
rect 35106 10724 35118 10727
rect 36446 10724 36452 10736
rect 35106 10696 36452 10724
rect 35106 10693 35118 10696
rect 35060 10687 35118 10693
rect 36446 10684 36452 10696
rect 36504 10684 36510 10736
rect 36538 10684 36544 10736
rect 36596 10684 36602 10736
rect 36906 10684 36912 10736
rect 36964 10724 36970 10736
rect 37728 10727 37786 10733
rect 36964 10696 37504 10724
rect 36964 10684 36970 10696
rect 34983 10628 35839 10656
rect 32585 10591 32643 10597
rect 32585 10557 32597 10591
rect 32631 10588 32643 10591
rect 32769 10591 32827 10597
rect 32769 10588 32781 10591
rect 32631 10560 32781 10588
rect 32631 10557 32643 10560
rect 32585 10551 32643 10557
rect 32769 10557 32781 10560
rect 32815 10557 32827 10591
rect 32769 10551 32827 10557
rect 32953 10591 33011 10597
rect 32953 10557 32965 10591
rect 32999 10588 33011 10591
rect 33962 10588 33968 10600
rect 32999 10560 33968 10588
rect 32999 10557 33011 10560
rect 32953 10551 33011 10557
rect 32784 10520 32812 10551
rect 33962 10548 33968 10560
rect 34020 10548 34026 10600
rect 35811 10588 35839 10628
rect 36354 10616 36360 10668
rect 36412 10616 36418 10668
rect 37476 10656 37504 10696
rect 37728 10693 37740 10727
rect 37774 10724 37786 10727
rect 38194 10724 38200 10736
rect 37774 10696 38200 10724
rect 37774 10693 37786 10696
rect 37728 10687 37786 10693
rect 38194 10684 38200 10696
rect 38252 10684 38258 10736
rect 38304 10724 38332 10764
rect 39209 10761 39221 10795
rect 39255 10792 39267 10795
rect 40494 10792 40500 10804
rect 39255 10764 40500 10792
rect 39255 10761 39267 10764
rect 39209 10755 39267 10761
rect 40494 10752 40500 10764
rect 40552 10792 40558 10804
rect 41233 10795 41291 10801
rect 41233 10792 41245 10795
rect 40552 10764 41245 10792
rect 40552 10752 40558 10764
rect 41233 10761 41245 10764
rect 41279 10761 41291 10795
rect 41233 10755 41291 10761
rect 42242 10752 42248 10804
rect 42300 10752 42306 10804
rect 43806 10752 43812 10804
rect 43864 10752 43870 10804
rect 45465 10795 45523 10801
rect 45465 10761 45477 10795
rect 45511 10792 45523 10795
rect 45830 10792 45836 10804
rect 45511 10764 45836 10792
rect 45511 10761 45523 10764
rect 45465 10755 45523 10761
rect 45830 10752 45836 10764
rect 45888 10752 45894 10804
rect 49602 10752 49608 10804
rect 49660 10792 49666 10804
rect 49660 10764 50292 10792
rect 49660 10752 49666 10764
rect 45646 10724 45652 10736
rect 38304 10696 41552 10724
rect 38930 10656 38936 10668
rect 37476 10628 38936 10656
rect 36814 10588 36820 10600
rect 35811 10560 36820 10588
rect 36814 10548 36820 10560
rect 36872 10548 36878 10600
rect 37476 10597 37504 10628
rect 38930 10616 38936 10628
rect 38988 10656 38994 10668
rect 38988 10628 39252 10656
rect 38988 10616 38994 10628
rect 37461 10591 37519 10597
rect 37461 10557 37473 10591
rect 37507 10557 37519 10591
rect 37461 10551 37519 10557
rect 39114 10548 39120 10600
rect 39172 10548 39178 10600
rect 39224 10588 39252 10628
rect 39298 10616 39304 10668
rect 39356 10616 39362 10668
rect 39761 10659 39819 10665
rect 39761 10656 39773 10659
rect 39408 10628 39773 10656
rect 39408 10588 39436 10628
rect 39761 10625 39773 10628
rect 39807 10625 39819 10659
rect 39761 10619 39819 10625
rect 40028 10659 40086 10665
rect 40028 10625 40040 10659
rect 40074 10656 40086 10659
rect 41322 10656 41328 10668
rect 40074 10628 41328 10656
rect 40074 10625 40086 10628
rect 40028 10619 40086 10625
rect 41322 10616 41328 10628
rect 41380 10616 41386 10668
rect 39224 10560 39436 10588
rect 33226 10520 33232 10532
rect 32784 10492 33232 10520
rect 33226 10480 33232 10492
rect 33284 10480 33290 10532
rect 33413 10523 33471 10529
rect 33413 10489 33425 10523
rect 33459 10520 33471 10523
rect 33594 10520 33600 10532
rect 33459 10492 33600 10520
rect 33459 10489 33471 10492
rect 33413 10483 33471 10489
rect 33594 10480 33600 10492
rect 33652 10480 33658 10532
rect 36173 10523 36231 10529
rect 36173 10489 36185 10523
rect 36219 10520 36231 10523
rect 37274 10520 37280 10532
rect 36219 10492 37280 10520
rect 36219 10489 36231 10492
rect 36173 10483 36231 10489
rect 37274 10480 37280 10492
rect 37332 10480 37338 10532
rect 41141 10523 41199 10529
rect 41141 10489 41153 10523
rect 41187 10520 41199 10523
rect 41524 10520 41552 10696
rect 42444 10696 45652 10724
rect 42444 10665 42472 10696
rect 42429 10659 42487 10665
rect 42429 10656 42441 10659
rect 41616 10628 42441 10656
rect 41616 10600 41644 10628
rect 42429 10625 42441 10628
rect 42475 10625 42487 10659
rect 42429 10619 42487 10625
rect 42696 10659 42754 10665
rect 42696 10625 42708 10659
rect 42742 10656 42754 10659
rect 43898 10656 43904 10668
rect 42742 10628 43904 10656
rect 42742 10625 42754 10628
rect 42696 10619 42754 10625
rect 43898 10616 43904 10628
rect 43956 10616 43962 10668
rect 44100 10665 44128 10696
rect 45646 10684 45652 10696
rect 45704 10724 45710 10736
rect 45741 10727 45799 10733
rect 45741 10724 45753 10727
rect 45704 10696 45753 10724
rect 45704 10684 45710 10696
rect 45741 10693 45753 10696
rect 45787 10693 45799 10727
rect 45741 10687 45799 10693
rect 46284 10727 46342 10733
rect 46284 10693 46296 10727
rect 46330 10724 46342 10727
rect 46474 10724 46480 10736
rect 46330 10696 46480 10724
rect 46330 10693 46342 10696
rect 46284 10687 46342 10693
rect 44085 10659 44143 10665
rect 44085 10625 44097 10659
rect 44131 10625 44143 10659
rect 44085 10619 44143 10625
rect 44352 10659 44410 10665
rect 44352 10625 44364 10659
rect 44398 10656 44410 10659
rect 44634 10656 44640 10668
rect 44398 10628 44640 10656
rect 44398 10625 44410 10628
rect 44352 10619 44410 10625
rect 44634 10616 44640 10628
rect 44692 10616 44698 10668
rect 45756 10656 45784 10687
rect 46474 10684 46480 10696
rect 46532 10684 46538 10736
rect 46658 10684 46664 10736
rect 46716 10724 46722 10736
rect 48222 10724 48228 10736
rect 46716 10696 48228 10724
rect 46716 10684 46722 10696
rect 48222 10684 48228 10696
rect 48280 10724 48286 10736
rect 49050 10724 49056 10736
rect 48280 10696 49056 10724
rect 48280 10684 48286 10696
rect 49050 10684 49056 10696
rect 49108 10684 49114 10736
rect 49878 10724 49884 10736
rect 49252 10696 49884 10724
rect 46017 10659 46075 10665
rect 46017 10656 46029 10659
rect 45756 10628 46029 10656
rect 46017 10625 46029 10628
rect 46063 10625 46075 10659
rect 46017 10619 46075 10625
rect 46106 10616 46112 10668
rect 46164 10656 46170 10668
rect 46676 10656 46704 10684
rect 46164 10628 46704 10656
rect 46164 10616 46170 10628
rect 41598 10548 41604 10600
rect 41656 10548 41662 10600
rect 41782 10548 41788 10600
rect 41840 10548 41846 10600
rect 47581 10591 47639 10597
rect 47581 10557 47593 10591
rect 47627 10557 47639 10591
rect 47581 10551 47639 10557
rect 47397 10523 47455 10529
rect 41187 10492 41414 10520
rect 41524 10492 42012 10520
rect 41187 10489 41199 10492
rect 41141 10483 41199 10489
rect 24995 10424 26464 10452
rect 24995 10421 25007 10424
rect 24949 10415 25007 10421
rect 26694 10412 26700 10464
rect 26752 10412 26758 10464
rect 28721 10455 28779 10461
rect 28721 10421 28733 10455
rect 28767 10452 28779 10455
rect 29086 10452 29092 10464
rect 28767 10424 29092 10452
rect 28767 10421 28779 10424
rect 28721 10415 28779 10421
rect 29086 10412 29092 10424
rect 29144 10412 29150 10464
rect 30745 10455 30803 10461
rect 30745 10421 30757 10455
rect 30791 10452 30803 10455
rect 30834 10452 30840 10464
rect 30791 10424 30840 10452
rect 30791 10421 30803 10424
rect 30745 10415 30803 10421
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 31846 10412 31852 10464
rect 31904 10412 31910 10464
rect 33042 10412 33048 10464
rect 33100 10452 33106 10464
rect 37642 10452 37648 10464
rect 33100 10424 37648 10452
rect 33100 10412 33106 10424
rect 37642 10412 37648 10424
rect 37700 10412 37706 10464
rect 38841 10455 38899 10461
rect 38841 10421 38853 10455
rect 38887 10452 38899 10455
rect 39574 10452 39580 10464
rect 38887 10424 39580 10452
rect 38887 10421 38899 10424
rect 38841 10415 38899 10421
rect 39574 10412 39580 10424
rect 39632 10412 39638 10464
rect 39669 10455 39727 10461
rect 39669 10421 39681 10455
rect 39715 10452 39727 10455
rect 40126 10452 40132 10464
rect 39715 10424 40132 10452
rect 39715 10421 39727 10424
rect 39669 10415 39727 10421
rect 40126 10412 40132 10424
rect 40184 10412 40190 10464
rect 41386 10452 41414 10492
rect 41874 10452 41880 10464
rect 41386 10424 41880 10452
rect 41874 10412 41880 10424
rect 41932 10412 41938 10464
rect 41984 10452 42012 10492
rect 47397 10489 47409 10523
rect 47443 10520 47455 10523
rect 47596 10520 47624 10551
rect 48314 10548 48320 10600
rect 48372 10588 48378 10600
rect 49252 10597 49280 10696
rect 49878 10684 49884 10696
rect 49936 10684 49942 10736
rect 50154 10684 50160 10736
rect 50212 10684 50218 10736
rect 49504 10659 49562 10665
rect 49504 10625 49516 10659
rect 49550 10656 49562 10659
rect 50172 10656 50200 10684
rect 49550 10628 50200 10656
rect 50264 10656 50292 10764
rect 50614 10752 50620 10804
rect 50672 10752 50678 10804
rect 50706 10752 50712 10804
rect 50764 10752 50770 10804
rect 51166 10752 51172 10804
rect 51224 10752 51230 10804
rect 51537 10795 51595 10801
rect 51276 10764 51488 10792
rect 51077 10727 51135 10733
rect 51077 10693 51089 10727
rect 51123 10724 51135 10727
rect 51276 10724 51304 10764
rect 51123 10696 51304 10724
rect 51123 10693 51135 10696
rect 51077 10687 51135 10693
rect 51460 10656 51488 10764
rect 51537 10761 51549 10795
rect 51583 10792 51595 10795
rect 52178 10792 52184 10804
rect 51583 10764 52184 10792
rect 51583 10761 51595 10764
rect 51537 10755 51595 10761
rect 52178 10752 52184 10764
rect 52236 10752 52242 10804
rect 54202 10752 54208 10804
rect 54260 10752 54266 10804
rect 55677 10795 55735 10801
rect 55677 10761 55689 10795
rect 55723 10792 55735 10795
rect 56870 10792 56876 10804
rect 55723 10764 56876 10792
rect 55723 10761 55735 10764
rect 55677 10755 55735 10761
rect 56870 10752 56876 10764
rect 56928 10752 56934 10804
rect 51810 10684 51816 10736
rect 51868 10724 51874 10736
rect 54220 10724 54248 10752
rect 51868 10696 54248 10724
rect 51868 10684 51874 10696
rect 51902 10656 51908 10668
rect 50264 10628 51304 10656
rect 51460 10628 51908 10656
rect 49550 10625 49562 10628
rect 49504 10619 49562 10625
rect 49237 10591 49295 10597
rect 49237 10588 49249 10591
rect 48372 10560 49249 10588
rect 48372 10548 48378 10560
rect 49237 10557 49249 10560
rect 49283 10557 49295 10591
rect 49237 10551 49295 10557
rect 51276 10520 51304 10628
rect 51902 10616 51908 10628
rect 51960 10616 51966 10668
rect 51997 10659 52055 10665
rect 51997 10625 52009 10659
rect 52043 10656 52055 10659
rect 52638 10656 52644 10668
rect 52043 10628 52644 10656
rect 52043 10625 52055 10628
rect 51997 10619 52055 10625
rect 52638 10616 52644 10628
rect 52696 10656 52702 10668
rect 52733 10659 52791 10665
rect 52733 10656 52745 10659
rect 52696 10628 52745 10656
rect 52696 10616 52702 10628
rect 52733 10625 52745 10628
rect 52779 10625 52791 10659
rect 52733 10619 52791 10625
rect 57514 10616 57520 10668
rect 57572 10616 57578 10668
rect 51350 10548 51356 10600
rect 51408 10588 51414 10600
rect 52181 10591 52239 10597
rect 51408 10560 52132 10588
rect 51408 10548 51414 10560
rect 52104 10520 52132 10560
rect 52181 10557 52193 10591
rect 52227 10588 52239 10591
rect 52362 10588 52368 10600
rect 52227 10560 52368 10588
rect 52227 10557 52239 10560
rect 52181 10551 52239 10557
rect 52362 10548 52368 10560
rect 52420 10548 52426 10600
rect 52546 10548 52552 10600
rect 52604 10588 52610 10600
rect 53285 10591 53343 10597
rect 53285 10588 53297 10591
rect 52604 10560 53297 10588
rect 52604 10548 52610 10560
rect 53285 10557 53297 10560
rect 53331 10557 53343 10591
rect 53285 10551 53343 10557
rect 54110 10548 54116 10600
rect 54168 10548 54174 10600
rect 54754 10548 54760 10600
rect 54812 10548 54818 10600
rect 55490 10548 55496 10600
rect 55548 10548 55554 10600
rect 56318 10548 56324 10600
rect 56376 10548 56382 10600
rect 56410 10548 56416 10600
rect 56468 10597 56474 10600
rect 56468 10591 56517 10597
rect 56468 10557 56471 10591
rect 56505 10557 56517 10591
rect 56468 10551 56517 10557
rect 56468 10548 56474 10551
rect 56594 10548 56600 10600
rect 56652 10548 56658 10600
rect 56778 10548 56784 10600
rect 56836 10588 56842 10600
rect 56873 10591 56931 10597
rect 56873 10588 56885 10591
rect 56836 10560 56885 10588
rect 56836 10548 56842 10560
rect 56873 10557 56885 10560
rect 56919 10557 56931 10591
rect 56873 10551 56931 10557
rect 57330 10548 57336 10600
rect 57388 10548 57394 10600
rect 58434 10548 58440 10600
rect 58492 10548 58498 10600
rect 54662 10520 54668 10532
rect 47443 10492 47624 10520
rect 47688 10492 48636 10520
rect 47443 10489 47455 10492
rect 47397 10483 47455 10489
rect 47688 10452 47716 10492
rect 41984 10424 47716 10452
rect 48222 10412 48228 10464
rect 48280 10412 48286 10464
rect 48498 10412 48504 10464
rect 48556 10412 48562 10464
rect 48608 10452 48636 10492
rect 50172 10492 51120 10520
rect 51276 10492 51948 10520
rect 52104 10492 54668 10520
rect 50172 10452 50200 10492
rect 48608 10424 50200 10452
rect 51092 10452 51120 10492
rect 51810 10452 51816 10464
rect 51092 10424 51816 10452
rect 51810 10412 51816 10424
rect 51868 10412 51874 10464
rect 51920 10452 51948 10492
rect 54662 10480 54668 10492
rect 54720 10480 54726 10532
rect 51994 10452 52000 10464
rect 51920 10424 52000 10452
rect 51994 10412 52000 10424
rect 52052 10412 52058 10464
rect 53466 10412 53472 10464
rect 53524 10412 53530 10464
rect 54202 10412 54208 10464
rect 54260 10412 54266 10464
rect 54938 10412 54944 10464
rect 54996 10412 55002 10464
rect 57882 10412 57888 10464
rect 57940 10412 57946 10464
rect 1104 10362 58880 10384
rect 1104 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 22616 10362
rect 22668 10310 22680 10362
rect 22732 10310 22744 10362
rect 22796 10310 22808 10362
rect 22860 10310 22872 10362
rect 22924 10310 37060 10362
rect 37112 10310 37124 10362
rect 37176 10310 37188 10362
rect 37240 10310 37252 10362
rect 37304 10310 37316 10362
rect 37368 10310 51504 10362
rect 51556 10310 51568 10362
rect 51620 10310 51632 10362
rect 51684 10310 51696 10362
rect 51748 10310 51760 10362
rect 51812 10310 58880 10362
rect 1104 10288 58880 10310
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 2740 10220 3464 10248
rect 2740 10208 2746 10220
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2130 10112 2136 10124
rect 1995 10084 2136 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10112 2283 10115
rect 2406 10112 2412 10124
rect 2271 10084 2412 10112
rect 2271 10081 2283 10084
rect 2225 10075 2283 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 3436 10112 3464 10220
rect 3510 10208 3516 10260
rect 3568 10208 3574 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 3752 10220 4721 10248
rect 3752 10208 3758 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 4948 10220 5580 10248
rect 4948 10208 4954 10220
rect 4522 10140 4528 10192
rect 4580 10180 4586 10192
rect 4908 10180 4936 10208
rect 4580 10152 4936 10180
rect 4580 10140 4586 10152
rect 5442 10140 5448 10192
rect 5500 10140 5506 10192
rect 5552 10180 5580 10220
rect 5810 10208 5816 10260
rect 5868 10208 5874 10260
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 6822 10248 6828 10260
rect 5960 10220 6828 10248
rect 5960 10208 5966 10220
rect 6454 10180 6460 10192
rect 5552 10152 6460 10180
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 5258 10112 5264 10124
rect 3436 10084 5264 10112
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 4246 10044 4252 10056
rect 4111 10016 4252 10044
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5460 10044 5488 10140
rect 6564 10124 6592 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 9030 10208 9036 10260
rect 9088 10208 9094 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 9766 10248 9772 10260
rect 9272 10220 9772 10248
rect 9272 10208 9278 10220
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12066 10248 12072 10260
rect 12023 10220 12072 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 12216 10220 12541 10248
rect 12216 10208 12222 10220
rect 12529 10217 12541 10220
rect 12575 10217 12587 10251
rect 13538 10248 13544 10260
rect 12529 10211 12587 10217
rect 13004 10220 13544 10248
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10180 6699 10183
rect 8662 10180 8668 10192
rect 6687 10152 8668 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 8662 10140 8668 10152
rect 8720 10180 8726 10192
rect 9048 10180 9076 10208
rect 8720 10152 9076 10180
rect 8720 10140 8726 10152
rect 9490 10140 9496 10192
rect 9548 10180 9554 10192
rect 12345 10183 12403 10189
rect 12345 10180 12357 10183
rect 9548 10152 12357 10180
rect 9548 10140 9554 10152
rect 12345 10149 12357 10152
rect 12391 10180 12403 10183
rect 13004 10180 13032 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 15010 10208 15016 10260
rect 15068 10248 15074 10260
rect 15068 10220 15700 10248
rect 15068 10208 15074 10220
rect 12391 10152 13032 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 5718 10072 5724 10124
rect 5776 10072 5782 10124
rect 5994 10072 6000 10124
rect 6052 10072 6058 10124
rect 6546 10072 6552 10124
rect 6604 10072 6610 10124
rect 11330 10072 11336 10124
rect 11388 10072 11394 10124
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 14458 10112 14464 10124
rect 13955 10084 14464 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 15473 10115 15531 10121
rect 14568 10084 15240 10112
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 4764 10016 5028 10044
rect 5460 10016 5641 10044
rect 4764 10004 4770 10016
rect 4617 9979 4675 9985
rect 4617 9945 4629 9979
rect 4663 9976 4675 9979
rect 4893 9979 4951 9985
rect 4893 9976 4905 9979
rect 4663 9948 4905 9976
rect 4663 9945 4675 9948
rect 4617 9939 4675 9945
rect 4893 9945 4905 9948
rect 4939 9945 4951 9979
rect 5000 9976 5028 10016
rect 5629 10013 5641 10016
rect 5675 10013 5687 10047
rect 5736 10044 5764 10072
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5736 10016 6101 10044
rect 5629 10007 5687 10013
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 10870 10004 10876 10056
rect 10928 10004 10934 10056
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 14148 10016 14381 10044
rect 14148 10004 14154 10016
rect 14369 10013 14381 10016
rect 14415 10044 14427 10047
rect 14568 10044 14596 10084
rect 15212 10053 15240 10084
rect 15473 10081 15485 10115
rect 15519 10112 15531 10115
rect 15672 10112 15700 10220
rect 15930 10208 15936 10260
rect 15988 10248 15994 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 15988 10220 16497 10248
rect 15988 10208 15994 10220
rect 15519 10084 15700 10112
rect 15749 10115 15807 10121
rect 15519 10081 15531 10084
rect 15473 10075 15531 10081
rect 15749 10081 15761 10115
rect 15795 10112 15807 10115
rect 15838 10112 15844 10124
rect 15795 10084 15844 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16408 10121 16436 10220
rect 16485 10217 16497 10220
rect 16531 10217 16543 10251
rect 16485 10211 16543 10217
rect 20530 10208 20536 10260
rect 20588 10208 20594 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 21082 10248 21088 10260
rect 20947 10220 21088 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 21082 10208 21088 10220
rect 21140 10208 21146 10260
rect 23845 10251 23903 10257
rect 23845 10217 23857 10251
rect 23891 10248 23903 10251
rect 24026 10248 24032 10260
rect 23891 10220 24032 10248
rect 23891 10217 23903 10220
rect 23845 10211 23903 10217
rect 24026 10208 24032 10220
rect 24084 10208 24090 10260
rect 24118 10208 24124 10260
rect 24176 10208 24182 10260
rect 24578 10248 24584 10260
rect 24504 10220 24584 10248
rect 19061 10183 19119 10189
rect 19061 10149 19073 10183
rect 19107 10149 19119 10183
rect 19061 10143 19119 10149
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10081 16451 10115
rect 19076 10112 19104 10143
rect 19978 10112 19984 10124
rect 19076 10084 19984 10112
rect 16393 10075 16451 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 24504 10121 24532 10220
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 24670 10208 24676 10260
rect 24728 10248 24734 10260
rect 32033 10251 32091 10257
rect 24728 10220 25268 10248
rect 24728 10208 24734 10220
rect 24489 10115 24547 10121
rect 24489 10081 24501 10115
rect 24535 10081 24547 10115
rect 24489 10075 24547 10081
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 25240 10112 25268 10220
rect 32033 10217 32045 10251
rect 32079 10248 32091 10251
rect 34882 10248 34888 10260
rect 32079 10220 34888 10248
rect 32079 10217 32091 10220
rect 32033 10211 32091 10217
rect 25409 10115 25467 10121
rect 25409 10112 25421 10115
rect 25240 10084 25421 10112
rect 25409 10081 25421 10084
rect 25455 10081 25467 10115
rect 25409 10075 25467 10081
rect 25682 10072 25688 10124
rect 25740 10072 25746 10124
rect 26510 10072 26516 10124
rect 26568 10112 26574 10124
rect 26973 10115 27031 10121
rect 26973 10112 26985 10115
rect 26568 10084 26985 10112
rect 26568 10072 26574 10084
rect 26973 10081 26985 10084
rect 27019 10112 27031 10115
rect 27430 10112 27436 10124
rect 27019 10084 27436 10112
rect 27019 10081 27031 10084
rect 26973 10075 27031 10081
rect 27430 10072 27436 10084
rect 27488 10072 27494 10124
rect 31110 10072 31116 10124
rect 31168 10112 31174 10124
rect 32140 10121 32168 10220
rect 34882 10208 34888 10220
rect 34940 10208 34946 10260
rect 35618 10208 35624 10260
rect 35676 10248 35682 10260
rect 35676 10220 36124 10248
rect 35676 10208 35682 10220
rect 33505 10183 33563 10189
rect 33505 10149 33517 10183
rect 33551 10180 33563 10183
rect 34330 10180 34336 10192
rect 33551 10152 34336 10180
rect 33551 10149 33563 10152
rect 33505 10143 33563 10149
rect 34330 10140 34336 10152
rect 34388 10140 34394 10192
rect 36096 10180 36124 10220
rect 36170 10208 36176 10260
rect 36228 10248 36234 10260
rect 36446 10248 36452 10260
rect 36228 10220 36452 10248
rect 36228 10208 36234 10220
rect 36446 10208 36452 10220
rect 36504 10208 36510 10260
rect 38565 10251 38623 10257
rect 38565 10217 38577 10251
rect 38611 10248 38623 10251
rect 38746 10248 38752 10260
rect 38611 10220 38752 10248
rect 38611 10217 38623 10220
rect 38565 10211 38623 10217
rect 38746 10208 38752 10220
rect 38804 10208 38810 10260
rect 39853 10251 39911 10257
rect 39853 10217 39865 10251
rect 39899 10248 39911 10251
rect 41782 10248 41788 10260
rect 39899 10220 41788 10248
rect 39899 10217 39911 10220
rect 39853 10211 39911 10217
rect 41782 10208 41788 10220
rect 41840 10208 41846 10260
rect 42797 10251 42855 10257
rect 42797 10217 42809 10251
rect 42843 10248 42855 10251
rect 44174 10248 44180 10260
rect 42843 10220 44180 10248
rect 42843 10217 42855 10220
rect 42797 10211 42855 10217
rect 44174 10208 44180 10220
rect 44232 10208 44238 10260
rect 46382 10248 46388 10260
rect 45940 10220 46388 10248
rect 44821 10183 44879 10189
rect 36096 10152 37136 10180
rect 32125 10115 32183 10121
rect 32125 10112 32137 10115
rect 31168 10084 32137 10112
rect 31168 10072 31174 10084
rect 32125 10081 32137 10084
rect 32171 10081 32183 10115
rect 32125 10075 32183 10081
rect 34238 10072 34244 10124
rect 34296 10072 34302 10124
rect 34348 10112 34376 10140
rect 35483 10115 35541 10121
rect 35483 10112 35495 10115
rect 34348 10084 35495 10112
rect 35483 10081 35495 10084
rect 35529 10081 35541 10115
rect 35483 10075 35541 10081
rect 35894 10072 35900 10124
rect 35952 10112 35958 10124
rect 36357 10115 36415 10121
rect 35952 10084 36216 10112
rect 35952 10072 35958 10084
rect 15378 10053 15384 10056
rect 14415 10016 14596 10044
rect 15197 10047 15255 10053
rect 14415 10013 14427 10016
rect 14369 10007 14427 10013
rect 15197 10013 15209 10047
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15356 10047 15384 10053
rect 15356 10013 15368 10047
rect 15356 10007 15384 10013
rect 15378 10004 15384 10007
rect 15436 10004 15442 10056
rect 16206 10004 16212 10056
rect 16264 10004 16270 10056
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 16632 10016 17049 10044
rect 16632 10004 16638 10016
rect 17037 10013 17049 10016
rect 17083 10013 17095 10047
rect 17037 10007 17095 10013
rect 17678 10004 17684 10056
rect 17736 10004 17742 10056
rect 20070 10004 20076 10056
rect 20128 10004 20134 10056
rect 22002 10044 22008 10056
rect 22060 10053 22066 10056
rect 21972 10016 22008 10044
rect 22002 10004 22008 10016
rect 22060 10007 22072 10053
rect 22060 10004 22066 10007
rect 22278 10004 22284 10056
rect 22336 10044 22342 10056
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22336 10016 22477 10044
rect 22336 10004 22342 10016
rect 22465 10013 22477 10016
rect 22511 10044 22523 10047
rect 23198 10044 23204 10056
rect 22511 10016 23204 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10044 24731 10047
rect 24854 10044 24860 10056
rect 24719 10016 24860 10044
rect 24719 10013 24731 10016
rect 24673 10007 24731 10013
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 25498 10004 25504 10056
rect 25556 10053 25562 10056
rect 25556 10047 25584 10053
rect 25572 10013 25584 10047
rect 25556 10007 25584 10013
rect 25556 10004 25562 10007
rect 26602 10004 26608 10056
rect 26660 10044 26666 10056
rect 26789 10047 26847 10053
rect 26789 10044 26801 10047
rect 26660 10016 26801 10044
rect 26660 10004 26666 10016
rect 26789 10013 26801 10016
rect 26835 10013 26847 10047
rect 26789 10007 26847 10013
rect 27985 10047 28043 10053
rect 27985 10013 27997 10047
rect 28031 10013 28043 10047
rect 27985 10007 28043 10013
rect 32392 10047 32450 10053
rect 32392 10013 32404 10047
rect 32438 10044 32450 10047
rect 32674 10044 32680 10056
rect 32438 10016 32680 10044
rect 32438 10013 32450 10016
rect 32392 10007 32450 10013
rect 5258 9976 5264 9988
rect 5000 9948 5264 9976
rect 4893 9939 4951 9945
rect 5258 9936 5264 9948
rect 5316 9976 5322 9988
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 5316 9948 5457 9976
rect 5316 9936 5322 9948
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 5445 9939 5503 9945
rect 12986 9936 12992 9988
rect 13044 9976 13050 9988
rect 13642 9979 13700 9985
rect 13642 9976 13654 9979
rect 13044 9948 13654 9976
rect 13044 9936 13050 9948
rect 13642 9945 13654 9948
rect 13688 9945 13700 9979
rect 13642 9939 13700 9945
rect 17948 9979 18006 9985
rect 17948 9945 17960 9979
rect 17994 9976 18006 9979
rect 18046 9976 18052 9988
rect 17994 9948 18052 9976
rect 17994 9945 18006 9948
rect 17948 9939 18006 9945
rect 18046 9936 18052 9948
rect 18104 9936 18110 9988
rect 22732 9979 22790 9985
rect 22732 9945 22744 9979
rect 22778 9976 22790 9979
rect 23014 9976 23020 9988
rect 22778 9948 23020 9976
rect 22778 9945 22790 9948
rect 22732 9939 22790 9945
rect 23014 9936 23020 9948
rect 23072 9936 23078 9988
rect 26329 9979 26387 9985
rect 26329 9945 26341 9979
rect 26375 9976 26387 9979
rect 26881 9979 26939 9985
rect 26881 9976 26893 9979
rect 26375 9948 26893 9976
rect 26375 9945 26387 9948
rect 26329 9939 26387 9945
rect 26881 9945 26893 9948
rect 26927 9945 26939 9979
rect 26881 9939 26939 9945
rect 10318 9868 10324 9920
rect 10376 9868 10382 9920
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9908 14611 9911
rect 15746 9908 15752 9920
rect 14599 9880 15752 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 19518 9868 19524 9920
rect 19576 9868 19582 9920
rect 19610 9868 19616 9920
rect 19668 9908 19674 9920
rect 26142 9908 26148 9920
rect 19668 9880 26148 9908
rect 19668 9868 19674 9880
rect 26142 9868 26148 9880
rect 26200 9868 26206 9920
rect 26234 9868 26240 9920
rect 26292 9908 26298 9920
rect 26421 9911 26479 9917
rect 26421 9908 26433 9911
rect 26292 9880 26433 9908
rect 26292 9868 26298 9880
rect 26421 9877 26433 9880
rect 26467 9877 26479 9911
rect 26421 9871 26479 9877
rect 27893 9911 27951 9917
rect 27893 9877 27905 9911
rect 27939 9908 27951 9911
rect 28000 9908 28028 10007
rect 32674 10004 32680 10016
rect 32732 10004 32738 10056
rect 33962 10004 33968 10056
rect 34020 10044 34026 10056
rect 34422 10044 34428 10056
rect 34020 10016 34428 10044
rect 34020 10004 34026 10016
rect 34422 10004 34428 10016
rect 34480 10004 34486 10056
rect 35342 10004 35348 10056
rect 35400 10004 35406 10056
rect 35618 10004 35624 10056
rect 35676 10004 35682 10056
rect 36188 10044 36216 10084
rect 36357 10081 36369 10115
rect 36403 10112 36415 10115
rect 36630 10112 36636 10124
rect 36403 10084 36636 10112
rect 36403 10081 36415 10084
rect 36357 10075 36415 10081
rect 36630 10072 36636 10084
rect 36688 10072 36694 10124
rect 37108 10121 37136 10152
rect 41524 10152 42196 10180
rect 41524 10124 41552 10152
rect 37093 10115 37151 10121
rect 37093 10081 37105 10115
rect 37139 10081 37151 10115
rect 37093 10075 37151 10081
rect 39022 10072 39028 10124
rect 39080 10072 39086 10124
rect 39206 10072 39212 10124
rect 39264 10072 39270 10124
rect 41322 10072 41328 10124
rect 41380 10072 41386 10124
rect 41506 10072 41512 10124
rect 41564 10072 41570 10124
rect 41874 10072 41880 10124
rect 41932 10072 41938 10124
rect 42168 10121 42196 10152
rect 44821 10149 44833 10183
rect 44867 10180 44879 10183
rect 45646 10180 45652 10192
rect 44867 10152 45652 10180
rect 44867 10149 44879 10152
rect 44821 10143 44879 10149
rect 45646 10140 45652 10152
rect 45704 10140 45710 10192
rect 42153 10115 42211 10121
rect 42153 10081 42165 10115
rect 42199 10081 42211 10115
rect 42153 10075 42211 10081
rect 42337 10115 42395 10121
rect 42337 10081 42349 10115
rect 42383 10112 42395 10115
rect 43162 10112 43168 10124
rect 42383 10084 43168 10112
rect 42383 10081 42395 10084
rect 42337 10075 42395 10081
rect 43162 10072 43168 10084
rect 43220 10072 43226 10124
rect 45186 10072 45192 10124
rect 45244 10112 45250 10124
rect 45557 10115 45615 10121
rect 45557 10112 45569 10115
rect 45244 10084 45569 10112
rect 45244 10072 45250 10084
rect 45557 10081 45569 10084
rect 45603 10112 45615 10115
rect 45940 10112 45968 10220
rect 46382 10208 46388 10220
rect 46440 10208 46446 10260
rect 46474 10208 46480 10260
rect 46532 10248 46538 10260
rect 48498 10248 48504 10260
rect 46532 10220 47072 10248
rect 46532 10208 46538 10220
rect 46106 10140 46112 10192
rect 46164 10140 46170 10192
rect 45603 10084 45968 10112
rect 46124 10112 46152 10140
rect 46571 10115 46629 10121
rect 46571 10112 46583 10115
rect 46124 10084 46583 10112
rect 45603 10081 45615 10084
rect 45557 10075 45615 10081
rect 46571 10081 46583 10084
rect 46617 10081 46629 10115
rect 46571 10075 46629 10081
rect 46728 10115 46786 10121
rect 46728 10081 46740 10115
rect 46774 10112 46786 10115
rect 47044 10112 47072 10220
rect 47136 10220 48504 10248
rect 47136 10189 47164 10220
rect 48498 10208 48504 10220
rect 48556 10208 48562 10260
rect 49050 10208 49056 10260
rect 49108 10248 49114 10260
rect 50430 10248 50436 10260
rect 49108 10220 50436 10248
rect 49108 10208 49114 10220
rect 50430 10208 50436 10220
rect 50488 10208 50494 10260
rect 50801 10251 50859 10257
rect 50801 10217 50813 10251
rect 50847 10248 50859 10251
rect 52454 10248 52460 10260
rect 50847 10220 52460 10248
rect 50847 10217 50859 10220
rect 50801 10211 50859 10217
rect 52454 10208 52460 10220
rect 52512 10208 52518 10260
rect 52638 10208 52644 10260
rect 52696 10208 52702 10260
rect 54110 10208 54116 10260
rect 54168 10208 54174 10260
rect 54202 10208 54208 10260
rect 54260 10208 54266 10260
rect 54941 10251 54999 10257
rect 54941 10217 54953 10251
rect 54987 10248 54999 10251
rect 55490 10248 55496 10260
rect 54987 10220 55496 10248
rect 54987 10217 54999 10220
rect 54941 10211 54999 10217
rect 55490 10208 55496 10220
rect 55548 10208 55554 10260
rect 47121 10183 47179 10189
rect 47121 10149 47133 10183
rect 47167 10149 47179 10183
rect 47121 10143 47179 10149
rect 51994 10140 52000 10192
rect 52052 10140 52058 10192
rect 46774 10084 47072 10112
rect 46774 10081 46786 10084
rect 46728 10075 46786 10081
rect 47762 10072 47768 10124
rect 47820 10112 47826 10124
rect 48222 10112 48228 10124
rect 47820 10084 48228 10112
rect 47820 10072 47826 10084
rect 48222 10072 48228 10084
rect 48280 10072 48286 10124
rect 51258 10072 51264 10124
rect 51316 10112 51322 10124
rect 52656 10121 52684 10208
rect 51721 10115 51779 10121
rect 51721 10112 51733 10115
rect 51316 10084 51733 10112
rect 51316 10072 51322 10084
rect 51721 10081 51733 10084
rect 51767 10081 51779 10115
rect 51721 10075 51779 10081
rect 52641 10115 52699 10121
rect 52641 10081 52653 10115
rect 52687 10081 52699 10115
rect 52641 10075 52699 10081
rect 36188 10016 36400 10044
rect 28252 9979 28310 9985
rect 28252 9945 28264 9979
rect 28298 9976 28310 9979
rect 28442 9976 28448 9988
rect 28298 9948 28448 9976
rect 28298 9945 28310 9948
rect 28252 9939 28310 9945
rect 28442 9936 28448 9948
rect 28500 9936 28506 9988
rect 30742 9936 30748 9988
rect 30800 9976 30806 9988
rect 30846 9979 30904 9985
rect 30846 9976 30858 9979
rect 30800 9948 30858 9976
rect 30800 9936 30806 9948
rect 30846 9945 30858 9948
rect 30892 9945 30904 9979
rect 30846 9939 30904 9945
rect 34057 9979 34115 9985
rect 34057 9945 34069 9979
rect 34103 9976 34115 9979
rect 34514 9976 34520 9988
rect 34103 9948 34520 9976
rect 34103 9945 34115 9948
rect 34057 9939 34115 9945
rect 34514 9936 34520 9948
rect 34572 9976 34578 9988
rect 36372 9976 36400 10016
rect 36538 10004 36544 10056
rect 36596 10004 36602 10056
rect 36814 10004 36820 10056
rect 36872 10044 36878 10056
rect 36909 10047 36967 10053
rect 36909 10044 36921 10047
rect 36872 10016 36921 10044
rect 36872 10004 36878 10016
rect 36909 10013 36921 10016
rect 36955 10044 36967 10047
rect 39224 10044 39252 10072
rect 36955 10016 39252 10044
rect 40977 10047 41035 10053
rect 36955 10013 36967 10016
rect 36909 10007 36967 10013
rect 40977 10013 40989 10047
rect 41023 10044 41035 10047
rect 41138 10044 41144 10056
rect 41023 10016 41144 10044
rect 41023 10013 41035 10016
rect 40977 10007 41035 10013
rect 41138 10004 41144 10016
rect 41196 10004 41202 10056
rect 41233 10047 41291 10053
rect 41233 10013 41245 10047
rect 41279 10044 41291 10047
rect 41598 10044 41604 10056
rect 41279 10016 41604 10044
rect 41279 10013 41291 10016
rect 41233 10007 41291 10013
rect 41598 10004 41604 10016
rect 41656 10004 41662 10056
rect 42429 10047 42487 10053
rect 42429 10013 42441 10047
rect 42475 10044 42487 10047
rect 42518 10044 42524 10056
rect 42475 10016 42524 10044
rect 42475 10013 42487 10016
rect 42429 10007 42487 10013
rect 42518 10004 42524 10016
rect 42576 10004 42582 10056
rect 43441 10047 43499 10053
rect 43441 10013 43453 10047
rect 43487 10013 43499 10047
rect 43441 10007 43499 10013
rect 36998 9976 37004 9988
rect 34572 9948 34836 9976
rect 36372 9948 37004 9976
rect 34572 9936 34578 9948
rect 28166 9908 28172 9920
rect 27939 9880 28172 9908
rect 27939 9877 27951 9880
rect 27893 9871 27951 9877
rect 28166 9868 28172 9880
rect 28224 9868 28230 9920
rect 29362 9868 29368 9920
rect 29420 9868 29426 9920
rect 29638 9868 29644 9920
rect 29696 9908 29702 9920
rect 29733 9911 29791 9917
rect 29733 9908 29745 9911
rect 29696 9880 29745 9908
rect 29696 9868 29702 9880
rect 29733 9877 29745 9880
rect 29779 9877 29791 9911
rect 29733 9871 29791 9877
rect 33594 9868 33600 9920
rect 33652 9868 33658 9920
rect 34698 9868 34704 9920
rect 34756 9868 34762 9920
rect 34808 9908 34836 9948
rect 36998 9936 37004 9948
rect 37056 9936 37062 9988
rect 37360 9979 37418 9985
rect 37360 9945 37372 9979
rect 37406 9976 37418 9979
rect 37550 9976 37556 9988
rect 37406 9948 37556 9976
rect 37406 9945 37418 9948
rect 37360 9939 37418 9945
rect 37550 9936 37556 9948
rect 37608 9936 37614 9988
rect 37642 9936 37648 9988
rect 37700 9976 37706 9988
rect 41506 9976 41512 9988
rect 37700 9948 41512 9976
rect 37700 9936 37706 9948
rect 41506 9936 41512 9948
rect 41564 9936 41570 9988
rect 41616 9976 41644 10004
rect 43456 9976 43484 10007
rect 46842 10004 46848 10056
rect 46900 10004 46906 10056
rect 47578 10004 47584 10056
rect 47636 10004 47642 10056
rect 49237 10047 49295 10053
rect 49237 10044 49249 10047
rect 48332 10016 49249 10044
rect 48332 9988 48360 10016
rect 49237 10013 49249 10016
rect 49283 10013 49295 10047
rect 49237 10007 49295 10013
rect 41616 9948 43484 9976
rect 43708 9979 43766 9985
rect 43708 9945 43720 9979
rect 43754 9976 43766 9979
rect 44082 9976 44088 9988
rect 43754 9948 44088 9976
rect 43754 9945 43766 9948
rect 43708 9939 43766 9945
rect 44082 9936 44088 9948
rect 44140 9936 44146 9988
rect 45373 9979 45431 9985
rect 45373 9945 45385 9979
rect 45419 9976 45431 9979
rect 46014 9976 46020 9988
rect 45419 9948 46020 9976
rect 45419 9945 45431 9948
rect 45373 9939 45431 9945
rect 46014 9936 46020 9948
rect 46072 9936 46078 9988
rect 47780 9948 48268 9976
rect 35618 9908 35624 9920
rect 34808 9880 35624 9908
rect 35618 9868 35624 9880
rect 35676 9868 35682 9920
rect 35802 9868 35808 9920
rect 35860 9908 35866 9920
rect 37458 9908 37464 9920
rect 35860 9880 37464 9908
rect 35860 9868 35866 9880
rect 37458 9868 37464 9880
rect 37516 9868 37522 9920
rect 38470 9868 38476 9920
rect 38528 9868 38534 9920
rect 38654 9868 38660 9920
rect 38712 9908 38718 9920
rect 38933 9911 38991 9917
rect 38933 9908 38945 9911
rect 38712 9880 38945 9908
rect 38712 9868 38718 9880
rect 38933 9877 38945 9880
rect 38979 9877 38991 9911
rect 38933 9871 38991 9877
rect 39114 9868 39120 9920
rect 39172 9908 39178 9920
rect 39669 9911 39727 9917
rect 39669 9908 39681 9911
rect 39172 9880 39681 9908
rect 39172 9868 39178 9880
rect 39669 9877 39681 9880
rect 39715 9908 39727 9911
rect 42794 9908 42800 9920
rect 39715 9880 42800 9908
rect 39715 9877 39727 9880
rect 39669 9871 39727 9877
rect 42794 9868 42800 9880
rect 42852 9868 42858 9920
rect 45002 9868 45008 9920
rect 45060 9868 45066 9920
rect 45462 9868 45468 9920
rect 45520 9868 45526 9920
rect 45925 9911 45983 9917
rect 45925 9877 45937 9911
rect 45971 9908 45983 9911
rect 47780 9908 47808 9948
rect 45971 9880 47808 9908
rect 45971 9877 45983 9880
rect 45925 9871 45983 9877
rect 47854 9868 47860 9920
rect 47912 9868 47918 9920
rect 48240 9908 48268 9948
rect 48314 9936 48320 9988
rect 48372 9936 48378 9988
rect 48992 9979 49050 9985
rect 48992 9945 49004 9979
rect 49038 9976 49050 9979
rect 49142 9976 49148 9988
rect 49038 9948 49148 9976
rect 49038 9945 49050 9948
rect 48992 9939 49050 9945
rect 49142 9936 49148 9948
rect 49200 9936 49206 9988
rect 49252 9976 49280 10007
rect 49970 10004 49976 10056
rect 50028 10004 50034 10056
rect 51442 10004 51448 10056
rect 51500 10004 51506 10056
rect 51626 10053 51632 10056
rect 51604 10047 51632 10053
rect 51604 10013 51616 10047
rect 51604 10007 51632 10013
rect 51626 10004 51632 10007
rect 51684 10004 51690 10056
rect 52457 10047 52515 10053
rect 52457 10013 52469 10047
rect 52503 10013 52515 10047
rect 52457 10007 52515 10013
rect 50338 9976 50344 9988
rect 49252 9948 50344 9976
rect 50338 9936 50344 9948
rect 50396 9936 50402 9988
rect 52472 9976 52500 10007
rect 52730 10004 52736 10056
rect 52788 10004 52794 10056
rect 53000 10047 53058 10053
rect 53000 10013 53012 10047
rect 53046 10044 53058 10047
rect 54220 10044 54248 10208
rect 54297 10115 54355 10121
rect 54297 10081 54309 10115
rect 54343 10081 54355 10115
rect 54297 10075 54355 10081
rect 53046 10016 54248 10044
rect 53046 10013 53058 10016
rect 53000 10007 53058 10013
rect 53466 9976 53472 9988
rect 52472 9948 53472 9976
rect 53466 9936 53472 9948
rect 53524 9936 53530 9988
rect 53834 9936 53840 9988
rect 53892 9976 53898 9988
rect 54312 9976 54340 10075
rect 56686 10072 56692 10124
rect 56744 10112 56750 10124
rect 56781 10115 56839 10121
rect 56781 10112 56793 10115
rect 56744 10084 56793 10112
rect 56744 10072 56750 10084
rect 56781 10081 56793 10084
rect 56827 10081 56839 10115
rect 56781 10075 56839 10081
rect 55122 10004 55128 10056
rect 55180 10044 55186 10056
rect 55309 10047 55367 10053
rect 55309 10044 55321 10047
rect 55180 10016 55321 10044
rect 55180 10004 55186 10016
rect 55309 10013 55321 10016
rect 55355 10044 55367 10047
rect 56704 10044 56732 10072
rect 58437 10047 58495 10053
rect 58437 10044 58449 10047
rect 55355 10016 58449 10044
rect 55355 10013 55367 10016
rect 55309 10007 55367 10013
rect 58437 10013 58449 10016
rect 58483 10013 58495 10047
rect 58437 10007 58495 10013
rect 53892 9948 54340 9976
rect 54481 9979 54539 9985
rect 53892 9936 53898 9948
rect 54481 9945 54493 9979
rect 54527 9976 54539 9979
rect 55398 9976 55404 9988
rect 54527 9948 55404 9976
rect 54527 9945 54539 9948
rect 54481 9939 54539 9945
rect 55398 9936 55404 9948
rect 55456 9936 55462 9988
rect 55576 9979 55634 9985
rect 55576 9945 55588 9979
rect 55622 9976 55634 9979
rect 56042 9976 56048 9988
rect 55622 9948 56048 9976
rect 55622 9945 55634 9948
rect 55576 9939 55634 9945
rect 56042 9936 56048 9948
rect 56100 9936 56106 9988
rect 57048 9979 57106 9985
rect 57048 9945 57060 9979
rect 57094 9976 57106 9979
rect 57606 9976 57612 9988
rect 57094 9948 57612 9976
rect 57094 9945 57106 9948
rect 57048 9939 57106 9945
rect 57606 9936 57612 9948
rect 57664 9936 57670 9988
rect 48406 9908 48412 9920
rect 48240 9880 48412 9908
rect 48406 9868 48412 9880
rect 48464 9868 48470 9920
rect 49326 9868 49332 9920
rect 49384 9868 49390 9920
rect 50430 9868 50436 9920
rect 50488 9908 50494 9920
rect 51442 9908 51448 9920
rect 50488 9880 51448 9908
rect 50488 9868 50494 9880
rect 51442 9868 51448 9880
rect 51500 9868 51506 9920
rect 54573 9911 54631 9917
rect 54573 9877 54585 9911
rect 54619 9908 54631 9911
rect 56410 9908 56416 9920
rect 54619 9880 56416 9908
rect 54619 9877 54631 9880
rect 54573 9871 54631 9877
rect 56410 9868 56416 9880
rect 56468 9868 56474 9920
rect 56686 9868 56692 9920
rect 56744 9868 56750 9920
rect 58158 9868 58164 9920
rect 58216 9868 58222 9920
rect 1104 9818 59040 9840
rect 1104 9766 15394 9818
rect 15446 9766 15458 9818
rect 15510 9766 15522 9818
rect 15574 9766 15586 9818
rect 15638 9766 15650 9818
rect 15702 9766 29838 9818
rect 29890 9766 29902 9818
rect 29954 9766 29966 9818
rect 30018 9766 30030 9818
rect 30082 9766 30094 9818
rect 30146 9766 44282 9818
rect 44334 9766 44346 9818
rect 44398 9766 44410 9818
rect 44462 9766 44474 9818
rect 44526 9766 44538 9818
rect 44590 9766 58726 9818
rect 58778 9766 58790 9818
rect 58842 9766 58854 9818
rect 58906 9766 58918 9818
rect 58970 9766 58982 9818
rect 59034 9766 59040 9818
rect 1104 9744 59040 9766
rect 4246 9664 4252 9716
rect 4304 9664 4310 9716
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 5353 9707 5411 9713
rect 5353 9704 5365 9707
rect 4856 9676 5365 9704
rect 4856 9664 4862 9676
rect 5353 9673 5365 9676
rect 5399 9673 5411 9707
rect 5353 9667 5411 9673
rect 5442 9664 5448 9716
rect 5500 9664 5506 9716
rect 12986 9664 12992 9716
rect 13044 9664 13050 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 25222 9704 25228 9716
rect 18288 9676 25228 9704
rect 18288 9664 18294 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 29454 9664 29460 9716
rect 29512 9664 29518 9716
rect 34698 9664 34704 9716
rect 34756 9704 34762 9716
rect 36170 9704 36176 9716
rect 34756 9676 36176 9704
rect 34756 9664 34762 9676
rect 36170 9664 36176 9676
rect 36228 9664 36234 9716
rect 36357 9707 36415 9713
rect 36357 9673 36369 9707
rect 36403 9704 36415 9707
rect 36630 9704 36636 9716
rect 36403 9676 36636 9704
rect 36403 9673 36415 9676
rect 36357 9667 36415 9673
rect 36630 9664 36636 9676
rect 36688 9664 36694 9716
rect 36998 9664 37004 9716
rect 37056 9704 37062 9716
rect 37826 9704 37832 9716
rect 37056 9676 37832 9704
rect 37056 9664 37062 9676
rect 37826 9664 37832 9676
rect 37884 9664 37890 9716
rect 39298 9704 39304 9716
rect 38672 9676 39304 9704
rect 2216 9639 2274 9645
rect 2216 9605 2228 9639
rect 2262 9636 2274 9639
rect 3050 9636 3056 9648
rect 2262 9608 3056 9636
rect 2262 9605 2274 9608
rect 2216 9599 2274 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4212 9608 4844 9636
rect 4212 9596 4218 9608
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2038 9568 2044 9580
rect 1995 9540 2044 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3344 9540 3525 9568
rect 3344 9444 3372 9540
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 3513 9531 3571 9537
rect 3804 9540 4445 9568
rect 3804 9444 3832 9540
rect 4433 9537 4445 9540
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 4816 9577 4844 9608
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 5166 9596 5172 9648
rect 5224 9596 5230 9648
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4724 9500 4752 9531
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 5460 9577 5488 9664
rect 38672 9648 38700 9676
rect 39298 9664 39304 9676
rect 39356 9704 39362 9716
rect 40957 9707 41015 9713
rect 39356 9676 40356 9704
rect 39356 9664 39362 9676
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 5868 9608 6377 9636
rect 5868 9596 5874 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 6917 9639 6975 9645
rect 6917 9605 6929 9639
rect 6963 9636 6975 9639
rect 8754 9636 8760 9648
rect 6963 9608 8760 9636
rect 6963 9605 6975 9608
rect 6917 9599 6975 9605
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 10220 9639 10278 9645
rect 10220 9605 10232 9639
rect 10266 9636 10278 9639
rect 10318 9636 10324 9648
rect 10266 9608 10324 9636
rect 10266 9605 10278 9608
rect 10220 9599 10278 9605
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 15188 9639 15246 9645
rect 13096 9608 14504 9636
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9568 9459 9571
rect 10042 9568 10048 9580
rect 9447 9540 10048 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 12618 9568 12624 9580
rect 12391 9540 12624 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13096 9577 13124 9608
rect 14476 9580 14504 9608
rect 15188 9605 15200 9639
rect 15234 9636 15246 9639
rect 15286 9636 15292 9648
rect 15234 9608 15292 9636
rect 15234 9605 15246 9608
rect 15188 9599 15246 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 17678 9596 17684 9648
rect 17736 9636 17742 9648
rect 19242 9636 19248 9648
rect 17736 9608 19248 9636
rect 17736 9596 17742 9608
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13170 9528 13176 9580
rect 13228 9568 13234 9580
rect 13337 9571 13395 9577
rect 13337 9568 13349 9571
rect 13228 9540 13349 9568
rect 13228 9528 13234 9540
rect 13337 9537 13349 9540
rect 13383 9537 13395 9571
rect 13337 9531 13395 9537
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14516 9540 14933 9568
rect 14516 9528 14522 9540
rect 14921 9537 14933 9540
rect 14967 9568 14979 9571
rect 17696 9568 17724 9596
rect 14967 9540 17724 9568
rect 17793 9571 17851 9577
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 17793 9537 17805 9571
rect 17839 9568 17851 9571
rect 17954 9568 17960 9580
rect 17839 9540 17960 9568
rect 17839 9537 17851 9540
rect 17793 9531 17851 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18064 9577 18092 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19420 9639 19478 9645
rect 19420 9605 19432 9639
rect 19466 9636 19478 9639
rect 19518 9636 19524 9648
rect 19466 9608 19524 9636
rect 19466 9605 19478 9608
rect 19420 9599 19478 9605
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 22278 9596 22284 9648
rect 22336 9596 22342 9648
rect 24213 9639 24271 9645
rect 24213 9605 24225 9639
rect 24259 9636 24271 9639
rect 25498 9636 25504 9648
rect 24259 9608 25504 9636
rect 24259 9605 24271 9608
rect 24213 9599 24271 9605
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 27062 9596 27068 9648
rect 27120 9636 27126 9648
rect 27341 9639 27399 9645
rect 27341 9636 27353 9639
rect 27120 9608 27353 9636
rect 27120 9596 27126 9608
rect 27341 9605 27353 9608
rect 27387 9605 27399 9639
rect 27341 9599 27399 9605
rect 28344 9639 28402 9645
rect 28344 9605 28356 9639
rect 28390 9636 28402 9639
rect 28534 9636 28540 9648
rect 28390 9608 28540 9636
rect 28390 9605 28402 9608
rect 28344 9599 28402 9605
rect 28534 9596 28540 9608
rect 28592 9596 28598 9648
rect 35434 9636 35440 9648
rect 34624 9608 35440 9636
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 18322 9528 18328 9580
rect 18380 9568 18386 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18380 9540 18521 9568
rect 18380 9528 18386 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 19153 9571 19211 9577
rect 19153 9537 19165 9571
rect 19199 9568 19211 9571
rect 19260 9568 19288 9596
rect 19199 9540 19288 9568
rect 22296 9568 22324 9596
rect 34624 9580 34652 9608
rect 35434 9596 35440 9608
rect 35492 9596 35498 9648
rect 37093 9639 37151 9645
rect 37093 9605 37105 9639
rect 37139 9636 37151 9639
rect 37918 9636 37924 9648
rect 37139 9608 37924 9636
rect 37139 9605 37151 9608
rect 37093 9599 37151 9605
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 22296 9540 22385 9568
rect 19199 9537 19211 9540
rect 19153 9531 19211 9537
rect 22373 9537 22385 9540
rect 22419 9537 22431 9571
rect 22373 9531 22431 9537
rect 22640 9571 22698 9577
rect 22640 9537 22652 9571
rect 22686 9568 22698 9571
rect 23014 9568 23020 9580
rect 22686 9540 23020 9568
rect 22686 9537 22698 9540
rect 22640 9531 22698 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 23474 9528 23480 9580
rect 23532 9568 23538 9580
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 23532 9540 24317 9568
rect 23532 9528 23538 9540
rect 24305 9537 24317 9540
rect 24351 9568 24363 9571
rect 26349 9571 26407 9577
rect 24351 9540 25544 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 25516 9512 25544 9540
rect 26349 9537 26361 9571
rect 26395 9568 26407 9571
rect 26510 9568 26516 9580
rect 26395 9540 26516 9568
rect 26395 9537 26407 9540
rect 26349 9531 26407 9537
rect 26510 9528 26516 9540
rect 26568 9528 26574 9580
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 29638 9568 29644 9580
rect 29595 9540 29644 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 29638 9528 29644 9540
rect 29696 9568 29702 9580
rect 29696 9540 29960 9568
rect 29696 9528 29702 9540
rect 4448 9472 4752 9500
rect 3326 9392 3332 9444
rect 3384 9392 3390 9444
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 3786 9432 3792 9444
rect 3743 9404 3792 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 3786 9392 3792 9404
rect 3844 9392 3850 9444
rect 4448 9376 4476 9472
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7616 9472 8217 9500
rect 7616 9460 7622 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 8938 9460 8944 9512
rect 8996 9460 9002 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9732 9472 9965 9500
rect 9732 9460 9738 9472
rect 9953 9469 9965 9472
rect 9999 9469 10011 9503
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 9953 9463 10011 9469
rect 11348 9472 12081 9500
rect 11348 9441 11376 9472
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 18601 9503 18659 9509
rect 18601 9469 18613 9503
rect 18647 9469 18659 9503
rect 18601 9463 18659 9469
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9401 11391 9435
rect 11333 9395 11391 9401
rect 4430 9324 4436 9376
rect 4488 9324 4494 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 6638 9364 6644 9376
rect 5500 9336 6644 9364
rect 5500 9324 5506 9336
rect 6638 9324 6644 9336
rect 6696 9364 6702 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6696 9336 7205 9364
rect 6696 9324 6702 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7650 9324 7656 9376
rect 7708 9324 7714 9376
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 8570 9364 8576 9376
rect 8435 9336 8576 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 10594 9364 10600 9376
rect 9815 9336 10600 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 11514 9324 11520 9376
rect 11572 9324 11578 9376
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14424 9336 14473 9364
rect 14424 9324 14430 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 14461 9327 14519 9333
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 15838 9364 15844 9376
rect 14875 9336 15844 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 16301 9367 16359 9373
rect 16301 9333 16313 9367
rect 16347 9364 16359 9367
rect 16574 9364 16580 9376
rect 16347 9336 16580 9364
rect 16347 9333 16359 9336
rect 16301 9327 16359 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16666 9324 16672 9376
rect 16724 9324 16730 9376
rect 18138 9324 18144 9376
rect 18196 9324 18202 9376
rect 18616 9364 18644 9463
rect 18782 9460 18788 9512
rect 18840 9460 18846 9512
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 20533 9435 20591 9441
rect 20533 9401 20545 9435
rect 20579 9432 20591 9435
rect 20640 9432 20668 9463
rect 24210 9460 24216 9512
rect 24268 9460 24274 9512
rect 24394 9460 24400 9512
rect 24452 9460 24458 9512
rect 25498 9460 25504 9512
rect 25556 9460 25562 9512
rect 26605 9503 26663 9509
rect 26605 9469 26617 9503
rect 26651 9500 26663 9503
rect 26694 9500 26700 9512
rect 26651 9472 26700 9500
rect 26651 9469 26663 9472
rect 26605 9463 26663 9469
rect 26694 9460 26700 9472
rect 26752 9500 26758 9512
rect 27893 9503 27951 9509
rect 27893 9500 27905 9503
rect 26752 9472 27905 9500
rect 26752 9460 26758 9472
rect 27893 9469 27905 9472
rect 27939 9500 27951 9503
rect 28074 9500 28080 9512
rect 27939 9472 28080 9500
rect 27939 9469 27951 9472
rect 27893 9463 27951 9469
rect 28074 9460 28080 9472
rect 28132 9460 28138 9512
rect 29733 9503 29791 9509
rect 29733 9469 29745 9503
rect 29779 9469 29791 9503
rect 29932 9500 29960 9540
rect 30558 9528 30564 9580
rect 30616 9577 30622 9580
rect 30616 9571 30644 9577
rect 30632 9537 30644 9571
rect 30616 9531 30644 9537
rect 32668 9571 32726 9577
rect 32668 9537 32680 9571
rect 32714 9568 32726 9571
rect 33134 9568 33140 9580
rect 32714 9540 33140 9568
rect 32714 9537 32726 9540
rect 32668 9531 32726 9537
rect 30616 9528 30622 9531
rect 33134 9528 33140 9540
rect 33192 9528 33198 9580
rect 34517 9571 34575 9577
rect 34517 9537 34529 9571
rect 34563 9568 34575 9571
rect 34606 9568 34612 9580
rect 34563 9540 34612 9568
rect 34563 9537 34575 9540
rect 34517 9531 34575 9537
rect 34606 9528 34612 9540
rect 34664 9528 34670 9580
rect 34790 9577 34796 9580
rect 34784 9531 34796 9577
rect 34790 9528 34796 9531
rect 34848 9528 34854 9580
rect 35158 9528 35164 9580
rect 35216 9568 35222 9580
rect 36265 9571 36323 9577
rect 36265 9568 36277 9571
rect 35216 9540 36277 9568
rect 35216 9528 35222 9540
rect 36265 9537 36277 9540
rect 36311 9537 36323 9571
rect 36265 9531 36323 9537
rect 30282 9500 30288 9512
rect 29932 9472 30288 9500
rect 29733 9463 29791 9469
rect 20579 9404 20668 9432
rect 23753 9435 23811 9441
rect 20579 9401 20591 9404
rect 20533 9395 20591 9401
rect 23753 9401 23765 9435
rect 23799 9432 23811 9435
rect 24228 9432 24256 9460
rect 23799 9404 24256 9432
rect 24857 9435 24915 9441
rect 23799 9401 23811 9404
rect 23753 9395 23811 9401
rect 24857 9401 24869 9435
rect 24903 9432 24915 9435
rect 25130 9432 25136 9444
rect 24903 9404 25136 9432
rect 24903 9401 24915 9404
rect 24857 9395 24915 9401
rect 25130 9392 25136 9404
rect 25188 9392 25194 9444
rect 19426 9364 19432 9376
rect 18616 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 21266 9324 21272 9376
rect 21324 9324 21330 9376
rect 23842 9324 23848 9376
rect 23900 9324 23906 9376
rect 25038 9324 25044 9376
rect 25096 9364 25102 9376
rect 25225 9367 25283 9373
rect 25225 9364 25237 9367
rect 25096 9336 25237 9364
rect 25096 9324 25102 9336
rect 25225 9333 25237 9336
rect 25271 9333 25283 9367
rect 29748 9364 29776 9463
rect 30282 9460 30288 9472
rect 30340 9460 30346 9512
rect 30466 9460 30472 9512
rect 30524 9460 30530 9512
rect 30745 9503 30803 9509
rect 30745 9469 30757 9503
rect 30791 9500 30803 9503
rect 31389 9503 31447 9509
rect 30791 9472 31340 9500
rect 30791 9469 30803 9472
rect 30745 9463 30803 9469
rect 30190 9392 30196 9444
rect 30248 9392 30254 9444
rect 31312 9432 31340 9472
rect 31389 9469 31401 9503
rect 31435 9500 31447 9503
rect 31938 9500 31944 9512
rect 31435 9472 31944 9500
rect 31435 9469 31447 9472
rect 31389 9463 31447 9469
rect 31938 9460 31944 9472
rect 31996 9460 32002 9512
rect 32122 9460 32128 9512
rect 32180 9500 32186 9512
rect 32401 9503 32459 9509
rect 32401 9500 32413 9503
rect 32180 9472 32413 9500
rect 32180 9460 32186 9472
rect 32401 9469 32413 9472
rect 32447 9469 32459 9503
rect 32401 9463 32459 9469
rect 36173 9503 36231 9509
rect 36173 9469 36185 9503
rect 36219 9500 36231 9503
rect 37108 9500 37136 9599
rect 37918 9596 37924 9608
rect 37976 9596 37982 9648
rect 38105 9639 38163 9645
rect 38105 9605 38117 9639
rect 38151 9636 38163 9639
rect 38654 9636 38660 9648
rect 38151 9608 38660 9636
rect 38151 9605 38163 9608
rect 38105 9599 38163 9605
rect 38654 9596 38660 9608
rect 38712 9596 38718 9648
rect 40328 9636 40356 9676
rect 40957 9673 40969 9707
rect 41003 9704 41015 9707
rect 41322 9704 41328 9716
rect 41003 9676 41328 9704
rect 41003 9673 41015 9676
rect 40957 9667 41015 9673
rect 40865 9639 40923 9645
rect 40865 9636 40877 9639
rect 40328 9608 40877 9636
rect 40865 9605 40877 9608
rect 40911 9605 40923 9639
rect 40865 9599 40923 9605
rect 37458 9528 37464 9580
rect 37516 9528 37522 9580
rect 38010 9528 38016 9580
rect 38068 9568 38074 9580
rect 38068 9540 38792 9568
rect 38068 9528 38074 9540
rect 36219 9472 37136 9500
rect 37476 9500 37504 9528
rect 38197 9503 38255 9509
rect 38197 9500 38209 9503
rect 37476 9472 38209 9500
rect 36219 9469 36231 9472
rect 36173 9463 36231 9469
rect 38197 9469 38209 9472
rect 38243 9500 38255 9503
rect 38562 9500 38568 9512
rect 38243 9472 38568 9500
rect 38243 9469 38255 9472
rect 38197 9463 38255 9469
rect 38562 9460 38568 9472
rect 38620 9460 38626 9512
rect 38764 9500 38792 9540
rect 39298 9528 39304 9580
rect 39356 9528 39362 9580
rect 39574 9528 39580 9580
rect 39632 9528 39638 9580
rect 40313 9571 40371 9577
rect 40313 9537 40325 9571
rect 40359 9568 40371 9571
rect 40972 9568 41000 9667
rect 41322 9664 41328 9676
rect 41380 9664 41386 9716
rect 41506 9664 41512 9716
rect 41564 9664 41570 9716
rect 41598 9664 41604 9716
rect 41656 9704 41662 9716
rect 42518 9704 42524 9716
rect 41656 9676 42524 9704
rect 41656 9664 41662 9676
rect 42518 9664 42524 9676
rect 42576 9704 42582 9716
rect 43901 9707 43959 9713
rect 43901 9704 43913 9707
rect 42576 9676 43913 9704
rect 42576 9664 42582 9676
rect 43901 9673 43913 9676
rect 43947 9704 43959 9707
rect 43990 9704 43996 9716
rect 43947 9676 43996 9704
rect 43947 9673 43959 9676
rect 43901 9667 43959 9673
rect 43990 9664 43996 9676
rect 44048 9664 44054 9716
rect 44082 9664 44088 9716
rect 44140 9664 44146 9716
rect 45189 9707 45247 9713
rect 45189 9673 45201 9707
rect 45235 9704 45247 9707
rect 45462 9704 45468 9716
rect 45235 9676 45468 9704
rect 45235 9673 45247 9676
rect 45189 9667 45247 9673
rect 41524 9636 41552 9664
rect 41969 9639 42027 9645
rect 41969 9636 41981 9639
rect 41524 9608 41981 9636
rect 41969 9605 41981 9608
rect 42015 9605 42027 9639
rect 41969 9599 42027 9605
rect 40359 9540 41000 9568
rect 44729 9571 44787 9577
rect 40359 9537 40371 9540
rect 40313 9531 40371 9537
rect 44729 9537 44741 9571
rect 44775 9568 44787 9571
rect 45002 9568 45008 9580
rect 44775 9540 45008 9568
rect 44775 9537 44787 9540
rect 44729 9531 44787 9537
rect 45002 9528 45008 9540
rect 45060 9528 45066 9580
rect 45204 9568 45232 9667
rect 45462 9664 45468 9676
rect 45520 9664 45526 9716
rect 46014 9664 46020 9716
rect 46072 9704 46078 9716
rect 46293 9707 46351 9713
rect 46293 9704 46305 9707
rect 46072 9676 46305 9704
rect 46072 9664 46078 9676
rect 46293 9673 46305 9676
rect 46339 9704 46351 9707
rect 46382 9704 46388 9716
rect 46339 9676 46388 9704
rect 46339 9673 46351 9676
rect 46293 9667 46351 9673
rect 46382 9664 46388 9676
rect 46440 9664 46446 9716
rect 46474 9664 46480 9716
rect 46532 9704 46538 9716
rect 46658 9704 46664 9716
rect 46532 9676 46664 9704
rect 46532 9664 46538 9676
rect 46658 9664 46664 9676
rect 46716 9664 46722 9716
rect 47029 9707 47087 9713
rect 47029 9673 47041 9707
rect 47075 9704 47087 9707
rect 47762 9704 47768 9716
rect 47075 9676 47768 9704
rect 47075 9673 47087 9676
rect 47029 9667 47087 9673
rect 47762 9664 47768 9676
rect 47820 9664 47826 9716
rect 53101 9707 53159 9713
rect 53101 9673 53113 9707
rect 53147 9704 53159 9707
rect 53466 9704 53472 9716
rect 53147 9676 53472 9704
rect 53147 9673 53159 9676
rect 53101 9667 53159 9673
rect 53466 9664 53472 9676
rect 53524 9664 53530 9716
rect 54662 9664 54668 9716
rect 54720 9704 54726 9716
rect 54720 9676 55076 9704
rect 54720 9664 54726 9676
rect 45281 9639 45339 9645
rect 45281 9605 45293 9639
rect 45327 9636 45339 9639
rect 46198 9636 46204 9648
rect 45327 9608 46204 9636
rect 45327 9605 45339 9608
rect 45281 9599 45339 9605
rect 46198 9596 46204 9608
rect 46256 9636 46262 9648
rect 46842 9636 46848 9648
rect 46256 9608 46848 9636
rect 46256 9596 46262 9608
rect 46842 9596 46848 9608
rect 46900 9596 46906 9648
rect 48584 9639 48642 9645
rect 48584 9605 48596 9639
rect 48630 9636 48642 9639
rect 49326 9636 49332 9648
rect 48630 9608 49332 9636
rect 48630 9605 48642 9608
rect 48584 9599 48642 9605
rect 49326 9596 49332 9608
rect 49384 9596 49390 9648
rect 54012 9639 54070 9645
rect 54012 9605 54024 9639
rect 54058 9636 54070 9639
rect 54938 9636 54944 9648
rect 54058 9608 54944 9636
rect 54058 9605 54070 9608
rect 54012 9599 54070 9605
rect 54938 9596 54944 9608
rect 54996 9596 55002 9648
rect 45204 9540 45600 9568
rect 39439 9503 39497 9509
rect 39439 9500 39451 9503
rect 38764 9472 39451 9500
rect 39439 9469 39451 9472
rect 39485 9469 39497 9503
rect 39439 9463 39497 9469
rect 40494 9460 40500 9512
rect 40552 9460 40558 9512
rect 40678 9460 40684 9512
rect 40736 9460 40742 9512
rect 45465 9503 45523 9509
rect 45465 9469 45477 9503
rect 45511 9469 45523 9503
rect 45572 9500 45600 9540
rect 45646 9528 45652 9580
rect 45704 9528 45710 9580
rect 46937 9571 46995 9577
rect 46937 9568 46949 9571
rect 46308 9540 46949 9568
rect 46308 9500 46336 9540
rect 46937 9537 46949 9540
rect 46983 9568 46995 9571
rect 47762 9568 47768 9580
rect 46983 9540 47768 9568
rect 46983 9537 46995 9540
rect 46937 9531 46995 9537
rect 47762 9528 47768 9540
rect 47820 9528 47826 9580
rect 47854 9528 47860 9580
rect 47912 9568 47918 9580
rect 48133 9571 48191 9577
rect 48133 9568 48145 9571
rect 47912 9540 48145 9568
rect 47912 9528 47918 9540
rect 48133 9537 48145 9540
rect 48179 9537 48191 9571
rect 48133 9531 48191 9537
rect 48314 9528 48320 9580
rect 48372 9528 48378 9580
rect 49694 9528 49700 9580
rect 49752 9568 49758 9580
rect 49789 9571 49847 9577
rect 49789 9568 49801 9571
rect 49752 9540 49801 9568
rect 49752 9528 49758 9540
rect 49789 9537 49801 9540
rect 49835 9537 49847 9571
rect 49789 9531 49847 9537
rect 51994 9528 52000 9580
rect 52052 9568 52058 9580
rect 53009 9571 53067 9577
rect 53009 9568 53021 9571
rect 52052 9540 53021 9568
rect 52052 9528 52058 9540
rect 53009 9537 53021 9540
rect 53055 9537 53067 9571
rect 53009 9531 53067 9537
rect 47121 9503 47179 9509
rect 47121 9500 47133 9503
rect 45572 9472 46336 9500
rect 46400 9472 47133 9500
rect 45465 9463 45523 9469
rect 34333 9435 34391 9441
rect 34333 9432 34345 9435
rect 31312 9404 31800 9432
rect 30834 9364 30840 9376
rect 29748 9336 30840 9364
rect 25225 9327 25283 9333
rect 30834 9324 30840 9336
rect 30892 9324 30898 9376
rect 31772 9373 31800 9404
rect 33704 9404 34345 9432
rect 31757 9367 31815 9373
rect 31757 9333 31769 9367
rect 31803 9364 31815 9367
rect 32030 9364 32036 9376
rect 31803 9336 32036 9364
rect 31803 9333 31815 9336
rect 31757 9327 31815 9333
rect 32030 9324 32036 9336
rect 32088 9324 32094 9376
rect 32398 9324 32404 9376
rect 32456 9364 32462 9376
rect 33704 9364 33732 9404
rect 34333 9401 34345 9404
rect 34379 9401 34391 9435
rect 34333 9395 34391 9401
rect 39853 9435 39911 9441
rect 39853 9401 39865 9435
rect 39899 9401 39911 9435
rect 39853 9395 39911 9401
rect 32456 9336 33732 9364
rect 32456 9324 32462 9336
rect 33778 9324 33784 9376
rect 33836 9324 33842 9376
rect 35894 9324 35900 9376
rect 35952 9324 35958 9376
rect 36722 9324 36728 9376
rect 36780 9324 36786 9376
rect 37642 9324 37648 9376
rect 37700 9324 37706 9376
rect 38657 9367 38715 9373
rect 38657 9333 38669 9367
rect 38703 9364 38715 9367
rect 39298 9364 39304 9376
rect 38703 9336 39304 9364
rect 38703 9333 38715 9336
rect 38657 9327 38715 9333
rect 39298 9324 39304 9336
rect 39356 9324 39362 9376
rect 39482 9324 39488 9376
rect 39540 9364 39546 9376
rect 39868 9364 39896 9395
rect 44818 9392 44824 9444
rect 44876 9392 44882 9444
rect 45480 9432 45508 9463
rect 45554 9432 45560 9444
rect 45480 9404 45560 9432
rect 45554 9392 45560 9404
rect 45612 9392 45618 9444
rect 46400 9376 46428 9472
rect 47121 9469 47133 9472
rect 47167 9469 47179 9503
rect 52181 9503 52239 9509
rect 52181 9500 52193 9503
rect 47121 9463 47179 9469
rect 51046 9472 52193 9500
rect 49697 9435 49755 9441
rect 49697 9401 49709 9435
rect 49743 9432 49755 9435
rect 51046 9432 51074 9472
rect 52181 9469 52193 9472
rect 52227 9469 52239 9503
rect 52181 9463 52239 9469
rect 52917 9503 52975 9509
rect 52917 9469 52929 9503
rect 52963 9469 52975 9503
rect 52917 9463 52975 9469
rect 49743 9404 51074 9432
rect 49743 9401 49755 9404
rect 49697 9395 49755 9401
rect 52932 9376 52960 9463
rect 53742 9460 53748 9512
rect 53800 9460 53806 9512
rect 55048 9500 55076 9676
rect 56042 9664 56048 9716
rect 56100 9664 56106 9716
rect 57241 9707 57299 9713
rect 57241 9673 57253 9707
rect 57287 9704 57299 9707
rect 57330 9704 57336 9716
rect 57287 9676 57336 9704
rect 57287 9673 57299 9676
rect 57241 9667 57299 9673
rect 57330 9664 57336 9676
rect 57388 9704 57394 9716
rect 57885 9707 57943 9713
rect 57885 9704 57897 9707
rect 57388 9676 57897 9704
rect 57388 9664 57394 9676
rect 57885 9673 57897 9676
rect 57931 9673 57943 9707
rect 57885 9667 57943 9673
rect 55493 9639 55551 9645
rect 55493 9605 55505 9639
rect 55539 9636 55551 9639
rect 56594 9636 56600 9648
rect 55539 9608 56600 9636
rect 55539 9605 55551 9608
rect 55493 9599 55551 9605
rect 56594 9596 56600 9608
rect 56652 9596 56658 9648
rect 55398 9528 55404 9580
rect 55456 9568 55462 9580
rect 55585 9571 55643 9577
rect 55585 9568 55597 9571
rect 55456 9540 55597 9568
rect 55456 9528 55462 9540
rect 55585 9537 55597 9540
rect 55631 9568 55643 9571
rect 56962 9568 56968 9580
rect 55631 9540 56968 9568
rect 55631 9537 55643 9540
rect 55585 9531 55643 9537
rect 56962 9528 56968 9540
rect 57020 9568 57026 9580
rect 57020 9540 57376 9568
rect 57020 9528 57026 9540
rect 57348 9512 57376 9540
rect 58158 9528 58164 9580
rect 58216 9568 58222 9580
rect 58437 9571 58495 9577
rect 58437 9568 58449 9571
rect 58216 9540 58449 9568
rect 58216 9528 58222 9540
rect 58437 9537 58449 9540
rect 58483 9537 58495 9571
rect 58437 9531 58495 9537
rect 55309 9503 55367 9509
rect 55309 9500 55321 9503
rect 55048 9472 55321 9500
rect 55309 9469 55321 9472
rect 55355 9469 55367 9503
rect 55309 9463 55367 9469
rect 56597 9503 56655 9509
rect 56597 9469 56609 9503
rect 56643 9469 56655 9503
rect 56597 9463 56655 9469
rect 55324 9432 55352 9463
rect 55582 9432 55588 9444
rect 55324 9404 55588 9432
rect 55582 9392 55588 9404
rect 55640 9392 55646 9444
rect 55953 9435 56011 9441
rect 55953 9401 55965 9435
rect 55999 9432 56011 9435
rect 56612 9432 56640 9463
rect 57330 9460 57336 9512
rect 57388 9460 57394 9512
rect 57422 9460 57428 9512
rect 57480 9460 57486 9512
rect 55999 9404 56640 9432
rect 55999 9401 56011 9404
rect 55953 9395 56011 9401
rect 39540 9336 39896 9364
rect 39540 9324 39546 9336
rect 41322 9324 41328 9376
rect 41380 9324 41386 9376
rect 46382 9324 46388 9376
rect 46440 9324 46446 9376
rect 46566 9324 46572 9376
rect 46624 9324 46630 9376
rect 47578 9324 47584 9376
rect 47636 9364 47642 9376
rect 47946 9364 47952 9376
rect 47636 9336 47952 9364
rect 47636 9324 47642 9336
rect 47946 9324 47952 9336
rect 48004 9324 48010 9376
rect 50338 9324 50344 9376
rect 50396 9364 50402 9376
rect 51077 9367 51135 9373
rect 51077 9364 51089 9367
rect 50396 9336 51089 9364
rect 50396 9324 50402 9336
rect 51077 9333 51089 9336
rect 51123 9333 51135 9367
rect 51077 9327 51135 9333
rect 51350 9324 51356 9376
rect 51408 9364 51414 9376
rect 51626 9364 51632 9376
rect 51408 9336 51632 9364
rect 51408 9324 51414 9336
rect 51626 9324 51632 9336
rect 51684 9324 51690 9376
rect 52914 9324 52920 9376
rect 52972 9324 52978 9376
rect 53469 9367 53527 9373
rect 53469 9333 53481 9367
rect 53515 9364 53527 9367
rect 54754 9364 54760 9376
rect 53515 9336 54760 9364
rect 53515 9333 53527 9336
rect 53469 9327 53527 9333
rect 54754 9324 54760 9336
rect 54812 9324 54818 9376
rect 55125 9367 55183 9373
rect 55125 9333 55137 9367
rect 55171 9364 55183 9367
rect 55306 9364 55312 9376
rect 55171 9336 55312 9364
rect 55171 9333 55183 9336
rect 55125 9327 55183 9333
rect 55306 9324 55312 9336
rect 55364 9324 55370 9376
rect 56870 9324 56876 9376
rect 56928 9324 56934 9376
rect 1104 9274 58880 9296
rect 1104 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 22616 9274
rect 22668 9222 22680 9274
rect 22732 9222 22744 9274
rect 22796 9222 22808 9274
rect 22860 9222 22872 9274
rect 22924 9222 37060 9274
rect 37112 9222 37124 9274
rect 37176 9222 37188 9274
rect 37240 9222 37252 9274
rect 37304 9222 37316 9274
rect 37368 9222 51504 9274
rect 51556 9222 51568 9274
rect 51620 9222 51632 9274
rect 51684 9222 51696 9274
rect 51748 9222 51760 9274
rect 51812 9222 58880 9274
rect 1104 9200 58880 9222
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6362 9160 6368 9172
rect 6144 9132 6368 9160
rect 6144 9120 6150 9132
rect 6362 9120 6368 9132
rect 6420 9160 6426 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 6420 9132 6469 9160
rect 6420 9120 6426 9132
rect 6457 9129 6469 9132
rect 6503 9129 6515 9163
rect 6457 9123 6515 9129
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7006 9160 7012 9172
rect 6963 9132 7012 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 7156 9132 7205 9160
rect 7156 9120 7162 9132
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 8938 9160 8944 9172
rect 8803 9132 8944 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 10413 9163 10471 9169
rect 10413 9129 10425 9163
rect 10459 9160 10471 9163
rect 10870 9160 10876 9172
rect 10459 9132 10876 9160
rect 10459 9129 10471 9132
rect 10413 9123 10471 9129
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11514 9120 11520 9172
rect 11572 9120 11578 9172
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16206 9160 16212 9172
rect 15979 9132 16212 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 18046 9120 18052 9172
rect 18104 9120 18110 9172
rect 18138 9120 18144 9172
rect 18196 9120 18202 9172
rect 19613 9163 19671 9169
rect 19613 9129 19625 9163
rect 19659 9160 19671 9163
rect 20070 9160 20076 9172
rect 19659 9132 20076 9160
rect 19659 9129 19671 9132
rect 19613 9123 19671 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 23014 9120 23020 9172
rect 23072 9160 23078 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 23072 9132 23305 9160
rect 23072 9120 23078 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 23293 9123 23351 9129
rect 23842 9120 23848 9172
rect 23900 9120 23906 9172
rect 25038 9120 25044 9172
rect 25096 9120 25102 9172
rect 26510 9120 26516 9172
rect 26568 9120 26574 9172
rect 28074 9120 28080 9172
rect 28132 9160 28138 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 28132 9132 29837 9160
rect 28132 9120 28138 9132
rect 29825 9129 29837 9132
rect 29871 9160 29883 9163
rect 31110 9160 31116 9172
rect 29871 9132 31116 9160
rect 29871 9129 29883 9132
rect 29825 9123 29883 9129
rect 31110 9120 31116 9132
rect 31168 9120 31174 9172
rect 31754 9120 31760 9172
rect 31812 9120 31818 9172
rect 33134 9120 33140 9172
rect 33192 9120 33198 9172
rect 33778 9120 33784 9172
rect 33836 9120 33842 9172
rect 34514 9120 34520 9172
rect 34572 9120 34578 9172
rect 36449 9163 36507 9169
rect 36449 9129 36461 9163
rect 36495 9160 36507 9163
rect 36538 9160 36544 9172
rect 36495 9132 36544 9160
rect 36495 9129 36507 9132
rect 36449 9123 36507 9129
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 10502 9092 10508 9104
rect 8904 9064 10508 9092
rect 8904 9052 8910 9064
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 11532 9092 11560 9120
rect 10888 9064 11560 9092
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 4522 9024 4528 9036
rect 4387 8996 4528 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 10888 9033 10916 9064
rect 11606 9052 11612 9104
rect 11664 9052 11670 9104
rect 10873 9027 10931 9033
rect 8588 8996 10364 9024
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3844 8928 3985 8956
rect 3844 8916 3850 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4264 8820 4292 8919
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 7374 8916 7380 8968
rect 7432 8916 7438 8968
rect 7650 8965 7656 8968
rect 7644 8956 7656 8965
rect 7611 8928 7656 8956
rect 7644 8919 7656 8928
rect 7650 8916 7656 8919
rect 7708 8916 7714 8968
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 8588 8888 8616 8996
rect 9766 8916 9772 8968
rect 9824 8916 9830 8968
rect 10336 8965 10364 8996
rect 10873 8993 10885 9027
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 9024 11023 9027
rect 11146 9024 11152 9036
rect 11011 8996 11152 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10980 8956 11008 8987
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 9024 16635 9027
rect 16684 9024 16712 9120
rect 16623 8996 16712 9024
rect 16761 9027 16819 9033
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 16761 8993 16773 9027
rect 16807 8993 16819 9027
rect 16761 8987 16819 8993
rect 16776 8956 16804 8987
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16908 8996 16957 9024
rect 16908 8984 16914 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 18156 9024 18184 9120
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 18156 8996 18613 9024
rect 16945 8987 17003 8993
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 9024 19579 9027
rect 19610 9024 19616 9036
rect 19567 8996 19616 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 19610 8984 19616 8996
rect 19668 9024 19674 9036
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 19668 8996 20177 9024
rect 19668 8984 19674 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 21266 8984 21272 9036
rect 21324 8984 21330 9036
rect 23860 9033 23888 9120
rect 25056 9033 25084 9120
rect 26421 9095 26479 9101
rect 25608 9064 25912 9092
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 8993 23903 9027
rect 23845 8987 23903 8993
rect 25041 9027 25099 9033
rect 25041 8993 25053 9027
rect 25087 8993 25099 9027
rect 25041 8987 25099 8993
rect 10367 8928 11008 8956
rect 16040 8928 16804 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 16040 8900 16068 8928
rect 6880 8860 8616 8888
rect 9125 8891 9183 8897
rect 6880 8848 6886 8860
rect 9125 8857 9137 8891
rect 9171 8857 9183 8891
rect 9125 8851 9183 8857
rect 4614 8820 4620 8832
rect 4264 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8820 4678 8832
rect 6454 8820 6460 8832
rect 4672 8792 6460 8820
rect 4672 8780 4678 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 9140 8820 9168 8851
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9272 8860 10824 8888
rect 9272 8848 9278 8860
rect 9490 8820 9496 8832
rect 8076 8792 9496 8820
rect 8076 8780 8082 8792
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 10686 8820 10692 8832
rect 10192 8792 10692 8820
rect 10192 8780 10198 8792
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10796 8829 10824 8860
rect 11330 8848 11336 8900
rect 11388 8888 11394 8900
rect 11425 8891 11483 8897
rect 11425 8888 11437 8891
rect 11388 8860 11437 8888
rect 11388 8848 11394 8860
rect 11425 8857 11437 8860
rect 11471 8857 11483 8891
rect 11425 8851 11483 8857
rect 11606 8848 11612 8900
rect 11664 8888 11670 8900
rect 11885 8891 11943 8897
rect 11885 8888 11897 8891
rect 11664 8860 11897 8888
rect 11664 8848 11670 8860
rect 11885 8857 11897 8860
rect 11931 8888 11943 8891
rect 15749 8891 15807 8897
rect 15749 8888 15761 8891
rect 11931 8860 15761 8888
rect 11931 8857 11943 8860
rect 11885 8851 11943 8857
rect 15749 8857 15761 8860
rect 15795 8888 15807 8891
rect 16022 8888 16028 8900
rect 15795 8860 16028 8888
rect 15795 8857 15807 8860
rect 15749 8851 15807 8857
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 16776 8888 16804 8928
rect 20073 8959 20131 8965
rect 20073 8925 20085 8959
rect 20119 8956 20131 8959
rect 21284 8956 21312 8984
rect 20119 8928 21312 8956
rect 22833 8959 22891 8965
rect 20119 8925 20131 8928
rect 20073 8919 20131 8925
rect 22833 8925 22845 8959
rect 22879 8956 22891 8959
rect 23658 8956 23664 8968
rect 22879 8928 23664 8956
rect 22879 8925 22891 8928
rect 22833 8919 22891 8925
rect 23658 8916 23664 8928
rect 23716 8956 23722 8968
rect 24394 8956 24400 8968
rect 23716 8928 24400 8956
rect 23716 8916 23722 8928
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 24854 8916 24860 8968
rect 24912 8956 24918 8968
rect 25608 8965 25636 9064
rect 25777 9027 25835 9033
rect 25777 8993 25789 9027
rect 25823 8993 25835 9027
rect 25777 8987 25835 8993
rect 25593 8959 25651 8965
rect 25593 8956 25605 8959
rect 24912 8928 25605 8956
rect 24912 8916 24918 8928
rect 25593 8925 25605 8928
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 19061 8891 19119 8897
rect 16776 8860 18920 8888
rect 10781 8823 10839 8829
rect 10781 8789 10793 8823
rect 10827 8820 10839 8823
rect 11790 8820 11796 8832
rect 10827 8792 11796 8820
rect 10827 8789 10839 8792
rect 10781 8783 10839 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 12342 8780 12348 8832
rect 12400 8780 12406 8832
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 16264 8792 17049 8820
rect 16264 8780 16270 8792
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 17402 8780 17408 8832
rect 17460 8780 17466 8832
rect 17957 8823 18015 8829
rect 17957 8789 17969 8823
rect 18003 8820 18015 8823
rect 18782 8820 18788 8832
rect 18003 8792 18788 8820
rect 18003 8789 18015 8792
rect 17957 8783 18015 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 18892 8820 18920 8860
rect 19061 8857 19073 8891
rect 19107 8888 19119 8891
rect 19794 8888 19800 8900
rect 19107 8860 19800 8888
rect 19107 8857 19119 8860
rect 19061 8851 19119 8857
rect 19794 8848 19800 8860
rect 19852 8888 19858 8900
rect 20346 8888 20352 8900
rect 19852 8860 20352 8888
rect 19852 8848 19858 8860
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 25792 8888 25820 8987
rect 25884 8956 25912 9064
rect 26421 9061 26433 9095
rect 26467 9061 26479 9095
rect 26421 9055 26479 9061
rect 26436 9024 26464 9055
rect 30190 9052 30196 9104
rect 30248 9092 30254 9104
rect 31772 9092 31800 9120
rect 30248 9064 31800 9092
rect 30248 9052 30254 9064
rect 27065 9027 27123 9033
rect 27065 9024 27077 9027
rect 26436 8996 27077 9024
rect 27065 8993 27077 8996
rect 27111 8993 27123 9027
rect 27065 8987 27123 8993
rect 28169 9027 28227 9033
rect 28169 8993 28181 9027
rect 28215 9024 28227 9027
rect 28902 9024 28908 9036
rect 28215 8996 28908 9024
rect 28215 8993 28227 8996
rect 28169 8987 28227 8993
rect 28902 8984 28908 8996
rect 28960 9024 28966 9036
rect 29181 9027 29239 9033
rect 29181 9024 29193 9027
rect 28960 8996 29193 9024
rect 28960 8984 28966 8996
rect 29181 8993 29193 8996
rect 29227 8993 29239 9027
rect 30653 9027 30711 9033
rect 30653 9024 30665 9027
rect 29181 8987 29239 8993
rect 30208 8996 30665 9024
rect 26053 8959 26111 8965
rect 26053 8956 26065 8959
rect 25884 8928 26065 8956
rect 26053 8925 26065 8928
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 26142 8916 26148 8968
rect 26200 8956 26206 8968
rect 28445 8959 28503 8965
rect 28445 8956 28457 8959
rect 26200 8928 28457 8956
rect 26200 8916 26206 8928
rect 28445 8925 28457 8928
rect 28491 8956 28503 8959
rect 30208 8956 30236 8996
rect 30653 8993 30665 8996
rect 30699 8993 30711 9027
rect 30653 8987 30711 8993
rect 33594 8984 33600 9036
rect 33652 9024 33658 9036
rect 33689 9027 33747 9033
rect 33689 9024 33701 9027
rect 33652 8996 33701 9024
rect 33652 8984 33658 8996
rect 33689 8993 33701 8996
rect 33735 8993 33747 9027
rect 33796 9024 33824 9120
rect 36464 9092 36492 9123
rect 36538 9120 36544 9132
rect 36596 9120 36602 9172
rect 37550 9120 37556 9172
rect 37608 9120 37614 9172
rect 37642 9120 37648 9172
rect 37700 9120 37706 9172
rect 37918 9120 37924 9172
rect 37976 9120 37982 9172
rect 38010 9120 38016 9172
rect 38068 9160 38074 9172
rect 38933 9163 38991 9169
rect 38933 9160 38945 9163
rect 38068 9132 38945 9160
rect 38068 9120 38074 9132
rect 38933 9129 38945 9132
rect 38979 9129 38991 9163
rect 38933 9123 38991 9129
rect 39206 9120 39212 9172
rect 39264 9160 39270 9172
rect 39301 9163 39359 9169
rect 39301 9160 39313 9163
rect 39264 9132 39313 9160
rect 39264 9120 39270 9132
rect 39301 9129 39313 9132
rect 39347 9160 39359 9163
rect 41966 9160 41972 9172
rect 39347 9132 41972 9160
rect 39347 9129 39359 9132
rect 39301 9123 39359 9129
rect 41966 9120 41972 9132
rect 42024 9120 42030 9172
rect 42245 9163 42303 9169
rect 42245 9129 42257 9163
rect 42291 9160 42303 9163
rect 42426 9160 42432 9172
rect 42291 9132 42432 9160
rect 42291 9129 42303 9132
rect 42245 9123 42303 9129
rect 42426 9120 42432 9132
rect 42484 9120 42490 9172
rect 43990 9120 43996 9172
rect 44048 9120 44054 9172
rect 45830 9120 45836 9172
rect 45888 9160 45894 9172
rect 46474 9160 46480 9172
rect 45888 9132 46480 9160
rect 45888 9120 45894 9132
rect 46474 9120 46480 9132
rect 46532 9120 46538 9172
rect 49142 9120 49148 9172
rect 49200 9160 49206 9172
rect 49329 9163 49387 9169
rect 49329 9160 49341 9163
rect 49200 9132 49341 9160
rect 49200 9120 49206 9132
rect 49329 9129 49341 9132
rect 49375 9129 49387 9163
rect 49329 9123 49387 9129
rect 49694 9120 49700 9172
rect 49752 9120 49758 9172
rect 50338 9120 50344 9172
rect 50396 9120 50402 9172
rect 52181 9163 52239 9169
rect 52181 9129 52193 9163
rect 52227 9160 52239 9163
rect 52546 9160 52552 9172
rect 52227 9132 52552 9160
rect 52227 9129 52239 9132
rect 52181 9123 52239 9129
rect 52546 9120 52552 9132
rect 52604 9120 52610 9172
rect 52641 9163 52699 9169
rect 52641 9129 52653 9163
rect 52687 9160 52699 9163
rect 52730 9160 52736 9172
rect 52687 9132 52736 9160
rect 52687 9129 52699 9132
rect 52641 9123 52699 9129
rect 52730 9120 52736 9132
rect 52788 9160 52794 9172
rect 53653 9163 53711 9169
rect 53653 9160 53665 9163
rect 52788 9132 53665 9160
rect 52788 9120 52794 9132
rect 53653 9129 53665 9132
rect 53699 9160 53711 9163
rect 53742 9160 53748 9172
rect 53699 9132 53748 9160
rect 53699 9129 53711 9132
rect 53653 9123 53711 9129
rect 53742 9120 53748 9132
rect 53800 9160 53806 9172
rect 55122 9160 55128 9172
rect 53800 9132 55128 9160
rect 53800 9120 53806 9132
rect 55122 9120 55128 9132
rect 55180 9120 55186 9172
rect 55306 9120 55312 9172
rect 55364 9120 55370 9172
rect 56229 9163 56287 9169
rect 56229 9129 56241 9163
rect 56275 9160 56287 9163
rect 56594 9160 56600 9172
rect 56275 9132 56600 9160
rect 56275 9129 56287 9132
rect 56229 9123 56287 9129
rect 56594 9120 56600 9132
rect 56652 9120 56658 9172
rect 56870 9120 56876 9172
rect 56928 9120 56934 9172
rect 57606 9120 57612 9172
rect 57664 9120 57670 9172
rect 35084 9064 36492 9092
rect 33873 9027 33931 9033
rect 33873 9024 33885 9027
rect 33796 8996 33885 9024
rect 33689 8987 33747 8993
rect 33873 8993 33885 8996
rect 33919 8993 33931 9027
rect 33873 8987 33931 8993
rect 28491 8928 30236 8956
rect 28491 8925 28503 8928
rect 28445 8919 28503 8925
rect 30282 8916 30288 8968
rect 30340 8956 30346 8968
rect 31481 8959 31539 8965
rect 31481 8956 31493 8959
rect 30340 8928 31493 8956
rect 30340 8916 30346 8928
rect 31481 8925 31493 8928
rect 31527 8925 31539 8959
rect 35084 8956 35112 9064
rect 35161 9027 35219 9033
rect 35161 8993 35173 9027
rect 35207 9024 35219 9027
rect 35207 8996 35848 9024
rect 35207 8993 35219 8996
rect 35161 8987 35219 8993
rect 35253 8959 35311 8965
rect 35253 8956 35265 8959
rect 35084 8928 35265 8956
rect 31481 8919 31539 8925
rect 35253 8925 35265 8928
rect 35299 8925 35311 8959
rect 35253 8919 35311 8925
rect 24872 8860 25820 8888
rect 24872 8832 24900 8860
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 29052 8860 30328 8888
rect 29052 8848 29058 8860
rect 19426 8820 19432 8832
rect 18892 8792 19432 8820
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19981 8823 20039 8829
rect 19981 8820 19993 8823
rect 19576 8792 19993 8820
rect 19576 8780 19582 8792
rect 19981 8789 19993 8792
rect 20027 8789 20039 8823
rect 19981 8783 20039 8789
rect 22462 8780 22468 8832
rect 22520 8820 22526 8832
rect 23109 8823 23167 8829
rect 23109 8820 23121 8823
rect 22520 8792 23121 8820
rect 22520 8780 22526 8792
rect 23109 8789 23121 8792
rect 23155 8820 23167 8823
rect 23198 8820 23204 8832
rect 23155 8792 23204 8820
rect 23155 8789 23167 8792
rect 23109 8783 23167 8789
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 24854 8780 24860 8832
rect 24912 8780 24918 8832
rect 25498 8780 25504 8832
rect 25556 8820 25562 8832
rect 25961 8823 26019 8829
rect 25961 8820 25973 8823
rect 25556 8792 25973 8820
rect 25556 8780 25562 8792
rect 25961 8789 25973 8792
rect 26007 8789 26019 8823
rect 25961 8783 26019 8789
rect 26694 8780 26700 8832
rect 26752 8820 26758 8832
rect 27433 8823 27491 8829
rect 27433 8820 27445 8823
rect 26752 8792 27445 8820
rect 26752 8780 26758 8792
rect 27433 8789 27445 8792
rect 27479 8789 27491 8823
rect 27433 8783 27491 8789
rect 28626 8780 28632 8832
rect 28684 8780 28690 8832
rect 29086 8780 29092 8832
rect 29144 8780 29150 8832
rect 30101 8823 30159 8829
rect 30101 8789 30113 8823
rect 30147 8820 30159 8823
rect 30190 8820 30196 8832
rect 30147 8792 30196 8820
rect 30147 8789 30159 8792
rect 30101 8783 30159 8789
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 30300 8820 30328 8860
rect 34514 8848 34520 8900
rect 34572 8888 34578 8900
rect 35158 8888 35164 8900
rect 34572 8860 35164 8888
rect 34572 8848 34578 8860
rect 35158 8848 35164 8860
rect 35216 8888 35222 8900
rect 35345 8891 35403 8897
rect 35345 8888 35357 8891
rect 35216 8860 35357 8888
rect 35216 8848 35222 8860
rect 35345 8857 35357 8860
rect 35391 8857 35403 8891
rect 35820 8888 35848 8996
rect 35894 8984 35900 9036
rect 35952 8984 35958 9036
rect 37660 9024 37688 9120
rect 37936 9092 37964 9120
rect 40405 9095 40463 9101
rect 40405 9092 40417 9095
rect 37936 9064 40417 9092
rect 40405 9061 40417 9064
rect 40451 9092 40463 9095
rect 40678 9092 40684 9104
rect 40451 9064 40684 9092
rect 40451 9061 40463 9064
rect 40405 9055 40463 9061
rect 40678 9052 40684 9064
rect 40736 9052 40742 9104
rect 42794 9052 42800 9104
rect 42852 9092 42858 9104
rect 46382 9092 46388 9104
rect 42852 9064 46388 9092
rect 42852 9052 42858 9064
rect 46382 9052 46388 9064
rect 46440 9052 46446 9104
rect 48317 9095 48375 9101
rect 48317 9061 48329 9095
rect 48363 9061 48375 9095
rect 48317 9055 48375 9061
rect 38105 9027 38163 9033
rect 38105 9024 38117 9027
rect 37660 8996 38117 9024
rect 38105 8993 38117 8996
rect 38151 8993 38163 9027
rect 38105 8987 38163 8993
rect 38381 9027 38439 9033
rect 38381 8993 38393 9027
rect 38427 9024 38439 9027
rect 38470 9024 38476 9036
rect 38427 8996 38476 9024
rect 38427 8993 38439 8996
rect 38381 8987 38439 8993
rect 38470 8984 38476 8996
rect 38528 8984 38534 9036
rect 38562 8984 38568 9036
rect 38620 9024 38626 9036
rect 40586 9024 40592 9036
rect 38620 8996 40592 9024
rect 38620 8984 38626 8996
rect 40586 8984 40592 8996
rect 40644 8984 40650 9036
rect 40696 9024 40724 9052
rect 44910 9024 44916 9036
rect 40696 8996 44916 9024
rect 44910 8984 44916 8996
rect 44968 9024 44974 9036
rect 47397 9027 47455 9033
rect 47397 9024 47409 9027
rect 44968 8996 47409 9024
rect 44968 8984 44974 8996
rect 47397 8993 47409 8996
rect 47443 9024 47455 9027
rect 47673 9027 47731 9033
rect 47673 9024 47685 9027
rect 47443 8996 47685 9024
rect 47443 8993 47455 8996
rect 47397 8987 47455 8993
rect 47673 8993 47685 8996
rect 47719 8993 47731 9027
rect 47673 8987 47731 8993
rect 37826 8916 37832 8968
rect 37884 8956 37890 8968
rect 39482 8956 39488 8968
rect 37884 8928 39488 8956
rect 37884 8916 37890 8928
rect 38396 8900 38424 8928
rect 39482 8916 39488 8928
rect 39540 8916 39546 8968
rect 43438 8916 43444 8968
rect 43496 8916 43502 8968
rect 45278 8916 45284 8968
rect 45336 8916 45342 8968
rect 36078 8888 36084 8900
rect 35820 8860 36084 8888
rect 35345 8851 35403 8857
rect 36078 8848 36084 8860
rect 36136 8848 36142 8900
rect 38378 8848 38384 8900
rect 38436 8848 38442 8900
rect 41966 8848 41972 8900
rect 42024 8848 42030 8900
rect 42150 8848 42156 8900
rect 42208 8848 42214 8900
rect 47688 8888 47716 8987
rect 47762 8984 47768 9036
rect 47820 9024 47826 9036
rect 47857 9027 47915 9033
rect 47857 9024 47869 9027
rect 47820 8996 47869 9024
rect 47820 8984 47826 8996
rect 47857 8993 47869 8996
rect 47903 8993 47915 9027
rect 48332 9024 48360 9055
rect 48685 9027 48743 9033
rect 48685 9024 48697 9027
rect 48332 8996 48697 9024
rect 47857 8987 47915 8993
rect 48685 8993 48697 8996
rect 48731 8993 48743 9027
rect 50356 9024 50384 9120
rect 53834 9052 53840 9104
rect 53892 9092 53898 9104
rect 54018 9092 54024 9104
rect 53892 9064 54024 9092
rect 53892 9052 53898 9064
rect 54018 9052 54024 9064
rect 54076 9052 54082 9104
rect 54662 9052 54668 9104
rect 54720 9052 54726 9104
rect 55324 9033 55352 9120
rect 55953 9095 56011 9101
rect 55953 9061 55965 9095
rect 55999 9092 56011 9095
rect 56410 9092 56416 9104
rect 55999 9064 56416 9092
rect 55999 9061 56011 9064
rect 55953 9055 56011 9061
rect 56410 9052 56416 9064
rect 56468 9052 56474 9104
rect 50801 9027 50859 9033
rect 50801 9024 50813 9027
rect 50356 8996 50813 9024
rect 48685 8987 48743 8993
rect 50801 8993 50813 8996
rect 50847 8993 50859 9027
rect 50801 8987 50859 8993
rect 55309 9027 55367 9033
rect 55309 8993 55321 9027
rect 55355 8993 55367 9027
rect 55309 8987 55367 8993
rect 56686 8984 56692 9036
rect 56744 9024 56750 9036
rect 56781 9027 56839 9033
rect 56781 9024 56793 9027
rect 56744 8996 56793 9024
rect 56744 8984 56750 8996
rect 56781 8993 56793 8996
rect 56827 8993 56839 9027
rect 56888 9024 56916 9120
rect 56965 9027 57023 9033
rect 56965 9024 56977 9027
rect 56888 8996 56977 9024
rect 56781 8987 56839 8993
rect 56965 8993 56977 8996
rect 57011 8993 57023 9027
rect 56965 8987 57023 8993
rect 47946 8916 47952 8968
rect 48004 8916 48010 8968
rect 51074 8965 51080 8968
rect 51068 8919 51080 8965
rect 51132 8956 51138 8968
rect 51132 8928 51168 8956
rect 51074 8916 51080 8919
rect 51132 8916 51138 8928
rect 58250 8916 58256 8968
rect 58308 8916 58314 8968
rect 52914 8888 52920 8900
rect 42812 8860 43300 8888
rect 47688 8860 52920 8888
rect 30466 8820 30472 8832
rect 30300 8792 30472 8820
rect 30466 8780 30472 8792
rect 30524 8780 30530 8832
rect 30561 8823 30619 8829
rect 30561 8789 30573 8823
rect 30607 8820 30619 8823
rect 30929 8823 30987 8829
rect 30929 8820 30941 8823
rect 30607 8792 30941 8820
rect 30607 8789 30619 8792
rect 30561 8783 30619 8789
rect 30929 8789 30941 8792
rect 30975 8789 30987 8823
rect 30929 8783 30987 8789
rect 31754 8780 31760 8832
rect 31812 8820 31818 8832
rect 31941 8823 31999 8829
rect 31941 8820 31953 8823
rect 31812 8792 31953 8820
rect 31812 8780 31818 8792
rect 31941 8789 31953 8792
rect 31987 8820 31999 8823
rect 32398 8820 32404 8832
rect 31987 8792 32404 8820
rect 31987 8789 31999 8792
rect 31941 8783 31999 8789
rect 32398 8780 32404 8792
rect 32456 8780 32462 8832
rect 35710 8780 35716 8832
rect 35768 8780 35774 8832
rect 41984 8820 42012 8848
rect 42812 8820 42840 8860
rect 41984 8792 42840 8820
rect 42886 8780 42892 8832
rect 42944 8780 42950 8832
rect 43272 8820 43300 8860
rect 52914 8848 52920 8860
rect 52972 8888 52978 8900
rect 56594 8888 56600 8900
rect 52972 8860 56600 8888
rect 52972 8848 52978 8860
rect 56594 8848 56600 8860
rect 56652 8848 56658 8900
rect 44637 8823 44695 8829
rect 44637 8820 44649 8823
rect 43272 8792 44649 8820
rect 44637 8789 44649 8792
rect 44683 8820 44695 8823
rect 45554 8820 45560 8832
rect 44683 8792 45560 8820
rect 44683 8789 44695 8792
rect 44637 8783 44695 8789
rect 45554 8780 45560 8792
rect 45612 8780 45618 8832
rect 57698 8780 57704 8832
rect 57756 8780 57762 8832
rect 1104 8730 59040 8752
rect 1104 8678 15394 8730
rect 15446 8678 15458 8730
rect 15510 8678 15522 8730
rect 15574 8678 15586 8730
rect 15638 8678 15650 8730
rect 15702 8678 29838 8730
rect 29890 8678 29902 8730
rect 29954 8678 29966 8730
rect 30018 8678 30030 8730
rect 30082 8678 30094 8730
rect 30146 8678 44282 8730
rect 44334 8678 44346 8730
rect 44398 8678 44410 8730
rect 44462 8678 44474 8730
rect 44526 8678 44538 8730
rect 44590 8678 58726 8730
rect 58778 8678 58790 8730
rect 58842 8678 58854 8730
rect 58906 8678 58918 8730
rect 58970 8678 58982 8730
rect 59034 8678 59040 8730
rect 1104 8656 59040 8678
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 7558 8576 7564 8628
rect 7616 8576 7622 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 9214 8616 9220 8628
rect 8067 8588 9220 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 11146 8616 11152 8628
rect 9539 8588 11152 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 18325 8619 18383 8625
rect 18325 8616 18337 8619
rect 18012 8588 18337 8616
rect 18012 8576 18018 8588
rect 18325 8585 18337 8588
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 18840 8588 20208 8616
rect 18840 8576 18846 8588
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 6362 8548 6368 8560
rect 6227 8520 6368 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 6362 8508 6368 8520
rect 6420 8548 6426 8560
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 6420 8520 6561 8548
rect 6420 8508 6426 8520
rect 6549 8517 6561 8520
rect 6595 8548 6607 8551
rect 6822 8548 6828 8560
rect 6595 8520 6828 8548
rect 6595 8517 6607 8520
rect 6549 8511 6607 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7929 8551 7987 8557
rect 7929 8517 7941 8551
rect 7975 8548 7987 8551
rect 8570 8548 8576 8560
rect 7975 8520 8576 8548
rect 7975 8517 7987 8520
rect 7929 8511 7987 8517
rect 8570 8508 8576 8520
rect 8628 8548 8634 8560
rect 8628 8520 9352 8548
rect 8628 8508 8634 8520
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7156 8452 7205 8480
rect 7156 8440 7162 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 8018 8480 8024 8492
rect 7193 8443 7251 8449
rect 7668 8452 8024 8480
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4540 8384 4997 8412
rect 4540 8356 4568 8384
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 4522 8304 4528 8356
rect 4580 8304 4586 8356
rect 7668 8344 7696 8452
rect 8018 8440 8024 8452
rect 8076 8480 8082 8492
rect 8481 8483 8539 8489
rect 8076 8452 8156 8480
rect 8076 8440 8082 8452
rect 7742 8372 7748 8424
rect 7800 8372 7806 8424
rect 8128 8421 8156 8452
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8662 8480 8668 8492
rect 8527 8452 8668 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8628 8384 8769 8412
rect 8628 8372 8634 8384
rect 8757 8381 8769 8384
rect 8803 8412 8815 8415
rect 8846 8412 8852 8424
rect 8803 8384 8852 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9324 8412 9352 8520
rect 11164 8520 11928 8548
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 11164 8489 11192 8520
rect 11900 8489 11928 8520
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16485 8551 16543 8557
rect 16485 8548 16497 8551
rect 16448 8520 16497 8548
rect 16448 8508 16454 8520
rect 16485 8517 16497 8520
rect 16531 8548 16543 8551
rect 18877 8551 18935 8557
rect 16531 8520 18552 8548
rect 16531 8517 16543 8520
rect 16485 8511 16543 8517
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 11931 8452 12357 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 17402 8440 17408 8492
rect 17460 8480 17466 8492
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17460 8452 17693 8480
rect 17460 8440 17466 8452
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 10275 8415 10333 8421
rect 10275 8412 10287 8415
rect 9324 8384 10287 8412
rect 10275 8381 10287 8384
rect 10321 8381 10333 8415
rect 10275 8375 10333 8381
rect 10410 8372 10416 8424
rect 10468 8372 10474 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10612 8384 10701 8412
rect 4632 8316 7696 8344
rect 7760 8344 7788 8372
rect 10612 8356 10640 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 11514 8412 11520 8424
rect 11379 8384 11520 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 11606 8372 11612 8424
rect 11664 8372 11670 8424
rect 12894 8372 12900 8424
rect 12952 8372 12958 8424
rect 17037 8415 17095 8421
rect 17037 8381 17049 8415
rect 17083 8412 17095 8415
rect 18524 8412 18552 8520
rect 18877 8517 18889 8551
rect 18923 8548 18935 8551
rect 19518 8548 19524 8560
rect 18923 8520 19524 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 19518 8508 19524 8520
rect 19576 8508 19582 8560
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 18831 8452 19901 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 19889 8449 19901 8452
rect 19935 8480 19947 8483
rect 20070 8480 20076 8492
rect 19935 8452 20076 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 17083 8384 18460 8412
rect 18524 8384 19073 8412
rect 17083 8381 17095 8384
rect 17037 8375 17095 8381
rect 7760 8316 9674 8344
rect 4632 8288 4660 8316
rect 4614 8236 4620 8288
rect 4672 8236 4678 8288
rect 4982 8236 4988 8288
rect 5040 8276 5046 8288
rect 5534 8276 5540 8288
rect 5040 8248 5540 8276
rect 5040 8236 5046 8248
rect 5534 8236 5540 8248
rect 5592 8276 5598 8288
rect 5813 8279 5871 8285
rect 5813 8276 5825 8279
rect 5592 8248 5825 8276
rect 5592 8236 5598 8248
rect 5813 8245 5825 8248
rect 5859 8276 5871 8279
rect 5902 8276 5908 8288
rect 5859 8248 5908 8276
rect 5859 8245 5871 8248
rect 5813 8239 5871 8245
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 9646 8276 9674 8316
rect 10594 8304 10600 8356
rect 10652 8304 10658 8356
rect 12253 8347 12311 8353
rect 12253 8313 12265 8347
rect 12299 8344 12311 8347
rect 12526 8344 12532 8356
rect 12299 8316 12532 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 17589 8347 17647 8353
rect 17589 8313 17601 8347
rect 17635 8344 17647 8347
rect 17954 8344 17960 8356
rect 17635 8316 17960 8344
rect 17635 8313 17647 8316
rect 17589 8307 17647 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18432 8353 18460 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 18417 8347 18475 8353
rect 18417 8313 18429 8347
rect 18463 8313 18475 8347
rect 19076 8344 19104 8375
rect 19242 8372 19248 8424
rect 19300 8372 19306 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19392 8384 19993 8412
rect 19392 8372 19398 8384
rect 19981 8381 19993 8384
rect 20027 8381 20039 8415
rect 20180 8412 20208 8588
rect 25222 8576 25228 8628
rect 25280 8576 25286 8628
rect 28442 8576 28448 8628
rect 28500 8576 28506 8628
rect 28626 8576 28632 8628
rect 28684 8576 28690 8628
rect 29086 8576 29092 8628
rect 29144 8616 29150 8628
rect 29917 8619 29975 8625
rect 29917 8616 29929 8619
rect 29144 8588 29929 8616
rect 29144 8576 29150 8588
rect 29917 8585 29929 8588
rect 29963 8616 29975 8619
rect 30374 8616 30380 8628
rect 29963 8588 30380 8616
rect 29963 8585 29975 8588
rect 29917 8579 29975 8585
rect 30374 8576 30380 8588
rect 30432 8576 30438 8628
rect 30742 8576 30748 8628
rect 30800 8576 30806 8628
rect 30834 8576 30840 8628
rect 30892 8576 30898 8628
rect 34790 8576 34796 8628
rect 34848 8616 34854 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 34848 8588 34897 8616
rect 34848 8576 34854 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 35710 8576 35716 8628
rect 35768 8576 35774 8628
rect 35897 8619 35955 8625
rect 35897 8585 35909 8619
rect 35943 8616 35955 8619
rect 36078 8616 36084 8628
rect 35943 8588 36084 8616
rect 35943 8585 35955 8588
rect 35897 8579 35955 8585
rect 36078 8576 36084 8588
rect 36136 8576 36142 8628
rect 42886 8576 42892 8628
rect 42944 8576 42950 8628
rect 48314 8576 48320 8628
rect 48372 8616 48378 8628
rect 48501 8619 48559 8625
rect 48501 8616 48513 8619
rect 48372 8588 48513 8616
rect 48372 8576 48378 8588
rect 48501 8585 48513 8588
rect 48547 8585 48559 8619
rect 48501 8579 48559 8585
rect 49970 8576 49976 8628
rect 50028 8616 50034 8628
rect 50157 8619 50215 8625
rect 50157 8616 50169 8619
rect 50028 8588 50169 8616
rect 50028 8576 50034 8588
rect 50157 8585 50169 8588
rect 50203 8585 50215 8619
rect 50157 8579 50215 8585
rect 50338 8576 50344 8628
rect 50396 8616 50402 8628
rect 51537 8619 51595 8625
rect 51537 8616 51549 8619
rect 50396 8588 51549 8616
rect 50396 8576 50402 8588
rect 51537 8585 51549 8588
rect 51583 8616 51595 8619
rect 52365 8619 52423 8625
rect 52365 8616 52377 8619
rect 51583 8588 52377 8616
rect 51583 8585 51595 8588
rect 51537 8579 51595 8585
rect 52365 8585 52377 8588
rect 52411 8616 52423 8619
rect 52730 8616 52736 8628
rect 52411 8588 52736 8616
rect 52411 8585 52423 8588
rect 52365 8579 52423 8585
rect 52730 8576 52736 8588
rect 52788 8576 52794 8628
rect 55766 8576 55772 8628
rect 55824 8616 55830 8628
rect 55861 8619 55919 8625
rect 55861 8616 55873 8619
rect 55824 8588 55873 8616
rect 55824 8576 55830 8588
rect 55861 8585 55873 8588
rect 55907 8585 55919 8619
rect 55861 8579 55919 8585
rect 20346 8508 20352 8560
rect 20404 8548 20410 8560
rect 25130 8548 25136 8560
rect 20404 8520 25136 8548
rect 20404 8508 20410 8520
rect 25130 8508 25136 8520
rect 25188 8508 25194 8560
rect 26544 8551 26602 8557
rect 26544 8517 26556 8551
rect 26590 8548 26602 8551
rect 26973 8551 27031 8557
rect 26973 8548 26985 8551
rect 26590 8520 26985 8548
rect 26590 8517 26602 8520
rect 26544 8511 26602 8517
rect 26973 8517 26985 8520
rect 27019 8517 27031 8551
rect 26973 8511 27031 8517
rect 26694 8440 26700 8492
rect 26752 8480 26758 8492
rect 26789 8483 26847 8489
rect 26789 8480 26801 8483
rect 26752 8452 26801 8480
rect 26752 8440 26758 8452
rect 26789 8449 26801 8452
rect 26835 8480 26847 8483
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 26835 8452 27905 8480
rect 26835 8449 26847 8452
rect 26789 8443 26847 8449
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 28644 8480 28672 8576
rect 28997 8483 29055 8489
rect 28997 8480 29009 8483
rect 28644 8452 29009 8480
rect 27893 8443 27951 8449
rect 28997 8449 29009 8452
rect 29043 8449 29055 8483
rect 28997 8443 29055 8449
rect 29362 8440 29368 8492
rect 29420 8440 29426 8492
rect 30190 8440 30196 8492
rect 30248 8440 30254 8492
rect 35529 8483 35587 8489
rect 35529 8449 35541 8483
rect 35575 8480 35587 8483
rect 35728 8480 35756 8576
rect 42788 8551 42846 8557
rect 42788 8517 42800 8551
rect 42834 8548 42846 8551
rect 42904 8548 42932 8576
rect 42834 8520 42932 8548
rect 42834 8517 42846 8520
rect 42788 8511 42846 8517
rect 45278 8508 45284 8560
rect 45336 8548 45342 8560
rect 50065 8551 50123 8557
rect 50065 8548 50077 8551
rect 45336 8520 50077 8548
rect 45336 8508 45342 8520
rect 50065 8517 50077 8520
rect 50111 8517 50123 8551
rect 50065 8511 50123 8517
rect 50525 8551 50583 8557
rect 50525 8517 50537 8551
rect 50571 8548 50583 8551
rect 51350 8548 51356 8560
rect 50571 8520 51356 8548
rect 50571 8517 50583 8520
rect 50525 8511 50583 8517
rect 38657 8483 38715 8489
rect 38657 8480 38669 8483
rect 35575 8452 35756 8480
rect 36556 8452 38669 8480
rect 35575 8449 35587 8452
rect 35529 8443 35587 8449
rect 23750 8412 23756 8424
rect 20180 8384 23756 8412
rect 19981 8375 20039 8381
rect 23750 8372 23756 8384
rect 23808 8372 23814 8424
rect 24026 8372 24032 8424
rect 24084 8372 24090 8424
rect 26878 8372 26884 8424
rect 26936 8412 26942 8424
rect 27525 8415 27583 8421
rect 27525 8412 27537 8415
rect 26936 8384 27537 8412
rect 26936 8372 26942 8384
rect 27525 8381 27537 8384
rect 27571 8381 27583 8415
rect 27525 8375 27583 8381
rect 31386 8372 31392 8424
rect 31444 8372 31450 8424
rect 22370 8344 22376 8356
rect 19076 8316 22376 8344
rect 18417 8307 18475 8313
rect 22370 8304 22376 8316
rect 22428 8304 22434 8356
rect 25332 8316 25544 8344
rect 10318 8276 10324 8288
rect 9646 8248 10324 8276
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 14093 8279 14151 8285
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 15102 8276 15108 8288
rect 14139 8248 15108 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 20162 8236 20168 8288
rect 20220 8276 20226 8288
rect 20625 8279 20683 8285
rect 20625 8276 20637 8279
rect 20220 8248 20637 8276
rect 20220 8236 20226 8248
rect 20625 8245 20637 8248
rect 20671 8245 20683 8279
rect 20625 8239 20683 8245
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23566 8276 23572 8288
rect 23523 8248 23572 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23566 8236 23572 8248
rect 23624 8236 23630 8288
rect 24670 8236 24676 8288
rect 24728 8276 24734 8288
rect 25332 8276 25360 8316
rect 24728 8248 25360 8276
rect 24728 8236 24734 8248
rect 25406 8236 25412 8288
rect 25464 8236 25470 8288
rect 25516 8276 25544 8316
rect 28902 8304 28908 8356
rect 28960 8344 28966 8356
rect 31846 8344 31852 8356
rect 28960 8316 31852 8344
rect 28960 8304 28966 8316
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 35986 8304 35992 8356
rect 36044 8344 36050 8356
rect 36081 8347 36139 8353
rect 36081 8344 36093 8347
rect 36044 8316 36093 8344
rect 36044 8304 36050 8316
rect 36081 8313 36093 8316
rect 36127 8313 36139 8347
rect 36081 8307 36139 8313
rect 28920 8276 28948 8304
rect 25516 8248 28948 8276
rect 32030 8236 32036 8288
rect 32088 8276 32094 8288
rect 34422 8276 34428 8288
rect 32088 8248 34428 8276
rect 32088 8236 32094 8248
rect 34422 8236 34428 8248
rect 34480 8276 34486 8288
rect 34517 8279 34575 8285
rect 34517 8276 34529 8279
rect 34480 8248 34529 8276
rect 34480 8236 34486 8248
rect 34517 8245 34529 8248
rect 34563 8276 34575 8279
rect 35342 8276 35348 8288
rect 34563 8248 35348 8276
rect 34563 8245 34575 8248
rect 34517 8239 34575 8245
rect 35342 8236 35348 8248
rect 35400 8276 35406 8288
rect 36556 8276 36584 8452
rect 38657 8449 38669 8452
rect 38703 8480 38715 8483
rect 39390 8480 39396 8492
rect 38703 8452 39396 8480
rect 38703 8449 38715 8452
rect 38657 8443 38715 8449
rect 39390 8440 39396 8452
rect 39448 8440 39454 8492
rect 42518 8440 42524 8492
rect 42576 8440 42582 8492
rect 42610 8440 42616 8492
rect 42668 8480 42674 8492
rect 45296 8480 45324 8508
rect 42668 8452 45324 8480
rect 42668 8440 42674 8452
rect 36630 8372 36636 8424
rect 36688 8372 36694 8424
rect 41414 8372 41420 8424
rect 41472 8372 41478 8424
rect 41598 8372 41604 8424
rect 41656 8372 41662 8424
rect 44545 8415 44603 8421
rect 44545 8381 44557 8415
rect 44591 8381 44603 8415
rect 44545 8375 44603 8381
rect 43901 8347 43959 8353
rect 43901 8313 43913 8347
rect 43947 8344 43959 8347
rect 44174 8344 44180 8356
rect 43947 8316 44180 8344
rect 43947 8313 43959 8316
rect 43901 8307 43959 8313
rect 44174 8304 44180 8316
rect 44232 8344 44238 8356
rect 44560 8344 44588 8375
rect 47578 8372 47584 8424
rect 47636 8372 47642 8424
rect 50080 8412 50108 8511
rect 51350 8508 51356 8520
rect 51408 8508 51414 8560
rect 57054 8508 57060 8560
rect 57112 8548 57118 8560
rect 57333 8551 57391 8557
rect 57333 8548 57345 8551
rect 57112 8520 57345 8548
rect 57112 8508 57118 8520
rect 57333 8517 57345 8520
rect 57379 8517 57391 8551
rect 57333 8511 57391 8517
rect 50617 8483 50675 8489
rect 50617 8449 50629 8483
rect 50663 8480 50675 8483
rect 51994 8480 52000 8492
rect 50663 8452 52000 8480
rect 50663 8449 50675 8452
rect 50617 8443 50675 8449
rect 51994 8440 52000 8452
rect 52052 8440 52058 8492
rect 52178 8440 52184 8492
rect 52236 8480 52242 8492
rect 53469 8483 53527 8489
rect 53469 8480 53481 8483
rect 52236 8452 53481 8480
rect 52236 8440 52242 8452
rect 53469 8449 53481 8452
rect 53515 8480 53527 8483
rect 55953 8483 56011 8489
rect 53515 8452 54524 8480
rect 53515 8449 53527 8452
rect 53469 8443 53527 8449
rect 50709 8415 50767 8421
rect 50709 8412 50721 8415
rect 50080 8384 50721 8412
rect 50709 8381 50721 8384
rect 50755 8412 50767 8415
rect 54018 8412 54024 8424
rect 50755 8384 54024 8412
rect 50755 8381 50767 8384
rect 50709 8375 50767 8381
rect 54018 8372 54024 8384
rect 54076 8372 54082 8424
rect 44232 8316 44588 8344
rect 51997 8347 52055 8353
rect 44232 8304 44238 8316
rect 51997 8313 52009 8347
rect 52043 8344 52055 8347
rect 52086 8344 52092 8356
rect 52043 8316 52092 8344
rect 52043 8313 52055 8316
rect 51997 8307 52055 8313
rect 52086 8304 52092 8316
rect 52144 8304 52150 8356
rect 52914 8304 52920 8356
rect 52972 8304 52978 8356
rect 53837 8347 53895 8353
rect 53837 8313 53849 8347
rect 53883 8344 53895 8347
rect 54496 8344 54524 8452
rect 55953 8449 55965 8483
rect 55999 8480 56011 8483
rect 56686 8480 56692 8492
rect 55999 8452 56692 8480
rect 55999 8449 56011 8452
rect 55953 8443 56011 8449
rect 56686 8440 56692 8452
rect 56744 8440 56750 8492
rect 57238 8440 57244 8492
rect 57296 8480 57302 8492
rect 57885 8483 57943 8489
rect 57885 8480 57897 8483
rect 57296 8452 57897 8480
rect 57296 8440 57302 8452
rect 57885 8449 57897 8452
rect 57931 8449 57943 8483
rect 57885 8443 57943 8449
rect 54570 8372 54576 8424
rect 54628 8372 54634 8424
rect 54757 8415 54815 8421
rect 54757 8381 54769 8415
rect 54803 8412 54815 8415
rect 55766 8412 55772 8424
rect 54803 8384 55772 8412
rect 54803 8381 54815 8384
rect 54757 8375 54815 8381
rect 55766 8372 55772 8384
rect 55824 8372 55830 8424
rect 56229 8415 56287 8421
rect 56229 8381 56241 8415
rect 56275 8381 56287 8415
rect 56229 8375 56287 8381
rect 55309 8347 55367 8353
rect 53883 8316 54055 8344
rect 54496 8316 55260 8344
rect 53883 8313 53895 8316
rect 53837 8307 53895 8313
rect 35400 8248 36584 8276
rect 35400 8236 35406 8248
rect 37458 8236 37464 8288
rect 37516 8276 37522 8288
rect 38378 8276 38384 8288
rect 37516 8248 38384 8276
rect 37516 8236 37522 8248
rect 38378 8236 38384 8248
rect 38436 8236 38442 8288
rect 40770 8236 40776 8288
rect 40828 8236 40834 8288
rect 41230 8236 41236 8288
rect 41288 8276 41294 8288
rect 42153 8279 42211 8285
rect 42153 8276 42165 8279
rect 41288 8248 42165 8276
rect 41288 8236 41294 8248
rect 42153 8245 42165 8248
rect 42199 8276 42211 8279
rect 43162 8276 43168 8288
rect 42199 8248 43168 8276
rect 42199 8245 42211 8248
rect 42153 8239 42211 8245
rect 43162 8236 43168 8248
rect 43220 8236 43226 8288
rect 43990 8236 43996 8288
rect 44048 8236 44054 8288
rect 48222 8236 48228 8288
rect 48280 8236 48286 8288
rect 51166 8236 51172 8288
rect 51224 8276 51230 8288
rect 53852 8276 53880 8307
rect 51224 8248 53880 8276
rect 51224 8236 51230 8248
rect 53926 8236 53932 8288
rect 53984 8236 53990 8288
rect 54027 8276 54055 8316
rect 54386 8276 54392 8288
rect 54027 8248 54392 8276
rect 54386 8236 54392 8248
rect 54444 8276 54450 8288
rect 54754 8276 54760 8288
rect 54444 8248 54760 8276
rect 54444 8236 54450 8248
rect 54754 8236 54760 8248
rect 54812 8236 54818 8288
rect 55232 8276 55260 8316
rect 55309 8313 55321 8347
rect 55355 8344 55367 8347
rect 55674 8344 55680 8356
rect 55355 8316 55680 8344
rect 55355 8313 55367 8316
rect 55309 8307 55367 8313
rect 55674 8304 55680 8316
rect 55732 8304 55738 8356
rect 56244 8344 56272 8375
rect 56594 8372 56600 8424
rect 56652 8412 56658 8424
rect 56652 8384 57284 8412
rect 56652 8372 56658 8384
rect 56873 8347 56931 8353
rect 56873 8344 56885 8347
rect 56244 8316 56885 8344
rect 56873 8313 56885 8316
rect 56919 8313 56931 8347
rect 57256 8344 57284 8384
rect 57422 8372 57428 8424
rect 57480 8372 57486 8424
rect 58434 8372 58440 8424
rect 58492 8372 58498 8424
rect 57440 8344 57468 8372
rect 57256 8316 57468 8344
rect 56873 8307 56931 8313
rect 55585 8279 55643 8285
rect 55585 8276 55597 8279
rect 55232 8248 55597 8276
rect 55585 8245 55597 8248
rect 55631 8276 55643 8279
rect 56226 8276 56232 8288
rect 55631 8248 56232 8276
rect 55631 8245 55643 8248
rect 55585 8239 55643 8245
rect 56226 8236 56232 8248
rect 56284 8236 56290 8288
rect 56778 8236 56784 8288
rect 56836 8236 56842 8288
rect 1104 8186 58880 8208
rect 1104 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 22616 8186
rect 22668 8134 22680 8186
rect 22732 8134 22744 8186
rect 22796 8134 22808 8186
rect 22860 8134 22872 8186
rect 22924 8134 37060 8186
rect 37112 8134 37124 8186
rect 37176 8134 37188 8186
rect 37240 8134 37252 8186
rect 37304 8134 37316 8186
rect 37368 8134 51504 8186
rect 51556 8134 51568 8186
rect 51620 8134 51632 8186
rect 51684 8134 51696 8186
rect 51748 8134 51760 8186
rect 51812 8134 58880 8186
rect 1104 8112 58880 8134
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 8018 8032 8024 8084
rect 8076 8032 8082 8084
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 11606 8072 11612 8084
rect 10376 8044 11612 8072
rect 10376 8032 10382 8044
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 12894 8072 12900 8084
rect 11931 8044 12900 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 14090 8072 14096 8084
rect 13955 8044 14096 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 3620 7976 3801 8004
rect 3620 7945 3648 7976
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 5721 8007 5779 8013
rect 5721 7973 5733 8007
rect 5767 7973 5779 8007
rect 7098 8004 7104 8016
rect 5721 7967 5779 7973
rect 6840 7976 7104 8004
rect 3605 7939 3663 7945
rect 3605 7905 3617 7939
rect 3651 7905 3663 7939
rect 3605 7899 3663 7905
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4479 7908 4813 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5736 7936 5764 7967
rect 5675 7908 5764 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 4816 7868 4844 7899
rect 6362 7896 6368 7948
rect 6420 7896 6426 7948
rect 6840 7945 6868 7976
rect 7098 7964 7104 7976
rect 7156 8004 7162 8016
rect 7760 8004 7788 8032
rect 13924 8004 13952 8035
rect 14090 8032 14096 8044
rect 14148 8072 14154 8084
rect 14826 8072 14832 8084
rect 14148 8044 14832 8072
rect 14148 8032 14154 8044
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19242 8072 19248 8084
rect 19107 8044 19248 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 19886 8032 19892 8084
rect 19944 8072 19950 8084
rect 20806 8072 20812 8084
rect 19944 8044 20812 8072
rect 19944 8032 19950 8044
rect 20806 8032 20812 8044
rect 20864 8032 20870 8084
rect 24118 8072 24124 8084
rect 22480 8044 24124 8072
rect 22480 8016 22508 8044
rect 24118 8032 24124 8044
rect 24176 8032 24182 8084
rect 29733 8075 29791 8081
rect 29733 8041 29745 8075
rect 29779 8072 29791 8075
rect 31386 8072 31392 8084
rect 29779 8044 31392 8072
rect 29779 8041 29791 8044
rect 29733 8035 29791 8041
rect 31386 8032 31392 8044
rect 31444 8032 31450 8084
rect 33597 8075 33655 8081
rect 33597 8041 33609 8075
rect 33643 8072 33655 8075
rect 34146 8072 34152 8084
rect 33643 8044 34152 8072
rect 33643 8041 33655 8044
rect 33597 8035 33655 8041
rect 34146 8032 34152 8044
rect 34204 8072 34210 8084
rect 34882 8072 34888 8084
rect 34204 8044 34888 8072
rect 34204 8032 34210 8044
rect 34882 8032 34888 8044
rect 34940 8032 34946 8084
rect 35158 8032 35164 8084
rect 35216 8072 35222 8084
rect 35253 8075 35311 8081
rect 35253 8072 35265 8075
rect 35216 8044 35265 8072
rect 35216 8032 35222 8044
rect 35253 8041 35265 8044
rect 35299 8041 35311 8075
rect 35253 8035 35311 8041
rect 40865 8075 40923 8081
rect 40865 8041 40877 8075
rect 40911 8072 40923 8075
rect 41414 8072 41420 8084
rect 40911 8044 41420 8072
rect 40911 8041 40923 8044
rect 40865 8035 40923 8041
rect 41414 8032 41420 8044
rect 41472 8032 41478 8084
rect 42794 8032 42800 8084
rect 42852 8032 42858 8084
rect 42981 8075 43039 8081
rect 42981 8041 42993 8075
rect 43027 8072 43039 8075
rect 43438 8072 43444 8084
rect 43027 8044 43444 8072
rect 43027 8041 43039 8044
rect 42981 8035 43039 8041
rect 43438 8032 43444 8044
rect 43496 8032 43502 8084
rect 45281 8075 45339 8081
rect 45281 8041 45293 8075
rect 45327 8072 45339 8075
rect 45830 8072 45836 8084
rect 45327 8044 45836 8072
rect 45327 8041 45339 8044
rect 45281 8035 45339 8041
rect 7156 7976 7788 8004
rect 12406 7976 13952 8004
rect 7156 7964 7162 7976
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 4816 7840 6868 7868
rect 6089 7803 6147 7809
rect 6089 7800 6101 7803
rect 4172 7772 6101 7800
rect 4172 7744 4200 7772
rect 6089 7769 6101 7772
rect 6135 7769 6147 7803
rect 6840 7800 6868 7840
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7064 7840 7389 7868
rect 7064 7828 7070 7840
rect 7377 7837 7389 7840
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8352 7840 8953 7868
rect 8352 7828 8358 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 9674 7868 9680 7880
rect 8987 7840 9680 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9674 7828 9680 7840
rect 9732 7868 9738 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 9732 7840 10517 7868
rect 9732 7828 9738 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 12406 7868 12434 7976
rect 17310 7964 17316 8016
rect 17368 7964 17374 8016
rect 20346 7964 20352 8016
rect 20404 8004 20410 8016
rect 20441 8007 20499 8013
rect 20441 8004 20453 8007
rect 20404 7976 20453 8004
rect 20404 7964 20410 7976
rect 20441 7973 20453 7976
rect 20487 7973 20499 8007
rect 20441 7967 20499 7973
rect 22462 7964 22468 8016
rect 22520 7964 22526 8016
rect 23109 8007 23167 8013
rect 23109 7973 23121 8007
rect 23155 8004 23167 8007
rect 23474 8004 23480 8016
rect 23155 7976 23480 8004
rect 23155 7973 23167 7976
rect 23109 7967 23167 7973
rect 23474 7964 23480 7976
rect 23532 7964 23538 8016
rect 24670 8004 24676 8016
rect 23768 7976 24676 8004
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7936 19303 7939
rect 19702 7936 19708 7948
rect 19291 7908 19708 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 20070 7945 20076 7948
rect 20048 7939 20076 7945
rect 20048 7905 20060 7939
rect 20048 7899 20076 7905
rect 20070 7896 20076 7899
rect 20128 7896 20134 7948
rect 20162 7896 20168 7948
rect 20220 7896 20226 7948
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7936 21143 7939
rect 21266 7936 21272 7948
rect 21131 7908 21272 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 21266 7896 21272 7908
rect 21324 7896 21330 7948
rect 22370 7896 22376 7948
rect 22428 7936 22434 7948
rect 22649 7939 22707 7945
rect 22649 7936 22661 7939
rect 22428 7908 22661 7936
rect 22428 7896 22434 7908
rect 22649 7905 22661 7908
rect 22695 7936 22707 7939
rect 23658 7936 23664 7948
rect 22695 7908 23664 7936
rect 22695 7905 22707 7908
rect 22649 7899 22707 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 11112 7840 12434 7868
rect 11112 7828 11118 7840
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 14734 7828 14740 7880
rect 14792 7828 14798 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17586 7868 17592 7880
rect 17267 7840 17592 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 17586 7828 17592 7840
rect 17644 7868 17650 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17644 7840 17693 7868
rect 17644 7828 17650 7840
rect 17681 7837 17693 7840
rect 17727 7868 17739 7871
rect 17727 7840 19334 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 8570 7800 8576 7812
rect 6840 7772 8576 7800
rect 6089 7763 6147 7769
rect 8570 7760 8576 7772
rect 8628 7760 8634 7812
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7800 8815 7803
rect 9186 7803 9244 7809
rect 9186 7800 9198 7803
rect 8803 7772 9198 7800
rect 8803 7769 8815 7772
rect 8757 7763 8815 7769
rect 9186 7769 9198 7772
rect 9232 7769 9244 7803
rect 9186 7763 9244 7769
rect 10226 7760 10232 7812
rect 10284 7800 10290 7812
rect 10772 7803 10830 7809
rect 10284 7772 10640 7800
rect 10284 7760 10290 7772
rect 10612 7744 10640 7772
rect 10772 7769 10784 7803
rect 10818 7800 10830 7803
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 10818 7772 11989 7800
rect 10818 7769 10830 7772
rect 10772 7763 10830 7769
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 12986 7800 12992 7812
rect 11977 7763 12035 7769
rect 12084 7772 12992 7800
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 4154 7692 4160 7744
rect 4212 7692 4218 7744
rect 4246 7692 4252 7744
rect 4304 7692 4310 7744
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5074 7732 5080 7744
rect 5031 7704 5080 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 6178 7692 6184 7744
rect 6236 7692 6242 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 12084 7732 12112 7772
rect 12986 7760 12992 7772
rect 13044 7760 13050 7812
rect 17494 7760 17500 7812
rect 17552 7760 17558 7812
rect 17954 7809 17960 7812
rect 17948 7800 17960 7809
rect 17915 7772 17960 7800
rect 17948 7763 17960 7772
rect 17954 7760 17960 7763
rect 18012 7760 18018 7812
rect 10652 7704 12112 7732
rect 10652 7692 10658 7704
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 14090 7692 14096 7744
rect 14148 7692 14154 7744
rect 15102 7692 15108 7744
rect 15160 7732 15166 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15160 7704 15853 7732
rect 15160 7692 15166 7704
rect 15841 7701 15853 7704
rect 15887 7732 15899 7735
rect 16206 7732 16212 7744
rect 15887 7704 16212 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 19306 7732 19334 7840
rect 19886 7828 19892 7880
rect 19944 7828 19950 7880
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20772 7840 20913 7868
rect 20772 7828 20778 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 23014 7828 23020 7880
rect 23072 7868 23078 7880
rect 23290 7868 23296 7880
rect 23072 7840 23296 7868
rect 23072 7828 23078 7840
rect 23290 7828 23296 7840
rect 23348 7868 23354 7880
rect 23768 7868 23796 7976
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 27522 8004 27528 8016
rect 24872 7976 27528 8004
rect 24872 7948 24900 7976
rect 27522 7964 27528 7976
rect 27580 8004 27586 8016
rect 27893 8007 27951 8013
rect 27893 8004 27905 8007
rect 27580 7976 27905 8004
rect 27580 7964 27586 7976
rect 27893 7973 27905 7976
rect 27939 7973 27951 8007
rect 27893 7967 27951 7973
rect 40586 7964 40592 8016
rect 40644 8004 40650 8016
rect 40773 8007 40831 8013
rect 40773 8004 40785 8007
rect 40644 7976 40785 8004
rect 40644 7964 40650 7976
rect 40773 7973 40785 7976
rect 40819 8004 40831 8007
rect 40819 7976 42656 8004
rect 40819 7973 40831 7976
rect 40773 7967 40831 7973
rect 24854 7896 24860 7948
rect 24912 7896 24918 7948
rect 25133 7939 25191 7945
rect 25133 7905 25145 7939
rect 25179 7936 25191 7939
rect 25406 7936 25412 7948
rect 25179 7908 25412 7936
rect 25179 7905 25191 7908
rect 25133 7899 25191 7905
rect 25406 7896 25412 7908
rect 25464 7896 25470 7948
rect 25777 7939 25835 7945
rect 25777 7905 25789 7939
rect 25823 7936 25835 7939
rect 26418 7936 26424 7948
rect 25823 7908 26424 7936
rect 25823 7905 25835 7908
rect 25777 7899 25835 7905
rect 26418 7896 26424 7908
rect 26476 7896 26482 7948
rect 31113 7939 31171 7945
rect 31113 7905 31125 7939
rect 31159 7936 31171 7939
rect 32122 7936 32128 7948
rect 31159 7908 32128 7936
rect 31159 7905 31171 7908
rect 31113 7899 31171 7905
rect 32122 7896 32128 7908
rect 32180 7896 32186 7948
rect 41524 7945 41552 7976
rect 42628 7948 42656 7976
rect 41509 7939 41567 7945
rect 41509 7905 41521 7939
rect 41555 7905 41567 7939
rect 41509 7899 41567 7905
rect 41966 7896 41972 7948
rect 42024 7936 42030 7948
rect 42245 7939 42303 7945
rect 42245 7936 42257 7939
rect 42024 7908 42257 7936
rect 42024 7896 42030 7908
rect 42245 7905 42257 7908
rect 42291 7905 42303 7939
rect 42245 7899 42303 7905
rect 42610 7896 42616 7948
rect 42668 7896 42674 7948
rect 42812 7936 42840 8032
rect 43070 7964 43076 8016
rect 43128 8004 43134 8016
rect 45296 8004 45324 8035
rect 45830 8032 45836 8044
rect 45888 8032 45894 8084
rect 46934 8032 46940 8084
rect 46992 8072 46998 8084
rect 47578 8072 47584 8084
rect 46992 8044 47584 8072
rect 46992 8032 46998 8044
rect 47578 8032 47584 8044
rect 47636 8032 47642 8084
rect 50430 8032 50436 8084
rect 50488 8072 50494 8084
rect 50488 8044 51074 8072
rect 50488 8032 50494 8044
rect 43128 7976 45324 8004
rect 51046 8004 51074 8044
rect 52730 8032 52736 8084
rect 52788 8072 52794 8084
rect 53193 8075 53251 8081
rect 53193 8072 53205 8075
rect 52788 8044 53205 8072
rect 52788 8032 52794 8044
rect 53193 8041 53205 8044
rect 53239 8072 53251 8075
rect 53561 8075 53619 8081
rect 53561 8072 53573 8075
rect 53239 8044 53573 8072
rect 53239 8041 53251 8044
rect 53193 8035 53251 8041
rect 53561 8041 53573 8044
rect 53607 8041 53619 8075
rect 53561 8035 53619 8041
rect 52178 8004 52184 8016
rect 51046 7976 52184 8004
rect 43128 7964 43134 7976
rect 52178 7964 52184 7976
rect 52236 7964 52242 8016
rect 43533 7939 43591 7945
rect 43533 7936 43545 7939
rect 42812 7908 43545 7936
rect 43533 7905 43545 7908
rect 43579 7905 43591 7939
rect 43533 7899 43591 7905
rect 43990 7896 43996 7948
rect 44048 7896 44054 7948
rect 48314 7896 48320 7948
rect 48372 7936 48378 7948
rect 49326 7936 49332 7948
rect 48372 7908 49332 7936
rect 48372 7896 48378 7908
rect 49326 7896 49332 7908
rect 49384 7936 49390 7948
rect 50798 7936 50804 7948
rect 49384 7908 50804 7936
rect 49384 7896 49390 7908
rect 50798 7896 50804 7908
rect 50856 7896 50862 7948
rect 53576 7936 53604 8035
rect 56594 8032 56600 8084
rect 56652 8032 56658 8084
rect 58069 8075 58127 8081
rect 58069 8041 58081 8075
rect 58115 8072 58127 8075
rect 58434 8072 58440 8084
rect 58115 8044 58440 8072
rect 58115 8041 58127 8044
rect 58069 8035 58127 8041
rect 58434 8032 58440 8044
rect 58492 8032 58498 8084
rect 53745 7939 53803 7945
rect 53745 7936 53757 7939
rect 53576 7908 53757 7936
rect 53745 7905 53757 7908
rect 53791 7936 53803 7939
rect 53791 7908 53880 7936
rect 53791 7905 53803 7908
rect 53745 7899 53803 7905
rect 23348 7840 23796 7868
rect 23348 7828 23354 7840
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 23992 7840 24409 7868
rect 23992 7828 23998 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 25222 7828 25228 7880
rect 25280 7868 25286 7880
rect 25869 7871 25927 7877
rect 25869 7868 25881 7871
rect 25280 7840 25881 7868
rect 25280 7828 25286 7840
rect 25869 7837 25881 7840
rect 25915 7837 25927 7871
rect 25869 7831 25927 7837
rect 31754 7828 31760 7880
rect 31812 7828 31818 7880
rect 33134 7828 33140 7880
rect 33192 7828 33198 7880
rect 36078 7828 36084 7880
rect 36136 7828 36142 7880
rect 36814 7828 36820 7880
rect 36872 7828 36878 7880
rect 37550 7828 37556 7880
rect 37608 7828 37614 7880
rect 38102 7828 38108 7880
rect 38160 7828 38166 7880
rect 39390 7828 39396 7880
rect 39448 7828 39454 7880
rect 41230 7828 41236 7880
rect 41288 7828 41294 7880
rect 41325 7871 41383 7877
rect 41325 7837 41337 7871
rect 41371 7868 41383 7871
rect 41414 7868 41420 7880
rect 41371 7840 41420 7868
rect 41371 7837 41383 7840
rect 41325 7831 41383 7837
rect 41414 7828 41420 7840
rect 41472 7868 41478 7880
rect 42061 7871 42119 7877
rect 42061 7868 42073 7871
rect 41472 7840 42073 7868
rect 41472 7828 41478 7840
rect 23477 7803 23535 7809
rect 23477 7769 23489 7803
rect 23523 7800 23535 7803
rect 24854 7800 24860 7812
rect 23523 7772 24860 7800
rect 23523 7769 23535 7772
rect 23477 7763 23535 7769
rect 24854 7760 24860 7772
rect 24912 7760 24918 7812
rect 25041 7803 25099 7809
rect 25041 7769 25053 7803
rect 25087 7800 25099 7803
rect 30868 7803 30926 7809
rect 25087 7772 25912 7800
rect 25087 7769 25099 7772
rect 25041 7763 25099 7769
rect 25884 7744 25912 7772
rect 30868 7769 30880 7803
rect 30914 7800 30926 7803
rect 31205 7803 31263 7809
rect 31205 7800 31217 7803
rect 30914 7772 31217 7800
rect 30914 7769 30926 7772
rect 30868 7763 30926 7769
rect 31205 7769 31217 7772
rect 31251 7769 31263 7803
rect 31205 7763 31263 7769
rect 35345 7803 35403 7809
rect 35345 7769 35357 7803
rect 35391 7800 35403 7803
rect 35894 7800 35900 7812
rect 35391 7772 35900 7800
rect 35391 7769 35403 7772
rect 35345 7763 35403 7769
rect 35894 7760 35900 7772
rect 35952 7760 35958 7812
rect 19794 7732 19800 7744
rect 19306 7704 19800 7732
rect 19794 7692 19800 7704
rect 19852 7732 19858 7744
rect 21450 7732 21456 7744
rect 19852 7704 21456 7732
rect 19852 7692 19858 7704
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 23569 7735 23627 7741
rect 23569 7701 23581 7735
rect 23615 7732 23627 7735
rect 24394 7732 24400 7744
rect 23615 7704 24400 7732
rect 23615 7701 23627 7704
rect 23569 7695 23627 7701
rect 24394 7692 24400 7704
rect 24452 7692 24458 7744
rect 25866 7692 25872 7744
rect 25924 7692 25930 7744
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 27157 7735 27215 7741
rect 27157 7732 27169 7735
rect 26752 7704 27169 7732
rect 26752 7692 26758 7704
rect 27157 7701 27169 7704
rect 27203 7701 27215 7735
rect 27157 7695 27215 7701
rect 32582 7692 32588 7744
rect 32640 7692 32646 7744
rect 35526 7692 35532 7744
rect 35584 7692 35590 7744
rect 36262 7692 36268 7744
rect 36320 7692 36326 7744
rect 36722 7692 36728 7744
rect 36780 7732 36786 7744
rect 37001 7735 37059 7741
rect 37001 7732 37013 7735
rect 36780 7704 37013 7732
rect 36780 7692 36786 7704
rect 37001 7701 37013 7704
rect 37047 7701 37059 7735
rect 37001 7695 37059 7701
rect 38746 7692 38752 7744
rect 38804 7692 38810 7744
rect 38838 7692 38844 7744
rect 38896 7692 38902 7744
rect 41690 7692 41696 7744
rect 41748 7692 41754 7744
rect 41984 7732 42012 7840
rect 42061 7837 42073 7840
rect 42107 7837 42119 7871
rect 42061 7831 42119 7837
rect 42153 7871 42211 7877
rect 42153 7837 42165 7871
rect 42199 7868 42211 7871
rect 42886 7868 42892 7880
rect 42199 7840 42892 7868
rect 42199 7837 42211 7840
rect 42153 7831 42211 7837
rect 42886 7828 42892 7840
rect 42944 7868 42950 7880
rect 43254 7868 43260 7880
rect 42944 7840 43260 7868
rect 42944 7828 42950 7840
rect 43254 7828 43260 7840
rect 43312 7828 43318 7880
rect 43441 7871 43499 7877
rect 43441 7837 43453 7871
rect 43487 7868 43499 7871
rect 44008 7868 44036 7896
rect 53852 7880 53880 7908
rect 43487 7840 44036 7868
rect 44545 7871 44603 7877
rect 43487 7837 43499 7840
rect 43441 7831 43499 7837
rect 44545 7837 44557 7871
rect 44591 7868 44603 7871
rect 44634 7868 44640 7880
rect 44591 7840 44640 7868
rect 44591 7837 44603 7840
rect 44545 7831 44603 7837
rect 44634 7828 44640 7840
rect 44692 7828 44698 7880
rect 48958 7828 48964 7880
rect 49016 7828 49022 7880
rect 50614 7828 50620 7880
rect 50672 7868 50678 7880
rect 50985 7871 51043 7877
rect 50985 7868 50997 7871
rect 50672 7840 50997 7868
rect 50672 7828 50678 7840
rect 50985 7837 50997 7840
rect 51031 7837 51043 7871
rect 50985 7831 51043 7837
rect 52270 7828 52276 7880
rect 52328 7828 52334 7880
rect 53834 7828 53840 7880
rect 53892 7828 53898 7880
rect 55950 7828 55956 7880
rect 56008 7828 56014 7880
rect 56410 7828 56416 7880
rect 56468 7868 56474 7880
rect 56689 7871 56747 7877
rect 56689 7868 56701 7871
rect 56468 7840 56701 7868
rect 56468 7828 56474 7840
rect 56689 7837 56701 7840
rect 56735 7837 56747 7871
rect 56689 7831 56747 7837
rect 56778 7828 56784 7880
rect 56836 7868 56842 7880
rect 56945 7871 57003 7877
rect 56945 7868 56957 7871
rect 56836 7840 56957 7868
rect 56836 7828 56842 7840
rect 56945 7837 56957 7840
rect 56991 7837 57003 7871
rect 56945 7831 57003 7837
rect 57422 7828 57428 7880
rect 57480 7868 57486 7880
rect 58345 7871 58403 7877
rect 58345 7868 58357 7871
rect 57480 7840 58357 7868
rect 57480 7828 57486 7840
rect 58345 7837 58357 7840
rect 58391 7837 58403 7871
rect 58345 7831 58403 7837
rect 48072 7803 48130 7809
rect 48072 7769 48084 7803
rect 48118 7800 48130 7803
rect 48409 7803 48467 7809
rect 48409 7800 48421 7803
rect 48118 7772 48421 7800
rect 48118 7769 48130 7772
rect 48072 7763 48130 7769
rect 48409 7769 48421 7772
rect 48455 7769 48467 7803
rect 48409 7763 48467 7769
rect 51258 7760 51264 7812
rect 51316 7800 51322 7812
rect 51721 7803 51779 7809
rect 51721 7800 51733 7803
rect 51316 7772 51733 7800
rect 51316 7760 51322 7772
rect 51721 7769 51733 7772
rect 51767 7769 51779 7803
rect 51721 7763 51779 7769
rect 54012 7803 54070 7809
rect 54012 7769 54024 7803
rect 54058 7800 54070 7803
rect 55309 7803 55367 7809
rect 55309 7800 55321 7803
rect 54058 7772 55321 7800
rect 54058 7769 54070 7772
rect 54012 7763 54070 7769
rect 55309 7769 55321 7772
rect 55355 7769 55367 7803
rect 55309 7763 55367 7769
rect 43346 7732 43352 7744
rect 41984 7704 43352 7732
rect 43346 7692 43352 7704
rect 43404 7692 43410 7744
rect 43898 7692 43904 7744
rect 43956 7692 43962 7744
rect 51626 7692 51632 7744
rect 51684 7692 51690 7744
rect 55125 7735 55183 7741
rect 55125 7701 55137 7735
rect 55171 7732 55183 7735
rect 55490 7732 55496 7744
rect 55171 7704 55496 7732
rect 55171 7701 55183 7704
rect 55125 7695 55183 7701
rect 55490 7692 55496 7704
rect 55548 7692 55554 7744
rect 1104 7642 59040 7664
rect 1104 7590 15394 7642
rect 15446 7590 15458 7642
rect 15510 7590 15522 7642
rect 15574 7590 15586 7642
rect 15638 7590 15650 7642
rect 15702 7590 29838 7642
rect 29890 7590 29902 7642
rect 29954 7590 29966 7642
rect 30018 7590 30030 7642
rect 30082 7590 30094 7642
rect 30146 7590 44282 7642
rect 44334 7590 44346 7642
rect 44398 7590 44410 7642
rect 44462 7590 44474 7642
rect 44526 7590 44538 7642
rect 44590 7590 58726 7642
rect 58778 7590 58790 7642
rect 58842 7590 58854 7642
rect 58906 7590 58918 7642
rect 58970 7590 58982 7642
rect 59034 7590 59040 7642
rect 1104 7568 59040 7590
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 5258 7528 5264 7540
rect 4304 7500 5264 7528
rect 4304 7488 4310 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 6840 7460 6868 7491
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8260 7500 8861 7528
rect 8260 7488 8266 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 9214 7488 9220 7540
rect 9272 7488 9278 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9355 7500 9873 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9861 7497 9873 7500
rect 9907 7528 9919 7531
rect 10410 7528 10416 7540
rect 9907 7500 10416 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 12250 7528 12256 7540
rect 10744 7500 12256 7528
rect 10744 7488 10750 7500
rect 12250 7488 12256 7500
rect 12308 7528 12314 7540
rect 12308 7500 12572 7528
rect 12308 7488 12314 7500
rect 7374 7460 7380 7472
rect 6420 7432 7380 7460
rect 6420 7420 6426 7432
rect 7374 7420 7380 7432
rect 7432 7460 7438 7472
rect 8294 7460 8300 7472
rect 7432 7432 8300 7460
rect 7432 7420 7438 7432
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 8481 7463 8539 7469
rect 8481 7429 8493 7463
rect 8527 7460 8539 7463
rect 8662 7460 8668 7472
rect 8527 7432 8668 7460
rect 8527 7429 8539 7432
rect 8481 7423 8539 7429
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 11793 7463 11851 7469
rect 11793 7429 11805 7463
rect 11839 7460 11851 7463
rect 11882 7460 11888 7472
rect 11839 7432 11888 7460
rect 11839 7429 11851 7432
rect 11793 7423 11851 7429
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 2400 7395 2458 7401
rect 2400 7361 2412 7395
rect 2446 7392 2458 7395
rect 3142 7392 3148 7404
rect 2446 7364 3148 7392
rect 2446 7361 2458 7364
rect 2400 7355 2458 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 7282 7392 7288 7404
rect 6043 7364 7288 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 9030 7392 9036 7404
rect 8159 7364 9036 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 12345 7395 12403 7401
rect 12345 7392 12357 7395
rect 9732 7364 12357 7392
rect 9732 7352 9738 7364
rect 12345 7361 12357 7364
rect 12391 7361 12403 7395
rect 12544 7392 12572 7500
rect 12894 7488 12900 7540
rect 12952 7488 12958 7540
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14550 7528 14556 7540
rect 14056 7500 14556 7528
rect 14056 7488 14062 7500
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14792 7500 14933 7528
rect 14792 7488 14798 7500
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 14921 7491 14979 7497
rect 17586 7488 17592 7540
rect 17644 7488 17650 7540
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7528 18935 7531
rect 19334 7528 19340 7540
rect 18923 7500 19340 7528
rect 18923 7497 18935 7500
rect 18877 7491 18935 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 20162 7528 20168 7540
rect 19475 7500 20168 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 23014 7528 23020 7540
rect 22066 7500 23020 7528
rect 12612 7463 12670 7469
rect 12612 7429 12624 7463
rect 12658 7460 12670 7463
rect 12912 7460 12940 7488
rect 12658 7432 12940 7460
rect 14461 7463 14519 7469
rect 12658 7429 12670 7432
rect 12612 7423 12670 7429
rect 14461 7429 14473 7463
rect 14507 7460 14519 7463
rect 15654 7460 15660 7472
rect 14507 7432 15660 7460
rect 14507 7429 14519 7432
rect 14461 7423 14519 7429
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 13814 7392 13820 7404
rect 12544 7364 13820 7392
rect 12345 7355 12403 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 17497 7395 17555 7401
rect 13924 7364 15976 7392
rect 2130 7284 2136 7336
rect 2188 7284 2194 7336
rect 3602 7284 3608 7336
rect 3660 7284 3666 7336
rect 5166 7333 5172 7336
rect 5144 7327 5172 7333
rect 5144 7293 5156 7327
rect 5144 7287 5172 7293
rect 5166 7284 5172 7287
rect 5224 7284 5230 7336
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 6086 7324 6092 7336
rect 5583 7296 6092 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 6178 7284 6184 7336
rect 6236 7284 6242 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 9122 7324 9128 7336
rect 8628 7296 9128 7324
rect 8628 7284 8634 7296
rect 9122 7284 9128 7296
rect 9180 7324 9186 7336
rect 9401 7327 9459 7333
rect 9401 7324 9413 7327
rect 9180 7296 9413 7324
rect 9180 7284 9186 7296
rect 9401 7293 9413 7296
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 10376 7296 10425 7324
rect 10376 7284 10382 7296
rect 10413 7293 10425 7296
rect 10459 7293 10471 7327
rect 13924 7324 13952 7364
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 10413 7287 10471 7293
rect 13648 7296 13952 7324
rect 14016 7296 14289 7324
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 3878 7188 3884 7200
rect 3559 7160 3884 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 5718 7188 5724 7200
rect 4387 7160 5724 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 10744 7160 11069 7188
rect 10744 7148 10750 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11514 7148 11520 7200
rect 11572 7188 11578 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 11572 7160 12081 7188
rect 11572 7148 11578 7160
rect 12069 7157 12081 7160
rect 12115 7188 12127 7191
rect 13648 7188 13676 7296
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 14016 7265 14044 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 15010 7284 15016 7336
rect 15068 7284 15074 7336
rect 15948 7268 15976 7364
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17604 7392 17632 7488
rect 22066 7460 22094 7500
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 23934 7488 23940 7540
rect 23992 7488 23998 7540
rect 24026 7488 24032 7540
rect 24084 7488 24090 7540
rect 24489 7531 24547 7537
rect 24489 7497 24501 7531
rect 24535 7528 24547 7531
rect 25866 7528 25872 7540
rect 24535 7500 25872 7528
rect 24535 7497 24547 7500
rect 24489 7491 24547 7497
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 30466 7488 30472 7540
rect 30524 7488 30530 7540
rect 30561 7531 30619 7537
rect 30561 7497 30573 7531
rect 30607 7528 30619 7531
rect 30834 7528 30840 7540
rect 30607 7500 30840 7528
rect 30607 7497 30619 7500
rect 30561 7491 30619 7497
rect 30834 7488 30840 7500
rect 30892 7488 30898 7540
rect 30929 7531 30987 7537
rect 30929 7497 30941 7531
rect 30975 7528 30987 7531
rect 31754 7528 31760 7540
rect 30975 7500 31760 7528
rect 30975 7497 30987 7500
rect 30929 7491 30987 7497
rect 31754 7488 31760 7500
rect 31812 7488 31818 7540
rect 32769 7531 32827 7537
rect 32769 7497 32781 7531
rect 32815 7528 32827 7531
rect 33134 7528 33140 7540
rect 32815 7500 33140 7528
rect 32815 7497 32827 7500
rect 32769 7491 32827 7497
rect 33134 7488 33140 7500
rect 33192 7488 33198 7540
rect 35158 7528 35164 7540
rect 34716 7500 35164 7528
rect 19628 7432 22094 7460
rect 17543 7364 17632 7392
rect 17764 7395 17822 7401
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17764 7361 17776 7395
rect 17810 7392 17822 7395
rect 18046 7392 18052 7404
rect 17810 7364 18052 7392
rect 17810 7361 17822 7364
rect 17764 7355 17822 7361
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19518 7392 19524 7404
rect 19383 7364 19524 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 17310 7284 17316 7336
rect 17368 7284 17374 7336
rect 18782 7284 18788 7336
rect 18840 7284 18846 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 19628 7333 19656 7432
rect 23566 7420 23572 7472
rect 23624 7420 23630 7472
rect 24670 7420 24676 7472
rect 24728 7420 24734 7472
rect 33962 7460 33968 7472
rect 33152 7432 33968 7460
rect 20248 7395 20306 7401
rect 20248 7361 20260 7395
rect 20294 7392 20306 7395
rect 20990 7392 20996 7404
rect 20294 7364 20996 7392
rect 20294 7361 20306 7364
rect 20248 7355 20306 7361
rect 20990 7352 20996 7364
rect 21048 7352 21054 7404
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 22462 7392 22468 7404
rect 21508 7364 22468 7392
rect 21508 7352 21514 7364
rect 22462 7352 22468 7364
rect 22520 7392 22526 7404
rect 22557 7395 22615 7401
rect 22557 7392 22569 7395
rect 22520 7364 22569 7392
rect 22520 7352 22526 7364
rect 22557 7361 22569 7364
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 22824 7395 22882 7401
rect 22824 7361 22836 7395
rect 22870 7392 22882 7395
rect 23584 7392 23612 7420
rect 22870 7364 23612 7392
rect 22870 7361 22882 7364
rect 22824 7355 22882 7361
rect 24394 7352 24400 7404
rect 24452 7352 24458 7404
rect 19613 7327 19671 7333
rect 19613 7324 19625 7327
rect 19300 7296 19625 7324
rect 19300 7284 19306 7296
rect 19613 7293 19625 7296
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 24688 7333 24716 7420
rect 25590 7352 25596 7404
rect 25648 7352 25654 7404
rect 25866 7352 25872 7404
rect 25924 7352 25930 7404
rect 26418 7352 26424 7404
rect 26476 7352 26482 7404
rect 33152 7401 33180 7432
rect 33962 7420 33968 7432
rect 34020 7460 34026 7472
rect 34716 7460 34744 7500
rect 35158 7488 35164 7500
rect 35216 7488 35222 7540
rect 35526 7488 35532 7540
rect 35584 7488 35590 7540
rect 35897 7531 35955 7537
rect 35897 7497 35909 7531
rect 35943 7528 35955 7531
rect 36630 7528 36636 7540
rect 35943 7500 36636 7528
rect 35943 7497 35955 7500
rect 35897 7491 35955 7497
rect 36630 7488 36636 7500
rect 36688 7488 36694 7540
rect 38933 7531 38991 7537
rect 38933 7497 38945 7531
rect 38979 7528 38991 7531
rect 39390 7528 39396 7540
rect 38979 7500 39396 7528
rect 38979 7497 38991 7500
rect 38933 7491 38991 7497
rect 39390 7488 39396 7500
rect 39448 7488 39454 7540
rect 41598 7488 41604 7540
rect 41656 7528 41662 7540
rect 41693 7531 41751 7537
rect 41693 7528 41705 7531
rect 41656 7500 41705 7528
rect 41656 7488 41662 7500
rect 41693 7497 41705 7500
rect 41739 7497 41751 7531
rect 41693 7491 41751 7497
rect 41966 7488 41972 7540
rect 42024 7488 42030 7540
rect 43346 7488 43352 7540
rect 43404 7528 43410 7540
rect 44361 7531 44419 7537
rect 43404 7500 44128 7528
rect 43404 7488 43410 7500
rect 34020 7432 34744 7460
rect 34784 7463 34842 7469
rect 34020 7420 34026 7432
rect 34784 7429 34796 7463
rect 34830 7460 34842 7463
rect 35544 7460 35572 7488
rect 34830 7432 35572 7460
rect 34830 7429 34842 7432
rect 34784 7423 34842 7429
rect 36170 7420 36176 7472
rect 36228 7460 36234 7472
rect 36449 7463 36507 7469
rect 36449 7460 36461 7463
rect 36228 7432 36461 7460
rect 36228 7420 36234 7432
rect 36449 7429 36461 7432
rect 36495 7429 36507 7463
rect 40580 7463 40638 7469
rect 36449 7423 36507 7429
rect 37660 7432 40356 7460
rect 37660 7404 37688 7432
rect 26605 7395 26663 7401
rect 26605 7361 26617 7395
rect 26651 7392 26663 7395
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 26651 7364 27353 7392
rect 26651 7361 26663 7364
rect 26605 7355 26663 7361
rect 27341 7361 27353 7364
rect 27387 7392 27399 7395
rect 27801 7395 27859 7401
rect 27801 7392 27813 7395
rect 27387 7364 27813 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 27801 7361 27813 7364
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 33137 7395 33195 7401
rect 33137 7361 33149 7395
rect 33183 7361 33195 7395
rect 33137 7355 33195 7361
rect 33229 7395 33287 7401
rect 33229 7361 33241 7395
rect 33275 7392 33287 7395
rect 34241 7395 34299 7401
rect 34241 7392 34253 7395
rect 33275 7364 34253 7392
rect 33275 7361 33287 7364
rect 33229 7355 33287 7361
rect 34241 7361 34253 7364
rect 34287 7361 34299 7395
rect 34241 7355 34299 7361
rect 19981 7327 20039 7333
rect 19981 7324 19993 7327
rect 19852 7296 19993 7324
rect 19852 7284 19858 7296
rect 19981 7293 19993 7296
rect 20027 7293 20039 7327
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 19981 7287 20039 7293
rect 22066 7296 22385 7324
rect 14001 7259 14059 7265
rect 14001 7256 14013 7259
rect 13872 7228 14013 7256
rect 13872 7216 13878 7228
rect 14001 7225 14013 7228
rect 14047 7225 14059 7259
rect 14001 7219 14059 7225
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 16025 7259 16083 7265
rect 16025 7256 16037 7259
rect 15988 7228 16037 7256
rect 15988 7216 15994 7228
rect 16025 7225 16037 7228
rect 16071 7256 16083 7259
rect 16071 7228 17540 7256
rect 16071 7225 16083 7228
rect 16025 7219 16083 7225
rect 12115 7160 13676 7188
rect 13725 7191 13783 7197
rect 12115 7157 12127 7160
rect 12069 7151 12127 7157
rect 13725 7157 13737 7191
rect 13771 7188 13783 7191
rect 13906 7188 13912 7200
rect 13771 7160 13912 7188
rect 13771 7157 13783 7160
rect 13725 7151 13783 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 16264 7160 16405 7188
rect 16264 7148 16270 7160
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 16669 7191 16727 7197
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 17034 7188 17040 7200
rect 16715 7160 17040 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 17512 7188 17540 7228
rect 18800 7188 18828 7284
rect 21361 7259 21419 7265
rect 21361 7225 21373 7259
rect 21407 7256 21419 7259
rect 22066 7256 22094 7296
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 24673 7327 24731 7333
rect 24673 7293 24685 7327
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 25682 7284 25688 7336
rect 25740 7333 25746 7336
rect 25740 7327 25789 7333
rect 25740 7293 25743 7327
rect 25777 7293 25789 7327
rect 26436 7324 26464 7352
rect 26789 7327 26847 7333
rect 26789 7324 26801 7327
rect 26436 7296 26801 7324
rect 25740 7287 25789 7293
rect 26789 7293 26801 7296
rect 26835 7293 26847 7327
rect 26789 7287 26847 7293
rect 25740 7284 25746 7287
rect 27062 7284 27068 7336
rect 27120 7324 27126 7336
rect 27433 7327 27491 7333
rect 27433 7324 27445 7327
rect 27120 7296 27445 7324
rect 27120 7284 27126 7296
rect 27433 7293 27445 7296
rect 27479 7293 27491 7327
rect 27433 7287 27491 7293
rect 27522 7284 27528 7336
rect 27580 7284 27586 7336
rect 28350 7284 28356 7336
rect 28408 7284 28414 7336
rect 29362 7284 29368 7336
rect 29420 7284 29426 7336
rect 30101 7327 30159 7333
rect 30101 7293 30113 7327
rect 30147 7324 30159 7327
rect 30190 7324 30196 7336
rect 30147 7296 30196 7324
rect 30147 7293 30159 7296
rect 30101 7287 30159 7293
rect 30190 7284 30196 7296
rect 30248 7284 30254 7336
rect 30377 7327 30435 7333
rect 30377 7293 30389 7327
rect 30423 7293 30435 7327
rect 30377 7287 30435 7293
rect 21407 7228 22094 7256
rect 21407 7225 21419 7228
rect 21361 7219 21419 7225
rect 26050 7216 26056 7268
rect 26108 7256 26114 7268
rect 26145 7259 26203 7265
rect 26145 7256 26157 7259
rect 26108 7228 26157 7256
rect 26108 7216 26114 7228
rect 26145 7225 26157 7228
rect 26191 7225 26203 7259
rect 27246 7256 27252 7268
rect 26145 7219 26203 7225
rect 26896 7228 27252 7256
rect 17512 7160 18828 7188
rect 18966 7148 18972 7200
rect 19024 7148 19030 7200
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 20772 7160 21833 7188
rect 20772 7148 20778 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 21821 7151 21879 7157
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 26896 7188 26924 7228
rect 27246 7216 27252 7228
rect 27304 7216 27310 7268
rect 27540 7256 27568 7284
rect 30392 7256 30420 7287
rect 30926 7284 30932 7336
rect 30984 7324 30990 7336
rect 32585 7327 32643 7333
rect 32585 7324 32597 7327
rect 30984 7296 32597 7324
rect 30984 7284 30990 7296
rect 32585 7293 32597 7296
rect 32631 7293 32643 7327
rect 32585 7287 32643 7293
rect 33321 7327 33379 7333
rect 33321 7293 33333 7327
rect 33367 7293 33379 7327
rect 33321 7287 33379 7293
rect 31205 7259 31263 7265
rect 31205 7256 31217 7259
rect 27540 7228 31217 7256
rect 31205 7225 31217 7228
rect 31251 7225 31263 7259
rect 32600 7256 32628 7287
rect 33336 7256 33364 7287
rect 33594 7284 33600 7336
rect 33652 7284 33658 7336
rect 32600 7228 33364 7256
rect 31205 7219 31263 7225
rect 24995 7160 26924 7188
rect 26973 7191 27031 7197
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 26973 7157 26985 7191
rect 27019 7188 27031 7191
rect 27614 7188 27620 7200
rect 27019 7160 27620 7188
rect 27019 7157 27031 7160
rect 26973 7151 27031 7157
rect 27614 7148 27620 7160
rect 27672 7148 27678 7200
rect 28721 7191 28779 7197
rect 28721 7157 28733 7191
rect 28767 7188 28779 7191
rect 29270 7188 29276 7200
rect 28767 7160 29276 7188
rect 28767 7157 28779 7160
rect 28721 7151 28779 7157
rect 29270 7148 29276 7160
rect 29328 7148 29334 7200
rect 29454 7148 29460 7200
rect 29512 7148 29518 7200
rect 34256 7188 34284 7355
rect 35066 7352 35072 7404
rect 35124 7392 35130 7404
rect 36357 7395 36415 7401
rect 36357 7392 36369 7395
rect 35124 7364 36369 7392
rect 35124 7352 35130 7364
rect 36357 7361 36369 7364
rect 36403 7361 36415 7395
rect 36357 7355 36415 7361
rect 37553 7395 37611 7401
rect 37553 7361 37565 7395
rect 37599 7392 37611 7395
rect 37642 7392 37648 7404
rect 37599 7364 37648 7392
rect 37599 7361 37611 7364
rect 37553 7355 37611 7361
rect 37642 7352 37648 7364
rect 37700 7352 37706 7404
rect 40328 7401 40356 7432
rect 40580 7429 40592 7463
rect 40626 7460 40638 7463
rect 40770 7460 40776 7472
rect 40626 7432 40776 7460
rect 40626 7429 40638 7432
rect 40580 7423 40638 7429
rect 40770 7420 40776 7432
rect 40828 7420 40834 7472
rect 44100 7460 44128 7500
rect 44361 7497 44373 7531
rect 44407 7528 44419 7531
rect 44634 7528 44640 7540
rect 44407 7500 44640 7528
rect 44407 7497 44419 7500
rect 44361 7491 44419 7497
rect 44634 7488 44640 7500
rect 44692 7488 44698 7540
rect 47762 7488 47768 7540
rect 47820 7488 47826 7540
rect 47857 7531 47915 7537
rect 47857 7497 47869 7531
rect 47903 7528 47915 7531
rect 48222 7528 48228 7540
rect 47903 7500 48228 7528
rect 47903 7497 47915 7500
rect 47857 7491 47915 7497
rect 48222 7488 48228 7500
rect 48280 7488 48286 7540
rect 48317 7531 48375 7537
rect 48317 7497 48329 7531
rect 48363 7528 48375 7531
rect 48958 7528 48964 7540
rect 48363 7500 48964 7528
rect 48363 7497 48375 7500
rect 48317 7491 48375 7497
rect 48958 7488 48964 7500
rect 49016 7488 49022 7540
rect 50798 7488 50804 7540
rect 50856 7528 50862 7540
rect 50856 7500 51074 7528
rect 50856 7488 50862 7500
rect 44821 7463 44879 7469
rect 44821 7460 44833 7463
rect 44100 7432 44833 7460
rect 44821 7429 44833 7432
rect 44867 7429 44879 7463
rect 47780 7460 47808 7488
rect 47946 7460 47952 7472
rect 47780 7432 47952 7460
rect 44821 7423 44879 7429
rect 47946 7420 47952 7432
rect 48004 7420 48010 7472
rect 48498 7420 48504 7472
rect 48556 7460 48562 7472
rect 48777 7463 48835 7469
rect 48777 7460 48789 7463
rect 48556 7432 48789 7460
rect 48556 7420 48562 7432
rect 48777 7429 48789 7432
rect 48823 7429 48835 7463
rect 51046 7460 51074 7500
rect 51626 7488 51632 7540
rect 51684 7528 51690 7540
rect 51721 7531 51779 7537
rect 51721 7528 51733 7531
rect 51684 7500 51733 7528
rect 51684 7488 51690 7500
rect 51721 7497 51733 7500
rect 51767 7497 51779 7531
rect 51721 7491 51779 7497
rect 52181 7531 52239 7537
rect 52181 7497 52193 7531
rect 52227 7528 52239 7531
rect 52270 7528 52276 7540
rect 52227 7500 52276 7528
rect 52227 7497 52239 7500
rect 52181 7491 52239 7497
rect 52270 7488 52276 7500
rect 52328 7488 52334 7540
rect 53834 7488 53840 7540
rect 53892 7488 53898 7540
rect 54849 7531 54907 7537
rect 54849 7497 54861 7531
rect 54895 7528 54907 7531
rect 55306 7528 55312 7540
rect 54895 7500 55312 7528
rect 54895 7497 54907 7500
rect 54849 7491 54907 7497
rect 55306 7488 55312 7500
rect 55364 7528 55370 7540
rect 56318 7528 56324 7540
rect 55364 7500 56324 7528
rect 55364 7488 55370 7500
rect 56318 7488 56324 7500
rect 56376 7488 56382 7540
rect 53852 7460 53880 7488
rect 51046 7432 51396 7460
rect 48777 7423 48835 7429
rect 37820 7395 37878 7401
rect 37820 7361 37832 7395
rect 37866 7392 37878 7395
rect 39025 7395 39083 7401
rect 39025 7392 39037 7395
rect 37866 7364 39037 7392
rect 37866 7361 37878 7364
rect 37820 7355 37878 7361
rect 39025 7361 39037 7364
rect 39071 7361 39083 7395
rect 39025 7355 39083 7361
rect 40313 7395 40371 7401
rect 40313 7361 40325 7395
rect 40359 7361 40371 7395
rect 40313 7355 40371 7361
rect 43070 7352 43076 7404
rect 43128 7352 43134 7404
rect 43162 7352 43168 7404
rect 43220 7401 43226 7404
rect 43220 7395 43269 7401
rect 43220 7361 43223 7395
rect 43257 7361 43269 7395
rect 43220 7355 43269 7361
rect 43220 7352 43226 7355
rect 43346 7352 43352 7404
rect 43404 7352 43410 7404
rect 44085 7395 44143 7401
rect 44085 7361 44097 7395
rect 44131 7392 44143 7395
rect 44729 7395 44787 7401
rect 44729 7392 44741 7395
rect 44131 7364 44741 7392
rect 44131 7361 44143 7364
rect 44085 7355 44143 7361
rect 44729 7361 44741 7364
rect 44775 7392 44787 7395
rect 45189 7395 45247 7401
rect 45189 7392 45201 7395
rect 44775 7364 45201 7392
rect 44775 7361 44787 7364
rect 44729 7355 44787 7361
rect 45189 7361 45201 7364
rect 45235 7361 45247 7395
rect 45189 7355 45247 7361
rect 48958 7352 48964 7404
rect 49016 7352 49022 7404
rect 49881 7395 49939 7401
rect 49881 7361 49893 7395
rect 49927 7392 49939 7395
rect 50706 7392 50712 7404
rect 49927 7364 50712 7392
rect 49927 7361 49939 7364
rect 49881 7355 49939 7361
rect 34514 7284 34520 7336
rect 34572 7284 34578 7336
rect 36541 7327 36599 7333
rect 36541 7324 36553 7327
rect 36372 7296 36553 7324
rect 36372 7268 36400 7296
rect 36541 7293 36553 7296
rect 36587 7324 36599 7327
rect 37001 7327 37059 7333
rect 37001 7324 37013 7327
rect 36587 7296 37013 7324
rect 36587 7293 36599 7296
rect 36541 7287 36599 7293
rect 37001 7293 37013 7296
rect 37047 7293 37059 7327
rect 37001 7287 37059 7293
rect 36354 7216 36360 7268
rect 36412 7216 36418 7268
rect 34698 7188 34704 7200
rect 34256 7160 34704 7188
rect 34698 7148 34704 7160
rect 34756 7148 34762 7200
rect 35618 7148 35624 7200
rect 35676 7188 35682 7200
rect 35989 7191 36047 7197
rect 35989 7188 36001 7191
rect 35676 7160 36001 7188
rect 35676 7148 35682 7160
rect 35989 7157 36001 7160
rect 36035 7157 36047 7191
rect 37016 7188 37044 7287
rect 39114 7284 39120 7336
rect 39172 7324 39178 7336
rect 39577 7327 39635 7333
rect 39577 7324 39589 7327
rect 39172 7296 39589 7324
rect 39172 7284 39178 7296
rect 39577 7293 39589 7296
rect 39623 7293 39635 7327
rect 39577 7287 39635 7293
rect 44174 7284 44180 7336
rect 44232 7324 44238 7336
rect 44269 7327 44327 7333
rect 44269 7324 44281 7327
rect 44232 7296 44281 7324
rect 44232 7284 44238 7296
rect 44269 7293 44281 7296
rect 44315 7293 44327 7327
rect 44269 7287 44327 7293
rect 44910 7284 44916 7336
rect 44968 7284 44974 7336
rect 45738 7284 45744 7336
rect 45796 7284 45802 7336
rect 46474 7284 46480 7336
rect 46532 7284 46538 7336
rect 46658 7284 46664 7336
rect 46716 7284 46722 7336
rect 47394 7284 47400 7336
rect 47452 7324 47458 7336
rect 47673 7327 47731 7333
rect 47673 7324 47685 7327
rect 47452 7296 47685 7324
rect 47452 7284 47458 7296
rect 47673 7293 47685 7296
rect 47719 7324 47731 7327
rect 48685 7327 48743 7333
rect 48685 7324 48697 7327
rect 47719 7296 48697 7324
rect 47719 7293 47731 7296
rect 47673 7287 47731 7293
rect 48685 7293 48697 7296
rect 48731 7324 48743 7327
rect 49896 7324 49924 7355
rect 50706 7352 50712 7364
rect 50764 7352 50770 7404
rect 51097 7395 51155 7401
rect 51097 7361 51109 7395
rect 51143 7392 51155 7395
rect 51258 7392 51264 7404
rect 51143 7364 51264 7392
rect 51143 7361 51155 7364
rect 51097 7355 51155 7361
rect 51258 7352 51264 7364
rect 51316 7352 51322 7404
rect 51368 7401 51396 7432
rect 53484 7432 53880 7460
rect 51353 7395 51411 7401
rect 51353 7361 51365 7395
rect 51399 7361 51411 7395
rect 51353 7355 51411 7361
rect 51813 7395 51871 7401
rect 51813 7361 51825 7395
rect 51859 7392 51871 7395
rect 51994 7392 52000 7404
rect 51859 7364 52000 7392
rect 51859 7361 51871 7364
rect 51813 7355 51871 7361
rect 51994 7352 52000 7364
rect 52052 7352 52058 7404
rect 53484 7401 53512 7432
rect 53926 7420 53932 7472
rect 53984 7420 53990 7472
rect 57330 7420 57336 7472
rect 57388 7460 57394 7472
rect 58253 7463 58311 7469
rect 58253 7460 58265 7463
rect 57388 7432 58265 7460
rect 57388 7420 57394 7432
rect 58253 7429 58265 7432
rect 58299 7429 58311 7463
rect 58253 7423 58311 7429
rect 53469 7395 53527 7401
rect 53469 7361 53481 7395
rect 53515 7361 53527 7395
rect 53469 7355 53527 7361
rect 53736 7395 53794 7401
rect 53736 7361 53748 7395
rect 53782 7392 53794 7395
rect 53944 7392 53972 7420
rect 53782 7364 53972 7392
rect 53782 7361 53794 7364
rect 53736 7355 53794 7361
rect 56226 7352 56232 7404
rect 56284 7352 56290 7404
rect 56318 7352 56324 7404
rect 56376 7401 56382 7404
rect 56376 7395 56425 7401
rect 56376 7361 56379 7395
rect 56413 7361 56425 7395
rect 56376 7355 56425 7361
rect 56376 7352 56382 7355
rect 56502 7352 56508 7404
rect 56560 7352 56566 7404
rect 57238 7352 57244 7404
rect 57296 7352 57302 7404
rect 58434 7352 58440 7404
rect 58492 7352 58498 7404
rect 48731 7296 49924 7324
rect 51629 7327 51687 7333
rect 48731 7293 48743 7296
rect 48685 7287 48743 7293
rect 51629 7293 51641 7327
rect 51675 7324 51687 7327
rect 51675 7296 52592 7324
rect 51675 7293 51687 7296
rect 51629 7287 51687 7293
rect 43625 7259 43683 7265
rect 43625 7225 43637 7259
rect 43671 7256 43683 7259
rect 43990 7256 43996 7268
rect 43671 7228 43996 7256
rect 43671 7225 43683 7228
rect 43625 7219 43683 7225
rect 43990 7216 43996 7228
rect 44048 7216 44054 7268
rect 45646 7216 45652 7268
rect 45704 7256 45710 7268
rect 45704 7228 47348 7256
rect 45704 7216 45710 7228
rect 38930 7188 38936 7200
rect 37016 7160 38936 7188
rect 35989 7151 36047 7157
rect 38930 7148 38936 7160
rect 38988 7148 38994 7200
rect 42429 7191 42487 7197
rect 42429 7157 42441 7191
rect 42475 7188 42487 7191
rect 45186 7188 45192 7200
rect 42475 7160 45192 7188
rect 42475 7157 42487 7160
rect 42429 7151 42487 7157
rect 45186 7148 45192 7160
rect 45244 7148 45250 7200
rect 45554 7148 45560 7200
rect 45612 7188 45618 7200
rect 47320 7197 47348 7228
rect 45925 7191 45983 7197
rect 45925 7188 45937 7191
rect 45612 7160 45937 7188
rect 45612 7148 45618 7160
rect 45925 7157 45937 7160
rect 45971 7157 45983 7191
rect 45925 7151 45983 7157
rect 47305 7191 47363 7197
rect 47305 7157 47317 7191
rect 47351 7188 47363 7191
rect 47578 7188 47584 7200
rect 47351 7160 47584 7188
rect 47351 7157 47363 7160
rect 47305 7151 47363 7157
rect 47578 7148 47584 7160
rect 47636 7148 47642 7200
rect 49421 7191 49479 7197
rect 49421 7157 49433 7191
rect 49467 7188 49479 7191
rect 49878 7188 49884 7200
rect 49467 7160 49884 7188
rect 49467 7157 49479 7160
rect 49421 7151 49479 7157
rect 49878 7148 49884 7160
rect 49936 7148 49942 7200
rect 49973 7191 50031 7197
rect 49973 7157 49985 7191
rect 50019 7188 50031 7191
rect 50614 7188 50620 7200
rect 50019 7160 50620 7188
rect 50019 7157 50031 7160
rect 49973 7151 50031 7157
rect 50614 7148 50620 7160
rect 50672 7148 50678 7200
rect 50706 7148 50712 7200
rect 50764 7188 50770 7200
rect 51644 7188 51672 7287
rect 52564 7265 52592 7296
rect 53282 7284 53288 7336
rect 53340 7284 53346 7336
rect 56781 7327 56839 7333
rect 56781 7324 56793 7327
rect 55232 7296 56793 7324
rect 52549 7259 52607 7265
rect 52549 7225 52561 7259
rect 52595 7256 52607 7259
rect 52595 7228 52868 7256
rect 52595 7225 52607 7228
rect 52549 7219 52607 7225
rect 50764 7160 51672 7188
rect 50764 7148 50770 7160
rect 52730 7148 52736 7200
rect 52788 7148 52794 7200
rect 52840 7188 52868 7228
rect 54202 7188 54208 7200
rect 52840 7160 54208 7188
rect 54202 7148 54208 7160
rect 54260 7148 54266 7200
rect 54754 7148 54760 7200
rect 54812 7188 54818 7200
rect 55232 7197 55260 7296
rect 56781 7293 56793 7296
rect 56827 7293 56839 7327
rect 56781 7287 56839 7293
rect 57330 7284 57336 7336
rect 57388 7324 57394 7336
rect 57425 7327 57483 7333
rect 57425 7324 57437 7327
rect 57388 7296 57437 7324
rect 57388 7284 57394 7296
rect 57425 7293 57437 7296
rect 57471 7293 57483 7327
rect 57425 7287 57483 7293
rect 55217 7191 55275 7197
rect 55217 7188 55229 7191
rect 54812 7160 55229 7188
rect 54812 7148 54818 7160
rect 55217 7157 55229 7160
rect 55263 7157 55275 7191
rect 55217 7151 55275 7157
rect 55585 7191 55643 7197
rect 55585 7157 55597 7191
rect 55631 7188 55643 7191
rect 56318 7188 56324 7200
rect 55631 7160 56324 7188
rect 55631 7157 55643 7160
rect 55585 7151 55643 7157
rect 56318 7148 56324 7160
rect 56376 7148 56382 7200
rect 56870 7148 56876 7200
rect 56928 7188 56934 7200
rect 57514 7188 57520 7200
rect 56928 7160 57520 7188
rect 56928 7148 56934 7160
rect 57514 7148 57520 7160
rect 57572 7188 57578 7200
rect 58069 7191 58127 7197
rect 58069 7188 58081 7191
rect 57572 7160 58081 7188
rect 57572 7148 57578 7160
rect 58069 7157 58081 7160
rect 58115 7157 58127 7191
rect 58069 7151 58127 7157
rect 1104 7098 58880 7120
rect 1104 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 22616 7098
rect 22668 7046 22680 7098
rect 22732 7046 22744 7098
rect 22796 7046 22808 7098
rect 22860 7046 22872 7098
rect 22924 7046 37060 7098
rect 37112 7046 37124 7098
rect 37176 7046 37188 7098
rect 37240 7046 37252 7098
rect 37304 7046 37316 7098
rect 37368 7046 51504 7098
rect 51556 7046 51568 7098
rect 51620 7046 51632 7098
rect 51684 7046 51696 7098
rect 51748 7046 51760 7098
rect 51812 7046 58880 7098
rect 1104 7024 58880 7046
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 3602 6984 3608 6996
rect 3467 6956 3608 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 9122 6944 9128 6996
rect 9180 6944 9186 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 12406 6956 13921 6984
rect 4614 6916 4620 6928
rect 4448 6888 4620 6916
rect 4448 6857 4476 6888
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 10045 6851 10103 6857
rect 10045 6817 10057 6851
rect 10091 6848 10103 6851
rect 11514 6848 11520 6860
rect 10091 6820 11520 6848
rect 10091 6817 10103 6820
rect 10045 6811 10103 6817
rect 11514 6808 11520 6820
rect 11572 6808 11578 6860
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6848 11943 6851
rect 12406 6848 12434 6956
rect 13909 6953 13921 6956
rect 13955 6953 13967 6987
rect 13909 6947 13967 6953
rect 11931 6820 12434 6848
rect 13924 6848 13952 6947
rect 17310 6944 17316 6996
rect 17368 6984 17374 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17368 6956 17509 6984
rect 17368 6944 17374 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 18046 6944 18052 6996
rect 18104 6984 18110 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 18104 6956 18429 6984
rect 18104 6944 18110 6956
rect 18417 6953 18429 6956
rect 18463 6953 18475 6987
rect 18417 6947 18475 6953
rect 19521 6987 19579 6993
rect 19521 6953 19533 6987
rect 19567 6984 19579 6987
rect 19794 6984 19800 6996
rect 19567 6956 19800 6984
rect 19567 6953 19579 6956
rect 19521 6947 19579 6953
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 20990 6944 20996 6996
rect 21048 6944 21054 6996
rect 22066 6956 24716 6984
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15838 6916 15844 6928
rect 15436 6888 15844 6916
rect 15436 6876 15442 6888
rect 15838 6876 15844 6888
rect 15896 6876 15902 6928
rect 22066 6916 22094 6956
rect 20272 6888 22094 6916
rect 24688 6916 24716 6956
rect 24854 6944 24860 6996
rect 24912 6984 24918 6996
rect 25041 6987 25099 6993
rect 25041 6984 25053 6987
rect 24912 6956 25053 6984
rect 24912 6944 24918 6956
rect 25041 6953 25053 6956
rect 25087 6984 25099 6987
rect 25682 6984 25688 6996
rect 25087 6956 25688 6984
rect 25087 6953 25099 6956
rect 25041 6947 25099 6953
rect 25682 6944 25688 6956
rect 25740 6944 25746 6996
rect 26694 6984 26700 6996
rect 25884 6956 26700 6984
rect 24946 6916 24952 6928
rect 24688 6888 24952 6916
rect 20272 6860 20300 6888
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 25884 6916 25912 6956
rect 26694 6944 26700 6956
rect 26752 6984 26758 6996
rect 27801 6987 27859 6993
rect 27801 6984 27813 6987
rect 26752 6956 27813 6984
rect 26752 6944 26758 6956
rect 27801 6953 27813 6956
rect 27847 6953 27859 6987
rect 27801 6947 27859 6953
rect 25424 6888 25912 6916
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 13924 6820 15117 6848
rect 11931 6817 11943 6820
rect 11885 6811 11943 6817
rect 15105 6817 15117 6820
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 15654 6808 15660 6860
rect 15712 6848 15718 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15712 6820 16037 6848
rect 15712 6808 15718 6820
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16025 6811 16083 6817
rect 18966 6808 18972 6860
rect 19024 6808 19030 6860
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 20254 6848 20260 6860
rect 19484 6820 20260 6848
rect 19484 6808 19490 6820
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 22094 6848 22100 6860
rect 21775 6820 22100 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22462 6808 22468 6860
rect 22520 6808 22526 6860
rect 24118 6808 24124 6860
rect 24176 6848 24182 6860
rect 25424 6848 25452 6888
rect 24176 6820 25452 6848
rect 24176 6808 24182 6820
rect 25498 6808 25504 6860
rect 25556 6808 25562 6860
rect 25884 6848 25912 6888
rect 25950 6851 26008 6857
rect 25950 6848 25962 6851
rect 25884 6820 25962 6848
rect 25950 6817 25962 6820
rect 25996 6817 26008 6851
rect 27816 6848 27844 6947
rect 29362 6944 29368 6996
rect 29420 6944 29426 6996
rect 33413 6987 33471 6993
rect 33413 6953 33425 6987
rect 33459 6984 33471 6987
rect 33594 6984 33600 6996
rect 33459 6956 33600 6984
rect 33459 6953 33471 6956
rect 33413 6947 33471 6953
rect 33594 6944 33600 6956
rect 33652 6944 33658 6996
rect 36173 6987 36231 6993
rect 36173 6953 36185 6987
rect 36219 6984 36231 6987
rect 36814 6984 36820 6996
rect 36219 6956 36820 6984
rect 36219 6953 36231 6956
rect 36173 6947 36231 6953
rect 36814 6944 36820 6956
rect 36872 6944 36878 6996
rect 37093 6987 37151 6993
rect 37093 6953 37105 6987
rect 37139 6984 37151 6987
rect 38102 6984 38108 6996
rect 37139 6956 38108 6984
rect 37139 6953 37151 6956
rect 37093 6947 37151 6953
rect 38102 6944 38108 6956
rect 38160 6944 38166 6996
rect 38194 6944 38200 6996
rect 38252 6984 38258 6996
rect 46385 6987 46443 6993
rect 38252 6956 38516 6984
rect 38252 6944 38258 6956
rect 33686 6876 33692 6928
rect 33744 6916 33750 6928
rect 33744 6888 34192 6916
rect 33744 6876 33750 6888
rect 34164 6860 34192 6888
rect 27890 6848 27896 6860
rect 27816 6820 27896 6848
rect 25950 6811 26008 6817
rect 27890 6808 27896 6820
rect 27948 6848 27954 6860
rect 27985 6851 28043 6857
rect 27985 6848 27997 6851
rect 27948 6820 27997 6848
rect 27948 6808 27954 6820
rect 27985 6817 27997 6820
rect 28031 6848 28043 6851
rect 28031 6820 28120 6848
rect 28031 6817 28043 6820
rect 27985 6811 28043 6817
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2130 6780 2136 6792
rect 2087 6752 2136 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2130 6740 2136 6752
rect 2188 6780 2194 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 2188 6752 4905 6780
rect 2188 6740 2194 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 5160 6783 5218 6789
rect 5160 6749 5172 6783
rect 5206 6749 5218 6783
rect 5160 6743 5218 6749
rect 2308 6715 2366 6721
rect 2308 6681 2320 6715
rect 2354 6712 2366 6715
rect 2958 6712 2964 6724
rect 2354 6684 2964 6712
rect 2354 6681 2366 6684
rect 2308 6675 2366 6681
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 3786 6604 3792 6656
rect 3844 6604 3850 6656
rect 4154 6604 4160 6656
rect 4212 6604 4218 6656
rect 4246 6604 4252 6656
rect 4304 6604 4310 6656
rect 4908 6644 4936 6743
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5184 6712 5212 6743
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 7708 6752 8401 6780
rect 7708 6740 7714 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 10778 6740 10784 6792
rect 10836 6740 10842 6792
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12400 6752 12541 6780
rect 12400 6740 12406 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12728 6752 14320 6780
rect 6380 6712 6408 6740
rect 5132 6684 5212 6712
rect 5276 6684 6408 6712
rect 6632 6715 6690 6721
rect 5132 6672 5138 6684
rect 5276 6644 5304 6684
rect 6632 6681 6644 6715
rect 6678 6712 6690 6715
rect 7837 6715 7895 6721
rect 7837 6712 7849 6715
rect 6678 6684 7849 6712
rect 6678 6681 6690 6684
rect 6632 6675 6690 6681
rect 7837 6681 7849 6684
rect 7883 6681 7895 6715
rect 7837 6675 7895 6681
rect 9030 6672 9036 6724
rect 9088 6712 9094 6724
rect 9585 6715 9643 6721
rect 9585 6712 9597 6715
rect 9088 6684 9597 6712
rect 9088 6672 9094 6684
rect 9585 6681 9597 6684
rect 9631 6712 9643 6715
rect 12728 6712 12756 6752
rect 12802 6721 12808 6724
rect 9631 6684 12756 6712
rect 9631 6681 9643 6684
rect 9585 6675 9643 6681
rect 12796 6675 12808 6721
rect 12802 6672 12808 6675
rect 12860 6672 12866 6724
rect 4908 6616 5304 6644
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 7742 6604 7748 6656
rect 7800 6604 7806 6656
rect 10134 6604 10140 6656
rect 10192 6604 10198 6656
rect 10870 6604 10876 6656
rect 10928 6604 10934 6656
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 13170 6644 13176 6656
rect 12483 6616 13176 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 14182 6604 14188 6656
rect 14240 6604 14246 6656
rect 14292 6644 14320 6752
rect 14826 6740 14832 6792
rect 14884 6740 14890 6792
rect 14918 6740 14924 6792
rect 14976 6789 14982 6792
rect 14976 6783 15025 6789
rect 14976 6749 14979 6783
rect 15013 6749 15025 6783
rect 14976 6743 15025 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16206 6780 16212 6792
rect 16163 6752 16212 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 14976 6740 14982 6743
rect 15194 6644 15200 6656
rect 14292 6616 15200 6644
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15856 6644 15884 6743
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 18138 6740 18144 6792
rect 18196 6740 18202 6792
rect 20533 6783 20591 6789
rect 20533 6749 20545 6783
rect 20579 6780 20591 6783
rect 20714 6780 20720 6792
rect 20579 6752 20720 6780
rect 20579 6749 20591 6752
rect 20533 6743 20591 6749
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 20916 6752 21557 6780
rect 16384 6715 16442 6721
rect 16384 6681 16396 6715
rect 16430 6712 16442 6715
rect 17589 6715 17647 6721
rect 17589 6712 17601 6715
rect 16430 6684 17601 6712
rect 16430 6681 16442 6684
rect 16384 6675 16442 6681
rect 17589 6681 17601 6684
rect 17635 6681 17647 6715
rect 17589 6675 17647 6681
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 20441 6715 20499 6721
rect 20441 6712 20453 6715
rect 19668 6684 20453 6712
rect 19668 6672 19674 6684
rect 20441 6681 20453 6684
rect 20487 6681 20499 6715
rect 20441 6675 20499 6681
rect 17034 6644 17040 6656
rect 15856 6616 17040 6644
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 19518 6604 19524 6656
rect 19576 6644 19582 6656
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 19576 6616 19809 6644
rect 19576 6604 19582 6616
rect 19797 6613 19809 6616
rect 19843 6644 19855 6647
rect 19886 6644 19892 6656
rect 19843 6616 19892 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 20916 6653 20944 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 21545 6743 21603 6749
rect 23860 6752 24409 6780
rect 21913 6715 21971 6721
rect 21913 6681 21925 6715
rect 21959 6712 21971 6715
rect 22462 6712 22468 6724
rect 21959 6684 22468 6712
rect 21959 6681 21971 6684
rect 21913 6675 21971 6681
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 22732 6715 22790 6721
rect 22732 6681 22744 6715
rect 22778 6712 22790 6715
rect 22922 6712 22928 6724
rect 22778 6684 22928 6712
rect 22778 6681 22790 6684
rect 22732 6675 22790 6681
rect 22922 6672 22928 6684
rect 22980 6672 22986 6724
rect 23860 6653 23888 6752
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 26050 6780 26056 6792
rect 24397 6743 24455 6749
rect 25240 6752 26056 6780
rect 25130 6712 25136 6724
rect 24228 6684 25136 6712
rect 20901 6647 20959 6653
rect 20901 6613 20913 6647
rect 20947 6613 20959 6647
rect 20901 6607 20959 6613
rect 23845 6647 23903 6653
rect 23845 6613 23857 6647
rect 23891 6613 23903 6647
rect 23845 6607 23903 6613
rect 23934 6604 23940 6656
rect 23992 6644 23998 6656
rect 24228 6653 24256 6684
rect 25130 6672 25136 6684
rect 25188 6712 25194 6724
rect 25240 6712 25268 6752
rect 26050 6740 26056 6752
rect 26108 6740 26114 6792
rect 28092 6780 28120 6820
rect 33962 6808 33968 6860
rect 34020 6808 34026 6860
rect 34146 6808 34152 6860
rect 34204 6808 34210 6860
rect 36446 6808 36452 6860
rect 36504 6848 36510 6860
rect 36814 6848 36820 6860
rect 36504 6820 36820 6848
rect 36504 6808 36510 6820
rect 36814 6808 36820 6820
rect 36872 6808 36878 6860
rect 38488 6848 38516 6956
rect 46385 6953 46397 6987
rect 46431 6984 46443 6987
rect 46658 6984 46664 6996
rect 46431 6956 46664 6984
rect 46431 6953 46443 6956
rect 46385 6947 46443 6953
rect 46658 6944 46664 6956
rect 46716 6944 46722 6996
rect 52549 6987 52607 6993
rect 52549 6953 52561 6987
rect 52595 6984 52607 6987
rect 53282 6984 53288 6996
rect 52595 6956 53288 6984
rect 52595 6953 52607 6956
rect 52549 6947 52607 6953
rect 53282 6944 53288 6956
rect 53340 6944 53346 6996
rect 55950 6944 55956 6996
rect 56008 6984 56014 6996
rect 56045 6987 56103 6993
rect 56045 6984 56057 6987
rect 56008 6956 56057 6984
rect 56008 6944 56014 6956
rect 56045 6953 56057 6956
rect 56091 6953 56103 6987
rect 56045 6947 56103 6953
rect 41693 6919 41751 6925
rect 41693 6885 41705 6919
rect 41739 6916 41751 6919
rect 41782 6916 41788 6928
rect 41739 6888 41788 6916
rect 41739 6885 41751 6888
rect 41693 6879 41751 6885
rect 41782 6876 41788 6888
rect 41840 6876 41846 6928
rect 51166 6876 51172 6928
rect 51224 6916 51230 6928
rect 51261 6919 51319 6925
rect 51261 6916 51273 6919
rect 51224 6888 51273 6916
rect 51224 6876 51230 6888
rect 51261 6885 51273 6888
rect 51307 6885 51319 6919
rect 51261 6879 51319 6885
rect 38657 6851 38715 6857
rect 38657 6848 38669 6851
rect 38488 6820 38669 6848
rect 38657 6817 38669 6820
rect 38703 6817 38715 6851
rect 38657 6811 38715 6817
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 28092 6752 29561 6780
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 31573 6783 31631 6789
rect 31573 6780 31585 6783
rect 29549 6743 29607 6749
rect 30944 6752 31585 6780
rect 25188 6684 25268 6712
rect 25188 6672 25194 6684
rect 25314 6672 25320 6724
rect 25372 6672 25378 6724
rect 26228 6715 26286 6721
rect 26228 6681 26240 6715
rect 26274 6712 26286 6715
rect 26970 6712 26976 6724
rect 26274 6684 26976 6712
rect 26274 6681 26286 6684
rect 26228 6675 26286 6681
rect 26970 6672 26976 6684
rect 27028 6672 27034 6724
rect 28258 6721 28264 6724
rect 28252 6675 28264 6721
rect 28258 6672 28264 6675
rect 28316 6672 28322 6724
rect 28350 6672 28356 6724
rect 28408 6672 28414 6724
rect 29454 6672 29460 6724
rect 29512 6712 29518 6724
rect 29794 6715 29852 6721
rect 29794 6712 29806 6715
rect 29512 6684 29806 6712
rect 29512 6672 29518 6684
rect 29794 6681 29806 6684
rect 29840 6681 29852 6715
rect 29794 6675 29852 6681
rect 24213 6647 24271 6653
rect 24213 6644 24225 6647
rect 23992 6616 24225 6644
rect 23992 6604 23998 6616
rect 24213 6613 24225 6616
rect 24259 6613 24271 6647
rect 24213 6607 24271 6613
rect 24394 6604 24400 6656
rect 24452 6644 24458 6656
rect 26326 6644 26332 6656
rect 24452 6616 26332 6644
rect 24452 6604 24458 6616
rect 26326 6604 26332 6616
rect 26384 6604 26390 6656
rect 27341 6647 27399 6653
rect 27341 6613 27353 6647
rect 27387 6644 27399 6647
rect 28368 6644 28396 6672
rect 30944 6653 30972 6752
rect 31573 6749 31585 6752
rect 31619 6749 31631 6783
rect 31573 6743 31631 6749
rect 32033 6783 32091 6789
rect 32033 6749 32045 6783
rect 32079 6780 32091 6783
rect 32122 6780 32128 6792
rect 32079 6752 32128 6780
rect 32079 6749 32091 6752
rect 32033 6743 32091 6749
rect 32122 6740 32128 6752
rect 32180 6780 32186 6792
rect 34514 6780 34520 6792
rect 32180 6752 34520 6780
rect 32180 6740 32186 6752
rect 34514 6740 34520 6752
rect 34572 6780 34578 6792
rect 34701 6783 34759 6789
rect 34701 6780 34713 6783
rect 34572 6752 34713 6780
rect 34572 6740 34578 6752
rect 34701 6749 34713 6752
rect 34747 6780 34759 6783
rect 37642 6780 37648 6792
rect 34747 6752 37648 6780
rect 34747 6749 34759 6752
rect 34701 6743 34759 6749
rect 37642 6740 37648 6752
rect 37700 6780 37706 6792
rect 38473 6783 38531 6789
rect 38473 6780 38485 6783
rect 37700 6752 38485 6780
rect 37700 6740 37706 6752
rect 38473 6749 38485 6752
rect 38519 6749 38531 6783
rect 38473 6743 38531 6749
rect 32300 6715 32358 6721
rect 32300 6681 32312 6715
rect 32346 6712 32358 6715
rect 32582 6712 32588 6724
rect 32346 6684 32588 6712
rect 32346 6681 32358 6684
rect 32300 6675 32358 6681
rect 32582 6672 32588 6684
rect 32640 6672 32646 6724
rect 34968 6715 35026 6721
rect 34968 6681 34980 6715
rect 35014 6712 35026 6715
rect 36262 6712 36268 6724
rect 35014 6684 36268 6712
rect 35014 6681 35026 6684
rect 34968 6675 35026 6681
rect 36262 6672 36268 6684
rect 36320 6672 36326 6724
rect 37550 6712 37556 6724
rect 36464 6684 37556 6712
rect 27387 6616 28396 6644
rect 30929 6647 30987 6653
rect 27387 6613 27399 6616
rect 27341 6607 27399 6613
rect 30929 6613 30941 6647
rect 30975 6613 30987 6647
rect 30929 6607 30987 6613
rect 31018 6604 31024 6656
rect 31076 6604 31082 6656
rect 33502 6604 33508 6656
rect 33560 6604 33566 6656
rect 33870 6604 33876 6656
rect 33928 6604 33934 6656
rect 36081 6647 36139 6653
rect 36081 6613 36093 6647
rect 36127 6644 36139 6647
rect 36464 6644 36492 6684
rect 37550 6672 37556 6684
rect 37608 6672 37614 6724
rect 38010 6672 38016 6724
rect 38068 6672 38074 6724
rect 38228 6715 38286 6721
rect 38228 6681 38240 6715
rect 38274 6712 38286 6715
rect 38562 6712 38568 6724
rect 38274 6684 38568 6712
rect 38274 6681 38286 6684
rect 38228 6675 38286 6681
rect 38562 6672 38568 6684
rect 38620 6672 38626 6724
rect 38672 6712 38700 6811
rect 38746 6808 38752 6860
rect 38804 6848 38810 6860
rect 38841 6851 38899 6857
rect 38841 6848 38853 6851
rect 38804 6820 38853 6848
rect 38804 6808 38810 6820
rect 38841 6817 38853 6820
rect 38887 6817 38899 6851
rect 43165 6851 43223 6857
rect 43165 6848 43177 6851
rect 38841 6811 38899 6817
rect 41386 6820 43177 6848
rect 38930 6740 38936 6792
rect 38988 6780 38994 6792
rect 39850 6780 39856 6792
rect 38988 6752 39856 6780
rect 38988 6740 38994 6752
rect 39850 6740 39856 6752
rect 39908 6780 39914 6792
rect 40037 6783 40095 6789
rect 40037 6780 40049 6783
rect 39908 6752 40049 6780
rect 39908 6740 39914 6752
rect 40037 6749 40049 6752
rect 40083 6749 40095 6783
rect 40037 6743 40095 6749
rect 40313 6783 40371 6789
rect 40313 6749 40325 6783
rect 40359 6780 40371 6783
rect 40954 6780 40960 6792
rect 40359 6752 40960 6780
rect 40359 6749 40371 6752
rect 40313 6743 40371 6749
rect 40954 6740 40960 6752
rect 41012 6780 41018 6792
rect 41386 6780 41414 6820
rect 43165 6817 43177 6820
rect 43211 6817 43223 6851
rect 43165 6811 43223 6817
rect 46569 6851 46627 6857
rect 46569 6817 46581 6851
rect 46615 6848 46627 6851
rect 46934 6848 46940 6860
rect 46615 6820 46940 6848
rect 46615 6817 46627 6820
rect 46569 6811 46627 6817
rect 41012 6752 41414 6780
rect 41012 6740 41018 6752
rect 41690 6740 41696 6792
rect 41748 6780 41754 6792
rect 42337 6783 42395 6789
rect 42337 6780 42349 6783
rect 41748 6752 42349 6780
rect 41748 6740 41754 6752
rect 42337 6749 42349 6752
rect 42383 6749 42395 6783
rect 43180 6780 43208 6811
rect 46934 6808 46940 6820
rect 46992 6808 46998 6860
rect 47118 6808 47124 6860
rect 47176 6848 47182 6860
rect 47213 6851 47271 6857
rect 47213 6848 47225 6851
rect 47176 6820 47225 6848
rect 47176 6808 47182 6820
rect 47213 6817 47225 6820
rect 47259 6817 47271 6851
rect 47213 6811 47271 6817
rect 47486 6808 47492 6860
rect 47544 6808 47550 6860
rect 47603 6808 47609 6860
rect 47661 6808 47667 6860
rect 48406 6808 48412 6860
rect 48464 6848 48470 6860
rect 48961 6851 49019 6857
rect 48961 6848 48973 6851
rect 48464 6820 48973 6848
rect 48464 6808 48470 6820
rect 48961 6817 48973 6820
rect 49007 6817 49019 6851
rect 48961 6811 49019 6817
rect 49050 6808 49056 6860
rect 49108 6808 49114 6860
rect 50614 6808 50620 6860
rect 50672 6857 50678 6860
rect 50672 6851 50721 6857
rect 50672 6817 50675 6851
rect 50709 6817 50721 6851
rect 50672 6811 50721 6817
rect 50672 6808 50678 6811
rect 51350 6808 51356 6860
rect 51408 6848 51414 6860
rect 51537 6851 51595 6857
rect 51537 6848 51549 6851
rect 51408 6820 51549 6848
rect 51408 6808 51414 6820
rect 51537 6817 51549 6820
rect 51583 6817 51595 6851
rect 51537 6811 51595 6817
rect 51813 6851 51871 6857
rect 51813 6817 51825 6851
rect 51859 6848 51871 6851
rect 52178 6848 52184 6860
rect 51859 6820 52184 6848
rect 51859 6817 51871 6820
rect 51813 6811 51871 6817
rect 52178 6808 52184 6820
rect 52236 6808 52242 6860
rect 54018 6808 54024 6860
rect 54076 6848 54082 6860
rect 54113 6851 54171 6857
rect 54113 6848 54125 6851
rect 54076 6820 54125 6848
rect 54076 6808 54082 6820
rect 54113 6817 54125 6820
rect 54159 6848 54171 6851
rect 55033 6851 55091 6857
rect 55033 6848 55045 6851
rect 54159 6820 55045 6848
rect 54159 6817 54171 6820
rect 54113 6811 54171 6817
rect 55033 6817 55045 6820
rect 55079 6817 55091 6851
rect 55033 6811 55091 6817
rect 55493 6851 55551 6857
rect 55493 6817 55505 6851
rect 55539 6848 55551 6851
rect 55582 6848 55588 6860
rect 55539 6820 55588 6848
rect 55539 6817 55551 6820
rect 55493 6811 55551 6817
rect 55582 6808 55588 6820
rect 55640 6808 55646 6860
rect 45002 6780 45008 6792
rect 43180 6752 45008 6780
rect 42337 6743 42395 6749
rect 45002 6740 45008 6752
rect 45060 6740 45066 6792
rect 45272 6783 45330 6789
rect 45272 6749 45284 6783
rect 45318 6780 45330 6783
rect 45554 6780 45560 6792
rect 45318 6752 45560 6780
rect 45318 6749 45330 6752
rect 45272 6743 45330 6749
rect 45554 6740 45560 6752
rect 45612 6740 45618 6792
rect 46750 6740 46756 6792
rect 46808 6740 46814 6792
rect 47762 6740 47768 6792
rect 47820 6740 47826 6792
rect 48332 6752 49924 6780
rect 40580 6715 40638 6721
rect 38672 6684 39712 6712
rect 36127 6616 36492 6644
rect 36127 6613 36139 6616
rect 36081 6607 36139 6613
rect 36538 6604 36544 6656
rect 36596 6604 36602 6656
rect 36633 6647 36691 6653
rect 36633 6613 36645 6647
rect 36679 6644 36691 6647
rect 36722 6644 36728 6656
rect 36679 6616 36728 6644
rect 36679 6613 36691 6616
rect 36633 6607 36691 6613
rect 36722 6604 36728 6616
rect 36780 6604 36786 6656
rect 36814 6604 36820 6656
rect 36872 6644 36878 6656
rect 38028 6644 38056 6672
rect 36872 6616 38056 6644
rect 36872 6604 36878 6616
rect 38102 6604 38108 6656
rect 38160 6644 38166 6656
rect 38654 6644 38660 6656
rect 38160 6616 38660 6644
rect 38160 6604 38166 6616
rect 38654 6604 38660 6616
rect 38712 6644 38718 6656
rect 38933 6647 38991 6653
rect 38933 6644 38945 6647
rect 38712 6616 38945 6644
rect 38712 6604 38718 6616
rect 38933 6613 38945 6616
rect 38979 6613 38991 6647
rect 38933 6607 38991 6613
rect 39301 6647 39359 6653
rect 39301 6613 39313 6647
rect 39347 6644 39359 6647
rect 39390 6644 39396 6656
rect 39347 6616 39396 6644
rect 39347 6613 39359 6616
rect 39301 6607 39359 6613
rect 39390 6604 39396 6616
rect 39448 6604 39454 6656
rect 39684 6653 39712 6684
rect 40580 6681 40592 6715
rect 40626 6712 40638 6715
rect 41785 6715 41843 6721
rect 41785 6712 41797 6715
rect 40626 6684 41797 6712
rect 40626 6681 40638 6684
rect 40580 6675 40638 6681
rect 41785 6681 41797 6684
rect 41831 6681 41843 6715
rect 41785 6675 41843 6681
rect 43432 6715 43490 6721
rect 43432 6681 43444 6715
rect 43478 6712 43490 6715
rect 43898 6712 43904 6724
rect 43478 6684 43904 6712
rect 43478 6681 43490 6684
rect 43432 6675 43490 6681
rect 43898 6672 43904 6684
rect 43956 6672 43962 6724
rect 43990 6672 43996 6724
rect 44048 6712 44054 6724
rect 48332 6712 48360 6752
rect 44048 6684 46796 6712
rect 44048 6672 44054 6684
rect 39669 6647 39727 6653
rect 39669 6613 39681 6647
rect 39715 6644 39727 6647
rect 43254 6644 43260 6656
rect 39715 6616 43260 6644
rect 39715 6613 39727 6616
rect 39669 6607 39727 6613
rect 43254 6604 43260 6616
rect 43312 6604 43318 6656
rect 44545 6647 44603 6653
rect 44545 6613 44557 6647
rect 44591 6644 44603 6647
rect 45738 6644 45744 6656
rect 44591 6616 45744 6644
rect 44591 6613 44603 6616
rect 44545 6607 44603 6613
rect 45738 6604 45744 6616
rect 45796 6604 45802 6656
rect 46768 6644 46796 6684
rect 48240 6684 48360 6712
rect 48409 6715 48467 6721
rect 47118 6644 47124 6656
rect 46768 6616 47124 6644
rect 47118 6604 47124 6616
rect 47176 6644 47182 6656
rect 48240 6644 48268 6684
rect 48409 6681 48421 6715
rect 48455 6712 48467 6715
rect 48869 6715 48927 6721
rect 48869 6712 48881 6715
rect 48455 6684 48881 6712
rect 48455 6681 48467 6684
rect 48409 6675 48467 6681
rect 48869 6681 48881 6684
rect 48915 6681 48927 6715
rect 48869 6675 48927 6681
rect 49896 6656 49924 6752
rect 49970 6740 49976 6792
rect 50028 6740 50034 6792
rect 50798 6740 50804 6792
rect 50856 6740 50862 6792
rect 51718 6789 51724 6792
rect 51675 6783 51724 6789
rect 51675 6749 51687 6783
rect 51721 6749 51724 6783
rect 51675 6743 51724 6749
rect 51718 6740 51724 6743
rect 51776 6740 51782 6792
rect 53834 6740 53840 6792
rect 53892 6780 53898 6792
rect 53929 6783 53987 6789
rect 53929 6780 53941 6783
rect 53892 6752 53941 6780
rect 53892 6740 53898 6752
rect 53929 6749 53941 6752
rect 53975 6749 53987 6783
rect 53929 6743 53987 6749
rect 54297 6783 54355 6789
rect 54297 6749 54309 6783
rect 54343 6780 54355 6783
rect 54343 6752 55168 6780
rect 54343 6749 54355 6752
rect 54297 6743 54355 6749
rect 53684 6715 53742 6721
rect 53684 6681 53696 6715
rect 53730 6712 53742 6715
rect 54202 6712 54208 6724
rect 53730 6684 54208 6712
rect 53730 6681 53742 6684
rect 53684 6675 53742 6681
rect 54202 6672 54208 6684
rect 54260 6672 54266 6724
rect 47176 6616 48268 6644
rect 47176 6604 47182 6616
rect 48314 6604 48320 6656
rect 48372 6644 48378 6656
rect 48501 6647 48559 6653
rect 48501 6644 48513 6647
rect 48372 6616 48513 6644
rect 48372 6604 48378 6616
rect 48501 6613 48513 6616
rect 48547 6613 48559 6647
rect 48501 6607 48559 6613
rect 49329 6647 49387 6653
rect 49329 6613 49341 6647
rect 49375 6644 49387 6647
rect 49418 6644 49424 6656
rect 49375 6616 49424 6644
rect 49375 6613 49387 6616
rect 49329 6607 49387 6613
rect 49418 6604 49424 6616
rect 49476 6604 49482 6656
rect 49878 6604 49884 6656
rect 49936 6644 49942 6656
rect 50433 6647 50491 6653
rect 50433 6644 50445 6647
rect 49936 6616 50445 6644
rect 49936 6604 49942 6616
rect 50433 6613 50445 6616
rect 50479 6644 50491 6647
rect 51166 6644 51172 6656
rect 50479 6616 51172 6644
rect 50479 6613 50491 6616
rect 50433 6607 50491 6613
rect 51166 6604 51172 6616
rect 51224 6604 51230 6656
rect 52454 6604 52460 6656
rect 52512 6604 52518 6656
rect 54386 6604 54392 6656
rect 54444 6604 54450 6656
rect 54570 6604 54576 6656
rect 54628 6644 54634 6656
rect 54757 6647 54815 6653
rect 54757 6644 54769 6647
rect 54628 6616 54769 6644
rect 54628 6604 54634 6616
rect 54757 6613 54769 6616
rect 54803 6613 54815 6647
rect 55140 6644 55168 6752
rect 56134 6740 56140 6792
rect 56192 6780 56198 6792
rect 56410 6780 56416 6792
rect 56192 6752 56416 6780
rect 56192 6740 56198 6752
rect 56410 6740 56416 6752
rect 56468 6740 56474 6792
rect 57422 6740 57428 6792
rect 57480 6780 57486 6792
rect 58437 6783 58495 6789
rect 58437 6780 58449 6783
rect 57480 6752 58449 6780
rect 57480 6740 57486 6752
rect 58437 6749 58449 6752
rect 58483 6749 58495 6783
rect 58437 6743 58495 6749
rect 55585 6715 55643 6721
rect 55585 6681 55597 6715
rect 55631 6712 55643 6715
rect 56502 6712 56508 6724
rect 55631 6684 56508 6712
rect 55631 6681 55643 6684
rect 55585 6675 55643 6681
rect 56502 6672 56508 6684
rect 56560 6672 56566 6724
rect 56680 6715 56738 6721
rect 56680 6681 56692 6715
rect 56726 6712 56738 6715
rect 57885 6715 57943 6721
rect 57885 6712 57897 6715
rect 56726 6684 57897 6712
rect 56726 6681 56738 6684
rect 56680 6675 56738 6681
rect 57885 6681 57897 6684
rect 57931 6681 57943 6715
rect 57885 6675 57943 6681
rect 55214 6644 55220 6656
rect 55140 6616 55220 6644
rect 54757 6607 54815 6613
rect 55214 6604 55220 6616
rect 55272 6644 55278 6656
rect 55677 6647 55735 6653
rect 55677 6644 55689 6647
rect 55272 6616 55689 6644
rect 55272 6604 55278 6616
rect 55677 6613 55689 6616
rect 55723 6644 55735 6647
rect 57054 6644 57060 6656
rect 55723 6616 57060 6644
rect 55723 6613 55735 6616
rect 55677 6607 55735 6613
rect 57054 6604 57060 6616
rect 57112 6604 57118 6656
rect 57790 6604 57796 6656
rect 57848 6604 57854 6656
rect 1104 6554 59040 6576
rect 1104 6502 15394 6554
rect 15446 6502 15458 6554
rect 15510 6502 15522 6554
rect 15574 6502 15586 6554
rect 15638 6502 15650 6554
rect 15702 6502 29838 6554
rect 29890 6502 29902 6554
rect 29954 6502 29966 6554
rect 30018 6502 30030 6554
rect 30082 6502 30094 6554
rect 30146 6502 44282 6554
rect 44334 6502 44346 6554
rect 44398 6502 44410 6554
rect 44462 6502 44474 6554
rect 44526 6502 44538 6554
rect 44590 6502 58726 6554
rect 58778 6502 58790 6554
rect 58842 6502 58854 6554
rect 58906 6502 58918 6554
rect 58970 6502 58982 6554
rect 59034 6502 59040 6554
rect 1104 6480 59040 6502
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 4212 6412 4537 6440
rect 4212 6400 4218 6412
rect 4525 6409 4537 6412
rect 4571 6440 4583 6443
rect 5166 6440 5172 6452
rect 4571 6412 5172 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 7098 6440 7104 6452
rect 6227 6412 7104 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7282 6400 7288 6452
rect 7340 6400 7346 6452
rect 7650 6400 7656 6452
rect 7708 6400 7714 6452
rect 7742 6400 7748 6452
rect 7800 6400 7806 6452
rect 10134 6400 10140 6452
rect 10192 6400 10198 6452
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6440 11115 6443
rect 11422 6440 11428 6452
rect 11103 6412 11428 6440
rect 11103 6409 11115 6412
rect 11057 6403 11115 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12802 6440 12808 6452
rect 12667 6412 12808 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13170 6400 13176 6452
rect 13228 6400 13234 6452
rect 13998 6440 14004 6452
rect 13740 6412 14004 6440
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 4338 6372 4344 6384
rect 2731 6344 4344 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 3786 6264 3792 6316
rect 3844 6264 3850 6316
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6564 6276 7205 6304
rect 6564 6248 6592 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 2314 6196 2320 6248
rect 2372 6196 2378 6248
rect 4062 6236 4068 6248
rect 2976 6208 4068 6236
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 2976 6168 3004 6208
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 6546 6196 6552 6248
rect 6604 6196 6610 6248
rect 7098 6196 7104 6248
rect 7156 6196 7162 6248
rect 7300 6236 7328 6400
rect 7760 6304 7788 6400
rect 9944 6375 10002 6381
rect 9944 6341 9956 6375
rect 9990 6372 10002 6375
rect 10152 6372 10180 6400
rect 9990 6344 10180 6372
rect 13081 6375 13139 6381
rect 9990 6341 10002 6344
rect 9944 6335 10002 6341
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13740 6372 13768 6412
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 16117 6443 16175 6449
rect 16117 6440 16129 6443
rect 14240 6412 16129 6440
rect 14240 6400 14246 6412
rect 16117 6409 16129 6412
rect 16163 6409 16175 6443
rect 16117 6403 16175 6409
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16908 6412 16957 6440
rect 16908 6400 16914 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 16945 6403 17003 6409
rect 17034 6400 17040 6452
rect 17092 6400 17098 6452
rect 17405 6443 17463 6449
rect 17405 6409 17417 6443
rect 17451 6440 17463 6443
rect 18138 6440 18144 6452
rect 17451 6412 18144 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 19242 6400 19248 6452
rect 19300 6400 19306 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 20441 6443 20499 6449
rect 20441 6440 20453 6443
rect 20312 6412 20453 6440
rect 20312 6400 20318 6412
rect 20441 6409 20453 6412
rect 20487 6409 20499 6443
rect 20441 6403 20499 6409
rect 22922 6400 22928 6452
rect 22980 6400 22986 6452
rect 24857 6443 24915 6449
rect 24857 6409 24869 6443
rect 24903 6440 24915 6443
rect 25590 6440 25596 6452
rect 24903 6412 25596 6440
rect 24903 6409 24915 6412
rect 24857 6403 24915 6409
rect 25590 6400 25596 6412
rect 25648 6400 25654 6452
rect 25869 6443 25927 6449
rect 25869 6409 25881 6443
rect 25915 6440 25927 6443
rect 26142 6440 26148 6452
rect 25915 6412 26148 6440
rect 25915 6409 25927 6412
rect 25869 6403 25927 6409
rect 13127 6344 13768 6372
rect 13808 6375 13866 6381
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13808 6341 13820 6375
rect 13854 6372 13866 6375
rect 14090 6372 14096 6384
rect 13854 6344 14096 6372
rect 13854 6341 13866 6344
rect 13808 6335 13866 6341
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 15746 6332 15752 6384
rect 15804 6372 15810 6384
rect 16209 6375 16267 6381
rect 16209 6372 16221 6375
rect 15804 6344 16221 6372
rect 15804 6332 15810 6344
rect 16209 6341 16221 6344
rect 16255 6341 16267 6375
rect 16209 6335 16267 6341
rect 17957 6375 18015 6381
rect 17957 6341 17969 6375
rect 18003 6372 18015 6375
rect 19260 6372 19288 6400
rect 18003 6344 19288 6372
rect 18003 6341 18015 6344
rect 17957 6335 18015 6341
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 7760 6276 8309 6304
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 12526 6304 12532 6316
rect 12115 6276 12532 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 15197 6307 15255 6313
rect 15197 6304 15209 6307
rect 13188 6276 15209 6304
rect 7745 6239 7803 6245
rect 7745 6236 7757 6239
rect 7300 6208 7757 6236
rect 7745 6205 7757 6208
rect 7791 6205 7803 6239
rect 7745 6199 7803 6205
rect 9214 6196 9220 6248
rect 9272 6196 9278 6248
rect 11900 6236 11928 6264
rect 13188 6236 13216 6276
rect 15197 6273 15209 6276
rect 15243 6273 15255 6307
rect 20714 6304 20720 6316
rect 15197 6267 15255 6273
rect 16316 6276 20720 6304
rect 11900 6208 13216 6236
rect 13262 6196 13268 6248
rect 13320 6196 13326 6248
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6205 13599 6239
rect 15212 6236 15240 6267
rect 16316 6245 16344 6276
rect 20714 6264 20720 6276
rect 20772 6304 20778 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20772 6276 20821 6304
rect 20772 6264 20778 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 23474 6264 23480 6316
rect 23532 6264 23538 6316
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15212 6208 16313 6236
rect 13541 6199 13599 6205
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 4985 6171 5043 6177
rect 4985 6168 4997 6171
rect 1995 6140 3004 6168
rect 3252 6140 4997 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2961 6103 3019 6109
rect 2961 6100 2973 6103
rect 1912 6072 2973 6100
rect 1912 6060 1918 6072
rect 2961 6069 2973 6072
rect 3007 6100 3019 6103
rect 3252 6100 3280 6140
rect 4985 6137 4997 6140
rect 5031 6168 5043 6171
rect 5353 6171 5411 6177
rect 5353 6168 5365 6171
rect 5031 6140 5365 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 5353 6137 5365 6140
rect 5399 6168 5411 6171
rect 6362 6168 6368 6180
rect 5399 6140 6368 6168
rect 5399 6137 5411 6140
rect 5353 6131 5411 6137
rect 6362 6128 6368 6140
rect 6420 6168 6426 6180
rect 6733 6171 6791 6177
rect 6733 6168 6745 6171
rect 6420 6140 6745 6168
rect 6420 6128 6426 6140
rect 6733 6137 6745 6140
rect 6779 6137 6791 6171
rect 13556 6168 13584 6199
rect 6733 6131 6791 6137
rect 12544 6140 13584 6168
rect 14921 6171 14979 6177
rect 12544 6112 12572 6140
rect 14921 6137 14933 6171
rect 14967 6168 14979 6171
rect 15010 6168 15016 6180
rect 14967 6140 15016 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 16482 6168 16488 6180
rect 15580 6140 16488 6168
rect 3007 6072 3280 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 4614 6100 4620 6112
rect 3384 6072 4620 6100
rect 3384 6060 3390 6072
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6100 5871 6103
rect 5902 6100 5908 6112
rect 5859 6072 5908 6100
rect 5859 6069 5871 6072
rect 5813 6063 5871 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 8662 6060 8668 6112
rect 8720 6060 8726 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 11790 6100 11796 6112
rect 9548 6072 11796 6100
rect 9548 6060 9554 6072
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6100 11943 6103
rect 12342 6100 12348 6112
rect 11931 6072 12348 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 12342 6060 12348 6072
rect 12400 6100 12406 6112
rect 12526 6100 12532 6112
rect 12400 6072 12532 6100
rect 12400 6060 12406 6072
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 12713 6103 12771 6109
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 12802 6100 12808 6112
rect 12759 6072 12808 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 15580 6109 15608 6140
rect 16482 6128 16488 6140
rect 16540 6168 16546 6180
rect 16776 6168 16804 6199
rect 18046 6196 18052 6248
rect 18104 6196 18110 6248
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 18196 6208 18797 6236
rect 18196 6196 18202 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 19300 6208 20085 6236
rect 19300 6196 19306 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 21910 6236 21916 6248
rect 20073 6199 20131 6205
rect 21192 6208 21916 6236
rect 19521 6171 19579 6177
rect 19521 6168 19533 6171
rect 16540 6140 16804 6168
rect 19352 6140 19533 6168
rect 16540 6128 16546 6140
rect 19352 6112 19380 6140
rect 19521 6137 19533 6140
rect 19567 6137 19579 6171
rect 19521 6131 19579 6137
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 13412 6072 15577 6100
rect 13412 6060 13418 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 15746 6060 15752 6112
rect 15804 6060 15810 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18782 6100 18788 6112
rect 18739 6072 18788 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 19334 6060 19340 6112
rect 19392 6060 19398 6112
rect 19426 6060 19432 6112
rect 19484 6060 19490 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 21192 6100 21220 6208
rect 21910 6196 21916 6208
rect 21968 6236 21974 6248
rect 21968 6208 23888 6236
rect 21968 6196 21974 6208
rect 21269 6171 21327 6177
rect 21269 6137 21281 6171
rect 21315 6168 21327 6171
rect 23860 6168 23888 6208
rect 23934 6196 23940 6248
rect 23992 6236 23998 6248
rect 26068 6245 26096 6412
rect 26142 6400 26148 6412
rect 26200 6400 26206 6452
rect 26237 6443 26295 6449
rect 26237 6409 26249 6443
rect 26283 6440 26295 6443
rect 26418 6440 26424 6452
rect 26283 6412 26424 6440
rect 26283 6409 26295 6412
rect 26237 6403 26295 6409
rect 26418 6400 26424 6412
rect 26476 6400 26482 6452
rect 26697 6443 26755 6449
rect 26697 6409 26709 6443
rect 26743 6440 26755 6443
rect 26878 6440 26884 6452
rect 26743 6412 26884 6440
rect 26743 6409 26755 6412
rect 26697 6403 26755 6409
rect 26878 6400 26884 6412
rect 26936 6400 26942 6452
rect 26970 6400 26976 6452
rect 27028 6400 27034 6452
rect 27890 6400 27896 6452
rect 27948 6400 27954 6452
rect 28169 6443 28227 6449
rect 28169 6409 28181 6443
rect 28215 6440 28227 6443
rect 28258 6440 28264 6452
rect 28215 6412 28264 6440
rect 28215 6409 28227 6412
rect 28169 6403 28227 6409
rect 28258 6400 28264 6412
rect 28316 6400 28322 6452
rect 30009 6443 30067 6449
rect 30009 6409 30021 6443
rect 30055 6440 30067 6443
rect 30190 6440 30196 6452
rect 30055 6412 30196 6440
rect 30055 6409 30067 6412
rect 30009 6403 30067 6409
rect 30190 6400 30196 6412
rect 30248 6400 30254 6452
rect 33686 6440 33692 6452
rect 31726 6412 33692 6440
rect 30377 6375 30435 6381
rect 26160 6344 30328 6372
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23992 6208 24225 6236
rect 23992 6196 23998 6208
rect 24213 6205 24225 6208
rect 24259 6205 24271 6239
rect 24213 6199 24271 6205
rect 26053 6239 26111 6245
rect 26053 6205 26065 6239
rect 26099 6205 26111 6239
rect 26053 6199 26111 6205
rect 26160 6180 26188 6344
rect 26326 6264 26332 6316
rect 26384 6304 26390 6316
rect 27062 6304 27068 6316
rect 26384 6276 27068 6304
rect 26384 6264 26390 6276
rect 27062 6264 27068 6276
rect 27120 6264 27126 6316
rect 27614 6264 27620 6316
rect 27672 6264 27678 6316
rect 29270 6264 29276 6316
rect 29328 6304 29334 6316
rect 29638 6304 29644 6316
rect 29328 6276 29644 6304
rect 29328 6264 29334 6276
rect 29638 6264 29644 6276
rect 29696 6264 29702 6316
rect 30300 6304 30328 6344
rect 30377 6341 30389 6375
rect 30423 6372 30435 6375
rect 30466 6372 30472 6384
rect 30423 6344 30472 6372
rect 30423 6341 30435 6344
rect 30377 6335 30435 6341
rect 30466 6332 30472 6344
rect 30524 6372 30530 6384
rect 31018 6372 31024 6384
rect 30524 6344 31024 6372
rect 30524 6332 30530 6344
rect 31018 6332 31024 6344
rect 31076 6332 31082 6384
rect 30300 6276 30604 6304
rect 28813 6239 28871 6245
rect 28813 6205 28825 6239
rect 28859 6236 28871 6239
rect 29365 6239 29423 6245
rect 28859 6208 28948 6236
rect 28859 6205 28871 6208
rect 28813 6199 28871 6205
rect 25409 6171 25467 6177
rect 25409 6168 25421 6171
rect 21315 6140 22048 6168
rect 23860 6140 25421 6168
rect 21315 6137 21327 6140
rect 21269 6131 21327 6137
rect 22020 6112 22048 6140
rect 25409 6137 25421 6140
rect 25455 6168 25467 6171
rect 26142 6168 26148 6180
rect 25455 6140 26148 6168
rect 25455 6137 25467 6140
rect 25409 6131 25467 6137
rect 26142 6128 26148 6140
rect 26200 6128 26206 6180
rect 28920 6177 28948 6208
rect 29365 6205 29377 6239
rect 29411 6205 29423 6239
rect 29365 6199 29423 6205
rect 29549 6239 29607 6245
rect 29549 6205 29561 6239
rect 29595 6205 29607 6239
rect 29549 6199 29607 6205
rect 28905 6171 28963 6177
rect 28905 6137 28917 6171
rect 28951 6137 28963 6171
rect 28905 6131 28963 6137
rect 21545 6103 21603 6109
rect 21545 6100 21557 6103
rect 19852 6072 21557 6100
rect 19852 6060 19858 6072
rect 21545 6069 21557 6072
rect 21591 6069 21603 6103
rect 21545 6063 21603 6069
rect 22002 6060 22008 6112
rect 22060 6060 22066 6112
rect 22370 6060 22376 6112
rect 22428 6100 22434 6112
rect 22649 6103 22707 6109
rect 22649 6100 22661 6103
rect 22428 6072 22661 6100
rect 22428 6060 22434 6072
rect 22649 6069 22661 6072
rect 22695 6069 22707 6103
rect 22649 6063 22707 6069
rect 23658 6060 23664 6112
rect 23716 6060 23722 6112
rect 29380 6100 29408 6199
rect 29564 6168 29592 6199
rect 30374 6196 30380 6248
rect 30432 6236 30438 6248
rect 30576 6245 30604 6276
rect 30469 6239 30527 6245
rect 30469 6236 30481 6239
rect 30432 6208 30481 6236
rect 30432 6196 30438 6208
rect 30469 6205 30481 6208
rect 30515 6205 30527 6239
rect 30469 6199 30527 6205
rect 30561 6239 30619 6245
rect 30561 6205 30573 6239
rect 30607 6236 30619 6239
rect 31021 6239 31079 6245
rect 31021 6236 31033 6239
rect 30607 6208 31033 6236
rect 30607 6205 30619 6208
rect 30561 6199 30619 6205
rect 31021 6205 31033 6208
rect 31067 6205 31079 6239
rect 31021 6199 31079 6205
rect 31389 6171 31447 6177
rect 31389 6168 31401 6171
rect 29564 6140 31401 6168
rect 31389 6137 31401 6140
rect 31435 6168 31447 6171
rect 31726 6168 31754 6412
rect 33686 6400 33692 6412
rect 33744 6400 33750 6452
rect 33781 6443 33839 6449
rect 33781 6409 33793 6443
rect 33827 6440 33839 6443
rect 35066 6440 35072 6452
rect 33827 6412 35072 6440
rect 33827 6409 33839 6412
rect 33781 6403 33839 6409
rect 35066 6400 35072 6412
rect 35124 6400 35130 6452
rect 35158 6400 35164 6452
rect 35216 6440 35222 6452
rect 35713 6443 35771 6449
rect 35216 6412 35664 6440
rect 35216 6400 35222 6412
rect 35636 6372 35664 6412
rect 35713 6409 35725 6443
rect 35759 6440 35771 6443
rect 36078 6440 36084 6452
rect 35759 6412 36084 6440
rect 35759 6409 35771 6412
rect 35713 6403 35771 6409
rect 36078 6400 36084 6412
rect 36136 6400 36142 6452
rect 36814 6400 36820 6452
rect 36872 6400 36878 6452
rect 38746 6440 38752 6452
rect 37660 6412 38752 6440
rect 36173 6375 36231 6381
rect 36173 6372 36185 6375
rect 35636 6344 36185 6372
rect 36173 6341 36185 6344
rect 36219 6372 36231 6375
rect 36538 6372 36544 6384
rect 36219 6344 36544 6372
rect 36219 6341 36231 6344
rect 36173 6335 36231 6341
rect 36538 6332 36544 6344
rect 36596 6332 36602 6384
rect 32122 6264 32128 6316
rect 32180 6264 32186 6316
rect 32392 6307 32450 6313
rect 32392 6273 32404 6307
rect 32438 6304 32450 6307
rect 32950 6304 32956 6316
rect 32438 6276 32956 6304
rect 32438 6273 32450 6276
rect 32392 6267 32450 6273
rect 32950 6264 32956 6276
rect 33008 6264 33014 6316
rect 34698 6264 34704 6316
rect 34756 6264 34762 6316
rect 35437 6307 35495 6313
rect 35437 6273 35449 6307
rect 35483 6304 35495 6307
rect 35986 6304 35992 6316
rect 35483 6276 35992 6304
rect 35483 6273 35495 6276
rect 35437 6267 35495 6273
rect 35986 6264 35992 6276
rect 36044 6304 36050 6316
rect 36081 6307 36139 6313
rect 36081 6304 36093 6307
rect 36044 6276 36093 6304
rect 36044 6264 36050 6276
rect 36081 6273 36093 6276
rect 36127 6273 36139 6307
rect 36081 6267 36139 6273
rect 36722 6264 36728 6316
rect 36780 6264 36786 6316
rect 37660 6313 37688 6412
rect 38746 6400 38752 6412
rect 38804 6400 38810 6452
rect 39298 6400 39304 6452
rect 39356 6440 39362 6452
rect 40037 6443 40095 6449
rect 40037 6440 40049 6443
rect 39356 6412 40049 6440
rect 39356 6400 39362 6412
rect 40037 6409 40049 6412
rect 40083 6409 40095 6443
rect 40037 6403 40095 6409
rect 41782 6400 41788 6452
rect 41840 6400 41846 6452
rect 42886 6400 42892 6452
rect 42944 6440 42950 6452
rect 43073 6443 43131 6449
rect 43073 6440 43085 6443
rect 42944 6412 43085 6440
rect 42944 6400 42950 6412
rect 43073 6409 43085 6412
rect 43119 6409 43131 6443
rect 43073 6403 43131 6409
rect 44269 6443 44327 6449
rect 44269 6409 44281 6443
rect 44315 6440 44327 6443
rect 44910 6440 44916 6452
rect 44315 6412 44916 6440
rect 44315 6409 44327 6412
rect 44269 6403 44327 6409
rect 44910 6400 44916 6412
rect 44968 6400 44974 6452
rect 45373 6443 45431 6449
rect 45373 6409 45385 6443
rect 45419 6440 45431 6443
rect 45462 6440 45468 6452
rect 45419 6412 45468 6440
rect 45419 6409 45431 6412
rect 45373 6403 45431 6409
rect 45462 6400 45468 6412
rect 45520 6400 45526 6452
rect 45833 6443 45891 6449
rect 45833 6409 45845 6443
rect 45879 6440 45891 6443
rect 46474 6440 46480 6452
rect 45879 6412 46480 6440
rect 45879 6409 45891 6412
rect 45833 6403 45891 6409
rect 46474 6400 46480 6412
rect 46532 6400 46538 6452
rect 47581 6443 47639 6449
rect 47581 6409 47593 6443
rect 47627 6409 47639 6443
rect 47581 6403 47639 6409
rect 37645 6307 37703 6313
rect 37645 6273 37657 6307
rect 37691 6273 37703 6307
rect 37645 6267 37703 6273
rect 39485 6307 39543 6313
rect 39485 6273 39497 6307
rect 39531 6304 39543 6307
rect 39945 6307 40003 6313
rect 39945 6304 39957 6307
rect 39531 6276 39957 6304
rect 39531 6273 39543 6276
rect 39485 6267 39543 6273
rect 39945 6273 39957 6276
rect 39991 6273 40003 6307
rect 41800 6304 41828 6400
rect 45020 6344 46060 6372
rect 45020 6316 45048 6344
rect 42429 6307 42487 6313
rect 42429 6304 42441 6307
rect 41800 6276 42441 6304
rect 39945 6267 40003 6273
rect 42429 6273 42441 6276
rect 42475 6273 42487 6307
rect 42429 6267 42487 6273
rect 45002 6264 45008 6316
rect 45060 6264 45066 6316
rect 45465 6307 45523 6313
rect 45465 6273 45477 6307
rect 45511 6304 45523 6307
rect 45646 6304 45652 6316
rect 45511 6276 45652 6304
rect 45511 6273 45523 6276
rect 45465 6267 45523 6273
rect 45646 6264 45652 6276
rect 45704 6264 45710 6316
rect 46032 6313 46060 6344
rect 47596 6316 47624 6403
rect 47670 6400 47676 6452
rect 47728 6440 47734 6452
rect 48041 6443 48099 6449
rect 48041 6440 48053 6443
rect 47728 6412 48053 6440
rect 47728 6400 47734 6412
rect 48041 6409 48053 6412
rect 48087 6440 48099 6443
rect 48409 6443 48467 6449
rect 48409 6440 48421 6443
rect 48087 6412 48421 6440
rect 48087 6409 48099 6412
rect 48041 6403 48099 6409
rect 48409 6409 48421 6412
rect 48455 6409 48467 6443
rect 48409 6403 48467 6409
rect 49418 6400 49424 6452
rect 49476 6400 49482 6452
rect 49970 6400 49976 6452
rect 50028 6400 50034 6452
rect 50798 6400 50804 6452
rect 50856 6440 50862 6452
rect 50856 6412 51074 6440
rect 50856 6400 50862 6412
rect 47946 6332 47952 6384
rect 48004 6332 48010 6384
rect 49436 6372 49464 6400
rect 49574 6375 49632 6381
rect 49574 6372 49586 6375
rect 49436 6344 49586 6372
rect 49574 6341 49586 6344
rect 49620 6341 49632 6375
rect 49574 6335 49632 6341
rect 46017 6307 46075 6313
rect 46017 6273 46029 6307
rect 46063 6273 46075 6307
rect 46017 6267 46075 6273
rect 46284 6307 46342 6313
rect 46284 6273 46296 6307
rect 46330 6304 46342 6307
rect 46566 6304 46572 6316
rect 46330 6276 46572 6304
rect 46330 6273 46342 6276
rect 46284 6267 46342 6273
rect 46566 6264 46572 6276
rect 46624 6264 46630 6316
rect 47578 6264 47584 6316
rect 47636 6264 47642 6316
rect 49326 6264 49332 6316
rect 49384 6264 49390 6316
rect 49988 6304 50016 6400
rect 51046 6372 51074 6412
rect 51166 6400 51172 6452
rect 51224 6440 51230 6452
rect 51994 6440 52000 6452
rect 51224 6412 52000 6440
rect 51224 6400 51230 6412
rect 51994 6400 52000 6412
rect 52052 6440 52058 6452
rect 52089 6443 52147 6449
rect 52089 6440 52101 6443
rect 52052 6412 52101 6440
rect 52052 6400 52058 6412
rect 52089 6409 52101 6412
rect 52135 6409 52147 6443
rect 52089 6403 52147 6409
rect 52454 6400 52460 6452
rect 52512 6440 52518 6452
rect 53101 6443 53159 6449
rect 53101 6440 53113 6443
rect 52512 6412 53113 6440
rect 52512 6400 52518 6412
rect 53101 6409 53113 6412
rect 53147 6409 53159 6443
rect 53101 6403 53159 6409
rect 54202 6400 54208 6452
rect 54260 6400 54266 6452
rect 54386 6400 54392 6452
rect 54444 6440 54450 6452
rect 54665 6443 54723 6449
rect 54665 6440 54677 6443
rect 54444 6412 54677 6440
rect 54444 6400 54450 6412
rect 54665 6409 54677 6412
rect 54711 6409 54723 6443
rect 54665 6403 54723 6409
rect 55582 6400 55588 6452
rect 55640 6400 55646 6452
rect 56137 6443 56195 6449
rect 56137 6409 56149 6443
rect 56183 6440 56195 6443
rect 56410 6440 56416 6452
rect 56183 6412 56416 6440
rect 56183 6409 56195 6412
rect 56137 6403 56195 6409
rect 56410 6400 56416 6412
rect 56468 6400 56474 6452
rect 57054 6400 57060 6452
rect 57112 6400 57118 6452
rect 57422 6400 57428 6452
rect 57480 6400 57486 6452
rect 57790 6400 57796 6452
rect 57848 6400 57854 6452
rect 52181 6375 52239 6381
rect 52181 6372 52193 6375
rect 51046 6344 52193 6372
rect 52181 6341 52193 6344
rect 52227 6372 52239 6375
rect 52730 6372 52736 6384
rect 52227 6344 52736 6372
rect 52227 6341 52239 6344
rect 52181 6335 52239 6341
rect 52730 6332 52736 6344
rect 52788 6332 52794 6384
rect 55600 6372 55628 6400
rect 56505 6375 56563 6381
rect 56505 6372 56517 6375
rect 55600 6344 56517 6372
rect 56505 6341 56517 6344
rect 56551 6341 56563 6375
rect 56505 6335 56563 6341
rect 49988 6276 50844 6304
rect 33778 6196 33784 6248
rect 33836 6236 33842 6248
rect 34422 6236 34428 6248
rect 33836 6208 34428 6236
rect 33836 6196 33842 6208
rect 34422 6196 34428 6208
rect 34480 6196 34486 6248
rect 34606 6245 34612 6248
rect 34584 6239 34612 6245
rect 34584 6205 34596 6239
rect 34584 6199 34612 6205
rect 34606 6196 34612 6199
rect 34664 6196 34670 6248
rect 35621 6239 35679 6245
rect 35621 6205 35633 6239
rect 35667 6205 35679 6239
rect 35621 6199 35679 6205
rect 31435 6140 31754 6168
rect 31435 6137 31447 6140
rect 31389 6131 31447 6137
rect 34882 6128 34888 6180
rect 34940 6168 34946 6180
rect 34977 6171 35035 6177
rect 34977 6168 34989 6171
rect 34940 6140 34989 6168
rect 34940 6128 34946 6140
rect 34977 6137 34989 6140
rect 35023 6137 35035 6171
rect 35636 6168 35664 6199
rect 35802 6196 35808 6248
rect 35860 6236 35866 6248
rect 36265 6239 36323 6245
rect 36265 6236 36277 6239
rect 35860 6208 36277 6236
rect 35860 6196 35866 6208
rect 36265 6205 36277 6208
rect 36311 6205 36323 6239
rect 36265 6199 36323 6205
rect 36740 6168 36768 6264
rect 37826 6196 37832 6248
rect 37884 6196 37890 6248
rect 38746 6245 38752 6248
rect 38565 6239 38623 6245
rect 38565 6236 38577 6239
rect 38120 6208 38577 6236
rect 35636 6140 36768 6168
rect 34977 6131 35035 6137
rect 30374 6100 30380 6112
rect 29380 6072 30380 6100
rect 30374 6060 30380 6072
rect 30432 6060 30438 6112
rect 33505 6103 33563 6109
rect 33505 6069 33517 6103
rect 33551 6100 33563 6103
rect 33686 6100 33692 6112
rect 33551 6072 33692 6100
rect 33551 6069 33563 6072
rect 33505 6063 33563 6069
rect 33686 6060 33692 6072
rect 33744 6060 33750 6112
rect 34992 6100 35020 6131
rect 38010 6128 38016 6180
rect 38068 6168 38074 6180
rect 38120 6168 38148 6208
rect 38565 6205 38577 6208
rect 38611 6205 38623 6239
rect 38565 6199 38623 6205
rect 38703 6239 38752 6245
rect 38703 6205 38715 6239
rect 38749 6205 38752 6239
rect 38703 6199 38752 6205
rect 38746 6196 38752 6199
rect 38804 6196 38810 6248
rect 38841 6239 38899 6245
rect 38841 6205 38853 6239
rect 38887 6236 38899 6239
rect 39022 6236 39028 6248
rect 38887 6208 39028 6236
rect 38887 6205 38899 6208
rect 38841 6199 38899 6205
rect 39022 6196 39028 6208
rect 39080 6196 39086 6248
rect 39850 6196 39856 6248
rect 39908 6236 39914 6248
rect 40129 6239 40187 6245
rect 40129 6236 40141 6239
rect 39908 6208 40141 6236
rect 39908 6196 39914 6208
rect 40129 6205 40141 6208
rect 40175 6205 40187 6239
rect 40129 6199 40187 6205
rect 45281 6239 45339 6245
rect 45281 6205 45293 6239
rect 45327 6236 45339 6239
rect 45327 6208 45416 6236
rect 45327 6205 45339 6208
rect 45281 6199 45339 6205
rect 38068 6140 38148 6168
rect 38068 6128 38074 6140
rect 38194 6128 38200 6180
rect 38252 6168 38258 6180
rect 38289 6171 38347 6177
rect 38289 6168 38301 6171
rect 38252 6140 38301 6168
rect 38252 6128 38258 6140
rect 38289 6137 38301 6140
rect 38335 6137 38347 6171
rect 38289 6131 38347 6137
rect 42610 6128 42616 6180
rect 42668 6168 42674 6180
rect 42668 6140 45048 6168
rect 42668 6128 42674 6140
rect 37458 6100 37464 6112
rect 34992 6072 37464 6100
rect 37458 6060 37464 6072
rect 37516 6060 37522 6112
rect 38378 6060 38384 6112
rect 38436 6100 38442 6112
rect 38838 6100 38844 6112
rect 38436 6072 38844 6100
rect 38436 6060 38442 6072
rect 38838 6060 38844 6072
rect 38896 6060 38902 6112
rect 39574 6060 39580 6112
rect 39632 6060 39638 6112
rect 44082 6060 44088 6112
rect 44140 6100 44146 6112
rect 45020 6109 45048 6140
rect 44637 6103 44695 6109
rect 44637 6100 44649 6103
rect 44140 6072 44649 6100
rect 44140 6060 44146 6072
rect 44637 6069 44649 6072
rect 44683 6069 44695 6103
rect 44637 6063 44695 6069
rect 45005 6103 45063 6109
rect 45005 6069 45017 6103
rect 45051 6100 45063 6103
rect 45388 6100 45416 6208
rect 47210 6196 47216 6248
rect 47268 6236 47274 6248
rect 48130 6236 48136 6248
rect 47268 6208 48136 6236
rect 47268 6196 47274 6208
rect 48130 6196 48136 6208
rect 48188 6196 48194 6248
rect 48961 6239 49019 6245
rect 48961 6205 48973 6239
rect 49007 6205 49019 6239
rect 48961 6199 49019 6205
rect 47397 6171 47455 6177
rect 47397 6137 47409 6171
rect 47443 6168 47455 6171
rect 48976 6168 49004 6199
rect 50816 6177 50844 6276
rect 51166 6264 51172 6316
rect 51224 6264 51230 6316
rect 51460 6276 52040 6304
rect 51460 6245 51488 6276
rect 52012 6248 52040 6276
rect 52546 6264 52552 6316
rect 52604 6304 52610 6316
rect 53193 6307 53251 6313
rect 53193 6304 53205 6307
rect 52604 6276 53205 6304
rect 52604 6264 52610 6276
rect 53193 6273 53205 6276
rect 53239 6273 53251 6307
rect 53193 6267 53251 6273
rect 53392 6276 54616 6304
rect 51261 6239 51319 6245
rect 51261 6205 51273 6239
rect 51307 6205 51319 6239
rect 51261 6199 51319 6205
rect 51445 6239 51503 6245
rect 51445 6205 51457 6239
rect 51491 6205 51503 6239
rect 51445 6199 51503 6205
rect 51905 6239 51963 6245
rect 51905 6205 51917 6239
rect 51951 6205 51963 6239
rect 51905 6199 51963 6205
rect 47443 6140 49004 6168
rect 50801 6171 50859 6177
rect 47443 6137 47455 6140
rect 47397 6131 47455 6137
rect 50801 6137 50813 6171
rect 50847 6137 50859 6171
rect 50801 6131 50859 6137
rect 51276 6112 51304 6199
rect 46658 6100 46664 6112
rect 45051 6072 46664 6100
rect 45051 6069 45063 6072
rect 45005 6063 45063 6069
rect 46658 6060 46664 6072
rect 46716 6100 46722 6112
rect 50246 6100 50252 6112
rect 46716 6072 50252 6100
rect 46716 6060 46722 6072
rect 50246 6060 50252 6072
rect 50304 6060 50310 6112
rect 50706 6060 50712 6112
rect 50764 6060 50770 6112
rect 51258 6060 51264 6112
rect 51316 6060 51322 6112
rect 51920 6100 51948 6199
rect 51994 6196 52000 6248
rect 52052 6196 52058 6248
rect 52086 6196 52092 6248
rect 52144 6236 52150 6248
rect 53392 6245 53420 6276
rect 53377 6239 53435 6245
rect 53377 6236 53389 6239
rect 52144 6208 53389 6236
rect 52144 6196 52150 6208
rect 53377 6205 53389 6208
rect 53423 6205 53435 6239
rect 53377 6199 53435 6205
rect 53561 6239 53619 6245
rect 53561 6205 53573 6239
rect 53607 6205 53619 6239
rect 53561 6199 53619 6205
rect 52549 6171 52607 6177
rect 52549 6137 52561 6171
rect 52595 6168 52607 6171
rect 53576 6168 53604 6199
rect 52595 6140 53604 6168
rect 52595 6137 52607 6140
rect 52549 6131 52607 6137
rect 52362 6100 52368 6112
rect 51920 6072 52368 6100
rect 52362 6060 52368 6072
rect 52420 6060 52426 6112
rect 52730 6060 52736 6112
rect 52788 6060 52794 6112
rect 54588 6109 54616 6276
rect 55306 6264 55312 6316
rect 55364 6264 55370 6316
rect 55490 6264 55496 6316
rect 55548 6264 55554 6316
rect 57808 6304 57836 6400
rect 58437 6307 58495 6313
rect 58437 6304 58449 6307
rect 57808 6276 58449 6304
rect 58437 6273 58449 6276
rect 58483 6273 58495 6307
rect 58437 6267 58495 6273
rect 56870 6196 56876 6248
rect 56928 6196 56934 6248
rect 56965 6239 57023 6245
rect 56965 6205 56977 6239
rect 57011 6236 57023 6239
rect 57330 6236 57336 6248
rect 57011 6208 57336 6236
rect 57011 6205 57023 6208
rect 56965 6199 57023 6205
rect 57330 6196 57336 6208
rect 57388 6236 57394 6248
rect 57885 6239 57943 6245
rect 57885 6236 57897 6239
rect 57388 6208 57897 6236
rect 57388 6196 57394 6208
rect 57885 6205 57897 6208
rect 57931 6205 57943 6239
rect 57885 6199 57943 6205
rect 54573 6103 54631 6109
rect 54573 6069 54585 6103
rect 54619 6100 54631 6103
rect 55398 6100 55404 6112
rect 54619 6072 55404 6100
rect 54619 6069 54631 6072
rect 54573 6063 54631 6069
rect 55398 6060 55404 6072
rect 55456 6060 55462 6112
rect 1104 6010 58880 6032
rect 1104 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 22616 6010
rect 22668 5958 22680 6010
rect 22732 5958 22744 6010
rect 22796 5958 22808 6010
rect 22860 5958 22872 6010
rect 22924 5958 37060 6010
rect 37112 5958 37124 6010
rect 37176 5958 37188 6010
rect 37240 5958 37252 6010
rect 37304 5958 37316 6010
rect 37368 5958 51504 6010
rect 51556 5958 51568 6010
rect 51620 5958 51632 6010
rect 51684 5958 51696 6010
rect 51748 5958 51760 6010
rect 51812 5958 58880 6010
rect 1104 5936 58880 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 2130 5896 2136 5908
rect 1964 5868 2136 5896
rect 1964 5769 1992 5868
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 8941 5899 8999 5905
rect 2372 5868 8800 5896
rect 2372 5856 2378 5868
rect 3326 5788 3332 5840
rect 3384 5788 3390 5840
rect 4448 5769 4476 5868
rect 6086 5788 6092 5840
rect 6144 5788 6150 5840
rect 6270 5788 6276 5840
rect 6328 5788 6334 5840
rect 8772 5837 8800 5868
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9214 5896 9220 5908
rect 8987 5868 9220 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9582 5896 9588 5908
rect 9508 5868 9588 5896
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9508 5828 9536 5868
rect 9582 5856 9588 5868
rect 9640 5896 9646 5908
rect 9640 5856 9674 5896
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10965 5899 11023 5905
rect 10965 5896 10977 5899
rect 10836 5868 10977 5896
rect 10836 5856 10842 5868
rect 10965 5865 10977 5868
rect 11011 5865 11023 5899
rect 10965 5859 11023 5865
rect 12986 5856 12992 5908
rect 13044 5856 13050 5908
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 13446 5896 13452 5908
rect 13127 5868 13452 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 14918 5896 14924 5908
rect 14783 5868 14924 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 17034 5896 17040 5908
rect 15252 5868 17040 5896
rect 15252 5856 15258 5868
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 19242 5856 19248 5908
rect 19300 5856 19306 5908
rect 22002 5856 22008 5908
rect 22060 5856 22066 5908
rect 24029 5899 24087 5905
rect 24029 5865 24041 5899
rect 24075 5896 24087 5899
rect 24118 5896 24124 5908
rect 24075 5868 24124 5896
rect 24075 5865 24087 5868
rect 24029 5859 24087 5865
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 26142 5856 26148 5908
rect 26200 5856 26206 5908
rect 27890 5856 27896 5908
rect 27948 5896 27954 5908
rect 29733 5899 29791 5905
rect 29733 5896 29745 5899
rect 27948 5868 29745 5896
rect 27948 5856 27954 5868
rect 29733 5865 29745 5868
rect 29779 5865 29791 5899
rect 29733 5859 29791 5865
rect 30374 5856 30380 5908
rect 30432 5856 30438 5908
rect 30926 5856 30932 5908
rect 30984 5896 30990 5908
rect 31110 5896 31116 5908
rect 30984 5868 31116 5896
rect 30984 5856 30990 5868
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 32950 5856 32956 5908
rect 33008 5856 33014 5908
rect 33502 5856 33508 5908
rect 33560 5856 33566 5908
rect 33686 5856 33692 5908
rect 33744 5856 33750 5908
rect 33870 5856 33876 5908
rect 33928 5896 33934 5908
rect 34425 5899 34483 5905
rect 34425 5896 34437 5899
rect 33928 5868 34437 5896
rect 33928 5856 33934 5868
rect 34425 5865 34437 5868
rect 34471 5896 34483 5899
rect 34606 5896 34612 5908
rect 34471 5868 34612 5896
rect 34471 5865 34483 5868
rect 34425 5859 34483 5865
rect 34606 5856 34612 5868
rect 34664 5856 34670 5908
rect 35345 5899 35403 5905
rect 35345 5865 35357 5899
rect 35391 5896 35403 5899
rect 35802 5896 35808 5908
rect 35391 5868 35808 5896
rect 35391 5865 35403 5868
rect 35345 5859 35403 5865
rect 35802 5856 35808 5868
rect 35860 5856 35866 5908
rect 37826 5856 37832 5908
rect 37884 5896 37890 5908
rect 38378 5896 38384 5908
rect 37884 5868 38384 5896
rect 37884 5856 37890 5868
rect 38378 5856 38384 5868
rect 38436 5856 38442 5908
rect 38608 5856 38614 5908
rect 38666 5896 38672 5908
rect 38841 5899 38899 5905
rect 38841 5896 38853 5899
rect 38666 5868 38853 5896
rect 38666 5856 38672 5868
rect 38841 5865 38853 5868
rect 38887 5865 38899 5899
rect 38841 5859 38899 5865
rect 39114 5856 39120 5908
rect 39172 5856 39178 5908
rect 45830 5856 45836 5908
rect 45888 5896 45894 5908
rect 46385 5899 46443 5905
rect 46385 5896 46397 5899
rect 45888 5868 46397 5896
rect 45888 5856 45894 5868
rect 46385 5865 46397 5868
rect 46431 5865 46443 5899
rect 46385 5859 46443 5865
rect 46566 5856 46572 5908
rect 46624 5896 46630 5908
rect 46937 5899 46995 5905
rect 46937 5896 46949 5899
rect 46624 5868 46949 5896
rect 46624 5856 46630 5868
rect 46937 5865 46949 5868
rect 46983 5865 46995 5899
rect 46937 5859 46995 5865
rect 47857 5899 47915 5905
rect 47857 5865 47869 5899
rect 47903 5896 47915 5899
rect 47946 5896 47952 5908
rect 47903 5868 47952 5896
rect 47903 5865 47915 5868
rect 47857 5859 47915 5865
rect 47946 5856 47952 5868
rect 48004 5856 48010 5908
rect 48130 5856 48136 5908
rect 48188 5896 48194 5908
rect 48225 5899 48283 5905
rect 48225 5896 48237 5899
rect 48188 5868 48237 5896
rect 48188 5856 48194 5868
rect 48225 5865 48237 5868
rect 48271 5865 48283 5899
rect 48225 5859 48283 5865
rect 8803 5800 9536 5828
rect 9646 5828 9674 5856
rect 12161 5831 12219 5837
rect 12161 5828 12173 5831
rect 9646 5800 12173 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 4614 5720 4620 5772
rect 4672 5720 4678 5772
rect 6288 5760 6316 5788
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6288 5732 6837 5760
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 9508 5769 9536 5800
rect 12161 5797 12173 5800
rect 12207 5828 12219 5831
rect 12207 5800 13768 5828
rect 12207 5797 12219 5800
rect 12161 5791 12219 5797
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 9364 5732 9413 5760
rect 9364 5720 9370 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4120 5664 5856 5692
rect 4120 5652 4126 5664
rect 2216 5627 2274 5633
rect 2216 5593 2228 5627
rect 2262 5624 2274 5627
rect 3050 5624 3056 5636
rect 2262 5596 3056 5624
rect 2262 5593 2274 5596
rect 2216 5587 2274 5593
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4798 5624 4804 5636
rect 4203 5596 4804 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4798 5584 4804 5596
rect 4856 5624 4862 5636
rect 5828 5633 5856 5664
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 6236 5664 6285 5692
rect 6236 5652 6242 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 7800 5664 8309 5692
rect 7800 5652 7806 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 9416 5692 9444 5723
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 13740 5769 13768 5800
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10100 5732 10333 5760
rect 10100 5720 10106 5732
rect 10321 5729 10333 5732
rect 10367 5760 10379 5763
rect 13725 5763 13783 5769
rect 10367 5732 11744 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 9416 5664 10517 5692
rect 8297 5655 8355 5661
rect 10505 5661 10517 5664
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 10870 5692 10876 5704
rect 10643 5664 10876 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11020 5664 11621 5692
rect 11020 5652 11026 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 5261 5627 5319 5633
rect 5261 5624 5273 5627
rect 4856 5596 5273 5624
rect 4856 5584 4862 5596
rect 5261 5593 5273 5596
rect 5307 5593 5319 5627
rect 5261 5587 5319 5593
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5624 5871 5627
rect 9309 5627 9367 5633
rect 5859 5596 7880 5624
rect 5859 5593 5871 5596
rect 5813 5587 5871 5593
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3752 5528 3801 5556
rect 3752 5516 3758 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4246 5516 4252 5568
rect 4304 5516 4310 5568
rect 4338 5516 4344 5568
rect 4396 5556 4402 5568
rect 6086 5556 6092 5568
rect 4396 5528 6092 5556
rect 4396 5516 4402 5528
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 7006 5516 7012 5568
rect 7064 5516 7070 5568
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 7745 5559 7803 5565
rect 7745 5556 7757 5559
rect 7248 5528 7757 5556
rect 7248 5516 7254 5528
rect 7745 5525 7757 5528
rect 7791 5525 7803 5559
rect 7852 5556 7880 5596
rect 9309 5593 9321 5627
rect 9355 5624 9367 5627
rect 11057 5627 11115 5633
rect 11057 5624 11069 5627
rect 9355 5596 11069 5624
rect 9355 5593 9367 5596
rect 9309 5587 9367 5593
rect 10520 5568 10548 5596
rect 11057 5593 11069 5596
rect 11103 5593 11115 5627
rect 11716 5624 11744 5732
rect 13725 5729 13737 5763
rect 13771 5729 13783 5763
rect 13725 5723 13783 5729
rect 13740 5692 13768 5723
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 13964 5732 14105 5760
rect 13964 5720 13970 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 14826 5692 14832 5704
rect 13740 5664 14832 5692
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 13354 5624 13360 5636
rect 11716 5596 13360 5624
rect 11057 5587 11115 5593
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 14936 5624 14964 5856
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 18288 5732 18429 5760
rect 18288 5720 18294 5732
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 22020 5760 22048 5856
rect 22833 5831 22891 5837
rect 22833 5797 22845 5831
rect 22879 5797 22891 5831
rect 22833 5791 22891 5797
rect 20680 5732 22048 5760
rect 20680 5720 20686 5732
rect 22370 5720 22376 5772
rect 22428 5720 22434 5772
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5760 22799 5763
rect 22848 5760 22876 5791
rect 26160 5769 26188 5856
rect 26789 5831 26847 5837
rect 26789 5797 26801 5831
rect 26835 5828 26847 5831
rect 26835 5800 27476 5828
rect 26835 5797 26847 5800
rect 26789 5791 26847 5797
rect 22787 5732 22876 5760
rect 23385 5763 23443 5769
rect 22787 5729 22799 5732
rect 22741 5723 22799 5729
rect 23385 5729 23397 5763
rect 23431 5729 23443 5763
rect 23385 5723 23443 5729
rect 26145 5763 26203 5769
rect 26145 5729 26157 5763
rect 26191 5729 26203 5763
rect 26145 5723 26203 5729
rect 15286 5652 15292 5704
rect 15344 5692 15350 5704
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15344 5664 15669 5692
rect 15344 5652 15350 5664
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16264 5664 16773 5692
rect 16264 5652 16270 5664
rect 16761 5661 16773 5664
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 17586 5652 17592 5704
rect 17644 5652 17650 5704
rect 18322 5652 18328 5704
rect 18380 5652 18386 5704
rect 21266 5652 21272 5704
rect 21324 5652 21330 5704
rect 22388 5692 22416 5720
rect 23400 5692 23428 5723
rect 26326 5720 26332 5772
rect 26384 5720 26390 5772
rect 27448 5769 27476 5800
rect 33520 5769 33548 5856
rect 27433 5763 27491 5769
rect 27433 5729 27445 5763
rect 27479 5729 27491 5763
rect 27433 5723 27491 5729
rect 33505 5763 33563 5769
rect 33505 5729 33517 5763
rect 33551 5729 33563 5763
rect 33704 5760 33732 5856
rect 38749 5831 38807 5837
rect 37568 5800 38700 5828
rect 33781 5763 33839 5769
rect 33781 5760 33793 5763
rect 33704 5732 33793 5760
rect 33505 5723 33563 5729
rect 33781 5729 33793 5732
rect 33827 5729 33839 5763
rect 33781 5723 33839 5729
rect 34422 5720 34428 5772
rect 34480 5760 34486 5772
rect 37568 5769 37596 5800
rect 37553 5763 37611 5769
rect 37553 5760 37565 5763
rect 34480 5732 37565 5760
rect 34480 5720 34486 5732
rect 37553 5729 37565 5732
rect 37599 5729 37611 5763
rect 37553 5723 37611 5729
rect 37734 5720 37740 5772
rect 37792 5760 37798 5772
rect 38105 5763 38163 5769
rect 38105 5760 38117 5763
rect 37792 5732 38117 5760
rect 37792 5720 37798 5732
rect 38105 5729 38117 5732
rect 38151 5729 38163 5763
rect 38672 5760 38700 5800
rect 38749 5797 38761 5831
rect 38795 5828 38807 5831
rect 39132 5828 39160 5856
rect 38795 5800 39160 5828
rect 38795 5797 38807 5800
rect 38749 5791 38807 5797
rect 39850 5788 39856 5840
rect 39908 5828 39914 5840
rect 45189 5831 45247 5837
rect 45189 5828 45201 5831
rect 39908 5800 45201 5828
rect 39908 5788 39914 5800
rect 45189 5797 45201 5800
rect 45235 5828 45247 5831
rect 45370 5828 45376 5840
rect 45235 5800 45376 5828
rect 45235 5797 45247 5800
rect 45189 5791 45247 5797
rect 45370 5788 45376 5800
rect 45428 5788 45434 5840
rect 39022 5760 39028 5772
rect 38672 5732 39028 5760
rect 38105 5723 38163 5729
rect 39022 5720 39028 5732
rect 39080 5720 39086 5772
rect 40862 5760 40868 5772
rect 39316 5732 40868 5760
rect 22388 5664 23428 5692
rect 24946 5652 24952 5704
rect 25004 5652 25010 5704
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 35437 5695 35495 5701
rect 35437 5661 35449 5695
rect 35483 5692 35495 5695
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 35483 5664 37841 5692
rect 35483 5661 35495 5664
rect 35437 5655 35495 5661
rect 37829 5661 37841 5664
rect 37875 5692 37887 5695
rect 39316 5692 39344 5732
rect 40862 5720 40868 5732
rect 40920 5720 40926 5772
rect 44082 5760 44088 5772
rect 43088 5732 44088 5760
rect 43088 5704 43116 5732
rect 44082 5720 44088 5732
rect 44140 5760 44146 5772
rect 44729 5763 44787 5769
rect 44729 5760 44741 5763
rect 44140 5732 44741 5760
rect 44140 5720 44146 5732
rect 44729 5729 44741 5732
rect 44775 5729 44787 5763
rect 44729 5723 44787 5729
rect 37875 5664 39344 5692
rect 37875 5661 37887 5664
rect 37829 5655 37887 5661
rect 39390 5652 39396 5704
rect 39448 5652 39454 5704
rect 40129 5695 40187 5701
rect 40129 5692 40141 5695
rect 39500 5664 40141 5692
rect 13495 5596 14964 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 19794 5624 19800 5636
rect 16540 5596 19800 5624
rect 16540 5584 16546 5596
rect 19794 5584 19800 5596
rect 19852 5584 19858 5636
rect 20380 5627 20438 5633
rect 20380 5593 20392 5627
rect 20426 5624 20438 5627
rect 20717 5627 20775 5633
rect 20717 5624 20729 5627
rect 20426 5596 20729 5624
rect 20426 5593 20438 5596
rect 20380 5587 20438 5593
rect 20717 5593 20729 5596
rect 20763 5593 20775 5627
rect 20717 5587 20775 5593
rect 23201 5627 23259 5633
rect 23201 5593 23213 5627
rect 23247 5624 23259 5627
rect 24210 5624 24216 5636
rect 23247 5596 24216 5624
rect 23247 5593 23259 5596
rect 23201 5587 23259 5593
rect 24210 5584 24216 5596
rect 24268 5584 24274 5636
rect 24302 5584 24308 5636
rect 24360 5584 24366 5636
rect 26421 5627 26479 5633
rect 26421 5624 26433 5627
rect 25332 5596 26433 5624
rect 9490 5556 9496 5568
rect 7852 5528 9496 5556
rect 7745 5519 7803 5525
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 10502 5516 10508 5568
rect 10560 5516 10566 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12621 5559 12679 5565
rect 12621 5556 12633 5559
rect 11848 5528 12633 5556
rect 11848 5516 11854 5528
rect 12621 5525 12633 5528
rect 12667 5556 12679 5559
rect 13262 5556 13268 5568
rect 12667 5528 13268 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13998 5556 14004 5568
rect 13587 5528 14004 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 15565 5559 15623 5565
rect 15565 5525 15577 5559
rect 15611 5556 15623 5559
rect 16022 5556 16028 5568
rect 15611 5528 16028 5556
rect 15611 5525 15623 5528
rect 15565 5519 15623 5525
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 16301 5559 16359 5565
rect 16301 5525 16313 5559
rect 16347 5556 16359 5559
rect 16666 5556 16672 5568
rect 16347 5528 16672 5556
rect 16347 5525 16359 5528
rect 16301 5519 16359 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 16945 5559 17003 5565
rect 16945 5525 16957 5559
rect 16991 5556 17003 5559
rect 17126 5556 17132 5568
rect 16991 5528 17132 5556
rect 16991 5525 17003 5528
rect 16945 5519 17003 5525
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 17678 5516 17684 5568
rect 17736 5516 17742 5568
rect 19058 5516 19064 5568
rect 19116 5516 19122 5568
rect 22097 5559 22155 5565
rect 22097 5525 22109 5559
rect 22143 5556 22155 5559
rect 22186 5556 22192 5568
rect 22143 5528 22192 5556
rect 22143 5525 22155 5528
rect 22097 5519 22155 5525
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 23293 5559 23351 5565
rect 23293 5525 23305 5559
rect 23339 5556 23351 5559
rect 24320 5556 24348 5584
rect 23339 5528 24348 5556
rect 23339 5525 23351 5528
rect 23293 5519 23351 5525
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 24854 5516 24860 5568
rect 24912 5556 24918 5568
rect 25332 5565 25360 5596
rect 26421 5593 26433 5596
rect 26467 5593 26479 5627
rect 26421 5587 26479 5593
rect 29730 5584 29736 5636
rect 29788 5624 29794 5636
rect 30285 5627 30343 5633
rect 30285 5624 30297 5627
rect 29788 5596 30297 5624
rect 29788 5584 29794 5596
rect 30285 5593 30297 5596
rect 30331 5593 30343 5627
rect 36814 5624 36820 5636
rect 30285 5587 30343 5593
rect 30760 5596 36820 5624
rect 25317 5559 25375 5565
rect 25317 5556 25329 5559
rect 24912 5528 25329 5556
rect 24912 5516 24918 5528
rect 25317 5525 25329 5528
rect 25363 5525 25375 5559
rect 25317 5519 25375 5525
rect 26878 5516 26884 5568
rect 26936 5516 26942 5568
rect 30650 5516 30656 5568
rect 30708 5556 30714 5568
rect 30760 5565 30788 5596
rect 36814 5584 36820 5596
rect 36872 5584 36878 5636
rect 37185 5627 37243 5633
rect 37185 5593 37197 5627
rect 37231 5624 37243 5627
rect 38381 5627 38439 5633
rect 37231 5596 37688 5624
rect 37231 5593 37243 5596
rect 37185 5587 37243 5593
rect 37660 5568 37688 5596
rect 38381 5593 38393 5627
rect 38427 5624 38439 5627
rect 38838 5624 38844 5636
rect 38427 5596 38844 5624
rect 38427 5593 38439 5596
rect 38381 5587 38439 5593
rect 38838 5584 38844 5596
rect 38896 5584 38902 5636
rect 39500 5624 39528 5664
rect 40129 5661 40141 5664
rect 40175 5661 40187 5695
rect 40129 5655 40187 5661
rect 41414 5652 41420 5704
rect 41472 5652 41478 5704
rect 41782 5652 41788 5704
rect 41840 5652 41846 5704
rect 42334 5652 42340 5704
rect 42392 5692 42398 5704
rect 42429 5695 42487 5701
rect 42429 5692 42441 5695
rect 42392 5664 42441 5692
rect 42392 5652 42398 5664
rect 42429 5661 42441 5664
rect 42475 5661 42487 5695
rect 42429 5655 42487 5661
rect 42978 5652 42984 5704
rect 43036 5652 43042 5704
rect 43070 5652 43076 5704
rect 43128 5652 43134 5704
rect 44174 5652 44180 5704
rect 44232 5692 44238 5704
rect 44361 5695 44419 5701
rect 44361 5692 44373 5695
rect 44232 5664 44373 5692
rect 44232 5652 44238 5664
rect 44361 5661 44373 5664
rect 44407 5661 44419 5695
rect 45388 5692 45416 5788
rect 47578 5720 47584 5772
rect 47636 5720 47642 5772
rect 48240 5760 48268 5859
rect 48590 5856 48596 5908
rect 48648 5896 48654 5908
rect 48685 5899 48743 5905
rect 48685 5896 48697 5899
rect 48648 5868 48697 5896
rect 48648 5856 48654 5868
rect 48685 5865 48697 5868
rect 48731 5896 48743 5899
rect 49050 5896 49056 5908
rect 48731 5868 49056 5896
rect 48731 5865 48743 5868
rect 48685 5859 48743 5865
rect 49050 5856 49056 5868
rect 49108 5856 49114 5908
rect 50706 5856 50712 5908
rect 50764 5856 50770 5908
rect 51258 5856 51264 5908
rect 51316 5896 51322 5908
rect 51629 5899 51687 5905
rect 51629 5896 51641 5899
rect 51316 5868 51641 5896
rect 51316 5856 51322 5868
rect 51629 5865 51641 5868
rect 51675 5865 51687 5899
rect 51629 5859 51687 5865
rect 51994 5856 52000 5908
rect 52052 5896 52058 5908
rect 52914 5896 52920 5908
rect 52052 5868 52920 5896
rect 52052 5856 52058 5868
rect 52914 5856 52920 5868
rect 52972 5856 52978 5908
rect 50724 5760 50752 5856
rect 50985 5763 51043 5769
rect 50985 5760 50997 5763
rect 48240 5732 48452 5760
rect 50724 5732 50997 5760
rect 45388 5664 48314 5692
rect 44361 5655 44419 5661
rect 38948 5596 39528 5624
rect 39945 5627 40003 5633
rect 30745 5559 30803 5565
rect 30745 5556 30757 5559
rect 30708 5528 30757 5556
rect 30708 5516 30714 5528
rect 30745 5525 30757 5528
rect 30791 5525 30803 5559
rect 30745 5519 30803 5525
rect 34146 5516 34152 5568
rect 34204 5556 34210 5568
rect 36906 5556 36912 5568
rect 34204 5528 36912 5556
rect 34204 5516 34210 5528
rect 36906 5516 36912 5528
rect 36964 5516 36970 5568
rect 37642 5516 37648 5568
rect 37700 5516 37706 5568
rect 38102 5516 38108 5568
rect 38160 5556 38166 5568
rect 38289 5559 38347 5565
rect 38289 5556 38301 5559
rect 38160 5528 38301 5556
rect 38160 5516 38166 5528
rect 38289 5525 38301 5528
rect 38335 5556 38347 5559
rect 38948 5556 38976 5596
rect 39945 5593 39957 5627
rect 39991 5593 40003 5627
rect 39945 5587 40003 5593
rect 38335 5528 38976 5556
rect 38335 5525 38347 5528
rect 38289 5519 38347 5525
rect 39390 5516 39396 5568
rect 39448 5556 39454 5568
rect 39960 5556 39988 5587
rect 42702 5584 42708 5636
rect 42760 5624 42766 5636
rect 42760 5596 46980 5624
rect 42760 5584 42766 5596
rect 39448 5528 39988 5556
rect 39448 5516 39454 5528
rect 40862 5516 40868 5568
rect 40920 5516 40926 5568
rect 41690 5516 41696 5568
rect 41748 5556 41754 5568
rect 42337 5559 42395 5565
rect 42337 5556 42349 5559
rect 41748 5528 42349 5556
rect 41748 5516 41754 5528
rect 42337 5525 42349 5528
rect 42383 5525 42395 5559
rect 42337 5519 42395 5525
rect 43622 5516 43628 5568
rect 43680 5556 43686 5568
rect 43809 5559 43867 5565
rect 43809 5556 43821 5559
rect 43680 5528 43821 5556
rect 43680 5516 43686 5528
rect 43809 5525 43821 5528
rect 43855 5525 43867 5559
rect 46952 5556 46980 5596
rect 47026 5584 47032 5636
rect 47084 5624 47090 5636
rect 47765 5627 47823 5633
rect 47765 5624 47777 5627
rect 47084 5596 47777 5624
rect 47084 5584 47090 5596
rect 47765 5593 47777 5596
rect 47811 5593 47823 5627
rect 47765 5587 47823 5593
rect 47210 5556 47216 5568
rect 46952 5528 47216 5556
rect 43809 5519 43867 5525
rect 47210 5516 47216 5528
rect 47268 5516 47274 5568
rect 48286 5556 48314 5664
rect 48424 5624 48452 5732
rect 50985 5729 50997 5732
rect 51031 5729 51043 5763
rect 50985 5723 51043 5729
rect 49697 5695 49755 5701
rect 49697 5661 49709 5695
rect 49743 5692 49755 5695
rect 49878 5692 49884 5704
rect 49743 5664 49884 5692
rect 49743 5661 49755 5664
rect 49697 5655 49755 5661
rect 49878 5652 49884 5664
rect 49936 5652 49942 5704
rect 50522 5652 50528 5704
rect 50580 5692 50586 5704
rect 50709 5695 50767 5701
rect 50709 5692 50721 5695
rect 50580 5664 50721 5692
rect 50580 5652 50586 5664
rect 50709 5661 50721 5664
rect 50755 5661 50767 5695
rect 50709 5655 50767 5661
rect 52012 5624 52040 5856
rect 52822 5652 52828 5704
rect 52880 5652 52886 5704
rect 53742 5652 53748 5704
rect 53800 5692 53806 5704
rect 54113 5695 54171 5701
rect 54113 5692 54125 5695
rect 53800 5664 54125 5692
rect 53800 5652 53806 5664
rect 54113 5661 54125 5664
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 54846 5652 54852 5704
rect 54904 5652 54910 5704
rect 55858 5652 55864 5704
rect 55916 5652 55922 5704
rect 55950 5652 55956 5704
rect 56008 5692 56014 5704
rect 56597 5695 56655 5701
rect 56597 5692 56609 5695
rect 56008 5664 56609 5692
rect 56008 5652 56014 5664
rect 56597 5661 56609 5664
rect 56643 5661 56655 5695
rect 56597 5655 56655 5661
rect 57330 5652 57336 5704
rect 57388 5652 57394 5704
rect 57790 5652 57796 5704
rect 57848 5692 57854 5704
rect 57885 5695 57943 5701
rect 57885 5692 57897 5695
rect 57848 5664 57897 5692
rect 57848 5652 57854 5664
rect 57885 5661 57897 5664
rect 57931 5661 57943 5695
rect 57885 5655 57943 5661
rect 48424 5596 52040 5624
rect 52362 5584 52368 5636
rect 52420 5624 52426 5636
rect 53285 5627 53343 5633
rect 53285 5624 53297 5627
rect 52420 5596 53297 5624
rect 52420 5584 52426 5596
rect 53285 5593 53297 5596
rect 53331 5624 53343 5627
rect 54478 5624 54484 5636
rect 53331 5596 54484 5624
rect 53331 5593 53343 5596
rect 53285 5587 53343 5593
rect 54478 5584 54484 5596
rect 54536 5624 54542 5636
rect 57701 5627 57759 5633
rect 57701 5624 57713 5627
rect 54536 5596 57713 5624
rect 54536 5584 54542 5596
rect 57701 5593 57713 5596
rect 57747 5593 57759 5627
rect 57701 5587 57759 5593
rect 48590 5556 48596 5568
rect 48286 5528 48596 5556
rect 48590 5516 48596 5528
rect 48648 5516 48654 5568
rect 48682 5516 48688 5568
rect 48740 5556 48746 5568
rect 49053 5559 49111 5565
rect 49053 5556 49065 5559
rect 48740 5528 49065 5556
rect 48740 5516 48746 5528
rect 49053 5525 49065 5528
rect 49099 5525 49111 5559
rect 49053 5519 49111 5525
rect 49786 5516 49792 5568
rect 49844 5556 49850 5568
rect 50157 5559 50215 5565
rect 50157 5556 50169 5559
rect 49844 5528 50169 5556
rect 49844 5516 49850 5528
rect 50157 5525 50169 5528
rect 50203 5525 50215 5559
rect 50157 5519 50215 5525
rect 51994 5516 52000 5568
rect 52052 5556 52058 5568
rect 52273 5559 52331 5565
rect 52273 5556 52285 5559
rect 52052 5528 52285 5556
rect 52052 5516 52058 5528
rect 52273 5525 52285 5528
rect 52319 5525 52331 5559
rect 52273 5519 52331 5525
rect 53558 5516 53564 5568
rect 53616 5516 53622 5568
rect 54202 5516 54208 5568
rect 54260 5556 54266 5568
rect 54297 5559 54355 5565
rect 54297 5556 54309 5559
rect 54260 5528 54309 5556
rect 54260 5516 54266 5528
rect 54297 5525 54309 5528
rect 54343 5525 54355 5559
rect 54297 5519 54355 5525
rect 54662 5516 54668 5568
rect 54720 5556 54726 5568
rect 55309 5559 55367 5565
rect 55309 5556 55321 5559
rect 54720 5528 55321 5556
rect 54720 5516 54726 5528
rect 55309 5525 55321 5528
rect 55355 5525 55367 5559
rect 55309 5519 55367 5525
rect 56042 5516 56048 5568
rect 56100 5516 56106 5568
rect 56778 5516 56784 5568
rect 56836 5516 56842 5568
rect 58158 5516 58164 5568
rect 58216 5556 58222 5568
rect 58529 5559 58587 5565
rect 58529 5556 58541 5559
rect 58216 5528 58541 5556
rect 58216 5516 58222 5528
rect 58529 5525 58541 5528
rect 58575 5525 58587 5559
rect 58529 5519 58587 5525
rect 1104 5466 59040 5488
rect 1104 5414 15394 5466
rect 15446 5414 15458 5466
rect 15510 5414 15522 5466
rect 15574 5414 15586 5466
rect 15638 5414 15650 5466
rect 15702 5414 29838 5466
rect 29890 5414 29902 5466
rect 29954 5414 29966 5466
rect 30018 5414 30030 5466
rect 30082 5414 30094 5466
rect 30146 5414 44282 5466
rect 44334 5414 44346 5466
rect 44398 5414 44410 5466
rect 44462 5414 44474 5466
rect 44526 5414 44538 5466
rect 44590 5414 58726 5466
rect 58778 5414 58790 5466
rect 58842 5414 58854 5466
rect 58906 5414 58918 5466
rect 58970 5414 58982 5466
rect 59034 5414 59040 5466
rect 1104 5392 59040 5414
rect 3050 5312 3056 5364
rect 3108 5312 3114 5364
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 4430 5352 4436 5364
rect 3660 5324 4436 5352
rect 3660 5312 3666 5324
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 5718 5312 5724 5364
rect 5776 5312 5782 5364
rect 6730 5352 6736 5364
rect 5920 5324 6736 5352
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 4525 5287 4583 5293
rect 4525 5284 4537 5287
rect 3936 5256 4537 5284
rect 3936 5244 3942 5256
rect 4525 5253 4537 5256
rect 4571 5284 4583 5287
rect 4614 5284 4620 5296
rect 4571 5256 4620 5284
rect 4571 5253 4583 5256
rect 4525 5247 4583 5253
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 1903 5188 5672 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 2958 5108 2964 5160
rect 3016 5108 3022 5160
rect 3694 5108 3700 5160
rect 3752 5108 3758 5160
rect 3786 5108 3792 5160
rect 3844 5108 3850 5160
rect 5074 5108 5080 5160
rect 5132 5108 5138 5160
rect 5644 5157 5672 5188
rect 5810 5176 5816 5228
rect 5868 5176 5874 5228
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5920 5148 5948 5324
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 10962 5352 10968 5364
rect 9447 5324 10968 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11977 5355 12035 5361
rect 11977 5352 11989 5355
rect 11204 5324 11989 5352
rect 11204 5312 11210 5324
rect 11977 5321 11989 5324
rect 12023 5321 12035 5355
rect 11977 5315 12035 5321
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 16114 5352 16120 5364
rect 15427 5324 16120 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 16114 5312 16120 5324
rect 16172 5312 16178 5364
rect 18230 5312 18236 5364
rect 18288 5312 18294 5364
rect 18322 5312 18328 5364
rect 18380 5312 18386 5364
rect 19702 5312 19708 5364
rect 19760 5312 19766 5364
rect 20073 5355 20131 5361
rect 20073 5321 20085 5355
rect 20119 5352 20131 5355
rect 21266 5352 21272 5364
rect 20119 5324 21272 5352
rect 20119 5321 20131 5324
rect 20073 5315 20131 5321
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 22373 5355 22431 5361
rect 22373 5321 22385 5355
rect 22419 5352 22431 5355
rect 23842 5352 23848 5364
rect 22419 5324 23848 5352
rect 22419 5321 22431 5324
rect 22373 5315 22431 5321
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 23934 5312 23940 5364
rect 23992 5312 23998 5364
rect 24302 5312 24308 5364
rect 24360 5312 24366 5364
rect 24394 5312 24400 5364
rect 24452 5312 24458 5364
rect 25409 5355 25467 5361
rect 25409 5321 25421 5355
rect 25455 5352 25467 5355
rect 25866 5352 25872 5364
rect 25455 5324 25872 5352
rect 25455 5321 25467 5324
rect 25409 5315 25467 5321
rect 25866 5312 25872 5324
rect 25924 5312 25930 5364
rect 26878 5352 26884 5364
rect 26712 5324 26884 5352
rect 8288 5287 8346 5293
rect 6380 5256 8064 5284
rect 6380 5228 6408 5256
rect 8036 5228 8064 5256
rect 8288 5253 8300 5287
rect 8334 5284 8346 5287
rect 8662 5284 8668 5296
rect 8334 5256 8668 5284
rect 8334 5253 8346 5256
rect 8288 5247 8346 5253
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 17120 5287 17178 5293
rect 13872 5256 17080 5284
rect 13872 5244 13878 5256
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6632 5219 6690 5225
rect 6632 5185 6644 5219
rect 6678 5216 6690 5219
rect 7006 5216 7012 5228
rect 6678 5188 7012 5216
rect 6678 5185 6690 5188
rect 6632 5179 6690 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9539 5188 9812 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 5675 5120 5948 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 4433 5083 4491 5089
rect 2240 5052 2774 5080
rect 2240 5021 2268 5052
rect 2225 5015 2283 5021
rect 2225 4981 2237 5015
rect 2271 4981 2283 5015
rect 2225 4975 2283 4981
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 2746 5012 2774 5052
rect 4433 5049 4445 5083
rect 4479 5080 4491 5083
rect 4479 5052 4752 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 4724 5024 4752 5052
rect 5718 5040 5724 5092
rect 5776 5080 5782 5092
rect 6380 5080 6408 5176
rect 9784 5160 9812 5188
rect 10502 5176 10508 5228
rect 10560 5225 10566 5228
rect 10560 5219 10588 5225
rect 10576 5185 10588 5219
rect 10560 5179 10588 5185
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11379 5188 11897 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 10560 5176 10566 5179
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 16022 5216 16028 5228
rect 13320 5188 16028 5216
rect 13320 5176 13326 5188
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 16224 5188 16865 5216
rect 16224 5160 16252 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 17052 5216 17080 5256
rect 17120 5253 17132 5287
rect 17166 5284 17178 5287
rect 17678 5284 17684 5296
rect 17166 5256 17684 5284
rect 17166 5253 17178 5256
rect 17120 5247 17178 5253
rect 17678 5244 17684 5256
rect 17736 5244 17742 5296
rect 19610 5284 19616 5296
rect 18616 5256 19616 5284
rect 17052 5188 17908 5216
rect 16853 5179 16911 5185
rect 9674 5108 9680 5160
rect 9732 5108 9738 5160
rect 9766 5108 9772 5160
rect 9824 5108 9830 5160
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 9876 5120 10425 5148
rect 5776 5052 6408 5080
rect 5776 5040 5782 5052
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 9876 5080 9904 5120
rect 10413 5117 10425 5120
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 11054 5148 11060 5160
rect 10735 5120 11060 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11054 5108 11060 5120
rect 11112 5108 11118 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11900 5120 12081 5148
rect 11900 5092 11928 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12894 5108 12900 5160
rect 12952 5108 12958 5160
rect 14274 5108 14280 5160
rect 14332 5108 14338 5160
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 14884 5120 15669 5148
rect 14884 5108 14890 5120
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 9364 5052 9904 5080
rect 10137 5083 10195 5089
rect 9364 5040 9370 5052
rect 10137 5049 10149 5083
rect 10183 5080 10195 5083
rect 10226 5080 10232 5092
rect 10183 5052 10232 5080
rect 10183 5049 10195 5052
rect 10137 5043 10195 5049
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 11882 5040 11888 5092
rect 11940 5040 11946 5092
rect 15672 5080 15700 5111
rect 16206 5108 16212 5160
rect 16264 5108 16270 5160
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 17880 5080 17908 5188
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 18616 5148 18644 5256
rect 19610 5244 19616 5256
rect 19668 5244 19674 5296
rect 19720 5284 19748 5312
rect 20441 5287 20499 5293
rect 20441 5284 20453 5287
rect 19720 5256 20453 5284
rect 20441 5253 20453 5256
rect 20487 5253 20499 5287
rect 20441 5247 20499 5253
rect 22732 5287 22790 5293
rect 22732 5253 22744 5287
rect 22778 5284 22790 5287
rect 23658 5284 23664 5296
rect 22778 5256 23664 5284
rect 22778 5253 22790 5256
rect 22732 5247 22790 5253
rect 23658 5244 23664 5256
rect 23716 5244 23722 5296
rect 26544 5287 26602 5293
rect 24228 5256 26464 5284
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5216 18751 5219
rect 19058 5216 19064 5228
rect 18739 5188 19064 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 19058 5176 19064 5188
rect 19116 5176 19122 5228
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19705 5219 19763 5225
rect 19705 5216 19717 5219
rect 19392 5188 19717 5216
rect 19392 5176 19398 5188
rect 19705 5185 19717 5188
rect 19751 5185 19763 5219
rect 19705 5179 19763 5185
rect 20162 5176 20168 5228
rect 20220 5216 20226 5228
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20220 5188 20545 5216
rect 20220 5176 20226 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 24228 5216 24256 5256
rect 25041 5219 25099 5225
rect 25041 5216 25053 5219
rect 20533 5179 20591 5185
rect 20732 5188 24256 5216
rect 24504 5188 25053 5216
rect 20732 5160 20760 5188
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 18012 5120 18797 5148
rect 18012 5108 18018 5120
rect 18785 5117 18797 5120
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 18877 5151 18935 5157
rect 18877 5117 18889 5151
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 19794 5148 19800 5160
rect 19567 5120 19800 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 18690 5080 18696 5092
rect 15672 5052 16896 5080
rect 17880 5052 18696 5080
rect 4338 5012 4344 5024
rect 2746 4984 4344 5012
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 4706 4972 4712 5024
rect 4764 4972 4770 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6730 5012 6736 5024
rect 6227 4984 6736 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10870 5012 10876 5024
rect 9732 4984 10876 5012
rect 9732 4972 9738 4984
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 12342 4972 12348 5024
rect 12400 4972 12406 5024
rect 13446 4972 13452 5024
rect 13504 5012 13510 5024
rect 14090 5012 14096 5024
rect 13504 4984 14096 5012
rect 13504 4972 13510 4984
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14608 4984 14933 5012
rect 14608 4972 14614 4984
rect 14921 4981 14933 4984
rect 14967 4981 14979 5015
rect 14921 4975 14979 4981
rect 15838 4972 15844 5024
rect 15896 4972 15902 5024
rect 16868 5012 16896 5052
rect 18690 5040 18696 5052
rect 18748 5040 18754 5092
rect 18892 5080 18920 5111
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 20349 5151 20407 5157
rect 20349 5117 20361 5151
rect 20395 5148 20407 5151
rect 20714 5148 20720 5160
rect 20395 5120 20720 5148
rect 20395 5117 20407 5120
rect 20349 5111 20407 5117
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 21082 5108 21088 5160
rect 21140 5108 21146 5160
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 24504 5157 24532 5188
rect 25041 5185 25053 5188
rect 25087 5185 25099 5219
rect 26436 5216 26464 5256
rect 26544 5253 26556 5287
rect 26590 5284 26602 5287
rect 26712 5284 26740 5324
rect 26878 5312 26884 5324
rect 26936 5312 26942 5364
rect 27246 5312 27252 5364
rect 27304 5312 27310 5364
rect 27890 5312 27896 5364
rect 27948 5352 27954 5364
rect 27985 5355 28043 5361
rect 27985 5352 27997 5355
rect 27948 5324 27997 5352
rect 27948 5312 27954 5324
rect 27985 5321 27997 5324
rect 28031 5352 28043 5355
rect 28442 5352 28448 5364
rect 28031 5324 28448 5352
rect 28031 5321 28043 5324
rect 27985 5315 28043 5321
rect 28442 5312 28448 5324
rect 28500 5352 28506 5364
rect 28721 5355 28779 5361
rect 28721 5352 28733 5355
rect 28500 5324 28733 5352
rect 28500 5312 28506 5324
rect 28721 5321 28733 5324
rect 28767 5321 28779 5355
rect 28721 5315 28779 5321
rect 35802 5312 35808 5364
rect 35860 5312 35866 5364
rect 36906 5312 36912 5364
rect 36964 5352 36970 5364
rect 40865 5355 40923 5361
rect 40865 5352 40877 5355
rect 36964 5324 40877 5352
rect 36964 5312 36970 5324
rect 40865 5321 40877 5324
rect 40911 5321 40923 5355
rect 40865 5315 40923 5321
rect 41049 5355 41107 5361
rect 41049 5321 41061 5355
rect 41095 5352 41107 5355
rect 41322 5352 41328 5364
rect 41095 5324 41328 5352
rect 41095 5321 41107 5324
rect 41049 5315 41107 5321
rect 27908 5284 27936 5312
rect 26590 5256 26740 5284
rect 26804 5256 27936 5284
rect 29457 5287 29515 5293
rect 26590 5253 26602 5256
rect 26544 5247 26602 5253
rect 26804 5225 26832 5256
rect 29457 5253 29469 5287
rect 29503 5284 29515 5287
rect 35820 5284 35848 5312
rect 37553 5287 37611 5293
rect 37553 5284 37565 5287
rect 29503 5256 30972 5284
rect 35820 5256 37565 5284
rect 29503 5253 29515 5256
rect 29457 5247 29515 5253
rect 26789 5219 26847 5225
rect 26436 5188 26740 5216
rect 25041 5179 25099 5185
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22152 5120 22477 5148
rect 22152 5108 22158 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 24489 5151 24547 5157
rect 24489 5148 24501 5151
rect 22465 5111 22523 5117
rect 23768 5120 24501 5148
rect 22370 5080 22376 5092
rect 18809 5052 22376 5080
rect 18809 5012 18837 5052
rect 22370 5040 22376 5052
rect 22428 5040 22434 5092
rect 23768 5024 23796 5120
rect 24489 5117 24501 5120
rect 24535 5117 24547 5151
rect 24489 5111 24547 5117
rect 24946 5108 24952 5160
rect 25004 5108 25010 5160
rect 26712 5148 26740 5188
rect 26789 5185 26801 5219
rect 26835 5185 26847 5219
rect 26789 5179 26847 5185
rect 27338 5176 27344 5228
rect 27396 5176 27402 5228
rect 27522 5176 27528 5228
rect 27580 5216 27586 5228
rect 29472 5216 29500 5247
rect 30944 5228 30972 5256
rect 37553 5253 37565 5256
rect 37599 5284 37611 5287
rect 37734 5284 37740 5296
rect 37599 5256 37740 5284
rect 37599 5253 37611 5256
rect 37553 5247 37611 5253
rect 37734 5244 37740 5256
rect 37792 5284 37798 5296
rect 37792 5256 38654 5284
rect 37792 5244 37798 5256
rect 27580 5188 29500 5216
rect 30193 5219 30251 5225
rect 27580 5176 27586 5188
rect 30193 5185 30205 5219
rect 30239 5216 30251 5219
rect 30558 5216 30564 5228
rect 30239 5188 30564 5216
rect 30239 5185 30251 5188
rect 30193 5179 30251 5185
rect 30558 5176 30564 5188
rect 30616 5176 30622 5228
rect 30926 5176 30932 5228
rect 30984 5176 30990 5228
rect 27157 5151 27215 5157
rect 26712 5120 27016 5148
rect 23845 5083 23903 5089
rect 23845 5049 23857 5083
rect 23891 5080 23903 5083
rect 24964 5080 24992 5108
rect 23891 5052 24992 5080
rect 26988 5080 27016 5120
rect 27157 5117 27169 5151
rect 27203 5148 27215 5151
rect 27430 5148 27436 5160
rect 27203 5120 27436 5148
rect 27203 5117 27215 5120
rect 27157 5111 27215 5117
rect 27430 5108 27436 5120
rect 27488 5148 27494 5160
rect 28353 5151 28411 5157
rect 28353 5148 28365 5151
rect 27488 5120 28365 5148
rect 27488 5108 27494 5120
rect 28353 5117 28365 5120
rect 28399 5117 28411 5151
rect 28353 5111 28411 5117
rect 30374 5108 30380 5160
rect 30432 5108 30438 5160
rect 31294 5148 31300 5160
rect 30484 5120 31300 5148
rect 30484 5080 30512 5120
rect 31294 5108 31300 5120
rect 31352 5108 31358 5160
rect 35986 5108 35992 5160
rect 36044 5148 36050 5160
rect 36357 5151 36415 5157
rect 36357 5148 36369 5151
rect 36044 5120 36369 5148
rect 36044 5108 36050 5120
rect 36357 5117 36369 5120
rect 36403 5117 36415 5151
rect 36357 5111 36415 5117
rect 38286 5108 38292 5160
rect 38344 5108 38350 5160
rect 33778 5080 33784 5092
rect 26988 5052 30512 5080
rect 31680 5052 33784 5080
rect 23891 5049 23903 5052
rect 23845 5043 23903 5049
rect 16868 4984 18837 5012
rect 20898 4972 20904 5024
rect 20956 4972 20962 5024
rect 21634 4972 21640 5024
rect 21692 4972 21698 5024
rect 23750 4972 23756 5024
rect 23808 4972 23814 5024
rect 27614 4972 27620 5024
rect 27672 5012 27678 5024
rect 27709 5015 27767 5021
rect 27709 5012 27721 5015
rect 27672 4984 27721 5012
rect 27672 4972 27678 4984
rect 27709 4981 27721 4984
rect 27755 4981 27767 5015
rect 27709 4975 27767 4981
rect 29454 4972 29460 5024
rect 29512 5012 29518 5024
rect 29549 5015 29607 5021
rect 29549 5012 29561 5015
rect 29512 4984 29561 5012
rect 29512 4972 29518 4984
rect 29549 4981 29561 4984
rect 29595 4981 29607 5015
rect 29549 4975 29607 4981
rect 31018 4972 31024 5024
rect 31076 4972 31082 5024
rect 31570 4972 31576 5024
rect 31628 5012 31634 5024
rect 31680 5021 31708 5052
rect 33778 5040 33784 5052
rect 33836 5040 33842 5092
rect 35710 5040 35716 5092
rect 35768 5080 35774 5092
rect 38626 5080 38654 5256
rect 39209 5151 39267 5157
rect 39209 5117 39221 5151
rect 39255 5148 39267 5151
rect 39482 5148 39488 5160
rect 39255 5120 39488 5148
rect 39255 5117 39267 5120
rect 39209 5111 39267 5117
rect 39482 5108 39488 5120
rect 39540 5108 39546 5160
rect 39666 5108 39672 5160
rect 39724 5148 39730 5160
rect 39853 5151 39911 5157
rect 39853 5148 39865 5151
rect 39724 5120 39865 5148
rect 39724 5108 39730 5120
rect 39853 5117 39865 5120
rect 39899 5117 39911 5151
rect 40880 5148 40908 5315
rect 41322 5312 41328 5324
rect 41380 5312 41386 5364
rect 41506 5312 41512 5364
rect 41564 5352 41570 5364
rect 43901 5355 43959 5361
rect 41564 5324 43024 5352
rect 41564 5312 41570 5324
rect 41874 5244 41880 5296
rect 41932 5284 41938 5296
rect 42061 5287 42119 5293
rect 42061 5284 42073 5287
rect 41932 5256 42073 5284
rect 41932 5244 41938 5256
rect 42061 5253 42073 5256
rect 42107 5253 42119 5287
rect 42996 5284 43024 5324
rect 43901 5321 43913 5355
rect 43947 5352 43959 5355
rect 44174 5352 44180 5364
rect 43947 5324 44180 5352
rect 43947 5321 43959 5324
rect 43901 5315 43959 5321
rect 44174 5312 44180 5324
rect 44232 5312 44238 5364
rect 46750 5312 46756 5364
rect 46808 5312 46814 5364
rect 51166 5312 51172 5364
rect 51224 5352 51230 5364
rect 53193 5355 53251 5361
rect 53193 5352 53205 5355
rect 51224 5324 53205 5352
rect 51224 5312 51230 5324
rect 53193 5321 53205 5324
rect 53239 5321 53251 5355
rect 53193 5315 53251 5321
rect 54662 5312 54668 5364
rect 54720 5312 54726 5364
rect 55033 5355 55091 5361
rect 55033 5321 55045 5355
rect 55079 5321 55091 5355
rect 55033 5315 55091 5321
rect 55125 5355 55183 5361
rect 55125 5321 55137 5355
rect 55171 5352 55183 5355
rect 55858 5352 55864 5364
rect 55171 5324 55864 5352
rect 55171 5321 55183 5324
rect 55125 5315 55183 5321
rect 43254 5284 43260 5296
rect 42996 5256 43260 5284
rect 42061 5247 42119 5253
rect 43254 5244 43260 5256
rect 43312 5284 43318 5296
rect 44361 5287 44419 5293
rect 44361 5284 44373 5287
rect 43312 5256 44373 5284
rect 43312 5244 43318 5256
rect 44361 5253 44373 5256
rect 44407 5284 44419 5287
rect 45097 5287 45155 5293
rect 45097 5284 45109 5287
rect 44407 5256 45109 5284
rect 44407 5253 44419 5256
rect 44361 5247 44419 5253
rect 45097 5253 45109 5256
rect 45143 5253 45155 5287
rect 45465 5287 45523 5293
rect 45465 5284 45477 5287
rect 45097 5247 45155 5253
rect 45204 5256 45477 5284
rect 41417 5219 41475 5225
rect 41417 5185 41429 5219
rect 41463 5216 41475 5219
rect 43073 5219 43131 5225
rect 43073 5216 43085 5219
rect 41463 5188 43085 5216
rect 41463 5185 41475 5188
rect 41417 5179 41475 5185
rect 43073 5185 43085 5188
rect 43119 5216 43131 5219
rect 43806 5216 43812 5228
rect 43119 5188 43812 5216
rect 43119 5185 43131 5188
rect 43073 5179 43131 5185
rect 43806 5176 43812 5188
rect 43864 5176 43870 5228
rect 44269 5219 44327 5225
rect 44269 5216 44281 5219
rect 44192 5188 44281 5216
rect 41693 5151 41751 5157
rect 41693 5148 41705 5151
rect 40880 5120 41705 5148
rect 39853 5111 39911 5117
rect 41693 5117 41705 5120
rect 41739 5117 41751 5151
rect 41693 5111 41751 5117
rect 41708 5080 41736 5111
rect 42426 5108 42432 5160
rect 42484 5108 42490 5160
rect 42886 5108 42892 5160
rect 42944 5148 42950 5160
rect 43717 5151 43775 5157
rect 43717 5148 43729 5151
rect 42944 5120 43729 5148
rect 42944 5108 42950 5120
rect 43717 5117 43729 5120
rect 43763 5117 43775 5151
rect 43717 5111 43775 5117
rect 42610 5080 42616 5092
rect 35768 5052 36676 5080
rect 38626 5052 38884 5080
rect 35768 5040 35774 5052
rect 36648 5024 36676 5052
rect 38856 5024 38884 5052
rect 40512 5052 41368 5080
rect 41708 5052 42616 5080
rect 31665 5015 31723 5021
rect 31665 5012 31677 5015
rect 31628 4984 31677 5012
rect 31628 4972 31634 4984
rect 31665 4981 31677 4984
rect 31711 4981 31723 5015
rect 31665 4975 31723 4981
rect 32398 4972 32404 5024
rect 32456 5012 32462 5024
rect 33413 5015 33471 5021
rect 33413 5012 33425 5015
rect 32456 4984 33425 5012
rect 32456 4972 32462 4984
rect 33413 4981 33425 4984
rect 33459 5012 33471 5015
rect 34882 5012 34888 5024
rect 33459 4984 34888 5012
rect 33459 4981 33471 4984
rect 33413 4975 33471 4981
rect 34882 4972 34888 4984
rect 34940 4972 34946 5024
rect 35802 4972 35808 5024
rect 35860 4972 35866 5024
rect 36630 4972 36636 5024
rect 36688 4972 36694 5024
rect 37734 4972 37740 5024
rect 37792 4972 37798 5024
rect 38562 4972 38568 5024
rect 38620 4972 38626 5024
rect 38838 4972 38844 5024
rect 38896 4972 38902 5024
rect 39298 4972 39304 5024
rect 39356 4972 39362 5024
rect 40034 4972 40040 5024
rect 40092 5012 40098 5024
rect 40512 5021 40540 5052
rect 40497 5015 40555 5021
rect 40497 5012 40509 5015
rect 40092 4984 40509 5012
rect 40092 4972 40098 4984
rect 40497 4981 40509 4984
rect 40543 4981 40555 5015
rect 41340 5012 41368 5052
rect 42610 5040 42616 5052
rect 42668 5040 42674 5092
rect 44192 5080 44220 5188
rect 44269 5185 44281 5188
rect 44315 5216 44327 5219
rect 45204 5216 45232 5256
rect 45465 5253 45477 5256
rect 45511 5253 45523 5287
rect 45465 5247 45523 5253
rect 49237 5287 49295 5293
rect 49237 5253 49249 5287
rect 49283 5284 49295 5287
rect 49602 5284 49608 5296
rect 49283 5256 49608 5284
rect 49283 5253 49295 5256
rect 49237 5247 49295 5253
rect 49602 5244 49608 5256
rect 49660 5244 49666 5296
rect 50985 5287 51043 5293
rect 50985 5253 50997 5287
rect 51031 5284 51043 5287
rect 51258 5284 51264 5296
rect 51031 5256 51264 5284
rect 51031 5253 51043 5256
rect 50985 5247 51043 5253
rect 44315 5188 45232 5216
rect 44315 5185 44327 5188
rect 44269 5179 44327 5185
rect 45278 5176 45284 5228
rect 45336 5176 45342 5228
rect 48705 5219 48763 5225
rect 48705 5185 48717 5219
rect 48751 5216 48763 5219
rect 48866 5216 48872 5228
rect 48751 5188 48872 5216
rect 48751 5185 48763 5188
rect 48705 5179 48763 5185
rect 48866 5176 48872 5188
rect 48924 5176 48930 5228
rect 48961 5219 49019 5225
rect 48961 5185 48973 5219
rect 49007 5216 49019 5219
rect 51000 5216 51028 5247
rect 51258 5244 51264 5256
rect 51316 5244 51322 5296
rect 55048 5284 55076 5315
rect 55858 5312 55864 5324
rect 55916 5312 55922 5364
rect 55950 5312 55956 5364
rect 56008 5312 56014 5364
rect 56134 5312 56140 5364
rect 56192 5352 56198 5364
rect 56192 5324 56548 5352
rect 56192 5312 56198 5324
rect 55968 5284 55996 5312
rect 55048 5256 55996 5284
rect 56042 5244 56048 5296
rect 56100 5284 56106 5296
rect 56238 5287 56296 5293
rect 56238 5284 56250 5287
rect 56100 5256 56250 5284
rect 56100 5244 56106 5256
rect 56238 5253 56250 5256
rect 56284 5253 56296 5287
rect 56238 5247 56296 5253
rect 56520 5228 56548 5324
rect 56686 5312 56692 5364
rect 56744 5352 56750 5364
rect 57517 5355 57575 5361
rect 57517 5352 57529 5355
rect 56744 5324 57529 5352
rect 56744 5312 56750 5324
rect 57517 5321 57529 5324
rect 57563 5321 57575 5355
rect 57517 5315 57575 5321
rect 57882 5312 57888 5364
rect 57940 5312 57946 5364
rect 51813 5219 51871 5225
rect 51813 5216 51825 5219
rect 49007 5188 51028 5216
rect 51092 5188 51825 5216
rect 49007 5185 49019 5188
rect 48961 5179 49019 5185
rect 51092 5160 51120 5188
rect 51813 5185 51825 5188
rect 51859 5216 51871 5219
rect 51902 5216 51908 5228
rect 51859 5188 51908 5216
rect 51859 5185 51871 5188
rect 51813 5179 51871 5185
rect 51902 5176 51908 5188
rect 51960 5176 51966 5228
rect 53282 5176 53288 5228
rect 53340 5176 53346 5228
rect 54018 5176 54024 5228
rect 54076 5216 54082 5228
rect 54573 5219 54631 5225
rect 54573 5216 54585 5219
rect 54076 5188 54585 5216
rect 54076 5176 54082 5188
rect 54573 5185 54585 5188
rect 54619 5216 54631 5219
rect 55214 5216 55220 5228
rect 54619 5188 55220 5216
rect 54619 5185 54631 5188
rect 54573 5179 54631 5185
rect 55214 5176 55220 5188
rect 55272 5176 55278 5228
rect 56502 5176 56508 5228
rect 56560 5176 56566 5228
rect 57701 5219 57759 5225
rect 57701 5185 57713 5219
rect 57747 5216 57759 5219
rect 57900 5216 57928 5312
rect 57747 5188 57928 5216
rect 57747 5185 57759 5188
rect 57701 5179 57759 5185
rect 44545 5151 44603 5157
rect 44545 5117 44557 5151
rect 44591 5117 44603 5151
rect 44545 5111 44603 5117
rect 42812 5052 44220 5080
rect 42812 5024 42840 5052
rect 41414 5012 41420 5024
rect 41340 4984 41420 5012
rect 40497 4975 40555 4981
rect 41414 4972 41420 4984
rect 41472 5012 41478 5024
rect 42702 5012 42708 5024
rect 41472 4984 42708 5012
rect 41472 4972 41478 4984
rect 42702 4972 42708 4984
rect 42760 4972 42766 5024
rect 42794 4972 42800 5024
rect 42852 4972 42858 5024
rect 43162 4972 43168 5024
rect 43220 4972 43226 5024
rect 44560 5012 44588 5111
rect 44726 5108 44732 5160
rect 44784 5148 44790 5160
rect 46017 5151 46075 5157
rect 46017 5148 46029 5151
rect 44784 5120 46029 5148
rect 44784 5108 44790 5120
rect 46017 5117 46029 5120
rect 46063 5117 46075 5151
rect 46017 5111 46075 5117
rect 47397 5151 47455 5157
rect 47397 5117 47409 5151
rect 47443 5117 47455 5151
rect 47397 5111 47455 5117
rect 47412 5080 47440 5111
rect 51074 5108 51080 5160
rect 51132 5108 51138 5160
rect 51350 5108 51356 5160
rect 51408 5148 51414 5160
rect 51629 5151 51687 5157
rect 51629 5148 51641 5151
rect 51408 5120 51641 5148
rect 51408 5108 51414 5120
rect 51629 5117 51641 5120
rect 51675 5117 51687 5151
rect 51629 5111 51687 5117
rect 52362 5108 52368 5160
rect 52420 5108 52426 5160
rect 53190 5108 53196 5160
rect 53248 5148 53254 5160
rect 53469 5151 53527 5157
rect 53469 5148 53481 5151
rect 53248 5120 53481 5148
rect 53248 5108 53254 5120
rect 53469 5117 53481 5120
rect 53515 5117 53527 5151
rect 53469 5111 53527 5117
rect 54478 5108 54484 5160
rect 54536 5108 54542 5160
rect 56686 5108 56692 5160
rect 56744 5148 56750 5160
rect 57149 5151 57207 5157
rect 57149 5148 57161 5151
rect 56744 5120 57161 5148
rect 56744 5108 56750 5120
rect 57149 5117 57161 5120
rect 57195 5117 57207 5151
rect 57149 5111 57207 5117
rect 57882 5108 57888 5160
rect 57940 5148 57946 5160
rect 58437 5151 58495 5157
rect 58437 5148 58449 5151
rect 57940 5120 58449 5148
rect 57940 5108 57946 5120
rect 58437 5117 58449 5120
rect 58483 5117 58495 5151
rect 58437 5111 58495 5117
rect 47581 5083 47639 5089
rect 47581 5080 47593 5083
rect 47412 5052 47593 5080
rect 47581 5049 47593 5052
rect 47627 5049 47639 5083
rect 47581 5043 47639 5049
rect 55122 5040 55128 5092
rect 55180 5080 55186 5092
rect 55180 5052 55444 5080
rect 55180 5040 55186 5052
rect 45005 5015 45063 5021
rect 45005 5012 45017 5015
rect 44560 4984 45017 5012
rect 45005 4981 45017 4984
rect 45051 5012 45063 5015
rect 46014 5012 46020 5024
rect 45051 4984 46020 5012
rect 45051 4981 45063 4984
rect 45005 4975 45063 4981
rect 46014 4972 46020 4984
rect 46072 4972 46078 5024
rect 46566 4972 46572 5024
rect 46624 4972 46630 5024
rect 50706 4972 50712 5024
rect 50764 5012 50770 5024
rect 51077 5015 51135 5021
rect 51077 5012 51089 5015
rect 50764 4984 51089 5012
rect 50764 4972 50770 4984
rect 51077 4981 51089 4984
rect 51123 4981 51135 5015
rect 51077 4975 51135 4981
rect 52914 4972 52920 5024
rect 52972 4972 52978 5024
rect 54113 5015 54171 5021
rect 54113 4981 54125 5015
rect 54159 5012 54171 5015
rect 55306 5012 55312 5024
rect 54159 4984 55312 5012
rect 54159 4981 54171 4984
rect 54113 4975 54171 4981
rect 55306 4972 55312 4984
rect 55364 4972 55370 5024
rect 55416 5012 55444 5052
rect 56597 5015 56655 5021
rect 56597 5012 56609 5015
rect 55416 4984 56609 5012
rect 56597 4981 56609 4984
rect 56643 4981 56655 5015
rect 56597 4975 56655 4981
rect 57698 4972 57704 5024
rect 57756 5012 57762 5024
rect 57885 5015 57943 5021
rect 57885 5012 57897 5015
rect 57756 4984 57897 5012
rect 57756 4972 57762 4984
rect 57885 4981 57897 4984
rect 57931 4981 57943 5015
rect 57885 4975 57943 4981
rect 1104 4922 58880 4944
rect 1104 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 22616 4922
rect 22668 4870 22680 4922
rect 22732 4870 22744 4922
rect 22796 4870 22808 4922
rect 22860 4870 22872 4922
rect 22924 4870 37060 4922
rect 37112 4870 37124 4922
rect 37176 4870 37188 4922
rect 37240 4870 37252 4922
rect 37304 4870 37316 4922
rect 37368 4870 51504 4922
rect 51556 4870 51568 4922
rect 51620 4870 51632 4922
rect 51684 4870 51696 4922
rect 51748 4870 51760 4922
rect 51812 4870 58880 4922
rect 1104 4848 58880 4870
rect 2130 4808 2136 4820
rect 1872 4780 2136 4808
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 1872 4681 1900 4780
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 3786 4808 3792 4820
rect 3283 4780 3792 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 7009 4811 7067 4817
rect 4540 4780 5856 4808
rect 3878 4740 3884 4752
rect 3804 4712 3884 4740
rect 3804 4681 3832 4712
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4430 4700 4436 4752
rect 4488 4700 4494 4752
rect 1857 4675 1915 4681
rect 1857 4672 1869 4675
rect 1728 4644 1869 4672
rect 1728 4632 1734 4644
rect 1857 4641 1869 4644
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 3789 4675 3847 4681
rect 3789 4641 3801 4675
rect 3835 4641 3847 4675
rect 4540 4672 4568 4780
rect 3789 4635 3847 4641
rect 3896 4644 4568 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 3896 4604 3924 4644
rect 4798 4632 4804 4684
rect 4856 4681 4862 4684
rect 4856 4675 4884 4681
rect 4872 4641 4884 4675
rect 4856 4635 4884 4641
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5828 4672 5856 4780
rect 7009 4777 7021 4811
rect 7055 4808 7067 4811
rect 7558 4808 7564 4820
rect 7055 4780 7564 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 11514 4808 11520 4820
rect 10888 4780 11520 4808
rect 10042 4740 10048 4752
rect 6380 4712 10048 4740
rect 6380 4681 6408 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5031 4644 5580 4672
rect 5828 4644 6377 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 4856 4632 4862 4635
rect 1811 4576 3924 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 2124 4539 2182 4545
rect 2124 4505 2136 4539
rect 2170 4536 2182 4539
rect 2314 4536 2320 4548
rect 2170 4508 2320 4536
rect 2170 4505 2182 4508
rect 2124 4499 2182 4505
rect 2314 4496 2320 4508
rect 2372 4496 2378 4548
rect 2682 4496 2688 4548
rect 2740 4536 2746 4548
rect 3421 4539 3479 4545
rect 3421 4536 3433 4539
rect 2740 4508 3433 4536
rect 2740 4496 2746 4508
rect 3421 4505 3433 4508
rect 3467 4505 3479 4539
rect 5552 4536 5580 4644
rect 6365 4641 6377 4644
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 8846 4672 8852 4684
rect 7515 4644 8852 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 10226 4672 10232 4684
rect 9171 4644 10232 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10594 4632 10600 4684
rect 10652 4632 10658 4684
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 5810 4604 5816 4616
rect 5675 4576 5816 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 6546 4604 6552 4616
rect 6052 4576 6552 4604
rect 6052 4564 6058 4576
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 7190 4604 7196 4616
rect 6687 4576 7196 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 7984 4576 8125 4604
rect 7984 4564 7990 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8220 4576 9674 4604
rect 5902 4536 5908 4548
rect 5552 4508 5908 4536
rect 3421 4499 3479 4505
rect 5902 4496 5908 4508
rect 5960 4496 5966 4548
rect 6086 4496 6092 4548
rect 6144 4536 6150 4548
rect 8220 4536 8248 4576
rect 6144 4508 8248 4536
rect 8757 4539 8815 4545
rect 6144 4496 6150 4508
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 9306 4536 9312 4548
rect 8803 4508 9312 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 9646 4536 9674 4576
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 10888 4613 10916 4780
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14148 4780 14933 4808
rect 14148 4768 14154 4780
rect 14921 4777 14933 4780
rect 14967 4808 14979 4811
rect 15010 4808 15016 4820
rect 14967 4780 15016 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 15010 4768 15016 4780
rect 15068 4808 15074 4820
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15068 4780 15761 4808
rect 15068 4768 15074 4780
rect 15749 4777 15761 4780
rect 15795 4808 15807 4811
rect 16206 4808 16212 4820
rect 15795 4780 16212 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 17586 4768 17592 4820
rect 17644 4768 17650 4820
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19760 4780 19809 4808
rect 19760 4768 19766 4780
rect 19797 4777 19809 4780
rect 19843 4808 19855 4811
rect 20622 4808 20628 4820
rect 19843 4780 20628 4808
rect 19843 4777 19855 4780
rect 19797 4771 19855 4777
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 23842 4768 23848 4820
rect 23900 4768 23906 4820
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 26237 4811 26295 4817
rect 24268 4780 26004 4808
rect 24268 4768 24274 4780
rect 10962 4700 10968 4752
rect 11020 4700 11026 4752
rect 11241 4743 11299 4749
rect 11241 4709 11253 4743
rect 11287 4740 11299 4743
rect 14645 4743 14703 4749
rect 11287 4712 11928 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 10980 4536 11008 4700
rect 11900 4681 11928 4712
rect 14645 4709 14657 4743
rect 14691 4740 14703 4743
rect 16298 4740 16304 4752
rect 14691 4712 16304 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 16298 4700 16304 4712
rect 16356 4700 16362 4752
rect 23477 4743 23535 4749
rect 23477 4709 23489 4743
rect 23523 4740 23535 4743
rect 23523 4712 23612 4740
rect 23523 4709 23535 4712
rect 23477 4703 23535 4709
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4641 11943 4675
rect 11885 4635 11943 4641
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12492 4644 12541 4672
rect 12492 4632 12498 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 16080 4644 18245 4672
rect 16080 4632 16086 4644
rect 18233 4641 18245 4644
rect 18279 4672 18291 4675
rect 21542 4672 21548 4684
rect 18279 4644 21548 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 21542 4632 21548 4644
rect 21600 4632 21606 4684
rect 23584 4681 23612 4712
rect 23569 4675 23627 4681
rect 23569 4641 23581 4675
rect 23615 4641 23627 4675
rect 23569 4635 23627 4641
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4604 13231 4607
rect 13262 4604 13268 4616
rect 13219 4576 13268 4604
rect 13219 4573 13231 4576
rect 13173 4567 13231 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 13906 4564 13912 4616
rect 13964 4564 13970 4616
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14056 4576 15117 4604
rect 14056 4564 14062 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 17034 4564 17040 4616
rect 17092 4604 17098 4616
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 17092 4576 17233 4604
rect 17092 4564 17098 4576
rect 17221 4573 17233 4576
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 18414 4564 18420 4616
rect 18472 4564 18478 4616
rect 20438 4564 20444 4616
rect 20496 4564 20502 4616
rect 21174 4564 21180 4616
rect 21232 4564 21238 4616
rect 21450 4564 21456 4616
rect 21508 4564 21514 4616
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 22186 4564 22192 4616
rect 22244 4604 22250 4616
rect 22353 4607 22411 4613
rect 22353 4604 22365 4607
rect 22244 4576 22365 4604
rect 22244 4564 22250 4576
rect 22353 4573 22365 4576
rect 22399 4573 22411 4607
rect 23860 4604 23888 4768
rect 24854 4740 24860 4752
rect 24596 4712 24860 4740
rect 24394 4632 24400 4684
rect 24452 4632 24458 4684
rect 24596 4681 24624 4712
rect 24854 4700 24860 4712
rect 24912 4700 24918 4752
rect 24581 4675 24639 4681
rect 24581 4641 24593 4675
rect 24627 4641 24639 4675
rect 25041 4675 25099 4681
rect 25041 4672 25053 4675
rect 24581 4635 24639 4641
rect 24688 4644 25053 4672
rect 24688 4604 24716 4644
rect 25041 4641 25053 4644
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25317 4675 25375 4681
rect 25317 4672 25329 4675
rect 25188 4644 25329 4672
rect 25188 4632 25194 4644
rect 25317 4641 25329 4644
rect 25363 4641 25375 4675
rect 25317 4635 25375 4641
rect 25455 4675 25513 4681
rect 25455 4641 25467 4675
rect 25501 4672 25513 4675
rect 25976 4672 26004 4780
rect 26237 4777 26249 4811
rect 26283 4808 26295 4811
rect 27338 4808 27344 4820
rect 26283 4780 27344 4808
rect 26283 4777 26295 4780
rect 26237 4771 26295 4777
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 28442 4768 28448 4820
rect 28500 4768 28506 4820
rect 30466 4808 30472 4820
rect 29748 4780 30472 4808
rect 25501 4644 26004 4672
rect 26697 4675 26755 4681
rect 25501 4641 25513 4644
rect 25455 4635 25513 4641
rect 26697 4641 26709 4675
rect 26743 4672 26755 4675
rect 27522 4672 27528 4684
rect 26743 4644 27528 4672
rect 26743 4641 26755 4644
rect 26697 4635 26755 4641
rect 27522 4632 27528 4644
rect 27580 4632 27586 4684
rect 29748 4681 29776 4780
rect 30466 4768 30472 4780
rect 30524 4768 30530 4820
rect 31294 4768 31300 4820
rect 31352 4808 31358 4820
rect 31352 4780 31754 4808
rect 31352 4768 31358 4780
rect 30190 4700 30196 4752
rect 30248 4700 30254 4752
rect 29733 4675 29791 4681
rect 29733 4641 29745 4675
rect 29779 4641 29791 4675
rect 30586 4675 30644 4681
rect 30586 4672 30598 4675
rect 29733 4635 29791 4641
rect 29840 4644 30598 4672
rect 23860 4576 24716 4604
rect 22353 4567 22411 4573
rect 25590 4564 25596 4616
rect 25648 4564 25654 4616
rect 27433 4607 27491 4613
rect 27433 4573 27445 4607
rect 27479 4604 27491 4607
rect 27706 4604 27712 4616
rect 27479 4576 27712 4604
rect 27479 4573 27491 4576
rect 27433 4567 27491 4573
rect 27706 4564 27712 4576
rect 27764 4564 27770 4616
rect 28074 4564 28080 4616
rect 28132 4564 28138 4616
rect 29362 4564 29368 4616
rect 29420 4564 29426 4616
rect 29549 4607 29607 4613
rect 29549 4573 29561 4607
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 9646 4508 11008 4536
rect 15289 4539 15347 4545
rect 15289 4505 15301 4539
rect 15335 4536 15347 4539
rect 16574 4536 16580 4548
rect 15335 4508 16580 4536
rect 15335 4505 15347 4508
rect 15289 4499 15347 4505
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 18690 4496 18696 4548
rect 18748 4536 18754 4548
rect 23750 4536 23756 4548
rect 18748 4508 23756 4536
rect 18748 4496 18754 4508
rect 23750 4496 23756 4508
rect 23808 4496 23814 4548
rect 3513 4471 3571 4477
rect 3513 4437 3525 4471
rect 3559 4468 3571 4471
rect 3602 4468 3608 4480
rect 3559 4440 3608 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8570 4468 8576 4480
rect 8067 4440 8576 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 9674 4428 9680 4480
rect 9732 4428 9738 4480
rect 10410 4428 10416 4480
rect 10468 4428 10474 4480
rect 10778 4428 10784 4480
rect 10836 4428 10842 4480
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 11333 4471 11391 4477
rect 11333 4468 11345 4471
rect 11296 4440 11345 4468
rect 11296 4428 11302 4440
rect 11333 4437 11345 4440
rect 11379 4437 11391 4471
rect 11333 4431 11391 4437
rect 12437 4471 12495 4477
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 12526 4468 12532 4480
rect 12483 4440 12532 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 13265 4471 13323 4477
rect 13265 4468 13277 4471
rect 13136 4440 13277 4468
rect 13136 4428 13142 4440
rect 13265 4437 13277 4440
rect 13311 4437 13323 4471
rect 13265 4431 13323 4437
rect 17954 4428 17960 4480
rect 18012 4428 18018 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 18095 4440 19073 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 19061 4437 19073 4440
rect 19107 4468 19119 4471
rect 19242 4468 19248 4480
rect 19107 4440 19248 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 19886 4428 19892 4480
rect 19944 4428 19950 4480
rect 20622 4428 20628 4480
rect 20680 4428 20686 4480
rect 22005 4471 22063 4477
rect 22005 4437 22017 4471
rect 22051 4468 22063 4471
rect 22186 4468 22192 4480
rect 22051 4440 22192 4468
rect 22051 4437 22063 4440
rect 22005 4431 22063 4437
rect 22186 4428 22192 4440
rect 22244 4428 22250 4480
rect 26786 4428 26792 4480
rect 26844 4428 26850 4480
rect 27522 4428 27528 4480
rect 27580 4428 27586 4480
rect 28721 4471 28779 4477
rect 28721 4437 28733 4471
rect 28767 4468 28779 4471
rect 28994 4468 29000 4480
rect 28767 4440 29000 4468
rect 28767 4437 28779 4440
rect 28721 4431 28779 4437
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 29564 4468 29592 4567
rect 29638 4564 29644 4616
rect 29696 4604 29702 4616
rect 29840 4604 29868 4644
rect 30586 4641 30598 4644
rect 30632 4641 30644 4675
rect 30586 4635 30644 4641
rect 30745 4675 30803 4681
rect 30745 4641 30757 4675
rect 30791 4672 30803 4675
rect 31570 4672 31576 4684
rect 30791 4644 31576 4672
rect 30791 4641 30803 4644
rect 30745 4635 30803 4641
rect 31570 4632 31576 4644
rect 31628 4632 31634 4684
rect 31726 4672 31754 4780
rect 33318 4768 33324 4820
rect 33376 4808 33382 4820
rect 33689 4811 33747 4817
rect 33689 4808 33701 4811
rect 33376 4780 33701 4808
rect 33376 4768 33382 4780
rect 33689 4777 33701 4780
rect 33735 4777 33747 4811
rect 33689 4771 33747 4777
rect 34422 4768 34428 4820
rect 34480 4768 34486 4820
rect 35710 4768 35716 4820
rect 35768 4768 35774 4820
rect 37829 4811 37887 4817
rect 37829 4777 37841 4811
rect 37875 4808 37887 4811
rect 38286 4808 38292 4820
rect 37875 4780 38292 4808
rect 37875 4777 37887 4780
rect 37829 4771 37887 4777
rect 38286 4768 38292 4780
rect 38344 4768 38350 4820
rect 38746 4808 38752 4820
rect 38396 4780 38752 4808
rect 32398 4700 32404 4752
rect 32456 4740 32462 4752
rect 32493 4743 32551 4749
rect 32493 4740 32505 4743
rect 32456 4712 32505 4740
rect 32456 4700 32462 4712
rect 32493 4709 32505 4712
rect 32539 4709 32551 4743
rect 32493 4703 32551 4709
rect 33042 4700 33048 4752
rect 33100 4740 33106 4752
rect 33597 4743 33655 4749
rect 33597 4740 33609 4743
rect 33100 4712 33609 4740
rect 33100 4700 33106 4712
rect 33597 4709 33609 4712
rect 33643 4740 33655 4743
rect 35728 4740 35756 4768
rect 38396 4740 38424 4780
rect 38746 4768 38752 4780
rect 38804 4768 38810 4820
rect 38838 4768 38844 4820
rect 38896 4808 38902 4820
rect 41785 4811 41843 4817
rect 38896 4780 41414 4808
rect 38896 4768 38902 4780
rect 33643 4712 35756 4740
rect 38028 4712 38424 4740
rect 38657 4743 38715 4749
rect 33643 4709 33655 4712
rect 33597 4703 33655 4709
rect 32033 4675 32091 4681
rect 32033 4672 32045 4675
rect 31726 4644 32045 4672
rect 32033 4641 32045 4644
rect 32079 4641 32091 4675
rect 32033 4635 32091 4641
rect 36906 4632 36912 4684
rect 36964 4672 36970 4684
rect 37185 4675 37243 4681
rect 37185 4672 37197 4675
rect 36964 4644 37197 4672
rect 36964 4632 36970 4644
rect 37185 4641 37197 4644
rect 37231 4641 37243 4675
rect 37185 4635 37243 4641
rect 29696 4576 29868 4604
rect 29696 4564 29702 4576
rect 30466 4564 30472 4616
rect 30524 4564 30530 4616
rect 31938 4564 31944 4616
rect 31996 4564 32002 4616
rect 33870 4564 33876 4616
rect 33928 4564 33934 4616
rect 34241 4607 34299 4613
rect 34241 4573 34253 4607
rect 34287 4573 34299 4607
rect 34241 4567 34299 4573
rect 31389 4539 31447 4545
rect 31389 4505 31401 4539
rect 31435 4536 31447 4539
rect 31849 4539 31907 4545
rect 31849 4536 31861 4539
rect 31435 4508 31861 4536
rect 31435 4505 31447 4508
rect 31389 4499 31447 4505
rect 31849 4505 31861 4508
rect 31895 4505 31907 4539
rect 34256 4536 34284 4567
rect 35526 4564 35532 4616
rect 35584 4564 35590 4616
rect 36262 4564 36268 4616
rect 36320 4564 36326 4616
rect 37461 4607 37519 4613
rect 37461 4573 37473 4607
rect 37507 4604 37519 4607
rect 38028 4604 38056 4712
rect 38657 4709 38669 4743
rect 38703 4740 38715 4743
rect 40126 4740 40132 4752
rect 38703 4712 40132 4740
rect 38703 4709 38715 4712
rect 38657 4703 38715 4709
rect 40126 4700 40132 4712
rect 40184 4700 40190 4752
rect 41386 4740 41414 4780
rect 41785 4777 41797 4811
rect 41831 4808 41843 4811
rect 42426 4808 42432 4820
rect 41831 4780 42432 4808
rect 41831 4777 41843 4780
rect 41785 4771 41843 4777
rect 42426 4768 42432 4780
rect 42484 4768 42490 4820
rect 48317 4811 48375 4817
rect 42536 4780 46060 4808
rect 42536 4740 42564 4780
rect 41386 4712 42564 4740
rect 43070 4700 43076 4752
rect 43128 4740 43134 4752
rect 44821 4743 44879 4749
rect 43128 4712 43300 4740
rect 43128 4700 43134 4712
rect 38105 4675 38163 4681
rect 38105 4641 38117 4675
rect 38151 4672 38163 4675
rect 40034 4672 40040 4684
rect 38151 4644 40040 4672
rect 38151 4641 38163 4644
rect 38105 4635 38163 4641
rect 40034 4632 40040 4644
rect 40092 4632 40098 4684
rect 42613 4675 42671 4681
rect 42613 4641 42625 4675
rect 42659 4672 42671 4675
rect 43162 4672 43168 4684
rect 42659 4644 43168 4672
rect 42659 4641 42671 4644
rect 42613 4635 42671 4641
rect 43162 4632 43168 4644
rect 43220 4632 43226 4684
rect 43272 4681 43300 4712
rect 44821 4709 44833 4743
rect 44867 4740 44879 4743
rect 45830 4740 45836 4752
rect 44867 4712 45836 4740
rect 44867 4709 44879 4712
rect 44821 4703 44879 4709
rect 43714 4681 43720 4684
rect 43257 4675 43315 4681
rect 43257 4641 43269 4675
rect 43303 4641 43315 4675
rect 43257 4635 43315 4641
rect 43671 4675 43720 4681
rect 43671 4641 43683 4675
rect 43717 4641 43720 4675
rect 43671 4635 43720 4641
rect 43714 4632 43720 4635
rect 43772 4632 43778 4684
rect 43809 4675 43867 4681
rect 43809 4641 43821 4675
rect 43855 4672 43867 4675
rect 44836 4672 44864 4703
rect 45830 4700 45836 4712
rect 45888 4700 45894 4752
rect 46032 4684 46060 4780
rect 48317 4777 48329 4811
rect 48363 4808 48375 4811
rect 49602 4808 49608 4820
rect 48363 4780 49608 4808
rect 48363 4777 48375 4780
rect 48317 4771 48375 4777
rect 49602 4768 49608 4780
rect 49660 4768 49666 4820
rect 51258 4808 51264 4820
rect 50172 4780 51264 4808
rect 47949 4743 48007 4749
rect 47949 4709 47961 4743
rect 47995 4740 48007 4743
rect 47995 4712 48452 4740
rect 47995 4709 48007 4712
rect 47949 4703 48007 4709
rect 43855 4644 44864 4672
rect 43855 4641 43867 4644
rect 43809 4635 43867 4641
rect 45370 4632 45376 4684
rect 45428 4672 45434 4684
rect 45557 4675 45615 4681
rect 45557 4672 45569 4675
rect 45428 4644 45569 4672
rect 45428 4632 45434 4644
rect 45557 4641 45569 4644
rect 45603 4641 45615 4675
rect 45557 4635 45615 4641
rect 46014 4632 46020 4684
rect 46072 4672 46078 4684
rect 48424 4681 48452 4712
rect 48866 4700 48872 4752
rect 48924 4740 48930 4752
rect 49053 4743 49111 4749
rect 49053 4740 49065 4743
rect 48924 4712 49065 4740
rect 48924 4700 48930 4712
rect 49053 4709 49065 4712
rect 49099 4709 49111 4743
rect 49053 4703 49111 4709
rect 50172 4681 50200 4780
rect 51258 4768 51264 4780
rect 51316 4768 51322 4820
rect 51537 4811 51595 4817
rect 51537 4777 51549 4811
rect 51583 4808 51595 4811
rect 52362 4808 52368 4820
rect 51583 4780 52368 4808
rect 51583 4777 51595 4780
rect 51537 4771 51595 4777
rect 52362 4768 52368 4780
rect 52420 4768 52426 4820
rect 53282 4768 53288 4820
rect 53340 4768 53346 4820
rect 55861 4811 55919 4817
rect 55861 4808 55873 4811
rect 53392 4780 55873 4808
rect 52270 4740 52276 4752
rect 51184 4712 52276 4740
rect 47121 4675 47179 4681
rect 47121 4672 47133 4675
rect 46072 4644 47133 4672
rect 46072 4632 46078 4644
rect 47121 4641 47133 4644
rect 47167 4672 47179 4675
rect 47397 4675 47455 4681
rect 47397 4672 47409 4675
rect 47167 4644 47409 4672
rect 47167 4641 47179 4644
rect 47121 4635 47179 4641
rect 47397 4641 47409 4644
rect 47443 4672 47455 4675
rect 48409 4675 48467 4681
rect 47443 4644 47716 4672
rect 47443 4641 47455 4644
rect 47397 4635 47455 4641
rect 37507 4576 38056 4604
rect 38197 4607 38255 4613
rect 37507 4573 37519 4576
rect 37461 4567 37519 4573
rect 38197 4573 38209 4607
rect 38243 4573 38255 4607
rect 38197 4567 38255 4573
rect 36170 4536 36176 4548
rect 34256 4508 36176 4536
rect 31849 4499 31907 4505
rect 36170 4496 36176 4508
rect 36228 4496 36234 4548
rect 38010 4496 38016 4548
rect 38068 4536 38074 4548
rect 38212 4536 38240 4567
rect 38654 4564 38660 4616
rect 38712 4604 38718 4616
rect 39301 4607 39359 4613
rect 39301 4604 39313 4607
rect 38712 4576 39313 4604
rect 38712 4564 38718 4576
rect 39301 4573 39313 4576
rect 39347 4573 39359 4607
rect 39301 4567 39359 4573
rect 40405 4607 40463 4613
rect 40405 4573 40417 4607
rect 40451 4604 40463 4607
rect 40954 4604 40960 4616
rect 40451 4576 40960 4604
rect 40451 4573 40463 4576
rect 40405 4567 40463 4573
rect 40954 4564 40960 4576
rect 41012 4564 41018 4616
rect 42426 4564 42432 4616
rect 42484 4564 42490 4616
rect 42794 4564 42800 4616
rect 42852 4564 42858 4616
rect 43530 4564 43536 4616
rect 43588 4564 43594 4616
rect 45462 4564 45468 4616
rect 45520 4604 45526 4616
rect 45833 4607 45891 4613
rect 45833 4604 45845 4607
rect 45520 4576 45845 4604
rect 45520 4564 45526 4576
rect 45833 4573 45845 4576
rect 45879 4573 45891 4607
rect 45833 4567 45891 4573
rect 46382 4564 46388 4616
rect 46440 4564 46446 4616
rect 46750 4564 46756 4616
rect 46808 4604 46814 4616
rect 47581 4607 47639 4613
rect 47581 4604 47593 4607
rect 46808 4576 47593 4604
rect 46808 4564 46814 4576
rect 47581 4573 47593 4576
rect 47627 4573 47639 4607
rect 47581 4567 47639 4573
rect 38068 4508 38240 4536
rect 40672 4539 40730 4545
rect 38068 4496 38074 4508
rect 40672 4505 40684 4539
rect 40718 4536 40730 4539
rect 40862 4536 40868 4548
rect 40718 4508 40868 4536
rect 40718 4505 40730 4508
rect 40672 4499 40730 4505
rect 40862 4496 40868 4508
rect 40920 4496 40926 4548
rect 41690 4496 41696 4548
rect 41748 4536 41754 4548
rect 44453 4539 44511 4545
rect 41748 4508 42840 4536
rect 41748 4496 41754 4508
rect 30190 4468 30196 4480
rect 29564 4440 30196 4468
rect 30190 4428 30196 4440
rect 30248 4428 30254 4480
rect 31478 4428 31484 4480
rect 31536 4428 31542 4480
rect 34974 4428 34980 4480
rect 35032 4428 35038 4480
rect 35710 4428 35716 4480
rect 35768 4428 35774 4480
rect 36630 4428 36636 4480
rect 36688 4428 36694 4480
rect 37369 4471 37427 4477
rect 37369 4437 37381 4471
rect 37415 4468 37427 4471
rect 38102 4468 38108 4480
rect 37415 4440 38108 4468
rect 37415 4437 37427 4440
rect 37369 4431 37427 4437
rect 38102 4428 38108 4440
rect 38160 4468 38166 4480
rect 38289 4471 38347 4477
rect 38289 4468 38301 4471
rect 38160 4440 38301 4468
rect 38160 4428 38166 4440
rect 38289 4437 38301 4440
rect 38335 4437 38347 4471
rect 38289 4431 38347 4437
rect 41874 4428 41880 4480
rect 41932 4428 41938 4480
rect 42812 4468 42840 4508
rect 44453 4505 44465 4539
rect 44499 4536 44511 4539
rect 45373 4539 45431 4545
rect 45373 4536 45385 4539
rect 44499 4508 45385 4536
rect 44499 4505 44511 4508
rect 44453 4499 44511 4505
rect 45373 4505 45385 4508
rect 45419 4505 45431 4539
rect 47688 4536 47716 4644
rect 48409 4641 48421 4675
rect 48455 4641 48467 4675
rect 48409 4635 48467 4641
rect 50157 4675 50215 4681
rect 50157 4641 50169 4675
rect 50203 4641 50215 4675
rect 50157 4635 50215 4641
rect 49050 4564 49056 4616
rect 49108 4604 49114 4616
rect 49697 4607 49755 4613
rect 49697 4604 49709 4607
rect 49108 4576 49709 4604
rect 49108 4564 49114 4576
rect 49697 4573 49709 4576
rect 49743 4573 49755 4607
rect 49697 4567 49755 4573
rect 50424 4607 50482 4613
rect 50424 4573 50436 4607
rect 50470 4604 50482 4607
rect 50706 4604 50712 4616
rect 50470 4576 50712 4604
rect 50470 4573 50482 4576
rect 50424 4567 50482 4573
rect 50706 4564 50712 4576
rect 50764 4564 50770 4616
rect 51184 4536 51212 4712
rect 52270 4700 52276 4712
rect 52328 4700 52334 4752
rect 52914 4700 52920 4752
rect 52972 4740 52978 4752
rect 53392 4740 53420 4780
rect 55861 4777 55873 4780
rect 55907 4777 55919 4811
rect 55861 4771 55919 4777
rect 52972 4712 53420 4740
rect 55125 4743 55183 4749
rect 52972 4700 52978 4712
rect 55125 4709 55137 4743
rect 55171 4709 55183 4743
rect 55125 4703 55183 4709
rect 55030 4632 55036 4684
rect 55088 4672 55094 4684
rect 55140 4672 55168 4703
rect 55398 4700 55404 4752
rect 55456 4740 55462 4752
rect 55456 4712 56272 4740
rect 55456 4700 55462 4712
rect 55088 4644 55168 4672
rect 55088 4632 55094 4644
rect 55214 4632 55220 4684
rect 55272 4672 55278 4684
rect 55490 4672 55496 4684
rect 55272 4644 55496 4672
rect 55272 4632 55278 4644
rect 55490 4632 55496 4644
rect 55548 4672 55554 4684
rect 56244 4681 56272 4712
rect 55585 4675 55643 4681
rect 55585 4672 55597 4675
rect 55548 4644 55597 4672
rect 55548 4632 55554 4644
rect 55585 4641 55597 4644
rect 55631 4641 55643 4675
rect 55585 4635 55643 4641
rect 56229 4675 56287 4681
rect 56229 4641 56241 4675
rect 56275 4641 56287 4675
rect 56229 4635 56287 4641
rect 56318 4632 56324 4684
rect 56376 4672 56382 4684
rect 56413 4675 56471 4681
rect 56413 4672 56425 4675
rect 56376 4644 56425 4672
rect 56376 4632 56382 4644
rect 56413 4641 56425 4644
rect 56459 4641 56471 4675
rect 56413 4635 56471 4641
rect 51534 4564 51540 4616
rect 51592 4604 51598 4616
rect 52181 4607 52239 4613
rect 52181 4604 52193 4607
rect 51592 4576 52193 4604
rect 51592 4564 51598 4576
rect 52181 4573 52193 4576
rect 52227 4573 52239 4607
rect 52181 4567 52239 4573
rect 52270 4564 52276 4616
rect 52328 4604 52334 4616
rect 52917 4607 52975 4613
rect 52917 4604 52929 4607
rect 52328 4576 52929 4604
rect 52328 4564 52334 4576
rect 52917 4573 52929 4576
rect 52963 4573 52975 4607
rect 52917 4567 52975 4573
rect 53101 4607 53159 4613
rect 53101 4573 53113 4607
rect 53147 4604 53159 4607
rect 53650 4604 53656 4616
rect 53147 4576 53656 4604
rect 53147 4573 53159 4576
rect 53101 4567 53159 4573
rect 53650 4564 53656 4576
rect 53708 4564 53714 4616
rect 53745 4607 53803 4613
rect 53745 4573 53757 4607
rect 53791 4604 53803 4607
rect 54012 4607 54070 4613
rect 53791 4576 53972 4604
rect 53791 4573 53803 4576
rect 53745 4567 53803 4573
rect 47688 4508 51212 4536
rect 45373 4499 45431 4505
rect 53944 4480 53972 4576
rect 54012 4573 54024 4607
rect 54058 4604 54070 4607
rect 55122 4604 55128 4616
rect 54058 4576 55128 4604
rect 54058 4573 54070 4576
rect 54012 4567 54070 4573
rect 55122 4564 55128 4576
rect 55180 4564 55186 4616
rect 58250 4564 58256 4616
rect 58308 4564 58314 4616
rect 54938 4496 54944 4548
rect 54996 4536 55002 4548
rect 55401 4539 55459 4545
rect 55401 4536 55413 4539
rect 54996 4508 55413 4536
rect 54996 4496 55002 4508
rect 55401 4505 55413 4508
rect 55447 4505 55459 4539
rect 55401 4499 55459 4505
rect 56134 4496 56140 4548
rect 56192 4536 56198 4548
rect 56505 4539 56563 4545
rect 56505 4536 56517 4539
rect 56192 4508 56517 4536
rect 56192 4496 56198 4508
rect 56505 4505 56517 4508
rect 56551 4505 56563 4539
rect 56505 4499 56563 4505
rect 57146 4496 57152 4548
rect 57204 4496 57210 4548
rect 43530 4468 43536 4480
rect 42812 4440 43536 4468
rect 43530 4428 43536 4440
rect 43588 4428 43594 4480
rect 45002 4428 45008 4480
rect 45060 4428 45066 4480
rect 45186 4428 45192 4480
rect 45244 4468 45250 4480
rect 45465 4471 45523 4477
rect 45465 4468 45477 4471
rect 45244 4440 45477 4468
rect 45244 4428 45250 4440
rect 45465 4437 45477 4440
rect 45511 4437 45523 4471
rect 45465 4431 45523 4437
rect 47489 4471 47547 4477
rect 47489 4437 47501 4471
rect 47535 4468 47547 4471
rect 47946 4468 47952 4480
rect 47535 4440 47952 4468
rect 47535 4437 47547 4440
rect 47489 4431 47547 4437
rect 47946 4428 47952 4440
rect 48004 4428 48010 4480
rect 49142 4428 49148 4480
rect 49200 4428 49206 4480
rect 50430 4428 50436 4480
rect 50488 4468 50494 4480
rect 51629 4471 51687 4477
rect 51629 4468 51641 4471
rect 50488 4440 51641 4468
rect 50488 4428 50494 4440
rect 51629 4437 51641 4440
rect 51675 4437 51687 4471
rect 51629 4431 51687 4437
rect 52362 4428 52368 4480
rect 52420 4428 52426 4480
rect 53466 4428 53472 4480
rect 53524 4468 53530 4480
rect 53561 4471 53619 4477
rect 53561 4468 53573 4471
rect 53524 4440 53573 4468
rect 53524 4428 53530 4440
rect 53561 4437 53573 4440
rect 53607 4437 53619 4471
rect 53561 4431 53619 4437
rect 53926 4428 53932 4480
rect 53984 4428 53990 4480
rect 56873 4471 56931 4477
rect 56873 4437 56885 4471
rect 56919 4468 56931 4471
rect 58066 4468 58072 4480
rect 56919 4440 58072 4468
rect 56919 4437 56931 4440
rect 56873 4431 56931 4437
rect 58066 4428 58072 4440
rect 58124 4428 58130 4480
rect 1104 4378 59040 4400
rect 1104 4326 15394 4378
rect 15446 4326 15458 4378
rect 15510 4326 15522 4378
rect 15574 4326 15586 4378
rect 15638 4326 15650 4378
rect 15702 4326 29838 4378
rect 29890 4326 29902 4378
rect 29954 4326 29966 4378
rect 30018 4326 30030 4378
rect 30082 4326 30094 4378
rect 30146 4326 44282 4378
rect 44334 4326 44346 4378
rect 44398 4326 44410 4378
rect 44462 4326 44474 4378
rect 44526 4326 44538 4378
rect 44590 4326 58726 4378
rect 58778 4326 58790 4378
rect 58842 4326 58854 4378
rect 58906 4326 58918 4378
rect 58970 4326 58982 4378
rect 59034 4326 59040 4378
rect 1104 4304 59040 4326
rect 2958 4224 2964 4276
rect 3016 4224 3022 4276
rect 3329 4267 3387 4273
rect 3329 4233 3341 4267
rect 3375 4264 3387 4267
rect 4246 4264 4252 4276
rect 3375 4236 4252 4264
rect 3375 4233 3387 4236
rect 3329 4227 3387 4233
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4396 4236 7420 4264
rect 4396 4224 4402 4236
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 6549 4199 6607 4205
rect 6549 4196 6561 4199
rect 2832 4168 6561 4196
rect 2832 4156 2838 4168
rect 6549 4165 6561 4168
rect 6595 4165 6607 4199
rect 6549 4159 6607 4165
rect 6638 4156 6644 4208
rect 6696 4196 6702 4208
rect 6825 4199 6883 4205
rect 6825 4196 6837 4199
rect 6696 4168 6837 4196
rect 6696 4156 6702 4168
rect 6825 4165 6837 4168
rect 6871 4196 6883 4199
rect 6914 4196 6920 4208
rect 6871 4168 6920 4196
rect 6871 4165 6883 4168
rect 6825 4159 6883 4165
rect 6914 4156 6920 4168
rect 6972 4156 6978 4208
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 4706 4128 4712 4140
rect 3467 4100 4712 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2133 4023 2191 4029
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 3605 4063 3663 4069
rect 2363 4032 3464 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2148 3992 2176 4023
rect 3234 3992 3240 4004
rect 2148 3964 3240 3992
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 3436 3992 3464 4032
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 4062 4060 4068 4072
rect 3651 4032 4068 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 4982 4060 4988 4072
rect 4203 4032 4988 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 5442 4020 5448 4072
rect 5500 4020 5506 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6086 4060 6092 4072
rect 5675 4032 6092 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6472 4060 6500 4088
rect 6227 4032 6500 4060
rect 6932 4060 6960 4156
rect 7392 4137 7420 4236
rect 8018 4224 8024 4276
rect 8076 4224 8082 4276
rect 8846 4224 8852 4276
rect 8904 4224 8910 4276
rect 9214 4224 9220 4276
rect 9272 4224 9278 4276
rect 9306 4224 9312 4276
rect 9364 4224 9370 4276
rect 9769 4267 9827 4273
rect 9769 4233 9781 4267
rect 9815 4233 9827 4267
rect 9769 4227 9827 4233
rect 8665 4199 8723 4205
rect 8665 4165 8677 4199
rect 8711 4196 8723 4199
rect 9784 4196 9812 4227
rect 10226 4224 10232 4276
rect 10284 4224 10290 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10468 4236 10701 4264
rect 10468 4224 10474 4236
rect 10689 4233 10701 4236
rect 10735 4233 10747 4267
rect 10689 4227 10747 4233
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 13446 4264 13452 4276
rect 12584 4236 13452 4264
rect 12584 4224 12590 4236
rect 13446 4224 13452 4236
rect 13504 4264 13510 4276
rect 13909 4267 13967 4273
rect 13909 4264 13921 4267
rect 13504 4236 13921 4264
rect 13504 4224 13510 4236
rect 13909 4233 13921 4236
rect 13955 4233 13967 4267
rect 13909 4227 13967 4233
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 15933 4267 15991 4273
rect 15933 4264 15945 4267
rect 15804 4236 15945 4264
rect 15804 4224 15810 4236
rect 15933 4233 15945 4236
rect 15979 4233 15991 4267
rect 15933 4227 15991 4233
rect 16114 4224 16120 4276
rect 16172 4224 16178 4276
rect 18233 4267 18291 4273
rect 18233 4233 18245 4267
rect 18279 4264 18291 4267
rect 18414 4264 18420 4276
rect 18279 4236 18420 4264
rect 18279 4233 18291 4236
rect 18233 4227 18291 4233
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 20162 4224 20168 4276
rect 20220 4224 20226 4276
rect 20257 4267 20315 4273
rect 20257 4233 20269 4267
rect 20303 4264 20315 4267
rect 20438 4264 20444 4276
rect 20303 4236 20444 4264
rect 20303 4233 20315 4236
rect 20257 4227 20315 4233
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 20622 4224 20628 4276
rect 20680 4264 20686 4276
rect 20717 4267 20775 4273
rect 20717 4264 20729 4267
rect 20680 4236 20729 4264
rect 20680 4224 20686 4236
rect 20717 4233 20729 4236
rect 20763 4233 20775 4267
rect 20717 4227 20775 4233
rect 20898 4224 20904 4276
rect 20956 4224 20962 4276
rect 21542 4224 21548 4276
rect 21600 4264 21606 4276
rect 24029 4267 24087 4273
rect 21600 4236 22094 4264
rect 21600 4224 21606 4236
rect 10597 4199 10655 4205
rect 10597 4196 10609 4199
rect 8711 4168 9812 4196
rect 9876 4168 10609 4196
rect 8711 4165 8723 4168
rect 8665 4159 8723 4165
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7834 4128 7840 4140
rect 7423 4100 7840 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 9214 4128 9220 4140
rect 8527 4100 9220 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 9214 4088 9220 4100
rect 9272 4128 9278 4140
rect 9876 4128 9904 4168
rect 10597 4165 10609 4168
rect 10643 4165 10655 4199
rect 16132 4196 16160 4224
rect 20916 4196 20944 4224
rect 16132 4168 18552 4196
rect 10597 4159 10655 4165
rect 9272 4100 9904 4128
rect 9272 4088 9278 4100
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 12084 4100 13461 4128
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 6932 4032 8309 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 3878 3992 3884 4004
rect 3436 3964 3884 3992
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 4522 3952 4528 4004
rect 4580 3952 4586 4004
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 6638 3992 6644 4004
rect 4755 3964 6644 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 8312 3992 8340 4023
rect 9490 4020 9496 4072
rect 9548 4020 9554 4072
rect 10870 4020 10876 4072
rect 10928 4020 10934 4072
rect 12084 4069 12112 4100
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 15988 4100 16160 4128
rect 15988 4088 15994 4100
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 10594 3992 10600 4004
rect 7944 3964 8248 3992
rect 8312 3964 10600 3992
rect 1489 3927 1547 3933
rect 1489 3893 1501 3927
rect 1535 3924 1547 3927
rect 1854 3924 1860 3936
rect 1535 3896 1860 3924
rect 1535 3893 1547 3896
rect 1489 3887 1547 3893
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 4540 3924 4568 3952
rect 7944 3924 7972 3964
rect 4540 3896 7972 3924
rect 8220 3924 8248 3964
rect 10594 3952 10600 3964
rect 10652 3992 10658 4004
rect 10962 3992 10968 4004
rect 10652 3964 10968 3992
rect 10652 3952 10658 3964
rect 10962 3952 10968 3964
rect 11020 3992 11026 4004
rect 11241 3995 11299 4001
rect 11241 3992 11253 3995
rect 11020 3964 11253 3992
rect 11020 3952 11026 3964
rect 11241 3961 11253 3964
rect 11287 3961 11299 3995
rect 11241 3955 11299 3961
rect 12084 3936 12112 4023
rect 12158 4020 12164 4072
rect 12216 4060 12222 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12216 4032 12449 4060
rect 12216 4020 12222 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 14200 3992 14228 4023
rect 14918 4020 14924 4072
rect 14976 4020 14982 4072
rect 16132 4069 16160 4100
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16264 4100 16865 4128
rect 16264 4088 16270 4100
rect 16853 4097 16865 4100
rect 16899 4128 16911 4131
rect 16942 4128 16948 4140
rect 16899 4100 16948 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17126 4137 17132 4140
rect 17120 4128 17132 4137
rect 17087 4100 17132 4128
rect 17120 4091 17132 4100
rect 17126 4088 17132 4091
rect 17184 4088 17190 4140
rect 18524 4128 18552 4168
rect 20640 4168 20944 4196
rect 18524 4100 18644 4128
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4060 15531 4063
rect 16025 4063 16083 4069
rect 16025 4060 16037 4063
rect 15519 4032 16037 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 16025 4029 16037 4032
rect 16071 4029 16083 4063
rect 16025 4023 16083 4029
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 15565 3995 15623 4001
rect 15565 3992 15577 3995
rect 14200 3964 15577 3992
rect 15565 3961 15577 3964
rect 15611 3961 15623 3995
rect 15565 3955 15623 3961
rect 10686 3924 10692 3936
rect 8220 3896 10692 3924
rect 10686 3884 10692 3896
rect 10744 3924 10750 3936
rect 10870 3924 10876 3936
rect 10744 3896 10876 3924
rect 10744 3884 10750 3896
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3924 11575 3927
rect 11882 3924 11888 3936
rect 11563 3896 11888 3924
rect 11563 3893 11575 3896
rect 11517 3887 11575 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12066 3884 12072 3936
rect 12124 3884 12130 3936
rect 14734 3884 14740 3936
rect 14792 3884 14798 3936
rect 16132 3924 16160 4023
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 17920 4032 18337 4060
rect 17920 4020 17926 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4029 18567 4063
rect 18616 4060 18644 4100
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 19518 4088 19524 4140
rect 19576 4088 19582 4140
rect 20640 4137 20668 4168
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4097 20683 4131
rect 22066 4128 22094 4236
rect 24029 4233 24041 4267
rect 24075 4264 24087 4267
rect 24302 4264 24308 4276
rect 24075 4236 24308 4264
rect 24075 4233 24087 4236
rect 24029 4227 24087 4233
rect 24302 4224 24308 4236
rect 24360 4264 24366 4276
rect 25777 4267 25835 4273
rect 25777 4264 25789 4267
rect 24360 4236 25789 4264
rect 24360 4224 24366 4236
rect 25777 4233 25789 4236
rect 25823 4233 25835 4267
rect 25777 4227 25835 4233
rect 27249 4267 27307 4273
rect 27249 4233 27261 4267
rect 27295 4264 27307 4267
rect 27522 4264 27528 4276
rect 27295 4236 27528 4264
rect 27295 4233 27307 4236
rect 27249 4227 27307 4233
rect 27522 4224 27528 4236
rect 27580 4224 27586 4276
rect 27614 4224 27620 4276
rect 27672 4224 27678 4276
rect 27706 4224 27712 4276
rect 27764 4224 27770 4276
rect 28442 4224 28448 4276
rect 28500 4224 28506 4276
rect 29362 4224 29368 4276
rect 29420 4264 29426 4276
rect 29733 4267 29791 4273
rect 29733 4264 29745 4267
rect 29420 4236 29745 4264
rect 29420 4224 29426 4236
rect 29733 4233 29745 4236
rect 29779 4233 29791 4267
rect 29733 4227 29791 4233
rect 30282 4224 30288 4276
rect 30340 4224 30346 4276
rect 30466 4224 30472 4276
rect 30524 4264 30530 4276
rect 31018 4264 31024 4276
rect 30524 4236 31024 4264
rect 30524 4224 30530 4236
rect 31018 4224 31024 4236
rect 31076 4224 31082 4276
rect 35069 4267 35127 4273
rect 35069 4233 35081 4267
rect 35115 4264 35127 4267
rect 35526 4264 35532 4276
rect 35115 4236 35532 4264
rect 35115 4233 35127 4236
rect 35069 4227 35127 4233
rect 35526 4224 35532 4236
rect 35584 4224 35590 4276
rect 35618 4224 35624 4276
rect 35676 4224 35682 4276
rect 35802 4224 35808 4276
rect 35860 4224 35866 4276
rect 35897 4267 35955 4273
rect 35897 4233 35909 4267
rect 35943 4264 35955 4267
rect 36262 4264 36268 4276
rect 35943 4236 36268 4264
rect 35943 4233 35955 4236
rect 35897 4227 35955 4233
rect 36262 4224 36268 4236
rect 36320 4224 36326 4276
rect 38194 4264 38200 4276
rect 37292 4236 38200 4264
rect 25869 4199 25927 4205
rect 23952 4168 24164 4196
rect 23952 4128 23980 4168
rect 22066 4100 23980 4128
rect 24136 4128 24164 4168
rect 25869 4165 25881 4199
rect 25915 4196 25927 4199
rect 27341 4199 27399 4205
rect 25915 4168 26924 4196
rect 25915 4165 25927 4168
rect 25869 4159 25927 4165
rect 26896 4128 26924 4168
rect 27341 4165 27353 4199
rect 27387 4196 27399 4199
rect 27632 4196 27660 4224
rect 27387 4168 27660 4196
rect 27387 4165 27399 4168
rect 27341 4159 27399 4165
rect 28077 4131 28135 4137
rect 24136 4100 24256 4128
rect 26896 4100 27936 4128
rect 20625 4091 20683 4097
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18616 4032 18981 4060
rect 18509 4023 18567 4029
rect 18969 4029 18981 4032
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 16390 3924 16396 3936
rect 16132 3896 16396 3924
rect 16390 3884 16396 3896
rect 16448 3924 16454 3936
rect 17494 3924 17500 3936
rect 16448 3896 17500 3924
rect 16448 3884 16454 3896
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 18524 3924 18552 4023
rect 19058 4020 19064 4072
rect 19116 4060 19122 4072
rect 19362 4063 19420 4069
rect 19362 4060 19374 4063
rect 19116 4032 19374 4060
rect 19116 4020 19122 4032
rect 19362 4029 19374 4032
rect 19408 4029 19420 4063
rect 19362 4023 19420 4029
rect 20809 4063 20867 4069
rect 20809 4029 20821 4063
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 23017 4063 23075 4069
rect 23017 4029 23029 4063
rect 23063 4060 23075 4063
rect 23474 4060 23480 4072
rect 23063 4032 23480 4060
rect 23063 4029 23075 4032
rect 23017 4023 23075 4029
rect 20824 3936 20852 4023
rect 22296 3992 22324 4023
rect 23474 4020 23480 4032
rect 23532 4020 23538 4072
rect 24228 4069 24256 4100
rect 23569 4063 23627 4069
rect 23569 4029 23581 4063
rect 23615 4060 23627 4063
rect 24121 4063 24179 4069
rect 24121 4060 24133 4063
rect 23615 4032 24133 4060
rect 23615 4029 23627 4032
rect 23569 4023 23627 4029
rect 24121 4029 24133 4032
rect 24167 4029 24179 4063
rect 24121 4023 24179 4029
rect 24213 4063 24271 4069
rect 24213 4029 24225 4063
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 25222 4020 25228 4072
rect 25280 4020 25286 4072
rect 26602 4020 26608 4072
rect 26660 4020 26666 4072
rect 26694 4020 26700 4072
rect 26752 4060 26758 4072
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 26752 4032 27169 4060
rect 26752 4020 26758 4032
rect 27157 4029 27169 4032
rect 27203 4060 27215 4063
rect 27430 4060 27436 4072
rect 27203 4032 27436 4060
rect 27203 4029 27215 4032
rect 27157 4023 27215 4029
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 27908 4001 27936 4100
rect 28077 4097 28089 4131
rect 28123 4097 28135 4131
rect 28077 4091 28135 4097
rect 28261 4131 28319 4137
rect 28261 4097 28273 4131
rect 28307 4128 28319 4131
rect 28460 4128 28488 4224
rect 29454 4156 29460 4208
rect 29512 4156 29518 4208
rect 30101 4199 30159 4205
rect 30101 4165 30113 4199
rect 30147 4196 30159 4199
rect 30300 4196 30328 4224
rect 30929 4199 30987 4205
rect 30929 4196 30941 4199
rect 30147 4168 30941 4196
rect 30147 4165 30159 4168
rect 30101 4159 30159 4165
rect 30929 4165 30941 4168
rect 30975 4165 30987 4199
rect 30929 4159 30987 4165
rect 35437 4199 35495 4205
rect 35437 4165 35449 4199
rect 35483 4196 35495 4199
rect 35636 4196 35664 4224
rect 35483 4168 35664 4196
rect 35483 4165 35495 4168
rect 35437 4159 35495 4165
rect 28307 4100 28488 4128
rect 28528 4131 28586 4137
rect 28307 4097 28319 4100
rect 28261 4091 28319 4097
rect 28528 4097 28540 4131
rect 28574 4128 28586 4131
rect 29472 4128 29500 4156
rect 28574 4100 29500 4128
rect 28574 4097 28586 4100
rect 28528 4091 28586 4097
rect 23661 3995 23719 4001
rect 23661 3992 23673 3995
rect 22296 3964 23673 3992
rect 23661 3961 23673 3964
rect 23707 3961 23719 3995
rect 23661 3955 23719 3961
rect 27893 3995 27951 4001
rect 27893 3961 27905 3995
rect 27939 3961 27951 3995
rect 27893 3955 27951 3961
rect 19334 3924 19340 3936
rect 18524 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 20806 3884 20812 3936
rect 20864 3884 20870 3936
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 22462 3924 22468 3936
rect 22152 3896 22468 3924
rect 22152 3884 22158 3896
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 22833 3927 22891 3933
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 23014 3924 23020 3936
rect 22879 3896 23020 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 24581 3927 24639 3933
rect 24581 3893 24593 3927
rect 24627 3924 24639 3927
rect 24854 3924 24860 3936
rect 24627 3896 24860 3924
rect 24627 3893 24639 3896
rect 24581 3887 24639 3893
rect 24854 3884 24860 3896
rect 24912 3884 24918 3936
rect 25498 3884 25504 3936
rect 25556 3884 25562 3936
rect 26050 3884 26056 3936
rect 26108 3884 26114 3936
rect 27154 3884 27160 3936
rect 27212 3924 27218 3936
rect 28092 3924 28120 4091
rect 30190 4088 30196 4140
rect 30248 4128 30254 4140
rect 30248 4100 30696 4128
rect 30248 4088 30254 4100
rect 30285 4063 30343 4069
rect 30285 4029 30297 4063
rect 30331 4029 30343 4063
rect 30285 4023 30343 4029
rect 29641 3995 29699 4001
rect 29641 3961 29653 3995
rect 29687 3992 29699 3995
rect 30190 3992 30196 4004
rect 29687 3964 30196 3992
rect 29687 3961 29699 3964
rect 29641 3955 29699 3961
rect 30190 3952 30196 3964
rect 30248 3952 30254 4004
rect 27212 3896 28120 3924
rect 30300 3924 30328 4023
rect 30558 3952 30564 4004
rect 30616 3952 30622 4004
rect 30668 3992 30696 4100
rect 31662 4088 31668 4140
rect 31720 4088 31726 4140
rect 35529 4131 35587 4137
rect 35529 4097 35541 4131
rect 35575 4128 35587 4131
rect 35820 4128 35848 4224
rect 37292 4196 37320 4236
rect 38194 4224 38200 4236
rect 38252 4224 38258 4276
rect 38654 4224 38660 4276
rect 38712 4224 38718 4276
rect 39025 4267 39083 4273
rect 39025 4233 39037 4267
rect 39071 4264 39083 4267
rect 39298 4264 39304 4276
rect 39071 4236 39304 4264
rect 39071 4233 39083 4236
rect 39025 4227 39083 4233
rect 39298 4224 39304 4236
rect 39356 4224 39362 4276
rect 39482 4224 39488 4276
rect 39540 4224 39546 4276
rect 39574 4224 39580 4276
rect 39632 4224 39638 4276
rect 41417 4267 41475 4273
rect 41417 4233 41429 4267
rect 41463 4264 41475 4267
rect 41690 4264 41696 4276
rect 41463 4236 41696 4264
rect 41463 4233 41475 4236
rect 41417 4227 41475 4233
rect 41690 4224 41696 4236
rect 41748 4224 41754 4276
rect 41877 4267 41935 4273
rect 41877 4233 41889 4267
rect 41923 4264 41935 4267
rect 42426 4264 42432 4276
rect 41923 4236 42432 4264
rect 41923 4233 41935 4236
rect 41877 4227 41935 4233
rect 42426 4224 42432 4236
rect 42484 4224 42490 4276
rect 42797 4267 42855 4273
rect 42797 4233 42809 4267
rect 42843 4264 42855 4267
rect 43162 4264 43168 4276
rect 42843 4236 43168 4264
rect 42843 4233 42855 4236
rect 42797 4227 42855 4233
rect 43162 4224 43168 4236
rect 43220 4224 43226 4276
rect 43257 4267 43315 4273
rect 43257 4233 43269 4267
rect 43303 4233 43315 4267
rect 43257 4227 43315 4233
rect 36280 4168 37320 4196
rect 37544 4199 37602 4205
rect 36280 4137 36308 4168
rect 37544 4165 37556 4199
rect 37590 4196 37602 4199
rect 37734 4196 37740 4208
rect 37590 4168 37740 4196
rect 37590 4165 37602 4168
rect 37544 4159 37602 4165
rect 37734 4156 37740 4168
rect 37792 4156 37798 4208
rect 39117 4199 39175 4205
rect 39117 4165 39129 4199
rect 39163 4196 39175 4199
rect 39592 4196 39620 4224
rect 39163 4168 39620 4196
rect 39163 4165 39175 4168
rect 39117 4159 39175 4165
rect 40954 4156 40960 4208
rect 41012 4196 41018 4208
rect 43272 4196 43300 4227
rect 44726 4224 44732 4276
rect 44784 4224 44790 4276
rect 45002 4224 45008 4276
rect 45060 4264 45066 4276
rect 45189 4267 45247 4273
rect 45189 4264 45201 4267
rect 45060 4236 45201 4264
rect 45060 4224 45066 4236
rect 45189 4233 45201 4236
rect 45235 4233 45247 4267
rect 45189 4227 45247 4233
rect 45557 4267 45615 4273
rect 45557 4233 45569 4267
rect 45603 4264 45615 4267
rect 46382 4264 46388 4276
rect 45603 4236 46388 4264
rect 45603 4233 45615 4236
rect 45557 4227 45615 4233
rect 46382 4224 46388 4236
rect 46440 4224 46446 4276
rect 48685 4267 48743 4273
rect 48685 4233 48697 4267
rect 48731 4264 48743 4267
rect 48774 4264 48780 4276
rect 48731 4236 48780 4264
rect 48731 4233 48743 4236
rect 48685 4227 48743 4233
rect 48774 4224 48780 4236
rect 48832 4224 48838 4276
rect 49050 4224 49056 4276
rect 49108 4224 49114 4276
rect 49513 4267 49571 4273
rect 49513 4233 49525 4267
rect 49559 4264 49571 4267
rect 49694 4264 49700 4276
rect 49559 4236 49700 4264
rect 49559 4233 49571 4236
rect 49513 4227 49571 4233
rect 49694 4224 49700 4236
rect 49752 4224 49758 4276
rect 50433 4267 50491 4273
rect 50433 4233 50445 4267
rect 50479 4264 50491 4267
rect 50982 4264 50988 4276
rect 50479 4236 50988 4264
rect 50479 4233 50491 4236
rect 50433 4227 50491 4233
rect 50982 4224 50988 4236
rect 51040 4224 51046 4276
rect 52270 4224 52276 4276
rect 52328 4224 52334 4276
rect 52730 4224 52736 4276
rect 52788 4224 52794 4276
rect 53101 4267 53159 4273
rect 53101 4233 53113 4267
rect 53147 4264 53159 4267
rect 55030 4264 55036 4276
rect 53147 4236 55036 4264
rect 53147 4233 53159 4236
rect 53101 4227 53159 4233
rect 55030 4224 55036 4236
rect 55088 4224 55094 4276
rect 55122 4224 55128 4276
rect 55180 4264 55186 4276
rect 55180 4236 56088 4264
rect 55180 4224 55186 4236
rect 51905 4199 51963 4205
rect 41012 4168 43024 4196
rect 43272 4168 43760 4196
rect 41012 4156 41018 4168
rect 35575 4100 35848 4128
rect 36265 4131 36323 4137
rect 35575 4097 35587 4100
rect 35529 4091 35587 4097
rect 36265 4097 36277 4131
rect 36311 4097 36323 4131
rect 36265 4091 36323 4097
rect 36906 4088 36912 4140
rect 36964 4128 36970 4140
rect 37001 4131 37059 4137
rect 37001 4128 37013 4131
rect 36964 4100 37013 4128
rect 36964 4088 36970 4100
rect 37001 4097 37013 4100
rect 37047 4097 37059 4131
rect 39758 4128 39764 4140
rect 37001 4091 37059 4097
rect 37108 4100 39764 4128
rect 31110 4020 31116 4072
rect 31168 4020 31174 4072
rect 31570 4020 31576 4072
rect 31628 4060 31634 4072
rect 32677 4063 32735 4069
rect 32677 4060 32689 4063
rect 31628 4032 32689 4060
rect 31628 4020 31634 4032
rect 32677 4029 32689 4032
rect 32723 4029 32735 4063
rect 32677 4023 32735 4029
rect 33134 4020 33140 4072
rect 33192 4060 33198 4072
rect 33413 4063 33471 4069
rect 33413 4060 33425 4063
rect 33192 4032 33425 4060
rect 33192 4020 33198 4032
rect 33413 4029 33425 4032
rect 33459 4029 33471 4063
rect 33413 4023 33471 4029
rect 34146 4020 34152 4072
rect 34204 4020 34210 4072
rect 34882 4020 34888 4072
rect 34940 4020 34946 4072
rect 35713 4063 35771 4069
rect 35713 4029 35725 4063
rect 35759 4029 35771 4063
rect 35713 4023 35771 4029
rect 32125 3995 32183 4001
rect 32125 3992 32137 3995
rect 30668 3964 32137 3992
rect 32125 3961 32137 3964
rect 32171 3961 32183 3995
rect 35728 3992 35756 4023
rect 36354 4020 36360 4072
rect 36412 4020 36418 4072
rect 36541 4063 36599 4069
rect 36541 4029 36553 4063
rect 36587 4060 36599 4063
rect 36630 4060 36636 4072
rect 36587 4032 36636 4060
rect 36587 4029 36599 4032
rect 36541 4023 36599 4029
rect 36556 3992 36584 4023
rect 36630 4020 36636 4032
rect 36688 4060 36694 4072
rect 37108 4060 37136 4100
rect 38948 4069 38976 4100
rect 39758 4088 39764 4100
rect 39816 4088 39822 4140
rect 40126 4088 40132 4140
rect 40184 4088 40190 4140
rect 41506 4088 41512 4140
rect 41564 4088 41570 4140
rect 41969 4131 42027 4137
rect 41969 4097 41981 4131
rect 42015 4128 42027 4131
rect 42794 4128 42800 4140
rect 42015 4100 42800 4128
rect 42015 4097 42027 4100
rect 41969 4091 42027 4097
rect 42794 4088 42800 4100
rect 42852 4088 42858 4140
rect 42889 4131 42947 4137
rect 42889 4097 42901 4131
rect 42935 4097 42947 4131
rect 42996 4128 43024 4168
rect 43622 4137 43628 4140
rect 43349 4131 43407 4137
rect 43349 4128 43361 4131
rect 42996 4100 43361 4128
rect 42889 4091 42947 4097
rect 43349 4097 43361 4100
rect 43395 4097 43407 4131
rect 43616 4128 43628 4137
rect 43583 4100 43628 4128
rect 43349 4091 43407 4097
rect 43616 4091 43628 4100
rect 36688 4032 37136 4060
rect 37277 4063 37335 4069
rect 36688 4020 36694 4032
rect 37277 4029 37289 4063
rect 37323 4029 37335 4063
rect 37277 4023 37335 4029
rect 38933 4063 38991 4069
rect 38933 4029 38945 4063
rect 38979 4029 38991 4063
rect 38933 4023 38991 4029
rect 35728 3964 36584 3992
rect 32125 3955 32183 3961
rect 30650 3924 30656 3936
rect 30300 3896 30656 3924
rect 27212 3884 27218 3896
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 31202 3884 31208 3936
rect 31260 3924 31266 3936
rect 31481 3927 31539 3933
rect 31481 3924 31493 3927
rect 31260 3896 31493 3924
rect 31260 3884 31266 3896
rect 31481 3893 31493 3896
rect 31527 3893 31539 3927
rect 31481 3887 31539 3893
rect 32858 3884 32864 3936
rect 32916 3884 32922 3936
rect 33226 3884 33232 3936
rect 33284 3924 33290 3936
rect 33597 3927 33655 3933
rect 33597 3924 33609 3927
rect 33284 3896 33609 3924
rect 33284 3884 33290 3896
rect 33597 3893 33609 3896
rect 33643 3893 33655 3927
rect 33597 3887 33655 3893
rect 34330 3884 34336 3936
rect 34388 3884 34394 3936
rect 35894 3884 35900 3936
rect 35952 3924 35958 3936
rect 36817 3927 36875 3933
rect 36817 3924 36829 3927
rect 35952 3896 36829 3924
rect 35952 3884 35958 3896
rect 36817 3893 36829 3896
rect 36863 3893 36875 3927
rect 37292 3924 37320 4023
rect 39022 4020 39028 4072
rect 39080 4060 39086 4072
rect 40865 4063 40923 4069
rect 40865 4060 40877 4063
rect 39080 4032 40877 4060
rect 39080 4020 39086 4032
rect 40865 4029 40877 4032
rect 40911 4029 40923 4063
rect 40865 4023 40923 4029
rect 41325 4063 41383 4069
rect 41325 4029 41337 4063
rect 41371 4060 41383 4063
rect 41414 4060 41420 4072
rect 41371 4032 41420 4060
rect 41371 4029 41383 4032
rect 41325 4023 41383 4029
rect 41414 4020 41420 4032
rect 41472 4020 41478 4072
rect 42705 4063 42763 4069
rect 42705 4029 42717 4063
rect 42751 4060 42763 4063
rect 42904 4060 42932 4091
rect 43254 4060 43260 4072
rect 42751 4032 42840 4060
rect 42904 4032 43260 4060
rect 42751 4029 42763 4032
rect 42705 4023 42763 4029
rect 40313 3995 40371 4001
rect 40313 3992 40325 3995
rect 38626 3964 40325 3992
rect 37642 3924 37648 3936
rect 37292 3896 37648 3924
rect 36817 3887 36875 3893
rect 37642 3884 37648 3896
rect 37700 3884 37706 3936
rect 38010 3884 38016 3936
rect 38068 3924 38074 3936
rect 38626 3924 38654 3964
rect 40313 3961 40325 3964
rect 40359 3961 40371 3995
rect 42812 3992 42840 4032
rect 43254 4020 43260 4032
rect 43312 4020 43318 4072
rect 43162 3992 43168 4004
rect 42812 3964 43168 3992
rect 40313 3955 40371 3961
rect 43162 3952 43168 3964
rect 43220 3952 43226 4004
rect 38068 3896 38654 3924
rect 38068 3884 38074 3896
rect 39574 3884 39580 3936
rect 39632 3884 39638 3936
rect 42058 3884 42064 3936
rect 42116 3924 42122 3936
rect 42153 3927 42211 3933
rect 42153 3924 42165 3927
rect 42116 3896 42165 3924
rect 42116 3884 42122 3896
rect 42153 3893 42165 3896
rect 42199 3893 42211 3927
rect 43364 3924 43392 4091
rect 43622 4088 43628 4091
rect 43680 4088 43686 4140
rect 43732 4128 43760 4168
rect 51905 4165 51917 4199
rect 51951 4196 51963 4199
rect 52748 4196 52776 4224
rect 53466 4196 53472 4208
rect 51951 4168 52776 4196
rect 52840 4168 53472 4196
rect 51951 4165 51963 4168
rect 51905 4159 51963 4165
rect 45097 4131 45155 4137
rect 43732 4100 45048 4128
rect 44910 4020 44916 4072
rect 44968 4020 44974 4072
rect 45020 4060 45048 4100
rect 45097 4097 45109 4131
rect 45143 4128 45155 4131
rect 46385 4131 46443 4137
rect 46385 4128 46397 4131
rect 45143 4100 46397 4128
rect 45143 4097 45155 4100
rect 45097 4091 45155 4097
rect 46385 4097 46397 4100
rect 46431 4097 46443 4131
rect 46385 4091 46443 4097
rect 48593 4131 48651 4137
rect 48593 4097 48605 4131
rect 48639 4128 48651 4131
rect 48682 4128 48688 4140
rect 48639 4100 48688 4128
rect 48639 4097 48651 4100
rect 48593 4091 48651 4097
rect 48682 4088 48688 4100
rect 48740 4088 48746 4140
rect 49786 4088 49792 4140
rect 49844 4088 49850 4140
rect 50341 4131 50399 4137
rect 50341 4097 50353 4131
rect 50387 4128 50399 4131
rect 51166 4128 51172 4140
rect 50387 4100 51172 4128
rect 50387 4097 50399 4100
rect 50341 4091 50399 4097
rect 51166 4088 51172 4100
rect 51224 4088 51230 4140
rect 51994 4088 52000 4140
rect 52052 4088 52058 4140
rect 52840 4128 52868 4168
rect 53466 4156 53472 4168
rect 53524 4156 53530 4208
rect 56060 4196 56088 4236
rect 56134 4224 56140 4276
rect 56192 4224 56198 4276
rect 56060 4168 58480 4196
rect 54202 4128 54208 4140
rect 52656 4100 52868 4128
rect 52932 4100 54208 4128
rect 46201 4063 46259 4069
rect 46201 4060 46213 4063
rect 45020 4032 46213 4060
rect 46201 4029 46213 4032
rect 46247 4029 46259 4063
rect 46201 4023 46259 4029
rect 46658 4020 46664 4072
rect 46716 4060 46722 4072
rect 46937 4063 46995 4069
rect 46937 4060 46949 4063
rect 46716 4032 46949 4060
rect 46716 4020 46722 4032
rect 46937 4029 46949 4032
rect 46983 4029 46995 4063
rect 46937 4023 46995 4029
rect 48130 4020 48136 4072
rect 48188 4020 48194 4072
rect 48409 4063 48467 4069
rect 48409 4029 48421 4063
rect 48455 4060 48467 4063
rect 49237 4063 49295 4069
rect 49237 4060 49249 4063
rect 48455 4032 49249 4060
rect 48455 4029 48467 4032
rect 48409 4023 48467 4029
rect 49237 4029 49249 4032
rect 49283 4029 49295 4063
rect 49237 4023 49295 4029
rect 49421 4063 49479 4069
rect 49421 4029 49433 4063
rect 49467 4060 49479 4063
rect 49804 4060 49832 4088
rect 49467 4032 49832 4060
rect 49467 4029 49479 4032
rect 49421 4023 49479 4029
rect 44928 3992 44956 4020
rect 46566 3992 46572 4004
rect 44928 3964 46572 3992
rect 46566 3952 46572 3964
rect 46624 3992 46630 4004
rect 47302 3992 47308 4004
rect 46624 3964 47308 3992
rect 46624 3952 46630 3964
rect 47302 3952 47308 3964
rect 47360 3992 47366 4004
rect 48424 3992 48452 4023
rect 47360 3964 48452 3992
rect 49252 3992 49280 4023
rect 50246 4020 50252 4072
rect 50304 4020 50310 4072
rect 51534 4060 51540 4072
rect 50448 4032 51540 4060
rect 49881 3995 49939 4001
rect 49252 3964 49372 3992
rect 47360 3952 47366 3964
rect 44266 3924 44272 3936
rect 43364 3896 44272 3924
rect 42153 3887 42211 3893
rect 44266 3884 44272 3896
rect 44324 3884 44330 3936
rect 44818 3884 44824 3936
rect 44876 3924 44882 3936
rect 45649 3927 45707 3933
rect 45649 3924 45661 3927
rect 44876 3896 45661 3924
rect 44876 3884 44882 3896
rect 45649 3893 45661 3896
rect 45695 3893 45707 3927
rect 45649 3887 45707 3893
rect 47578 3884 47584 3936
rect 47636 3884 47642 3936
rect 47762 3884 47768 3936
rect 47820 3924 47826 3936
rect 49234 3924 49240 3936
rect 47820 3896 49240 3924
rect 47820 3884 47826 3896
rect 49234 3884 49240 3896
rect 49292 3884 49298 3936
rect 49344 3924 49372 3964
rect 49881 3961 49893 3995
rect 49927 3992 49939 3995
rect 50448 3992 50476 4032
rect 51534 4020 51540 4032
rect 51592 4020 51598 4072
rect 51721 4063 51779 4069
rect 51721 4029 51733 4063
rect 51767 4029 51779 4063
rect 51721 4023 51779 4029
rect 51813 4063 51871 4069
rect 51813 4029 51825 4063
rect 51859 4060 51871 4063
rect 52012 4060 52040 4088
rect 51859 4032 52040 4060
rect 51859 4029 51871 4032
rect 51813 4023 51871 4029
rect 49927 3964 50476 3992
rect 50801 3995 50859 4001
rect 49927 3961 49939 3964
rect 49881 3955 49939 3961
rect 50801 3961 50813 3995
rect 50847 3992 50859 3995
rect 51350 3992 51356 4004
rect 50847 3964 51356 3992
rect 50847 3961 50859 3964
rect 50801 3955 50859 3961
rect 51350 3952 51356 3964
rect 51408 3952 51414 4004
rect 51736 3992 51764 4023
rect 52656 3992 52684 4100
rect 52730 4020 52736 4072
rect 52788 4060 52794 4072
rect 52825 4063 52883 4069
rect 52825 4060 52837 4063
rect 52788 4032 52837 4060
rect 52788 4020 52794 4032
rect 52825 4029 52837 4032
rect 52871 4029 52883 4063
rect 52825 4023 52883 4029
rect 51736 3964 52684 3992
rect 51169 3927 51227 3933
rect 51169 3924 51181 3927
rect 49344 3896 51181 3924
rect 51169 3893 51181 3896
rect 51215 3924 51227 3927
rect 51736 3924 51764 3964
rect 51215 3896 51764 3924
rect 52932 3924 52960 4100
rect 54202 4088 54208 4100
rect 54260 4128 54266 4140
rect 54481 4131 54539 4137
rect 54260 4100 54432 4128
rect 54260 4088 54266 4100
rect 53009 4063 53067 4069
rect 53009 4029 53021 4063
rect 53055 4060 53067 4063
rect 53282 4060 53288 4072
rect 53055 4032 53288 4060
rect 53055 4029 53067 4032
rect 53009 4023 53067 4029
rect 53282 4020 53288 4032
rect 53340 4060 53346 4072
rect 54018 4060 54024 4072
rect 53340 4032 54024 4060
rect 53340 4020 53346 4032
rect 54018 4020 54024 4032
rect 54076 4020 54082 4072
rect 54113 4063 54171 4069
rect 54113 4029 54125 4063
rect 54159 4029 54171 4063
rect 54113 4023 54171 4029
rect 54297 4063 54355 4069
rect 54297 4029 54309 4063
rect 54343 4029 54355 4063
rect 54404 4060 54432 4100
rect 54481 4097 54493 4131
rect 54527 4128 54539 4131
rect 54662 4128 54668 4140
rect 54527 4100 54668 4128
rect 54527 4097 54539 4100
rect 54481 4091 54539 4097
rect 54662 4088 54668 4100
rect 54720 4088 54726 4140
rect 55306 4088 55312 4140
rect 55364 4137 55370 4140
rect 55364 4131 55392 4137
rect 55380 4097 55392 4131
rect 55364 4091 55392 4097
rect 57701 4131 57759 4137
rect 57701 4097 57713 4131
rect 57747 4128 57759 4131
rect 57974 4128 57980 4140
rect 57747 4100 57980 4128
rect 57747 4097 57759 4100
rect 57701 4091 57759 4097
rect 55364 4088 55370 4091
rect 57974 4088 57980 4100
rect 58032 4088 58038 4140
rect 58452 4137 58480 4168
rect 58437 4131 58495 4137
rect 58437 4097 58449 4131
rect 58483 4097 58495 4131
rect 58437 4091 58495 4097
rect 55217 4063 55275 4069
rect 55217 4060 55229 4063
rect 54404 4032 55229 4060
rect 54297 4023 54355 4029
rect 55217 4029 55229 4032
rect 55263 4029 55275 4063
rect 55217 4023 55275 4029
rect 55493 4063 55551 4069
rect 55493 4029 55505 4063
rect 55539 4060 55551 4063
rect 56042 4060 56048 4072
rect 55539 4032 56048 4060
rect 55539 4029 55551 4032
rect 55493 4023 55551 4029
rect 53469 3995 53527 4001
rect 53469 3961 53481 3995
rect 53515 3992 53527 3995
rect 54128 3992 54156 4023
rect 53515 3964 54156 3992
rect 53515 3961 53527 3964
rect 53469 3955 53527 3961
rect 53098 3924 53104 3936
rect 52932 3896 53104 3924
rect 51215 3893 51227 3896
rect 51169 3887 51227 3893
rect 53098 3884 53104 3896
rect 53156 3884 53162 3936
rect 53374 3884 53380 3936
rect 53432 3924 53438 3936
rect 53561 3927 53619 3933
rect 53561 3924 53573 3927
rect 53432 3896 53573 3924
rect 53432 3884 53438 3896
rect 53561 3893 53573 3896
rect 53607 3893 53619 3927
rect 54312 3924 54340 4023
rect 56042 4020 56048 4032
rect 56100 4020 56106 4072
rect 57241 4063 57299 4069
rect 57241 4029 57253 4063
rect 57287 4060 57299 4063
rect 58342 4060 58348 4072
rect 57287 4032 58348 4060
rect 57287 4029 57299 4032
rect 57241 4023 57299 4029
rect 58342 4020 58348 4032
rect 58400 4020 58406 4072
rect 54754 3952 54760 4004
rect 54812 3992 54818 4004
rect 54941 3995 54999 4001
rect 54941 3992 54953 3995
rect 54812 3964 54953 3992
rect 54812 3952 54818 3964
rect 54941 3961 54953 3964
rect 54987 3961 54999 3995
rect 54941 3955 54999 3961
rect 56134 3952 56140 4004
rect 56192 3992 56198 4004
rect 58434 3992 58440 4004
rect 56192 3964 58440 3992
rect 56192 3952 56198 3964
rect 58434 3952 58440 3964
rect 58492 3952 58498 4004
rect 55582 3924 55588 3936
rect 54312 3896 55588 3924
rect 53561 3887 53619 3893
rect 55582 3884 55588 3896
rect 55640 3924 55646 3936
rect 57885 3927 57943 3933
rect 57885 3924 57897 3927
rect 55640 3896 57897 3924
rect 55640 3884 55646 3896
rect 57885 3893 57897 3896
rect 57931 3893 57943 3927
rect 57885 3887 57943 3893
rect 1104 3834 58880 3856
rect 1104 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 22616 3834
rect 22668 3782 22680 3834
rect 22732 3782 22744 3834
rect 22796 3782 22808 3834
rect 22860 3782 22872 3834
rect 22924 3782 37060 3834
rect 37112 3782 37124 3834
rect 37176 3782 37188 3834
rect 37240 3782 37252 3834
rect 37304 3782 37316 3834
rect 37368 3782 51504 3834
rect 51556 3782 51568 3834
rect 51620 3782 51632 3834
rect 51684 3782 51696 3834
rect 51748 3782 51760 3834
rect 51812 3782 58880 3834
rect 1104 3760 58880 3782
rect 3234 3680 3240 3732
rect 3292 3680 3298 3732
rect 3878 3680 3884 3732
rect 3936 3680 3942 3732
rect 4798 3680 4804 3732
rect 4856 3680 4862 3732
rect 4982 3680 4988 3732
rect 5040 3680 5046 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 5500 3692 7144 3720
rect 5500 3680 5506 3692
rect 3602 3544 3608 3596
rect 3660 3544 3666 3596
rect 4522 3544 4528 3596
rect 4580 3544 4586 3596
rect 4614 3544 4620 3596
rect 4672 3544 4678 3596
rect 4816 3584 4844 3680
rect 5810 3612 5816 3664
rect 5868 3612 5874 3664
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 4816 3556 5457 3584
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5828 3584 5856 3612
rect 5675 3556 5856 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1670 3516 1676 3528
rect 1627 3488 1676 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 1854 3525 1860 3528
rect 1848 3516 1860 3525
rect 1815 3488 1860 3516
rect 1848 3479 1860 3488
rect 1854 3476 1860 3479
rect 1912 3476 1918 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4632 3516 4660 3544
rect 4387 3488 4660 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 3436 3448 3464 3479
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5718 3476 5724 3528
rect 5776 3518 5782 3528
rect 5813 3519 5871 3525
rect 5813 3518 5825 3519
rect 5776 3490 5825 3518
rect 5776 3476 5782 3490
rect 5813 3485 5825 3490
rect 5859 3485 5871 3519
rect 7116 3516 7144 3692
rect 9766 3680 9772 3732
rect 9824 3680 9830 3732
rect 10778 3720 10784 3732
rect 10244 3692 10784 3720
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 10244 3652 10272 3692
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11020 3692 11192 3720
rect 11020 3680 11026 3692
rect 9723 3624 10272 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 7432 3556 7757 3584
rect 7432 3544 7438 3556
rect 7745 3553 7757 3556
rect 7791 3553 7803 3587
rect 11164 3584 11192 3692
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11425 3723 11483 3729
rect 11425 3720 11437 3723
rect 11388 3692 11437 3720
rect 11388 3680 11394 3692
rect 11425 3689 11437 3692
rect 11471 3689 11483 3723
rect 11425 3683 11483 3689
rect 11808 3692 13584 3720
rect 11808 3593 11836 3692
rect 11882 3612 11888 3664
rect 11940 3652 11946 3664
rect 11940 3624 12020 3652
rect 11940 3612 11946 3624
rect 11992 3593 12020 3624
rect 12342 3612 12348 3664
rect 12400 3612 12406 3664
rect 12434 3612 12440 3664
rect 12492 3612 12498 3664
rect 13556 3652 13584 3692
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13964 3692 14105 3720
rect 13964 3680 13970 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 14734 3680 14740 3732
rect 14792 3680 14798 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 16393 3723 16451 3729
rect 16393 3720 16405 3723
rect 14976 3692 16405 3720
rect 14976 3680 14982 3692
rect 16393 3689 16405 3692
rect 16439 3689 16451 3723
rect 16393 3683 16451 3689
rect 13556 3624 14688 3652
rect 11793 3587 11851 3593
rect 11793 3584 11805 3587
rect 11164 3556 11805 3584
rect 7745 3547 7803 3553
rect 11793 3553 11805 3556
rect 11839 3553 11851 3587
rect 11793 3547 11851 3553
rect 11977 3587 12035 3593
rect 11977 3553 11989 3587
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 7282 3516 7288 3528
rect 7116 3488 7288 3516
rect 5813 3479 5871 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 5258 3448 5264 3460
rect 3436 3420 5264 3448
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6058 3451 6116 3457
rect 6058 3448 6070 3451
rect 5960 3420 6070 3448
rect 5960 3408 5966 3420
rect 6058 3417 6070 3420
rect 6104 3417 6116 3451
rect 6058 3411 6116 3417
rect 6270 3408 6276 3460
rect 6328 3448 6334 3460
rect 6328 3420 7052 3448
rect 6328 3408 6334 3420
rect 2958 3340 2964 3392
rect 3016 3340 3022 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 5718 3380 5724 3392
rect 4304 3352 5724 3380
rect 4304 3340 4310 3352
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 7024 3380 7052 3420
rect 7190 3380 7196 3392
rect 7024 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 9140 3380 9168 3479
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 10882 3519 10940 3525
rect 10882 3516 10894 3519
rect 9732 3488 10894 3516
rect 9732 3476 9738 3488
rect 10882 3485 10894 3488
rect 10928 3485 10940 3519
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 10882 3479 10940 3485
rect 10980 3488 11161 3516
rect 10980 3460 11008 3488
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 12360 3516 12388 3612
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14660 3593 14688 3624
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 11655 3488 12388 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 12526 3476 12532 3528
rect 12584 3476 12590 3528
rect 12796 3519 12854 3525
rect 12796 3485 12808 3519
rect 12842 3516 12854 3519
rect 13078 3516 13084 3528
rect 12842 3488 13084 3516
rect 12842 3485 12854 3488
rect 12796 3479 12854 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14461 3519 14519 3525
rect 14461 3516 14473 3519
rect 14424 3488 14473 3516
rect 14424 3476 14430 3488
rect 14461 3485 14473 3488
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 10962 3408 10968 3460
rect 11020 3448 11026 3460
rect 12544 3448 12572 3476
rect 11020 3420 12572 3448
rect 11020 3408 11026 3420
rect 11146 3380 11152 3392
rect 9140 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 12069 3383 12127 3389
rect 12069 3349 12081 3383
rect 12115 3380 12127 3383
rect 12250 3380 12256 3392
rect 12115 3352 12256 3380
rect 12115 3349 12127 3352
rect 12069 3343 12127 3349
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3380 13967 3383
rect 13998 3380 14004 3392
rect 13955 3352 14004 3380
rect 13955 3349 13967 3352
rect 13909 3343 13967 3349
rect 13998 3340 14004 3352
rect 14056 3380 14062 3392
rect 14292 3380 14320 3476
rect 14056 3352 14320 3380
rect 14660 3380 14688 3547
rect 14752 3448 14780 3680
rect 15010 3544 15016 3596
rect 15068 3544 15074 3596
rect 15028 3516 15056 3544
rect 15746 3516 15752 3528
rect 15028 3488 15752 3516
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 15258 3451 15316 3457
rect 15258 3448 15270 3451
rect 14752 3420 15270 3448
rect 15258 3417 15270 3420
rect 15304 3417 15316 3451
rect 16408 3448 16436 3683
rect 16482 3680 16488 3732
rect 16540 3680 16546 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 19337 3723 19395 3729
rect 17000 3692 19104 3720
rect 17000 3680 17006 3692
rect 17494 3652 17500 3664
rect 17144 3624 17500 3652
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 17144 3593 17172 3624
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 17681 3655 17739 3661
rect 17681 3621 17693 3655
rect 17727 3652 17739 3655
rect 17862 3652 17868 3664
rect 17727 3624 17868 3652
rect 17727 3621 17739 3624
rect 17681 3615 17739 3621
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16724 3556 16957 3584
rect 16724 3544 16730 3556
rect 16945 3553 16957 3556
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 16850 3476 16856 3528
rect 16908 3476 16914 3528
rect 16666 3448 16672 3460
rect 16408 3420 16672 3448
rect 15258 3411 15316 3417
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 17512 3448 17540 3612
rect 19076 3593 19104 3692
rect 19337 3689 19349 3723
rect 19383 3720 19395 3723
rect 19518 3720 19524 3732
rect 19383 3692 19524 3720
rect 19383 3689 19395 3692
rect 19337 3683 19395 3689
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 20993 3723 21051 3729
rect 20993 3689 21005 3723
rect 21039 3720 21051 3723
rect 21174 3720 21180 3732
rect 21039 3692 21180 3720
rect 21039 3689 21051 3692
rect 20993 3683 21051 3689
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24213 3723 24271 3729
rect 24213 3720 24225 3723
rect 23532 3692 24225 3720
rect 23532 3680 23538 3692
rect 24213 3689 24225 3692
rect 24259 3720 24271 3723
rect 25130 3720 25136 3732
rect 24259 3692 25136 3720
rect 24259 3689 24271 3692
rect 24213 3683 24271 3689
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 27617 3723 27675 3729
rect 27617 3689 27629 3723
rect 27663 3720 27675 3723
rect 28074 3720 28080 3732
rect 27663 3692 28080 3720
rect 27663 3689 27675 3692
rect 27617 3683 27675 3689
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 29730 3680 29736 3732
rect 29788 3680 29794 3732
rect 32953 3723 33011 3729
rect 32953 3689 32965 3723
rect 32999 3720 33011 3723
rect 33318 3720 33324 3732
rect 32999 3692 33324 3720
rect 32999 3689 33011 3692
rect 32953 3683 33011 3689
rect 33318 3680 33324 3692
rect 33376 3720 33382 3732
rect 34146 3720 34152 3732
rect 33376 3692 34152 3720
rect 33376 3680 33382 3692
rect 34146 3680 34152 3692
rect 34204 3680 34210 3732
rect 34425 3723 34483 3729
rect 34425 3689 34437 3723
rect 34471 3720 34483 3723
rect 34882 3720 34888 3732
rect 34471 3692 34888 3720
rect 34471 3689 34483 3692
rect 34425 3683 34483 3689
rect 34882 3680 34888 3692
rect 34940 3680 34946 3732
rect 39022 3680 39028 3732
rect 39080 3680 39086 3732
rect 39301 3723 39359 3729
rect 39301 3689 39313 3723
rect 39347 3720 39359 3723
rect 39390 3720 39396 3732
rect 39347 3692 39396 3720
rect 39347 3689 39359 3692
rect 39301 3683 39359 3689
rect 39390 3680 39396 3692
rect 39448 3680 39454 3732
rect 39574 3680 39580 3732
rect 39632 3680 39638 3732
rect 40037 3723 40095 3729
rect 40037 3689 40049 3723
rect 40083 3720 40095 3723
rect 40402 3720 40408 3732
rect 40083 3692 40408 3720
rect 40083 3689 40095 3692
rect 40037 3683 40095 3689
rect 40402 3680 40408 3692
rect 40460 3680 40466 3732
rect 41782 3680 41788 3732
rect 41840 3680 41846 3732
rect 41966 3680 41972 3732
rect 42024 3720 42030 3732
rect 42024 3692 42564 3720
rect 42024 3680 42030 3692
rect 19061 3587 19119 3593
rect 19061 3553 19073 3587
rect 19107 3584 19119 3587
rect 39592 3584 39620 3680
rect 41690 3612 41696 3664
rect 41748 3652 41754 3664
rect 41984 3652 42012 3680
rect 41748 3624 42012 3652
rect 41748 3612 41754 3624
rect 19107 3556 19656 3584
rect 19107 3553 19119 3556
rect 19061 3547 19119 3553
rect 18782 3476 18788 3528
rect 18840 3525 18846 3528
rect 18840 3516 18852 3525
rect 18840 3488 18885 3516
rect 18840 3479 18852 3488
rect 18840 3476 18846 3479
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19628 3525 19656 3556
rect 35728 3556 37688 3584
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19484 3488 19533 3516
rect 19484 3476 19490 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 19702 3516 19708 3528
rect 19659 3488 19708 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 19886 3525 19892 3528
rect 19880 3516 19892 3525
rect 19847 3488 19892 3516
rect 19880 3479 19892 3488
rect 19886 3476 19892 3479
rect 19944 3476 19950 3528
rect 22186 3476 22192 3528
rect 22244 3525 22250 3528
rect 22244 3479 22256 3525
rect 22244 3476 22250 3479
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22833 3519 22891 3525
rect 22833 3516 22845 3519
rect 22520 3488 22845 3516
rect 22520 3476 22526 3488
rect 22833 3485 22845 3488
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23100 3519 23158 3525
rect 23100 3485 23112 3519
rect 23146 3485 23158 3519
rect 23100 3479 23158 3485
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 25498 3516 25504 3528
rect 24811 3488 25504 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 20806 3448 20812 3460
rect 17512 3420 20812 3448
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 16390 3380 16396 3392
rect 14660 3352 16396 3380
rect 14056 3340 14062 3352
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 21082 3340 21088 3392
rect 21140 3340 21146 3392
rect 22848 3380 22876 3479
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 23124 3448 23152 3479
rect 24780 3448 24808 3479
rect 25498 3476 25504 3488
rect 25556 3516 25562 3528
rect 26237 3519 26295 3525
rect 26237 3516 26249 3519
rect 25556 3488 26249 3516
rect 25556 3476 25562 3488
rect 26237 3485 26249 3488
rect 26283 3485 26295 3519
rect 26237 3479 26295 3485
rect 26504 3519 26562 3525
rect 26504 3485 26516 3519
rect 26550 3516 26562 3519
rect 26786 3516 26792 3528
rect 26550 3488 26792 3516
rect 26550 3485 26562 3488
rect 26504 3479 26562 3485
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 27982 3476 27988 3528
rect 28040 3516 28046 3528
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 28040 3488 28457 3516
rect 28040 3476 28046 3488
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 28810 3476 28816 3528
rect 28868 3476 28874 3528
rect 29086 3476 29092 3528
rect 29144 3516 29150 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29144 3488 29561 3516
rect 29144 3476 29150 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 29917 3519 29975 3525
rect 29917 3485 29929 3519
rect 29963 3516 29975 3519
rect 31573 3519 31631 3525
rect 31573 3516 31585 3519
rect 29963 3488 31585 3516
rect 29963 3485 29975 3488
rect 29917 3479 29975 3485
rect 31573 3485 31585 3488
rect 31619 3516 31631 3519
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 31619 3488 33057 3516
rect 31619 3485 31631 3488
rect 31573 3479 31631 3485
rect 33045 3485 33057 3488
rect 33091 3516 33103 3519
rect 34698 3516 34704 3528
rect 33091 3488 34704 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 34698 3476 34704 3488
rect 34756 3516 34762 3528
rect 35728 3516 35756 3556
rect 37660 3525 37688 3556
rect 38764 3556 39620 3584
rect 39669 3587 39727 3593
rect 34756 3488 35756 3516
rect 36357 3519 36415 3525
rect 34756 3476 34762 3488
rect 36357 3485 36369 3519
rect 36403 3516 36415 3519
rect 37645 3519 37703 3525
rect 36403 3488 36860 3516
rect 36403 3485 36415 3488
rect 36357 3479 36415 3485
rect 23072 3420 23152 3448
rect 23216 3420 24808 3448
rect 23072 3408 23078 3420
rect 23216 3380 23244 3420
rect 24854 3408 24860 3460
rect 24912 3448 24918 3460
rect 25010 3451 25068 3457
rect 25010 3448 25022 3451
rect 24912 3420 25022 3448
rect 24912 3408 24918 3420
rect 25010 3417 25022 3420
rect 25056 3417 25068 3451
rect 25010 3411 25068 3417
rect 25590 3408 25596 3460
rect 25648 3408 25654 3460
rect 29365 3451 29423 3457
rect 29365 3417 29377 3451
rect 29411 3448 29423 3451
rect 30162 3451 30220 3457
rect 30162 3448 30174 3451
rect 29411 3420 30174 3448
rect 29411 3417 29423 3420
rect 29365 3411 29423 3417
rect 30162 3417 30174 3420
rect 30208 3417 30220 3451
rect 30162 3411 30220 3417
rect 31840 3451 31898 3457
rect 31840 3417 31852 3451
rect 31886 3448 31898 3451
rect 32858 3448 32864 3460
rect 31886 3420 32864 3448
rect 31886 3417 31898 3420
rect 31840 3411 31898 3417
rect 32858 3408 32864 3420
rect 32916 3408 32922 3460
rect 33312 3451 33370 3457
rect 33312 3417 33324 3451
rect 33358 3448 33370 3451
rect 33594 3448 33600 3460
rect 33358 3420 33600 3448
rect 33358 3417 33370 3420
rect 33312 3411 33370 3417
rect 33594 3408 33600 3420
rect 33652 3408 33658 3460
rect 34968 3451 35026 3457
rect 34968 3417 34980 3451
rect 35014 3448 35026 3451
rect 35710 3448 35716 3460
rect 35014 3420 35716 3448
rect 35014 3417 35026 3420
rect 34968 3411 35026 3417
rect 35710 3408 35716 3420
rect 35768 3408 35774 3460
rect 22848 3352 23244 3380
rect 24673 3383 24731 3389
rect 24673 3349 24685 3383
rect 24719 3380 24731 3383
rect 25608 3380 25636 3408
rect 24719 3352 25636 3380
rect 26145 3383 26203 3389
rect 24719 3349 24731 3352
rect 24673 3343 24731 3349
rect 26145 3349 26157 3383
rect 26191 3380 26203 3383
rect 26602 3380 26608 3392
rect 26191 3352 26608 3380
rect 26191 3349 26203 3352
rect 26145 3343 26203 3349
rect 26602 3340 26608 3352
rect 26660 3340 26666 3392
rect 27890 3340 27896 3392
rect 27948 3340 27954 3392
rect 31297 3383 31355 3389
rect 31297 3349 31309 3383
rect 31343 3380 31355 3383
rect 31938 3380 31944 3392
rect 31343 3352 31944 3380
rect 31343 3349 31355 3352
rect 31297 3343 31355 3349
rect 31938 3340 31944 3352
rect 31996 3340 32002 3392
rect 36081 3383 36139 3389
rect 36081 3349 36093 3383
rect 36127 3380 36139 3383
rect 36372 3380 36400 3479
rect 36832 3392 36860 3488
rect 37645 3485 37657 3519
rect 37691 3516 37703 3519
rect 37734 3516 37740 3528
rect 37691 3488 37740 3516
rect 37691 3485 37703 3488
rect 37645 3479 37703 3485
rect 37734 3476 37740 3488
rect 37792 3476 37798 3528
rect 37912 3519 37970 3525
rect 37912 3485 37924 3519
rect 37958 3516 37970 3519
rect 38764 3516 38792 3556
rect 39669 3553 39681 3587
rect 39715 3584 39727 3587
rect 39758 3584 39764 3596
rect 39715 3556 39764 3584
rect 39715 3553 39727 3556
rect 39669 3547 39727 3553
rect 39758 3544 39764 3556
rect 39816 3584 39822 3596
rect 39816 3556 40540 3584
rect 39816 3544 39822 3556
rect 37958 3488 38792 3516
rect 37958 3485 37970 3488
rect 37912 3479 37970 3485
rect 39114 3476 39120 3528
rect 39172 3476 39178 3528
rect 39850 3476 39856 3528
rect 39908 3476 39914 3528
rect 40405 3519 40463 3525
rect 40405 3485 40417 3519
rect 40451 3485 40463 3519
rect 40405 3479 40463 3485
rect 37090 3408 37096 3460
rect 37148 3408 37154 3460
rect 40420 3392 40448 3479
rect 36127 3352 36400 3380
rect 36127 3349 36139 3352
rect 36081 3343 36139 3349
rect 36814 3340 36820 3392
rect 36872 3340 36878 3392
rect 40402 3340 40408 3392
rect 40460 3340 40466 3392
rect 40512 3380 40540 3556
rect 42334 3544 42340 3596
rect 42392 3544 42398 3596
rect 42536 3593 42564 3692
rect 42886 3680 42892 3732
rect 42944 3680 42950 3732
rect 43162 3680 43168 3732
rect 43220 3720 43226 3732
rect 43346 3720 43352 3732
rect 43220 3692 43352 3720
rect 43220 3680 43226 3692
rect 43346 3680 43352 3692
rect 43404 3720 43410 3732
rect 44542 3720 44548 3732
rect 43404 3692 44548 3720
rect 43404 3680 43410 3692
rect 44542 3680 44548 3692
rect 44600 3680 44606 3732
rect 46385 3723 46443 3729
rect 46385 3689 46397 3723
rect 46431 3720 46443 3723
rect 46658 3720 46664 3732
rect 46431 3692 46664 3720
rect 46431 3689 46443 3692
rect 46385 3683 46443 3689
rect 46658 3680 46664 3692
rect 46716 3680 46722 3732
rect 48958 3680 48964 3732
rect 49016 3680 49022 3732
rect 49329 3723 49387 3729
rect 49329 3689 49341 3723
rect 49375 3720 49387 3723
rect 49878 3720 49884 3732
rect 49375 3692 49884 3720
rect 49375 3689 49387 3692
rect 49329 3683 49387 3689
rect 49878 3680 49884 3692
rect 49936 3680 49942 3732
rect 52730 3680 52736 3732
rect 52788 3720 52794 3732
rect 52914 3720 52920 3732
rect 52788 3692 52920 3720
rect 52788 3680 52794 3692
rect 52914 3680 52920 3692
rect 52972 3680 52978 3732
rect 53190 3680 53196 3732
rect 53248 3680 53254 3732
rect 53926 3720 53932 3732
rect 53300 3692 53932 3720
rect 48976 3652 49004 3680
rect 49605 3655 49663 3661
rect 49605 3652 49617 3655
rect 48976 3624 49617 3652
rect 49605 3621 49617 3624
rect 49651 3621 49663 3655
rect 49605 3615 49663 3621
rect 49712 3624 51212 3652
rect 42521 3587 42579 3593
rect 42521 3553 42533 3587
rect 42567 3553 42579 3587
rect 42521 3547 42579 3553
rect 40672 3519 40730 3525
rect 40672 3485 40684 3519
rect 40718 3516 40730 3519
rect 41874 3516 41880 3528
rect 40718 3488 41880 3516
rect 40718 3485 40730 3488
rect 40672 3479 40730 3485
rect 41874 3476 41880 3488
rect 41932 3476 41938 3528
rect 42242 3476 42248 3528
rect 42300 3476 42306 3528
rect 42536 3516 42564 3547
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45005 3587 45063 3593
rect 45005 3584 45017 3587
rect 44324 3556 45017 3584
rect 44324 3544 44330 3556
rect 45005 3553 45017 3556
rect 45051 3553 45063 3587
rect 49712 3584 49740 3624
rect 45005 3547 45063 3553
rect 48976 3556 49740 3584
rect 44013 3519 44071 3525
rect 42536 3488 43944 3516
rect 41138 3408 41144 3460
rect 41196 3448 41202 3460
rect 43806 3448 43812 3460
rect 41196 3420 43812 3448
rect 41196 3408 41202 3420
rect 43806 3408 43812 3420
rect 43864 3408 43870 3460
rect 43916 3448 43944 3488
rect 44013 3485 44025 3519
rect 44059 3516 44071 3519
rect 44818 3516 44824 3528
rect 44059 3488 44824 3516
rect 44059 3485 44071 3488
rect 44013 3479 44071 3485
rect 44818 3476 44824 3488
rect 44876 3476 44882 3528
rect 45020 3516 45048 3547
rect 46477 3519 46535 3525
rect 46477 3516 46489 3519
rect 45020 3488 46489 3516
rect 46477 3485 46489 3488
rect 46523 3516 46535 3519
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 46523 3488 47961 3516
rect 46523 3485 46535 3488
rect 46477 3479 46535 3485
rect 47949 3485 47961 3488
rect 47995 3516 48007 3519
rect 48498 3516 48504 3528
rect 47995 3488 48504 3516
rect 47995 3485 48007 3488
rect 47949 3479 48007 3485
rect 48498 3476 48504 3488
rect 48556 3516 48562 3528
rect 48976 3516 49004 3556
rect 50246 3544 50252 3596
rect 50304 3584 50310 3596
rect 50801 3587 50859 3593
rect 50801 3584 50813 3587
rect 50304 3556 50813 3584
rect 50304 3544 50310 3556
rect 50801 3553 50813 3556
rect 50847 3553 50859 3587
rect 50801 3547 50859 3553
rect 51184 3528 51212 3624
rect 53300 3593 53328 3692
rect 53926 3680 53932 3692
rect 53984 3720 53990 3732
rect 56502 3720 56508 3732
rect 53984 3692 56508 3720
rect 53984 3680 53990 3692
rect 54665 3655 54723 3661
rect 54665 3621 54677 3655
rect 54711 3652 54723 3655
rect 54846 3652 54852 3664
rect 54711 3624 54852 3652
rect 54711 3621 54723 3624
rect 54665 3615 54723 3621
rect 54846 3612 54852 3624
rect 54904 3612 54910 3664
rect 54938 3612 54944 3664
rect 54996 3612 55002 3664
rect 55582 3612 55588 3664
rect 55640 3612 55646 3664
rect 53285 3587 53343 3593
rect 53285 3553 53297 3587
rect 53331 3553 53343 3587
rect 53285 3547 53343 3553
rect 48556 3488 49004 3516
rect 48556 3476 48562 3488
rect 49142 3476 49148 3528
rect 49200 3476 49206 3528
rect 49789 3519 49847 3525
rect 49789 3485 49801 3519
rect 49835 3485 49847 3519
rect 49789 3479 49847 3485
rect 44910 3448 44916 3460
rect 43916 3420 44916 3448
rect 44910 3408 44916 3420
rect 44968 3408 44974 3460
rect 45272 3451 45330 3457
rect 45272 3417 45284 3451
rect 45318 3448 45330 3451
rect 45462 3448 45468 3460
rect 45318 3420 45468 3448
rect 45318 3417 45330 3420
rect 45272 3411 45330 3417
rect 45462 3408 45468 3420
rect 45520 3408 45526 3460
rect 46744 3451 46802 3457
rect 46744 3417 46756 3451
rect 46790 3448 46802 3451
rect 47578 3448 47584 3460
rect 46790 3420 47584 3448
rect 46790 3417 46802 3420
rect 46744 3411 46802 3417
rect 47578 3408 47584 3420
rect 47636 3408 47642 3460
rect 48216 3451 48274 3457
rect 48216 3417 48228 3451
rect 48262 3448 48274 3451
rect 49160 3448 49188 3476
rect 48262 3420 49188 3448
rect 48262 3417 48274 3420
rect 48216 3411 48274 3417
rect 41690 3380 41696 3392
rect 40512 3352 41696 3380
rect 41690 3340 41696 3352
rect 41748 3340 41754 3392
rect 41874 3340 41880 3392
rect 41932 3340 41938 3392
rect 46106 3340 46112 3392
rect 46164 3380 46170 3392
rect 47670 3380 47676 3392
rect 46164 3352 47676 3380
rect 46164 3340 46170 3352
rect 47670 3340 47676 3352
rect 47728 3340 47734 3392
rect 47857 3383 47915 3389
rect 47857 3349 47869 3383
rect 47903 3380 47915 3383
rect 48774 3380 48780 3392
rect 47903 3352 48780 3380
rect 47903 3349 47915 3352
rect 47857 3343 47915 3349
rect 48774 3340 48780 3352
rect 48832 3340 48838 3392
rect 49804 3380 49832 3479
rect 50522 3476 50528 3528
rect 50580 3476 50586 3528
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 51813 3519 51871 3525
rect 51813 3516 51825 3519
rect 51224 3488 51825 3516
rect 51224 3476 51230 3488
rect 51813 3485 51825 3488
rect 51859 3516 51871 3519
rect 53300 3516 53328 3547
rect 54294 3544 54300 3596
rect 54352 3584 54358 3596
rect 55401 3587 55459 3593
rect 55401 3584 55413 3587
rect 54352 3556 55413 3584
rect 54352 3544 54358 3556
rect 55401 3553 55413 3556
rect 55447 3553 55459 3587
rect 55401 3547 55459 3553
rect 51859 3488 53328 3516
rect 51859 3485 51871 3488
rect 51813 3479 51871 3485
rect 53374 3476 53380 3528
rect 53432 3476 53438 3528
rect 53558 3525 53564 3528
rect 53552 3516 53564 3525
rect 53519 3488 53564 3516
rect 53552 3479 53564 3488
rect 53558 3476 53564 3479
rect 53616 3476 53622 3528
rect 55600 3525 55628 3612
rect 56244 3593 56272 3692
rect 56502 3680 56508 3692
rect 56560 3680 56566 3732
rect 57701 3723 57759 3729
rect 57701 3689 57713 3723
rect 57747 3720 57759 3723
rect 57882 3720 57888 3732
rect 57747 3692 57888 3720
rect 57747 3689 57759 3692
rect 57701 3683 57759 3689
rect 57882 3680 57888 3692
rect 57940 3680 57946 3732
rect 57609 3655 57667 3661
rect 57609 3621 57621 3655
rect 57655 3652 57667 3655
rect 57790 3652 57796 3664
rect 57655 3624 57796 3652
rect 57655 3621 57667 3624
rect 57609 3615 57667 3621
rect 57790 3612 57796 3624
rect 57848 3612 57854 3664
rect 56229 3587 56287 3593
rect 56229 3553 56241 3587
rect 56275 3553 56287 3587
rect 56229 3547 56287 3553
rect 58158 3544 58164 3596
rect 58216 3544 58222 3596
rect 58253 3587 58311 3593
rect 58253 3553 58265 3587
rect 58299 3553 58311 3587
rect 58253 3547 58311 3553
rect 54757 3519 54815 3525
rect 54757 3485 54769 3519
rect 54803 3485 54815 3519
rect 54757 3479 54815 3485
rect 55585 3519 55643 3525
rect 55585 3485 55597 3519
rect 55631 3485 55643 3519
rect 55585 3479 55643 3485
rect 56496 3519 56554 3525
rect 56496 3485 56508 3519
rect 56542 3516 56554 3519
rect 57698 3516 57704 3528
rect 56542 3488 57704 3516
rect 56542 3485 56554 3488
rect 56496 3479 56554 3485
rect 52080 3451 52138 3457
rect 52080 3417 52092 3451
rect 52126 3448 52138 3451
rect 53392 3448 53420 3476
rect 52126 3420 53420 3448
rect 52126 3417 52138 3420
rect 52080 3411 52138 3417
rect 54202 3408 54208 3460
rect 54260 3408 54266 3460
rect 54772 3448 54800 3479
rect 57698 3476 57704 3488
rect 57756 3476 57762 3528
rect 58066 3476 58072 3528
rect 58124 3476 58130 3528
rect 56594 3448 56600 3460
rect 54772 3420 56600 3448
rect 56594 3408 56600 3420
rect 56652 3408 56658 3460
rect 56686 3408 56692 3460
rect 56744 3408 56750 3460
rect 57422 3408 57428 3460
rect 57480 3448 57486 3460
rect 58268 3448 58296 3547
rect 57480 3420 58296 3448
rect 57480 3408 57486 3420
rect 54220 3380 54248 3408
rect 49804 3352 54248 3380
rect 55490 3340 55496 3392
rect 55548 3380 55554 3392
rect 55677 3383 55735 3389
rect 55677 3380 55689 3383
rect 55548 3352 55689 3380
rect 55548 3340 55554 3352
rect 55677 3349 55689 3352
rect 55723 3349 55735 3383
rect 55677 3343 55735 3349
rect 56045 3383 56103 3389
rect 56045 3349 56057 3383
rect 56091 3380 56103 3383
rect 56704 3380 56732 3408
rect 56091 3352 56732 3380
rect 56091 3349 56103 3352
rect 56045 3343 56103 3349
rect 57698 3340 57704 3392
rect 57756 3380 57762 3392
rect 58526 3380 58532 3392
rect 57756 3352 58532 3380
rect 57756 3340 57762 3352
rect 58526 3340 58532 3352
rect 58584 3340 58590 3392
rect 1104 3290 59040 3312
rect 1104 3238 15394 3290
rect 15446 3238 15458 3290
rect 15510 3238 15522 3290
rect 15574 3238 15586 3290
rect 15638 3238 15650 3290
rect 15702 3238 29838 3290
rect 29890 3238 29902 3290
rect 29954 3238 29966 3290
rect 30018 3238 30030 3290
rect 30082 3238 30094 3290
rect 30146 3238 44282 3290
rect 44334 3238 44346 3290
rect 44398 3238 44410 3290
rect 44462 3238 44474 3290
rect 44526 3238 44538 3290
rect 44590 3238 58726 3290
rect 58778 3238 58790 3290
rect 58842 3238 58854 3290
rect 58906 3238 58918 3290
rect 58970 3238 58982 3290
rect 59034 3238 59040 3290
rect 1104 3216 59040 3238
rect 2774 3136 2780 3188
rect 2832 3136 2838 3188
rect 2866 3136 2872 3188
rect 2924 3136 2930 3188
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 5074 3176 5080 3188
rect 4295 3148 5080 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3176 5503 3179
rect 5491 3148 6776 3176
rect 5491 3145 5503 3148
rect 5445 3139 5503 3145
rect 1578 3068 1584 3120
rect 1636 3068 1642 3120
rect 2884 3108 2912 3136
rect 3114 3111 3172 3117
rect 3114 3108 3126 3111
rect 1688 3080 2820 3108
rect 2884 3080 3126 3108
rect 1688 3052 1716 3080
rect 1670 3000 1676 3052
rect 1728 3000 1734 3052
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2222 3040 2228 3052
rect 1995 3012 2228 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2792 3040 2820 3080
rect 3114 3077 3126 3080
rect 3160 3077 3172 3111
rect 3114 3071 3172 3077
rect 3252 3080 5580 3108
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2792 3012 2881 3040
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 3252 3040 3280 3080
rect 2869 3003 2927 3009
rect 2976 3012 3280 3040
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2976 2972 3004 3012
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 5552 2984 5580 3080
rect 5810 3068 5816 3120
rect 5868 3108 5874 3120
rect 5868 3080 6408 3108
rect 5868 3068 5874 3080
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5776 3012 5917 3040
rect 5776 3000 5782 3012
rect 5905 3009 5917 3012
rect 5951 3040 5963 3043
rect 5994 3040 6000 3052
rect 5951 3012 6000 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 6380 3049 6408 3080
rect 6638 3049 6644 3052
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6632 3040 6644 3049
rect 6599 3012 6644 3040
rect 6365 3003 6423 3009
rect 6632 3003 6644 3012
rect 2179 2944 3004 2972
rect 4893 2975 4951 2981
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 4893 2941 4905 2975
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 4908 2904 4936 2935
rect 5534 2932 5540 2984
rect 5592 2932 5598 2984
rect 5994 2904 6000 2916
rect 4908 2876 6000 2904
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 4617 2839 4675 2845
rect 4617 2805 4629 2839
rect 4663 2836 4675 2839
rect 5626 2836 5632 2848
rect 4663 2808 5632 2836
rect 4663 2805 4675 2808
rect 4617 2799 4675 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 6104 2836 6132 3003
rect 6638 3000 6644 3003
rect 6696 3000 6702 3052
rect 6748 3040 6776 3148
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7340 3148 7757 3176
rect 7340 3136 7346 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 7984 3148 8217 3176
rect 7984 3136 7990 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 11974 3136 11980 3188
rect 12032 3136 12038 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12124 3148 12173 3176
rect 12124 3136 12130 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 14277 3179 14335 3185
rect 14277 3145 14289 3179
rect 14323 3176 14335 3179
rect 15378 3176 15384 3188
rect 14323 3148 15384 3176
rect 14323 3145 14335 3148
rect 14277 3139 14335 3145
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 16390 3136 16396 3188
rect 16448 3136 16454 3188
rect 16758 3136 16764 3188
rect 16816 3136 16822 3188
rect 18046 3136 18052 3188
rect 18104 3136 18110 3188
rect 20806 3136 20812 3188
rect 20864 3136 20870 3188
rect 21450 3136 21456 3188
rect 21508 3176 21514 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21508 3148 21833 3176
rect 21508 3136 21514 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 22189 3179 22247 3185
rect 22189 3145 22201 3179
rect 22235 3176 22247 3179
rect 22278 3176 22284 3188
rect 22235 3148 22284 3176
rect 22235 3145 22247 3148
rect 22189 3139 22247 3145
rect 22278 3136 22284 3148
rect 22336 3136 22342 3188
rect 22925 3179 22983 3185
rect 22925 3145 22937 3179
rect 22971 3176 22983 3179
rect 23106 3176 23112 3188
rect 22971 3148 23112 3176
rect 22971 3145 22983 3148
rect 22925 3139 22983 3145
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 25280 3148 25513 3176
rect 25280 3136 25286 3148
rect 25501 3145 25513 3148
rect 25547 3145 25559 3179
rect 25501 3139 25559 3145
rect 25961 3179 26019 3185
rect 25961 3145 25973 3179
rect 26007 3176 26019 3179
rect 26050 3176 26056 3188
rect 26007 3148 26056 3176
rect 26007 3145 26019 3148
rect 25961 3139 26019 3145
rect 26050 3136 26056 3148
rect 26108 3136 26114 3188
rect 26234 3136 26240 3188
rect 26292 3136 26298 3188
rect 26697 3179 26755 3185
rect 26697 3145 26709 3179
rect 26743 3176 26755 3179
rect 27062 3176 27068 3188
rect 26743 3148 27068 3176
rect 26743 3145 26755 3148
rect 26697 3139 26755 3145
rect 27062 3136 27068 3148
rect 27120 3136 27126 3188
rect 27890 3136 27896 3188
rect 27948 3136 27954 3188
rect 28810 3136 28816 3188
rect 28868 3176 28874 3188
rect 30377 3179 30435 3185
rect 30377 3176 30389 3179
rect 28868 3148 30389 3176
rect 28868 3136 28874 3148
rect 30377 3145 30389 3148
rect 30423 3145 30435 3179
rect 30377 3139 30435 3145
rect 30745 3179 30803 3185
rect 30745 3145 30757 3179
rect 30791 3176 30803 3179
rect 31478 3176 31484 3188
rect 30791 3148 31484 3176
rect 30791 3145 30803 3148
rect 30745 3139 30803 3145
rect 31478 3136 31484 3148
rect 31536 3136 31542 3188
rect 31570 3136 31576 3188
rect 31628 3136 31634 3188
rect 32490 3136 32496 3188
rect 32548 3136 32554 3188
rect 32861 3179 32919 3185
rect 32861 3145 32873 3179
rect 32907 3176 32919 3179
rect 33134 3176 33140 3188
rect 32907 3148 33140 3176
rect 32907 3145 32919 3148
rect 32861 3139 32919 3145
rect 33134 3136 33140 3148
rect 33192 3136 33198 3188
rect 33226 3136 33232 3188
rect 33284 3136 33290 3188
rect 33321 3179 33379 3185
rect 33321 3145 33333 3179
rect 33367 3176 33379 3179
rect 34330 3176 34336 3188
rect 33367 3148 34336 3176
rect 33367 3145 33379 3148
rect 33321 3139 33379 3145
rect 34330 3136 34336 3148
rect 34388 3136 34394 3188
rect 35986 3136 35992 3188
rect 36044 3136 36050 3188
rect 36265 3179 36323 3185
rect 36265 3145 36277 3179
rect 36311 3176 36323 3179
rect 36354 3176 36360 3188
rect 36311 3148 36360 3176
rect 36311 3145 36323 3148
rect 36265 3139 36323 3145
rect 36354 3136 36360 3148
rect 36412 3136 36418 3188
rect 36906 3136 36912 3188
rect 36964 3176 36970 3188
rect 37277 3179 37335 3185
rect 37277 3176 37289 3179
rect 36964 3148 37289 3176
rect 36964 3136 36970 3148
rect 37277 3145 37289 3148
rect 37323 3145 37335 3179
rect 37277 3139 37335 3145
rect 39393 3179 39451 3185
rect 39393 3145 39405 3179
rect 39439 3176 39451 3179
rect 39666 3176 39672 3188
rect 39439 3148 39672 3176
rect 39439 3145 39451 3148
rect 39393 3139 39451 3145
rect 39666 3136 39672 3148
rect 39724 3136 39730 3188
rect 39850 3136 39856 3188
rect 39908 3176 39914 3188
rect 40129 3179 40187 3185
rect 40129 3176 40141 3179
rect 39908 3148 40141 3176
rect 39908 3136 39914 3148
rect 40129 3145 40141 3148
rect 40175 3145 40187 3179
rect 40129 3139 40187 3145
rect 41785 3179 41843 3185
rect 41785 3145 41797 3179
rect 41831 3145 41843 3179
rect 41785 3139 41843 3145
rect 42061 3179 42119 3185
rect 42061 3145 42073 3179
rect 42107 3176 42119 3179
rect 42150 3176 42156 3188
rect 42107 3148 42156 3176
rect 42107 3145 42119 3148
rect 42061 3139 42119 3145
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 10962 3108 10968 3120
rect 8076 3080 10968 3108
rect 8076 3068 8082 3080
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 6748 3012 8125 3040
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 9600 3049 9628 3080
rect 10962 3068 10968 3080
rect 11020 3108 11026 3120
rect 15504 3111 15562 3117
rect 11020 3080 11376 3108
rect 11020 3068 11026 3080
rect 9318 3043 9376 3049
rect 9318 3040 9330 3043
rect 8628 3012 9330 3040
rect 8628 3000 8634 3012
rect 9318 3009 9330 3012
rect 9364 3009 9376 3043
rect 9318 3003 9376 3009
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 11077 3043 11135 3049
rect 11077 3009 11089 3043
rect 11123 3040 11135 3043
rect 11238 3040 11244 3052
rect 11123 3012 11244 3040
rect 11123 3009 11135 3012
rect 11077 3003 11135 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11348 3049 11376 3080
rect 12544 3080 13584 3108
rect 12544 3052 12572 3080
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3009 11391 3043
rect 11333 3003 11391 3009
rect 11790 3000 11796 3052
rect 11848 3000 11854 3052
rect 12526 3000 12532 3052
rect 12584 3000 12590 3052
rect 13262 3000 13268 3052
rect 13320 3049 13326 3052
rect 13556 3049 13584 3080
rect 15504 3077 15516 3111
rect 15550 3108 15562 3111
rect 15838 3108 15844 3120
rect 15550 3080 15844 3108
rect 15550 3077 15562 3080
rect 15504 3071 15562 3077
rect 15838 3068 15844 3080
rect 15896 3068 15902 3120
rect 17954 3108 17960 3120
rect 17328 3080 17960 3108
rect 13320 3040 13332 3049
rect 13541 3043 13599 3049
rect 13320 3012 13365 3040
rect 13320 3003 13332 3012
rect 13541 3009 13553 3043
rect 13587 3009 13599 3043
rect 15194 3040 15200 3052
rect 13541 3003 13599 3009
rect 14752 3012 15200 3040
rect 13320 3000 13326 3003
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2972 13783 2975
rect 14752 2972 14780 3012
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 15746 3049 15752 3052
rect 15742 3003 15752 3049
rect 15804 3040 15810 3052
rect 15933 3043 15991 3049
rect 15804 3012 15842 3040
rect 15746 3000 15752 3003
rect 15804 3000 15810 3012
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 13771 2944 14320 2972
rect 13771 2941 13783 2944
rect 13725 2935 13783 2941
rect 7929 2907 7987 2913
rect 7929 2904 7941 2907
rect 7300 2876 7941 2904
rect 7300 2836 7328 2876
rect 7929 2873 7941 2876
rect 7975 2873 7987 2907
rect 7929 2867 7987 2873
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 11388 2876 12434 2904
rect 11388 2864 11394 2876
rect 6104 2808 7328 2836
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2836 10011 2839
rect 11146 2836 11152 2848
rect 9999 2808 11152 2836
rect 9999 2805 10011 2808
rect 9953 2799 10011 2805
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12406 2836 12434 2876
rect 12894 2836 12900 2848
rect 12406 2808 12900 2836
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 14292 2836 14320 2944
rect 14384 2944 14780 2972
rect 14384 2913 14412 2944
rect 14369 2907 14427 2913
rect 14369 2873 14381 2907
rect 14415 2873 14427 2907
rect 15948 2904 15976 3003
rect 16132 2972 16160 3003
rect 16942 3000 16948 3052
rect 17000 3000 17006 3052
rect 17328 2972 17356 3080
rect 17954 3068 17960 3080
rect 18012 3108 18018 3120
rect 18417 3111 18475 3117
rect 18417 3108 18429 3111
rect 18012 3080 18429 3108
rect 18012 3068 18018 3080
rect 18417 3077 18429 3080
rect 18463 3077 18475 3111
rect 18417 3071 18475 3077
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3040 17463 3043
rect 17862 3040 17868 3052
rect 17451 3012 17868 3040
rect 17451 3009 17463 3012
rect 17405 3003 17463 3009
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 20036 3012 20085 3040
rect 20036 3000 20042 3012
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 16132 2944 17356 2972
rect 17957 2975 18015 2981
rect 17957 2941 17969 2975
rect 18003 2972 18015 2975
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18003 2944 18521 2972
rect 18003 2941 18015 2944
rect 17957 2935 18015 2941
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 18690 2932 18696 2984
rect 18748 2932 18754 2984
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18840 2944 19073 2972
rect 18840 2932 18846 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 15948 2876 16896 2904
rect 14369 2867 14427 2873
rect 16298 2836 16304 2848
rect 14292 2808 16304 2836
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 16868 2836 16896 2876
rect 18874 2836 18880 2848
rect 16868 2808 18880 2836
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 20824 2836 20852 3136
rect 25869 3111 25927 3117
rect 22066 3080 22784 3108
rect 21450 3000 21456 3052
rect 21508 3040 21514 3052
rect 22066 3040 22094 3080
rect 22756 3049 22784 3080
rect 25869 3077 25881 3111
rect 25915 3108 25927 3111
rect 26252 3108 26280 3136
rect 27908 3108 27936 3136
rect 25915 3080 26280 3108
rect 26528 3080 27936 3108
rect 25915 3077 25927 3080
rect 25869 3071 25927 3077
rect 21508 3012 22094 3040
rect 22741 3043 22799 3049
rect 21508 3000 21514 3012
rect 22741 3009 22753 3043
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 23124 3012 24164 3040
rect 21082 2932 21088 2984
rect 21140 2932 21146 2984
rect 21637 2975 21695 2981
rect 21637 2941 21649 2975
rect 21683 2972 21695 2975
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 21683 2944 22293 2972
rect 21683 2941 21695 2944
rect 21637 2935 21695 2941
rect 22281 2941 22293 2944
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 23124 2972 23152 3012
rect 22511 2944 23152 2972
rect 23201 2975 23259 2981
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 23201 2941 23213 2975
rect 23247 2941 23259 2975
rect 23201 2935 23259 2941
rect 21100 2904 21128 2932
rect 22186 2904 22192 2916
rect 21100 2876 22192 2904
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 22480 2836 22508 2935
rect 23216 2904 23244 2935
rect 24026 2932 24032 2984
rect 24084 2932 24090 2984
rect 24136 2972 24164 3012
rect 25038 3000 25044 3052
rect 25096 3000 25102 3052
rect 26528 3049 26556 3080
rect 28994 3068 29000 3120
rect 29052 3108 29058 3120
rect 29150 3111 29208 3117
rect 29150 3108 29162 3111
rect 29052 3080 29162 3108
rect 29052 3068 29058 3080
rect 29150 3077 29162 3080
rect 29196 3077 29208 3111
rect 29150 3071 29208 3077
rect 26513 3043 26571 3049
rect 26513 3009 26525 3043
rect 26559 3009 26571 3043
rect 26513 3003 26571 3009
rect 27341 3043 27399 3049
rect 27341 3009 27353 3043
rect 27387 3040 27399 3043
rect 28074 3040 28080 3052
rect 27387 3012 28080 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 28442 3000 28448 3052
rect 28500 3040 28506 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28500 3012 28917 3040
rect 28500 3000 28506 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 30837 3043 30895 3049
rect 30837 3009 30849 3043
rect 30883 3040 30895 3043
rect 31205 3043 31263 3049
rect 31205 3040 31217 3043
rect 30883 3012 31217 3040
rect 30883 3009 30895 3012
rect 30837 3003 30895 3009
rect 31205 3009 31217 3012
rect 31251 3009 31263 3043
rect 31205 3003 31263 3009
rect 26145 2975 26203 2981
rect 26145 2972 26157 2975
rect 24136 2944 26157 2972
rect 26145 2941 26157 2944
rect 26191 2972 26203 2975
rect 26694 2972 26700 2984
rect 26191 2944 26700 2972
rect 26191 2941 26203 2944
rect 26145 2935 26203 2941
rect 26694 2932 26700 2944
rect 26752 2932 26758 2984
rect 27062 2932 27068 2984
rect 27120 2972 27126 2984
rect 27617 2975 27675 2981
rect 27617 2972 27629 2975
rect 27120 2944 27629 2972
rect 27120 2932 27126 2944
rect 27617 2941 27629 2944
rect 27663 2941 27675 2975
rect 27617 2935 27675 2941
rect 30926 2932 30932 2984
rect 30984 2932 30990 2984
rect 24578 2904 24584 2916
rect 23216 2876 24584 2904
rect 24578 2864 24584 2876
rect 24636 2864 24642 2916
rect 30285 2907 30343 2913
rect 30285 2873 30297 2907
rect 30331 2904 30343 2907
rect 31588 2904 31616 3136
rect 32401 3111 32459 3117
rect 32401 3077 32413 3111
rect 32447 3108 32459 3111
rect 33244 3108 33272 3136
rect 32447 3080 33272 3108
rect 32447 3077 32459 3080
rect 32401 3071 32459 3077
rect 33410 3068 33416 3120
rect 33468 3068 33474 3120
rect 33594 3068 33600 3120
rect 33652 3108 33658 3120
rect 33873 3111 33931 3117
rect 33873 3108 33885 3111
rect 33652 3080 33885 3108
rect 33652 3068 33658 3080
rect 33873 3077 33885 3080
rect 33919 3077 33931 3111
rect 33873 3071 33931 3077
rect 34876 3111 34934 3117
rect 34876 3077 34888 3111
rect 34922 3108 34934 3111
rect 34974 3108 34980 3120
rect 34922 3080 34980 3108
rect 34922 3077 34934 3080
rect 34876 3071 34934 3077
rect 34974 3068 34980 3080
rect 35032 3068 35038 3120
rect 35342 3068 35348 3120
rect 35400 3108 35406 3120
rect 37090 3108 37096 3120
rect 35400 3080 37096 3108
rect 35400 3068 35406 3080
rect 37090 3068 37096 3080
rect 37148 3068 37154 3120
rect 37734 3068 37740 3120
rect 37792 3108 37798 3120
rect 41800 3108 41828 3139
rect 42150 3136 42156 3148
rect 42208 3136 42214 3188
rect 42794 3136 42800 3188
rect 42852 3176 42858 3188
rect 45373 3179 45431 3185
rect 45373 3176 45385 3179
rect 42852 3148 45385 3176
rect 42852 3136 42858 3148
rect 45373 3145 45385 3148
rect 45419 3145 45431 3179
rect 45373 3139 45431 3145
rect 47029 3179 47087 3185
rect 47029 3145 47041 3179
rect 47075 3176 47087 3179
rect 47210 3176 47216 3188
rect 47075 3148 47216 3176
rect 47075 3145 47087 3148
rect 47029 3139 47087 3145
rect 47210 3136 47216 3148
rect 47268 3136 47274 3188
rect 47397 3179 47455 3185
rect 47397 3145 47409 3179
rect 47443 3176 47455 3179
rect 48130 3176 48136 3188
rect 47443 3148 48136 3176
rect 47443 3145 47455 3148
rect 47397 3139 47455 3145
rect 48130 3136 48136 3148
rect 48188 3136 48194 3188
rect 49881 3179 49939 3185
rect 48240 3148 48728 3176
rect 37792 3080 40448 3108
rect 41800 3080 42656 3108
rect 37792 3068 37798 3080
rect 34609 3043 34667 3049
rect 34609 3009 34621 3043
rect 34655 3040 34667 3043
rect 34698 3040 34704 3052
rect 34655 3012 34704 3040
rect 34655 3009 34667 3012
rect 34609 3003 34667 3009
rect 34698 3000 34704 3012
rect 34756 3000 34762 3052
rect 36814 3000 36820 3052
rect 36872 3000 36878 3052
rect 38028 3049 38056 3080
rect 40420 3052 40448 3080
rect 38013 3043 38071 3049
rect 38013 3009 38025 3043
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 38280 3043 38338 3049
rect 38280 3009 38292 3043
rect 38326 3040 38338 3043
rect 38562 3040 38568 3052
rect 38326 3012 38568 3040
rect 38326 3009 38338 3012
rect 38280 3003 38338 3009
rect 38562 3000 38568 3012
rect 38620 3000 38626 3052
rect 40402 3000 40408 3052
rect 40460 3000 40466 3052
rect 40672 3043 40730 3049
rect 40672 3009 40684 3043
rect 40718 3040 40730 3043
rect 40954 3040 40960 3052
rect 40718 3012 40960 3040
rect 40718 3009 40730 3012
rect 40672 3003 40730 3009
rect 40954 3000 40960 3012
rect 41012 3000 41018 3052
rect 42628 3049 42656 3080
rect 44634 3068 44640 3120
rect 44692 3108 44698 3120
rect 44692 3080 46428 3108
rect 44692 3068 44698 3080
rect 41877 3043 41935 3049
rect 41877 3009 41889 3043
rect 41923 3009 41935 3043
rect 41877 3003 41935 3009
rect 42613 3043 42671 3049
rect 42613 3009 42625 3043
rect 42659 3040 42671 3043
rect 42978 3040 42984 3052
rect 42659 3012 42984 3040
rect 42659 3009 42671 3012
rect 42613 3003 42671 3009
rect 31849 2975 31907 2981
rect 31849 2941 31861 2975
rect 31895 2972 31907 2975
rect 31938 2972 31944 2984
rect 31895 2944 31944 2972
rect 31895 2941 31907 2944
rect 31849 2935 31907 2941
rect 31938 2932 31944 2944
rect 31996 2932 32002 2984
rect 32309 2975 32367 2981
rect 32309 2941 32321 2975
rect 32355 2972 32367 2975
rect 33042 2972 33048 2984
rect 32355 2944 33048 2972
rect 32355 2941 32367 2944
rect 32309 2935 32367 2941
rect 33042 2932 33048 2944
rect 33100 2972 33106 2984
rect 33137 2975 33195 2981
rect 33137 2972 33149 2975
rect 33100 2944 33149 2972
rect 33100 2932 33106 2944
rect 33137 2941 33149 2944
rect 33183 2941 33195 2975
rect 33137 2935 33195 2941
rect 34425 2975 34483 2981
rect 34425 2941 34437 2975
rect 34471 2941 34483 2975
rect 34425 2935 34483 2941
rect 30331 2876 31616 2904
rect 33781 2907 33839 2913
rect 30331 2873 30343 2876
rect 30285 2867 30343 2873
rect 33781 2873 33793 2907
rect 33827 2904 33839 2907
rect 34440 2904 34468 2935
rect 36354 2932 36360 2984
rect 36412 2972 36418 2984
rect 37829 2975 37887 2981
rect 37829 2972 37841 2975
rect 36412 2944 37841 2972
rect 36412 2932 36418 2944
rect 37829 2941 37841 2944
rect 37875 2941 37887 2975
rect 37829 2935 37887 2941
rect 39482 2932 39488 2984
rect 39540 2932 39546 2984
rect 41892 2972 41920 3003
rect 42978 3000 42984 3012
rect 43036 3000 43042 3052
rect 45094 3000 45100 3052
rect 45152 3000 45158 3052
rect 46290 3000 46296 3052
rect 46348 3000 46354 3052
rect 46400 3040 46428 3080
rect 47578 3068 47584 3120
rect 47636 3068 47642 3120
rect 47670 3068 47676 3120
rect 47728 3108 47734 3120
rect 48240 3108 48268 3148
rect 47728 3080 48268 3108
rect 47728 3068 47734 3080
rect 48314 3068 48320 3120
rect 48372 3068 48378 3120
rect 46400 3012 47072 3040
rect 42794 2972 42800 2984
rect 41892 2944 42800 2972
rect 42794 2932 42800 2944
rect 42852 2932 42858 2984
rect 42889 2975 42947 2981
rect 42889 2941 42901 2975
rect 42935 2941 42947 2975
rect 42889 2935 42947 2941
rect 33827 2876 34468 2904
rect 33827 2873 33839 2876
rect 33781 2867 33839 2873
rect 35986 2864 35992 2916
rect 36044 2904 36050 2916
rect 36814 2904 36820 2916
rect 36044 2876 36820 2904
rect 36044 2864 36050 2876
rect 36814 2864 36820 2876
rect 36872 2864 36878 2916
rect 41966 2864 41972 2916
rect 42024 2904 42030 2916
rect 42904 2904 42932 2935
rect 43622 2932 43628 2984
rect 43680 2972 43686 2984
rect 44085 2975 44143 2981
rect 44085 2972 44097 2975
rect 43680 2944 44097 2972
rect 43680 2932 43686 2944
rect 44085 2941 44097 2944
rect 44131 2941 44143 2975
rect 44085 2935 44143 2941
rect 45925 2975 45983 2981
rect 45925 2941 45937 2975
rect 45971 2941 45983 2975
rect 45925 2935 45983 2941
rect 42024 2876 42932 2904
rect 42024 2864 42030 2876
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 45940 2904 45968 2935
rect 46566 2932 46572 2984
rect 46624 2972 46630 2984
rect 46753 2975 46811 2981
rect 46753 2972 46765 2975
rect 46624 2944 46765 2972
rect 46624 2932 46630 2944
rect 46753 2941 46765 2944
rect 46799 2941 46811 2975
rect 46753 2935 46811 2941
rect 46937 2975 46995 2981
rect 46937 2941 46949 2975
rect 46983 2941 46995 2975
rect 47044 2972 47072 3012
rect 47210 3000 47216 3052
rect 47268 3040 47274 3052
rect 48332 3040 48360 3068
rect 48498 3040 48504 3052
rect 48556 3049 48562 3052
rect 47268 3012 48360 3040
rect 48466 3012 48504 3040
rect 47268 3000 47274 3012
rect 48498 3000 48504 3012
rect 48556 3003 48566 3049
rect 48700 3040 48728 3148
rect 49881 3145 49893 3179
rect 49927 3176 49939 3179
rect 50522 3176 50528 3188
rect 49927 3148 50528 3176
rect 49927 3145 49939 3148
rect 49881 3139 49939 3145
rect 50522 3136 50528 3148
rect 50580 3136 50586 3188
rect 50982 3136 50988 3188
rect 51040 3136 51046 3188
rect 51166 3136 51172 3188
rect 51224 3136 51230 3188
rect 51276 3148 55168 3176
rect 48768 3111 48826 3117
rect 48768 3077 48780 3111
rect 48814 3108 48826 3111
rect 50430 3108 50436 3120
rect 48814 3080 50436 3108
rect 48814 3077 48826 3080
rect 48768 3071 48826 3077
rect 50430 3068 50436 3080
rect 50488 3068 50494 3120
rect 51184 3108 51212 3136
rect 51092 3080 51212 3108
rect 51092 3049 51120 3080
rect 50525 3043 50583 3049
rect 50525 3040 50537 3043
rect 48700 3012 50537 3040
rect 50525 3009 50537 3012
rect 50571 3009 50583 3043
rect 50525 3003 50583 3009
rect 50801 3043 50859 3049
rect 50801 3009 50813 3043
rect 50847 3009 50859 3043
rect 50801 3003 50859 3009
rect 51084 3043 51142 3049
rect 51084 3009 51096 3043
rect 51130 3009 51142 3043
rect 51276 3040 51304 3148
rect 55140 3117 55168 3148
rect 55674 3136 55680 3188
rect 55732 3136 55738 3188
rect 56134 3136 56140 3188
rect 56192 3136 56198 3188
rect 56502 3136 56508 3188
rect 56560 3136 56566 3188
rect 56686 3136 56692 3188
rect 56744 3176 56750 3188
rect 57885 3179 57943 3185
rect 57885 3176 57897 3179
rect 56744 3148 57897 3176
rect 56744 3136 56750 3148
rect 57885 3145 57897 3148
rect 57931 3145 57943 3179
rect 57885 3139 57943 3145
rect 55125 3111 55183 3117
rect 52564 3080 53788 3108
rect 51084 3003 51142 3009
rect 51184 3012 51304 3040
rect 51344 3043 51402 3049
rect 48556 3000 48562 3003
rect 48133 2975 48191 2981
rect 48133 2972 48145 2975
rect 47044 2944 48145 2972
rect 46937 2935 46995 2941
rect 48133 2941 48145 2944
rect 48179 2941 48191 2975
rect 50816 2972 50844 3003
rect 51184 2972 51212 3012
rect 51344 3009 51356 3043
rect 51390 3040 51402 3043
rect 52362 3040 52368 3052
rect 51390 3012 52368 3040
rect 51390 3009 51402 3012
rect 51344 3003 51402 3009
rect 52362 3000 52368 3012
rect 52420 3000 52426 3052
rect 50816 2944 51212 2972
rect 48133 2935 48191 2941
rect 43036 2876 45968 2904
rect 46952 2904 46980 2935
rect 48314 2904 48320 2916
rect 46952 2876 48320 2904
rect 43036 2864 43042 2876
rect 48314 2864 48320 2876
rect 48372 2864 48378 2916
rect 51074 2904 51080 2916
rect 49436 2876 51080 2904
rect 20824 2808 22508 2836
rect 23750 2796 23756 2848
rect 23808 2796 23814 2848
rect 46477 2839 46535 2845
rect 46477 2805 46489 2839
rect 46523 2836 46535 2839
rect 47762 2836 47768 2848
rect 46523 2808 47768 2836
rect 46523 2805 46535 2808
rect 46477 2799 46535 2805
rect 47762 2796 47768 2808
rect 47820 2796 47826 2848
rect 47854 2796 47860 2848
rect 47912 2836 47918 2848
rect 49436 2836 49464 2876
rect 51074 2864 51080 2876
rect 51132 2864 51138 2916
rect 52564 2904 52592 3080
rect 53098 3000 53104 3052
rect 53156 3000 53162 3052
rect 53190 3000 53196 3052
rect 53248 3000 53254 3052
rect 53653 3043 53711 3049
rect 53653 3040 53665 3043
rect 53300 3012 53665 3040
rect 53006 2932 53012 2984
rect 53064 2932 53070 2984
rect 53300 2904 53328 3012
rect 53653 3009 53665 3012
rect 53699 3009 53711 3043
rect 53760 3040 53788 3080
rect 55125 3077 55137 3111
rect 55171 3077 55183 3111
rect 55692 3108 55720 3136
rect 55692 3080 55996 3108
rect 55125 3071 55183 3077
rect 55968 3049 55996 3080
rect 55953 3043 56011 3049
rect 53760 3012 55720 3040
rect 53653 3003 53711 3009
rect 53558 2932 53564 2984
rect 53616 2972 53622 2984
rect 55692 2981 55720 3012
rect 55953 3009 55965 3043
rect 55999 3009 56011 3043
rect 55953 3003 56011 3009
rect 56321 3043 56379 3049
rect 56321 3009 56333 3043
rect 56367 3040 56379 3043
rect 56520 3040 56548 3136
rect 56588 3111 56646 3117
rect 56588 3077 56600 3111
rect 56634 3108 56646 3111
rect 56778 3108 56784 3120
rect 56634 3080 56784 3108
rect 56634 3077 56646 3080
rect 56588 3071 56646 3077
rect 56778 3068 56784 3080
rect 56836 3068 56842 3120
rect 56367 3012 56548 3040
rect 56367 3009 56379 3012
rect 56321 3003 56379 3009
rect 54113 2975 54171 2981
rect 54113 2972 54125 2975
rect 53616 2944 54125 2972
rect 53616 2932 53622 2944
rect 54113 2941 54125 2944
rect 54159 2941 54171 2975
rect 54113 2935 54171 2941
rect 55677 2975 55735 2981
rect 55677 2941 55689 2975
rect 55723 2941 55735 2975
rect 55677 2935 55735 2941
rect 58250 2932 58256 2984
rect 58308 2932 58314 2984
rect 58437 2975 58495 2981
rect 58437 2941 58449 2975
rect 58483 2941 58495 2975
rect 58437 2935 58495 2941
rect 52012 2876 52592 2904
rect 52840 2876 53328 2904
rect 47912 2808 49464 2836
rect 47912 2796 47918 2808
rect 49970 2796 49976 2848
rect 50028 2796 50034 2848
rect 51350 2796 51356 2848
rect 51408 2836 51414 2848
rect 52012 2836 52040 2876
rect 52840 2848 52868 2876
rect 53742 2864 53748 2916
rect 53800 2864 53806 2916
rect 54386 2864 54392 2916
rect 54444 2904 54450 2916
rect 57701 2907 57759 2913
rect 54444 2876 56272 2904
rect 54444 2864 54450 2876
rect 51408 2808 52040 2836
rect 52457 2839 52515 2845
rect 51408 2796 51414 2808
rect 52457 2805 52469 2839
rect 52503 2836 52515 2839
rect 52822 2836 52828 2848
rect 52503 2808 52828 2836
rect 52503 2805 52515 2808
rect 52457 2799 52515 2805
rect 52822 2796 52828 2808
rect 52880 2796 52886 2848
rect 53561 2839 53619 2845
rect 53561 2805 53573 2839
rect 53607 2836 53619 2839
rect 53760 2836 53788 2864
rect 53607 2808 53788 2836
rect 56244 2836 56272 2876
rect 57701 2873 57713 2907
rect 57747 2904 57759 2907
rect 58268 2904 58296 2932
rect 57747 2876 58296 2904
rect 57747 2873 57759 2876
rect 57701 2867 57759 2873
rect 58452 2836 58480 2935
rect 56244 2808 58480 2836
rect 53607 2805 53619 2808
rect 53561 2799 53619 2805
rect 1104 2746 58880 2768
rect 1104 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 22616 2746
rect 22668 2694 22680 2746
rect 22732 2694 22744 2746
rect 22796 2694 22808 2746
rect 22860 2694 22872 2746
rect 22924 2694 37060 2746
rect 37112 2694 37124 2746
rect 37176 2694 37188 2746
rect 37240 2694 37252 2746
rect 37304 2694 37316 2746
rect 37368 2694 51504 2746
rect 51556 2694 51568 2746
rect 51620 2694 51632 2746
rect 51684 2694 51696 2746
rect 51748 2694 51760 2746
rect 51812 2694 58880 2746
rect 1104 2672 58880 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2682 2632 2688 2644
rect 2179 2604 2688 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 4430 2632 4436 2644
rect 2915 2604 4436 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5258 2592 5264 2644
rect 5316 2592 5322 2644
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 9766 2632 9772 2644
rect 6227 2604 9772 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 11790 2632 11796 2644
rect 9907 2604 11796 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 16942 2632 16948 2644
rect 12483 2604 16948 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 18874 2592 18880 2644
rect 18932 2592 18938 2644
rect 20165 2635 20223 2641
rect 20165 2601 20177 2635
rect 20211 2632 20223 2635
rect 21450 2632 21456 2644
rect 20211 2604 21456 2632
rect 20211 2601 20223 2604
rect 20165 2595 20223 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 22097 2635 22155 2641
rect 22097 2601 22109 2635
rect 22143 2632 22155 2635
rect 22370 2632 22376 2644
rect 22143 2604 22376 2632
rect 22143 2601 22155 2604
rect 22097 2595 22155 2601
rect 22370 2592 22376 2604
rect 22428 2592 22434 2644
rect 24121 2635 24179 2641
rect 24121 2601 24133 2635
rect 24167 2632 24179 2635
rect 25038 2632 25044 2644
rect 24167 2604 25044 2632
rect 24167 2601 24179 2604
rect 24121 2595 24179 2601
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 25317 2635 25375 2641
rect 25317 2601 25329 2635
rect 25363 2632 25375 2635
rect 27154 2632 27160 2644
rect 25363 2604 27160 2632
rect 25363 2601 25375 2604
rect 25317 2595 25375 2601
rect 27154 2592 27160 2604
rect 27212 2592 27218 2644
rect 27893 2635 27951 2641
rect 27893 2601 27905 2635
rect 27939 2632 27951 2635
rect 29086 2632 29092 2644
rect 27939 2604 29092 2632
rect 27939 2601 27951 2604
rect 27893 2595 27951 2601
rect 29086 2592 29092 2604
rect 29144 2592 29150 2644
rect 30377 2635 30435 2641
rect 30377 2601 30389 2635
rect 30423 2632 30435 2635
rect 31662 2632 31668 2644
rect 30423 2604 31668 2632
rect 30423 2601 30435 2604
rect 30377 2595 30435 2601
rect 31662 2592 31668 2604
rect 31720 2592 31726 2644
rect 34054 2592 34060 2644
rect 34112 2632 34118 2644
rect 34241 2635 34299 2641
rect 34241 2632 34253 2635
rect 34112 2604 34253 2632
rect 34112 2592 34118 2604
rect 34241 2601 34253 2604
rect 34287 2601 34299 2635
rect 34241 2595 34299 2601
rect 36170 2592 36176 2644
rect 36228 2592 36234 2644
rect 39114 2592 39120 2644
rect 39172 2632 39178 2644
rect 39393 2635 39451 2641
rect 39393 2632 39405 2635
rect 39172 2604 39405 2632
rect 39172 2592 39178 2604
rect 39393 2601 39405 2604
rect 39439 2601 39451 2635
rect 39393 2595 39451 2601
rect 40954 2592 40960 2644
rect 41012 2632 41018 2644
rect 41325 2635 41383 2641
rect 41325 2632 41337 2635
rect 41012 2604 41337 2632
rect 41012 2592 41018 2604
rect 41325 2601 41337 2604
rect 41371 2601 41383 2635
rect 41325 2595 41383 2601
rect 42794 2592 42800 2644
rect 42852 2632 42858 2644
rect 43901 2635 43959 2641
rect 43901 2632 43913 2635
rect 42852 2604 43913 2632
rect 42852 2592 42858 2604
rect 43901 2601 43913 2604
rect 43947 2601 43959 2635
rect 43901 2595 43959 2601
rect 45189 2635 45247 2641
rect 45189 2601 45201 2635
rect 45235 2632 45247 2635
rect 45278 2632 45284 2644
rect 45235 2604 45284 2632
rect 45235 2601 45247 2604
rect 45189 2595 45247 2601
rect 45278 2592 45284 2604
rect 45336 2592 45342 2644
rect 47026 2592 47032 2644
rect 47084 2592 47090 2644
rect 47394 2592 47400 2644
rect 47452 2592 47458 2644
rect 48314 2592 48320 2644
rect 48372 2632 48378 2644
rect 49053 2635 49111 2641
rect 49053 2632 49065 2635
rect 48372 2604 49065 2632
rect 48372 2592 48378 2604
rect 49053 2601 49065 2604
rect 49099 2601 49111 2635
rect 49053 2595 49111 2601
rect 49970 2592 49976 2644
rect 50028 2592 50034 2644
rect 51166 2592 51172 2644
rect 51224 2632 51230 2644
rect 51629 2635 51687 2641
rect 51629 2632 51641 2635
rect 51224 2604 51641 2632
rect 51224 2592 51230 2604
rect 51629 2601 51641 2604
rect 51675 2601 51687 2635
rect 51629 2595 51687 2601
rect 54202 2592 54208 2644
rect 54260 2592 54266 2644
rect 56873 2635 56931 2641
rect 56873 2601 56885 2635
rect 56919 2632 56931 2635
rect 57330 2632 57336 2644
rect 56919 2604 57336 2632
rect 56919 2601 56931 2604
rect 56873 2595 56931 2601
rect 57330 2592 57336 2604
rect 57388 2592 57394 2644
rect 57790 2592 57796 2644
rect 57848 2592 57854 2644
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 3068 2536 6377 2564
rect 3068 2505 3096 2536
rect 6365 2533 6377 2536
rect 6411 2533 6423 2567
rect 6365 2527 6423 2533
rect 16574 2524 16580 2576
rect 16632 2564 16638 2576
rect 16761 2567 16819 2573
rect 16761 2564 16773 2567
rect 16632 2536 16773 2564
rect 16632 2524 16638 2536
rect 16761 2533 16773 2536
rect 16807 2533 16819 2567
rect 16761 2527 16819 2533
rect 40494 2524 40500 2576
rect 40552 2564 40558 2576
rect 49988 2564 50016 2592
rect 57808 2564 57836 2592
rect 40552 2536 42932 2564
rect 40552 2524 40558 2536
rect 3053 2499 3111 2505
rect 3053 2465 3065 2499
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3384 2468 4261 2496
rect 3384 2456 3390 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 6454 2456 6460 2508
rect 6512 2496 6518 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6512 2468 6837 2496
rect 6512 2456 6518 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 6914 2456 6920 2508
rect 6972 2456 6978 2508
rect 12986 2496 12992 2508
rect 9324 2468 12992 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1596 2360 1624 2391
rect 2314 2388 2320 2440
rect 2372 2388 2378 2440
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3200 2400 3801 2428
rect 3200 2388 3206 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 4948 2400 5457 2428
rect 4948 2388 4954 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5675 2400 6914 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 3878 2360 3884 2372
rect 1596 2332 3884 2360
rect 3878 2320 3884 2332
rect 3936 2320 3942 2372
rect 5902 2320 5908 2372
rect 5960 2320 5966 2372
rect 6730 2320 6736 2372
rect 6788 2320 6794 2372
rect 3605 2295 3663 2301
rect 3605 2261 3617 2295
rect 3651 2292 3663 2295
rect 5920 2292 5948 2320
rect 3651 2264 5948 2292
rect 6886 2292 6914 2400
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 9324 2437 9352 2468
rect 12986 2456 12992 2468
rect 13044 2456 13050 2508
rect 13449 2499 13507 2505
rect 13449 2465 13461 2499
rect 13495 2496 13507 2499
rect 13814 2496 13820 2508
rect 13495 2468 13820 2496
rect 13495 2465 13507 2468
rect 13449 2459 13507 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15344 2468 15577 2496
rect 15344 2456 15350 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 16724 2468 17264 2496
rect 16724 2456 16730 2468
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7248 2400 7389 2428
rect 7248 2388 7254 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2428 13967 2431
rect 13998 2428 14004 2440
rect 13955 2400 14004 2428
rect 13955 2397 13967 2400
rect 13909 2391 13967 2397
rect 8573 2363 8631 2369
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 8846 2360 8852 2372
rect 8619 2332 8852 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 10410 2320 10416 2372
rect 10468 2320 10474 2372
rect 11900 2360 11928 2391
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 14458 2388 14464 2440
rect 14516 2388 14522 2440
rect 15194 2388 15200 2440
rect 15252 2388 15258 2440
rect 15378 2388 15384 2440
rect 15436 2428 15442 2440
rect 17236 2437 17264 2468
rect 17310 2456 17316 2508
rect 17368 2496 17374 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17368 2468 17693 2496
rect 17368 2456 17374 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22649 2499 22707 2505
rect 22649 2496 22661 2499
rect 22152 2468 22661 2496
rect 22152 2456 22158 2468
rect 22649 2465 22661 2468
rect 22695 2465 22707 2499
rect 22649 2459 22707 2465
rect 28718 2456 28724 2508
rect 28776 2456 28782 2508
rect 34054 2456 34060 2508
rect 34112 2496 34118 2508
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 34112 2468 35173 2496
rect 34112 2456 34118 2468
rect 35161 2465 35173 2468
rect 35207 2465 35219 2499
rect 35161 2459 35219 2465
rect 37182 2456 37188 2508
rect 37240 2496 37246 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 37240 2468 37749 2496
rect 37240 2456 37246 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 39022 2456 39028 2508
rect 39080 2496 39086 2508
rect 40313 2499 40371 2505
rect 40313 2496 40325 2499
rect 39080 2468 40325 2496
rect 39080 2456 39086 2468
rect 40313 2465 40325 2468
rect 40359 2465 40371 2499
rect 40313 2459 40371 2465
rect 41969 2499 42027 2505
rect 41969 2465 41981 2499
rect 42015 2496 42027 2499
rect 42058 2496 42064 2508
rect 42015 2468 42064 2496
rect 42015 2465 42027 2468
rect 41969 2459 42027 2465
rect 42058 2456 42064 2468
rect 42116 2456 42122 2508
rect 42904 2505 42932 2536
rect 46860 2536 50016 2564
rect 56704 2536 57836 2564
rect 42889 2499 42947 2505
rect 42889 2465 42901 2499
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 15436 2400 16957 2428
rect 15436 2388 15442 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 19061 2431 19119 2437
rect 19061 2397 19073 2431
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 19659 2400 20944 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 14274 2360 14280 2372
rect 11900 2332 14280 2360
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 15013 2363 15071 2369
rect 15013 2329 15025 2363
rect 15059 2360 15071 2363
rect 19076 2360 19104 2391
rect 15059 2332 19104 2360
rect 15059 2329 15071 2332
rect 15013 2323 15071 2329
rect 20438 2320 20444 2372
rect 20496 2320 20502 2372
rect 20916 2360 20944 2400
rect 20990 2388 20996 2440
rect 21048 2428 21054 2440
rect 21453 2431 21511 2437
rect 21453 2428 21465 2431
rect 21048 2400 21465 2428
rect 21048 2388 21054 2400
rect 21453 2397 21465 2400
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 21634 2388 21640 2440
rect 21692 2428 21698 2440
rect 21913 2431 21971 2437
rect 21913 2428 21925 2431
rect 21692 2400 21925 2428
rect 21692 2388 21698 2400
rect 21913 2397 21925 2400
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 22186 2388 22192 2440
rect 22244 2388 22250 2440
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23808 2400 23949 2428
rect 23808 2388 23814 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 26050 2428 26056 2440
rect 24811 2400 26056 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 26050 2388 26056 2400
rect 26108 2388 26114 2440
rect 26602 2388 26608 2440
rect 26660 2388 26666 2440
rect 27341 2431 27399 2437
rect 27341 2397 27353 2431
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 22646 2360 22652 2372
rect 20916 2332 22652 2360
rect 22646 2320 22652 2332
rect 22704 2320 22710 2372
rect 25590 2320 25596 2372
rect 25648 2320 25654 2372
rect 27356 2360 27384 2391
rect 28166 2388 28172 2440
rect 28224 2388 28230 2440
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2428 29883 2431
rect 31202 2428 31208 2440
rect 29871 2400 31208 2428
rect 29871 2397 29883 2400
rect 29825 2391 29883 2397
rect 31202 2388 31208 2400
rect 31260 2388 31266 2440
rect 31849 2431 31907 2437
rect 31849 2397 31861 2431
rect 31895 2428 31907 2431
rect 31938 2428 31944 2440
rect 31895 2400 31944 2428
rect 31895 2397 31907 2400
rect 31849 2391 31907 2397
rect 31938 2388 31944 2400
rect 31996 2388 32002 2440
rect 33318 2388 33324 2440
rect 33376 2388 33382 2440
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 29362 2360 29368 2372
rect 27356 2332 29368 2360
rect 29362 2320 29368 2332
rect 29420 2320 29426 2372
rect 30466 2320 30472 2372
rect 30524 2360 30530 2372
rect 30653 2363 30711 2369
rect 30653 2360 30665 2363
rect 30524 2332 30665 2360
rect 30524 2320 30530 2332
rect 30653 2329 30665 2332
rect 30699 2329 30711 2363
rect 30653 2323 30711 2329
rect 32030 2320 32036 2372
rect 32088 2360 32094 2372
rect 32309 2363 32367 2369
rect 32309 2360 32321 2363
rect 32088 2332 32321 2360
rect 32088 2320 32094 2332
rect 32309 2329 32321 2332
rect 32355 2329 32367 2363
rect 32309 2323 32367 2329
rect 32950 2320 32956 2372
rect 33008 2360 33014 2372
rect 33612 2360 33640 2391
rect 34790 2388 34796 2440
rect 34848 2388 34854 2440
rect 34882 2388 34888 2440
rect 34940 2428 34946 2440
rect 36725 2431 36783 2437
rect 36725 2428 36737 2431
rect 34940 2400 36737 2428
rect 34940 2388 34946 2400
rect 36725 2397 36737 2400
rect 36771 2397 36783 2431
rect 36725 2391 36783 2397
rect 36814 2388 36820 2440
rect 36872 2428 36878 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36872 2400 37289 2428
rect 36872 2388 36878 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37918 2388 37924 2440
rect 37976 2428 37982 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 37976 2400 38761 2428
rect 37976 2388 37982 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 39666 2388 39672 2440
rect 39724 2428 39730 2440
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 39724 2400 39865 2428
rect 39724 2388 39730 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39853 2391 39911 2397
rect 40218 2388 40224 2440
rect 40276 2428 40282 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 40276 2400 42441 2428
rect 40276 2388 40282 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 44174 2388 44180 2440
rect 44232 2428 44238 2440
rect 44453 2431 44511 2437
rect 44453 2428 44465 2431
rect 44232 2400 44465 2428
rect 44232 2388 44238 2400
rect 44453 2397 44465 2400
rect 44499 2397 44511 2431
rect 44453 2391 44511 2397
rect 45005 2431 45063 2437
rect 45005 2397 45017 2431
rect 45051 2397 45063 2431
rect 45005 2391 45063 2397
rect 33008 2332 33640 2360
rect 33008 2320 33014 2332
rect 9674 2292 9680 2304
rect 6886 2264 9680 2292
rect 3651 2261 3663 2264
rect 3605 2255 3663 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 45020 2292 45048 2391
rect 46658 2388 46664 2440
rect 46716 2388 46722 2440
rect 46860 2437 46888 2536
rect 48682 2456 48688 2508
rect 48740 2496 48746 2508
rect 50617 2499 50675 2505
rect 50617 2496 50629 2499
rect 48740 2468 50629 2496
rect 48740 2456 48746 2468
rect 50617 2465 50629 2468
rect 50663 2465 50675 2499
rect 50617 2459 50675 2465
rect 46845 2431 46903 2437
rect 46845 2397 46857 2431
rect 46891 2397 46903 2431
rect 46845 2391 46903 2397
rect 48774 2388 48780 2440
rect 48832 2428 48838 2440
rect 49605 2431 49663 2437
rect 49605 2428 49617 2431
rect 48832 2400 49617 2428
rect 48832 2388 48838 2400
rect 49605 2397 49617 2400
rect 49651 2397 49663 2431
rect 49605 2391 49663 2397
rect 50154 2388 50160 2440
rect 50212 2388 50218 2440
rect 51074 2388 51080 2440
rect 51132 2428 51138 2440
rect 52181 2431 52239 2437
rect 52181 2428 52193 2431
rect 51132 2400 52193 2428
rect 51132 2388 51138 2400
rect 52181 2397 52193 2400
rect 52227 2397 52239 2431
rect 52181 2391 52239 2397
rect 52638 2388 52644 2440
rect 52696 2428 52702 2440
rect 53929 2431 53987 2437
rect 53929 2428 53941 2431
rect 52696 2400 53941 2428
rect 52696 2388 52702 2400
rect 53929 2397 53941 2400
rect 53975 2397 53987 2431
rect 53929 2391 53987 2397
rect 54754 2388 54760 2440
rect 54812 2388 54818 2440
rect 56704 2437 56732 2536
rect 57422 2456 57428 2508
rect 57480 2456 57486 2508
rect 57606 2456 57612 2508
rect 57664 2456 57670 2508
rect 58434 2456 58440 2508
rect 58492 2456 58498 2508
rect 56689 2431 56747 2437
rect 56689 2397 56701 2431
rect 56735 2397 56747 2431
rect 56689 2391 56747 2397
rect 57238 2388 57244 2440
rect 57296 2388 57302 2440
rect 57333 2431 57391 2437
rect 57333 2397 57345 2431
rect 57379 2428 57391 2431
rect 57624 2428 57652 2456
rect 57379 2400 57652 2428
rect 57379 2397 57391 2400
rect 57333 2391 57391 2397
rect 45278 2320 45284 2372
rect 45336 2360 45342 2372
rect 45557 2363 45615 2369
rect 45557 2360 45569 2363
rect 45336 2332 45569 2360
rect 45336 2320 45342 2332
rect 45557 2329 45569 2332
rect 45603 2329 45615 2363
rect 45557 2323 45615 2329
rect 46934 2320 46940 2372
rect 46992 2360 46998 2372
rect 47765 2363 47823 2369
rect 47765 2360 47777 2363
rect 46992 2332 47777 2360
rect 46992 2320 46998 2332
rect 47765 2329 47777 2332
rect 47811 2329 47823 2363
rect 47765 2323 47823 2329
rect 52086 2320 52092 2372
rect 52144 2360 52150 2372
rect 52917 2363 52975 2369
rect 52917 2360 52929 2363
rect 52144 2332 52929 2360
rect 52144 2320 52150 2332
rect 52917 2329 52929 2332
rect 52963 2329 52975 2363
rect 52917 2323 52975 2329
rect 53650 2320 53656 2372
rect 53708 2320 53714 2372
rect 55214 2320 55220 2372
rect 55272 2360 55278 2372
rect 55493 2363 55551 2369
rect 55493 2360 55505 2363
rect 55272 2332 55505 2360
rect 55272 2320 55278 2332
rect 55493 2329 55505 2332
rect 55539 2329 55551 2363
rect 55493 2323 55551 2329
rect 47578 2292 47584 2304
rect 45020 2264 47584 2292
rect 47578 2252 47584 2264
rect 47636 2252 47642 2304
rect 53668 2292 53696 2320
rect 57885 2295 57943 2301
rect 57885 2292 57897 2295
rect 53668 2264 57897 2292
rect 57885 2261 57897 2264
rect 57931 2261 57943 2295
rect 57885 2255 57943 2261
rect 1104 2202 59040 2224
rect 1104 2150 15394 2202
rect 15446 2150 15458 2202
rect 15510 2150 15522 2202
rect 15574 2150 15586 2202
rect 15638 2150 15650 2202
rect 15702 2150 29838 2202
rect 29890 2150 29902 2202
rect 29954 2150 29966 2202
rect 30018 2150 30030 2202
rect 30082 2150 30094 2202
rect 30146 2150 44282 2202
rect 44334 2150 44346 2202
rect 44398 2150 44410 2202
rect 44462 2150 44474 2202
rect 44526 2150 44538 2202
rect 44590 2150 58726 2202
rect 58778 2150 58790 2202
rect 58842 2150 58854 2202
rect 58906 2150 58918 2202
rect 58970 2150 58982 2202
rect 59034 2150 59040 2202
rect 1104 2128 59040 2150
rect 2314 2048 2320 2100
rect 2372 2088 2378 2100
rect 6362 2088 6368 2100
rect 2372 2060 6368 2088
rect 2372 2048 2378 2060
rect 6362 2048 6368 2060
rect 6420 2048 6426 2100
rect 14458 2048 14464 2100
rect 14516 2088 14522 2100
rect 19610 2088 19616 2100
rect 14516 2060 19616 2088
rect 14516 2048 14522 2060
rect 19610 2048 19616 2060
rect 19668 2048 19674 2100
<< via1 >>
rect 8172 27718 8224 27770
rect 8236 27718 8288 27770
rect 8300 27718 8352 27770
rect 8364 27718 8416 27770
rect 8428 27718 8480 27770
rect 22616 27718 22668 27770
rect 22680 27718 22732 27770
rect 22744 27718 22796 27770
rect 22808 27718 22860 27770
rect 22872 27718 22924 27770
rect 37060 27718 37112 27770
rect 37124 27718 37176 27770
rect 37188 27718 37240 27770
rect 37252 27718 37304 27770
rect 37316 27718 37368 27770
rect 51504 27718 51556 27770
rect 51568 27718 51620 27770
rect 51632 27718 51684 27770
rect 51696 27718 51748 27770
rect 51760 27718 51812 27770
rect 15394 27174 15446 27226
rect 15458 27174 15510 27226
rect 15522 27174 15574 27226
rect 15586 27174 15638 27226
rect 15650 27174 15702 27226
rect 29838 27174 29890 27226
rect 29902 27174 29954 27226
rect 29966 27174 30018 27226
rect 30030 27174 30082 27226
rect 30094 27174 30146 27226
rect 44282 27174 44334 27226
rect 44346 27174 44398 27226
rect 44410 27174 44462 27226
rect 44474 27174 44526 27226
rect 44538 27174 44590 27226
rect 58726 27174 58778 27226
rect 58790 27174 58842 27226
rect 58854 27174 58906 27226
rect 58918 27174 58970 27226
rect 58982 27174 59034 27226
rect 8172 26630 8224 26682
rect 8236 26630 8288 26682
rect 8300 26630 8352 26682
rect 8364 26630 8416 26682
rect 8428 26630 8480 26682
rect 22616 26630 22668 26682
rect 22680 26630 22732 26682
rect 22744 26630 22796 26682
rect 22808 26630 22860 26682
rect 22872 26630 22924 26682
rect 37060 26630 37112 26682
rect 37124 26630 37176 26682
rect 37188 26630 37240 26682
rect 37252 26630 37304 26682
rect 37316 26630 37368 26682
rect 51504 26630 51556 26682
rect 51568 26630 51620 26682
rect 51632 26630 51684 26682
rect 51696 26630 51748 26682
rect 51760 26630 51812 26682
rect 15394 26086 15446 26138
rect 15458 26086 15510 26138
rect 15522 26086 15574 26138
rect 15586 26086 15638 26138
rect 15650 26086 15702 26138
rect 29838 26086 29890 26138
rect 29902 26086 29954 26138
rect 29966 26086 30018 26138
rect 30030 26086 30082 26138
rect 30094 26086 30146 26138
rect 44282 26086 44334 26138
rect 44346 26086 44398 26138
rect 44410 26086 44462 26138
rect 44474 26086 44526 26138
rect 44538 26086 44590 26138
rect 58726 26086 58778 26138
rect 58790 26086 58842 26138
rect 58854 26086 58906 26138
rect 58918 26086 58970 26138
rect 58982 26086 59034 26138
rect 8172 25542 8224 25594
rect 8236 25542 8288 25594
rect 8300 25542 8352 25594
rect 8364 25542 8416 25594
rect 8428 25542 8480 25594
rect 22616 25542 22668 25594
rect 22680 25542 22732 25594
rect 22744 25542 22796 25594
rect 22808 25542 22860 25594
rect 22872 25542 22924 25594
rect 37060 25542 37112 25594
rect 37124 25542 37176 25594
rect 37188 25542 37240 25594
rect 37252 25542 37304 25594
rect 37316 25542 37368 25594
rect 51504 25542 51556 25594
rect 51568 25542 51620 25594
rect 51632 25542 51684 25594
rect 51696 25542 51748 25594
rect 51760 25542 51812 25594
rect 15394 24998 15446 25050
rect 15458 24998 15510 25050
rect 15522 24998 15574 25050
rect 15586 24998 15638 25050
rect 15650 24998 15702 25050
rect 29838 24998 29890 25050
rect 29902 24998 29954 25050
rect 29966 24998 30018 25050
rect 30030 24998 30082 25050
rect 30094 24998 30146 25050
rect 44282 24998 44334 25050
rect 44346 24998 44398 25050
rect 44410 24998 44462 25050
rect 44474 24998 44526 25050
rect 44538 24998 44590 25050
rect 58726 24998 58778 25050
rect 58790 24998 58842 25050
rect 58854 24998 58906 25050
rect 58918 24998 58970 25050
rect 58982 24998 59034 25050
rect 8172 24454 8224 24506
rect 8236 24454 8288 24506
rect 8300 24454 8352 24506
rect 8364 24454 8416 24506
rect 8428 24454 8480 24506
rect 22616 24454 22668 24506
rect 22680 24454 22732 24506
rect 22744 24454 22796 24506
rect 22808 24454 22860 24506
rect 22872 24454 22924 24506
rect 37060 24454 37112 24506
rect 37124 24454 37176 24506
rect 37188 24454 37240 24506
rect 37252 24454 37304 24506
rect 37316 24454 37368 24506
rect 51504 24454 51556 24506
rect 51568 24454 51620 24506
rect 51632 24454 51684 24506
rect 51696 24454 51748 24506
rect 51760 24454 51812 24506
rect 15394 23910 15446 23962
rect 15458 23910 15510 23962
rect 15522 23910 15574 23962
rect 15586 23910 15638 23962
rect 15650 23910 15702 23962
rect 29838 23910 29890 23962
rect 29902 23910 29954 23962
rect 29966 23910 30018 23962
rect 30030 23910 30082 23962
rect 30094 23910 30146 23962
rect 44282 23910 44334 23962
rect 44346 23910 44398 23962
rect 44410 23910 44462 23962
rect 44474 23910 44526 23962
rect 44538 23910 44590 23962
rect 58726 23910 58778 23962
rect 58790 23910 58842 23962
rect 58854 23910 58906 23962
rect 58918 23910 58970 23962
rect 58982 23910 59034 23962
rect 15200 23647 15252 23656
rect 15200 23613 15209 23647
rect 15209 23613 15243 23647
rect 15243 23613 15252 23647
rect 15200 23604 15252 23613
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 18144 23604 18196 23656
rect 18236 23647 18288 23656
rect 18236 23613 18245 23647
rect 18245 23613 18279 23647
rect 18279 23613 18288 23647
rect 18236 23604 18288 23613
rect 47584 23647 47636 23656
rect 47584 23613 47593 23647
rect 47593 23613 47627 23647
rect 47627 23613 47636 23647
rect 47584 23604 47636 23613
rect 53288 23647 53340 23656
rect 53288 23613 53297 23647
rect 53297 23613 53331 23647
rect 53331 23613 53340 23647
rect 53288 23604 53340 23613
rect 54024 23647 54076 23656
rect 54024 23613 54033 23647
rect 54033 23613 54067 23647
rect 54067 23613 54076 23647
rect 54024 23604 54076 23613
rect 14556 23511 14608 23520
rect 14556 23477 14565 23511
rect 14565 23477 14599 23511
rect 14599 23477 14608 23511
rect 14556 23468 14608 23477
rect 16212 23468 16264 23520
rect 17408 23511 17460 23520
rect 17408 23477 17417 23511
rect 17417 23477 17451 23511
rect 17451 23477 17460 23511
rect 17408 23468 17460 23477
rect 18880 23511 18932 23520
rect 18880 23477 18889 23511
rect 18889 23477 18923 23511
rect 18923 23477 18932 23511
rect 18880 23468 18932 23477
rect 46848 23511 46900 23520
rect 46848 23477 46857 23511
rect 46857 23477 46891 23511
rect 46891 23477 46900 23511
rect 46848 23468 46900 23477
rect 48136 23468 48188 23520
rect 48228 23511 48280 23520
rect 48228 23477 48237 23511
rect 48237 23477 48271 23511
rect 48271 23477 48280 23511
rect 48228 23468 48280 23477
rect 49332 23468 49384 23520
rect 54484 23536 54536 23588
rect 52736 23511 52788 23520
rect 52736 23477 52745 23511
rect 52745 23477 52779 23511
rect 52779 23477 52788 23511
rect 52736 23468 52788 23477
rect 53472 23511 53524 23520
rect 53472 23477 53481 23511
rect 53481 23477 53515 23511
rect 53515 23477 53524 23511
rect 53472 23468 53524 23477
rect 8172 23366 8224 23418
rect 8236 23366 8288 23418
rect 8300 23366 8352 23418
rect 8364 23366 8416 23418
rect 8428 23366 8480 23418
rect 22616 23366 22668 23418
rect 22680 23366 22732 23418
rect 22744 23366 22796 23418
rect 22808 23366 22860 23418
rect 22872 23366 22924 23418
rect 37060 23366 37112 23418
rect 37124 23366 37176 23418
rect 37188 23366 37240 23418
rect 37252 23366 37304 23418
rect 37316 23366 37368 23418
rect 51504 23366 51556 23418
rect 51568 23366 51620 23418
rect 51632 23366 51684 23418
rect 51696 23366 51748 23418
rect 51760 23366 51812 23418
rect 18236 23264 18288 23316
rect 42524 23264 42576 23316
rect 46848 23264 46900 23316
rect 15108 23128 15160 23180
rect 20444 23196 20496 23248
rect 52552 23264 52604 23316
rect 54024 23264 54076 23316
rect 48596 23196 48648 23248
rect 48136 23128 48188 23180
rect 6644 23103 6696 23112
rect 6644 23069 6653 23103
rect 6653 23069 6687 23103
rect 6687 23069 6696 23103
rect 6644 23060 6696 23069
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 14372 23035 14424 23044
rect 14372 23001 14406 23035
rect 14406 23001 14424 23035
rect 14372 22992 14424 23001
rect 17408 23060 17460 23112
rect 17960 23060 18012 23112
rect 20352 23103 20404 23112
rect 20352 23069 20361 23103
rect 20361 23069 20395 23103
rect 20395 23069 20404 23103
rect 20352 23060 20404 23069
rect 22284 23060 22336 23112
rect 23572 23103 23624 23112
rect 23572 23069 23581 23103
rect 23581 23069 23615 23103
rect 23615 23069 23624 23103
rect 23572 23060 23624 23069
rect 34060 23103 34112 23112
rect 34060 23069 34069 23103
rect 34069 23069 34103 23103
rect 34103 23069 34112 23103
rect 34060 23060 34112 23069
rect 36452 23103 36504 23112
rect 36452 23069 36461 23103
rect 36461 23069 36495 23103
rect 36495 23069 36504 23103
rect 36452 23060 36504 23069
rect 40408 23103 40460 23112
rect 40408 23069 40417 23103
rect 40417 23069 40451 23103
rect 40451 23069 40460 23103
rect 40408 23060 40460 23069
rect 45560 23103 45612 23112
rect 45560 23069 45569 23103
rect 45569 23069 45603 23103
rect 45603 23069 45612 23103
rect 45560 23060 45612 23069
rect 16764 22992 16816 23044
rect 35808 22992 35860 23044
rect 42708 22992 42760 23044
rect 6092 22967 6144 22976
rect 6092 22933 6101 22967
rect 6101 22933 6135 22967
rect 6135 22933 6144 22967
rect 6092 22924 6144 22933
rect 11060 22924 11112 22976
rect 16304 22924 16356 22976
rect 18052 22967 18104 22976
rect 18052 22933 18061 22967
rect 18061 22933 18095 22967
rect 18095 22933 18104 22967
rect 18052 22924 18104 22933
rect 19248 22924 19300 22976
rect 19800 22967 19852 22976
rect 19800 22933 19809 22967
rect 19809 22933 19843 22967
rect 19843 22933 19852 22967
rect 19800 22924 19852 22933
rect 22192 22967 22244 22976
rect 22192 22933 22201 22967
rect 22201 22933 22235 22967
rect 22235 22933 22244 22967
rect 22192 22924 22244 22933
rect 23204 22924 23256 22976
rect 33416 22967 33468 22976
rect 33416 22933 33425 22967
rect 33425 22933 33459 22967
rect 33459 22933 33468 22967
rect 33416 22924 33468 22933
rect 34244 22924 34296 22976
rect 35992 22924 36044 22976
rect 39856 22967 39908 22976
rect 39856 22933 39865 22967
rect 39865 22933 39899 22967
rect 39899 22933 39908 22967
rect 39856 22924 39908 22933
rect 45008 22967 45060 22976
rect 45008 22933 45017 22967
rect 45017 22933 45051 22967
rect 45051 22933 45060 22967
rect 45008 22924 45060 22933
rect 46204 22967 46256 22976
rect 46204 22933 46213 22967
rect 46213 22933 46247 22967
rect 46247 22933 46256 22967
rect 46204 22924 46256 22933
rect 48044 22924 48096 22976
rect 48228 22924 48280 22976
rect 49148 23060 49200 23112
rect 51540 23103 51592 23112
rect 51540 23069 51549 23103
rect 51549 23069 51583 23103
rect 51583 23069 51592 23103
rect 51540 23060 51592 23069
rect 51908 23103 51960 23112
rect 51908 23069 51917 23103
rect 51917 23069 51951 23103
rect 51951 23069 51960 23103
rect 51908 23060 51960 23069
rect 55220 23060 55272 23112
rect 56600 23103 56652 23112
rect 56600 23069 56609 23103
rect 56609 23069 56643 23103
rect 56643 23069 56652 23103
rect 56600 23060 56652 23069
rect 49056 22992 49108 23044
rect 52736 22992 52788 23044
rect 54208 22992 54260 23044
rect 49976 22924 50028 22976
rect 50068 22924 50120 22976
rect 50252 22924 50304 22976
rect 55128 22924 55180 22976
rect 56048 22967 56100 22976
rect 56048 22933 56057 22967
rect 56057 22933 56091 22967
rect 56091 22933 56100 22967
rect 56048 22924 56100 22933
rect 15394 22822 15446 22874
rect 15458 22822 15510 22874
rect 15522 22822 15574 22874
rect 15586 22822 15638 22874
rect 15650 22822 15702 22874
rect 29838 22822 29890 22874
rect 29902 22822 29954 22874
rect 29966 22822 30018 22874
rect 30030 22822 30082 22874
rect 30094 22822 30146 22874
rect 44282 22822 44334 22874
rect 44346 22822 44398 22874
rect 44410 22822 44462 22874
rect 44474 22822 44526 22874
rect 44538 22822 44590 22874
rect 58726 22822 58778 22874
rect 58790 22822 58842 22874
rect 58854 22822 58906 22874
rect 58918 22822 58970 22874
rect 58982 22822 59034 22874
rect 12164 22720 12216 22772
rect 14096 22652 14148 22704
rect 14556 22652 14608 22704
rect 15200 22720 15252 22772
rect 17132 22720 17184 22772
rect 17960 22720 18012 22772
rect 18144 22763 18196 22772
rect 18144 22729 18153 22763
rect 18153 22729 18187 22763
rect 18187 22729 18196 22763
rect 18144 22720 18196 22729
rect 18880 22720 18932 22772
rect 20352 22720 20404 22772
rect 22192 22720 22244 22772
rect 23572 22720 23624 22772
rect 36452 22720 36504 22772
rect 38660 22720 38712 22772
rect 39856 22720 39908 22772
rect 46204 22720 46256 22772
rect 47584 22720 47636 22772
rect 48136 22720 48188 22772
rect 13636 22627 13688 22636
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 15476 22627 15528 22636
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 16764 22652 16816 22704
rect 3700 22559 3752 22568
rect 3700 22525 3709 22559
rect 3709 22525 3743 22559
rect 3743 22525 3752 22559
rect 3700 22516 3752 22525
rect 4436 22559 4488 22568
rect 4436 22525 4445 22559
rect 4445 22525 4479 22559
rect 4479 22525 4488 22559
rect 4436 22516 4488 22525
rect 7104 22559 7156 22568
rect 7104 22525 7113 22559
rect 7113 22525 7147 22559
rect 7147 22525 7156 22559
rect 7104 22516 7156 22525
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 10048 22559 10100 22568
rect 10048 22525 10057 22559
rect 10057 22525 10091 22559
rect 10091 22525 10100 22559
rect 10048 22516 10100 22525
rect 10692 22559 10744 22568
rect 10692 22525 10701 22559
rect 10701 22525 10735 22559
rect 10735 22525 10744 22559
rect 10692 22516 10744 22525
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 15292 22516 15344 22568
rect 16120 22559 16172 22568
rect 16120 22525 16129 22559
rect 16129 22525 16163 22559
rect 16163 22525 16172 22559
rect 16120 22516 16172 22525
rect 4896 22491 4948 22500
rect 4896 22457 4905 22491
rect 4905 22457 4939 22491
rect 4939 22457 4948 22491
rect 4896 22448 4948 22457
rect 9956 22448 10008 22500
rect 3056 22423 3108 22432
rect 3056 22389 3065 22423
rect 3065 22389 3099 22423
rect 3099 22389 3108 22423
rect 3056 22380 3108 22389
rect 3884 22423 3936 22432
rect 3884 22389 3893 22423
rect 3893 22389 3927 22423
rect 3927 22389 3936 22423
rect 3884 22380 3936 22389
rect 5724 22380 5776 22432
rect 9220 22423 9272 22432
rect 9220 22389 9229 22423
rect 9229 22389 9263 22423
rect 9263 22389 9272 22423
rect 9220 22380 9272 22389
rect 10140 22380 10192 22432
rect 10876 22380 10928 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 12624 22423 12676 22432
rect 12624 22389 12633 22423
rect 12633 22389 12667 22423
rect 12667 22389 12676 22423
rect 12624 22380 12676 22389
rect 16580 22448 16632 22500
rect 17960 22584 18012 22636
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 19524 22559 19576 22568
rect 19524 22525 19533 22559
rect 19533 22525 19567 22559
rect 19567 22525 19576 22559
rect 19524 22516 19576 22525
rect 20628 22584 20680 22636
rect 32036 22652 32088 22704
rect 22376 22584 22428 22636
rect 33784 22584 33836 22636
rect 34336 22584 34388 22636
rect 20444 22559 20496 22568
rect 20444 22525 20453 22559
rect 20453 22525 20487 22559
rect 20487 22525 20496 22559
rect 20444 22516 20496 22525
rect 13820 22380 13872 22432
rect 20720 22559 20772 22568
rect 20720 22525 20729 22559
rect 20729 22525 20763 22559
rect 20763 22525 20772 22559
rect 20720 22516 20772 22525
rect 20812 22448 20864 22500
rect 23388 22516 23440 22568
rect 26332 22559 26384 22568
rect 26332 22525 26341 22559
rect 26341 22525 26375 22559
rect 26375 22525 26384 22559
rect 26332 22516 26384 22525
rect 27896 22516 27948 22568
rect 29184 22559 29236 22568
rect 29184 22525 29193 22559
rect 29193 22525 29227 22559
rect 29227 22525 29236 22559
rect 29184 22516 29236 22525
rect 31576 22559 31628 22568
rect 31576 22525 31585 22559
rect 31585 22525 31619 22559
rect 31619 22525 31628 22559
rect 31576 22516 31628 22525
rect 31668 22516 31720 22568
rect 24860 22448 24912 22500
rect 26792 22491 26844 22500
rect 26792 22457 26801 22491
rect 26801 22457 26835 22491
rect 26835 22457 26844 22491
rect 26792 22448 26844 22457
rect 23296 22423 23348 22432
rect 23296 22389 23305 22423
rect 23305 22389 23339 22423
rect 23339 22389 23348 22423
rect 23296 22380 23348 22389
rect 25596 22380 25648 22432
rect 27712 22380 27764 22432
rect 27804 22380 27856 22432
rect 28172 22380 28224 22432
rect 28632 22423 28684 22432
rect 28632 22389 28641 22423
rect 28641 22389 28675 22423
rect 28675 22389 28684 22423
rect 28632 22380 28684 22389
rect 30564 22423 30616 22432
rect 30564 22389 30573 22423
rect 30573 22389 30607 22423
rect 30607 22389 30616 22423
rect 30564 22380 30616 22389
rect 31024 22423 31076 22432
rect 31024 22389 31033 22423
rect 31033 22389 31067 22423
rect 31067 22389 31076 22423
rect 31024 22380 31076 22389
rect 33048 22380 33100 22432
rect 33324 22559 33376 22568
rect 33324 22525 33333 22559
rect 33333 22525 33367 22559
rect 33367 22525 33376 22559
rect 33324 22516 33376 22525
rect 33968 22516 34020 22568
rect 35256 22448 35308 22500
rect 37464 22516 37516 22568
rect 38568 22559 38620 22568
rect 38568 22525 38577 22559
rect 38577 22525 38611 22559
rect 38611 22525 38620 22559
rect 38568 22516 38620 22525
rect 40592 22559 40644 22568
rect 40592 22525 40601 22559
rect 40601 22525 40635 22559
rect 40635 22525 40644 22559
rect 40592 22516 40644 22525
rect 42064 22559 42116 22568
rect 42064 22525 42073 22559
rect 42073 22525 42107 22559
rect 42107 22525 42116 22559
rect 42064 22516 42116 22525
rect 42432 22559 42484 22568
rect 42432 22525 42441 22559
rect 42441 22525 42475 22559
rect 42475 22525 42484 22559
rect 42432 22516 42484 22525
rect 42708 22516 42760 22568
rect 43444 22516 43496 22568
rect 45008 22584 45060 22636
rect 49976 22652 50028 22704
rect 48872 22627 48924 22636
rect 48872 22593 48881 22627
rect 48881 22593 48915 22627
rect 48915 22593 48924 22627
rect 48872 22584 48924 22593
rect 49148 22627 49200 22636
rect 49148 22593 49157 22627
rect 49157 22593 49191 22627
rect 49191 22593 49200 22627
rect 49148 22584 49200 22593
rect 50068 22627 50120 22636
rect 50068 22593 50077 22627
rect 50077 22593 50111 22627
rect 50111 22593 50120 22627
rect 50068 22584 50120 22593
rect 51080 22652 51132 22704
rect 50252 22584 50304 22636
rect 51172 22584 51224 22636
rect 34244 22380 34296 22432
rect 34428 22380 34480 22432
rect 37556 22380 37608 22432
rect 38936 22380 38988 22432
rect 39212 22380 39264 22432
rect 40776 22423 40828 22432
rect 40776 22389 40785 22423
rect 40785 22389 40819 22423
rect 40819 22389 40828 22423
rect 40776 22380 40828 22389
rect 41512 22423 41564 22432
rect 41512 22389 41521 22423
rect 41521 22389 41555 22423
rect 41555 22389 41564 22423
rect 41512 22380 41564 22389
rect 43628 22380 43680 22432
rect 45284 22423 45336 22432
rect 45284 22389 45293 22423
rect 45293 22389 45327 22423
rect 45327 22389 45336 22423
rect 45284 22380 45336 22389
rect 48228 22516 48280 22568
rect 51540 22763 51592 22772
rect 51540 22729 51549 22763
rect 51549 22729 51583 22763
rect 51583 22729 51592 22763
rect 51540 22720 51592 22729
rect 53288 22720 53340 22772
rect 53472 22720 53524 22772
rect 56600 22763 56652 22772
rect 56600 22729 56609 22763
rect 56609 22729 56643 22763
rect 56643 22729 56652 22763
rect 56600 22720 56652 22729
rect 53288 22584 53340 22636
rect 56048 22652 56100 22704
rect 55220 22627 55272 22636
rect 55220 22593 55229 22627
rect 55229 22593 55263 22627
rect 55263 22593 55272 22627
rect 55220 22584 55272 22593
rect 53932 22559 53984 22568
rect 53932 22525 53941 22559
rect 53941 22525 53975 22559
rect 53975 22525 53984 22559
rect 53932 22516 53984 22525
rect 54024 22516 54076 22568
rect 49424 22491 49476 22500
rect 49424 22457 49433 22491
rect 49433 22457 49467 22491
rect 49467 22457 49476 22491
rect 49424 22448 49476 22457
rect 46664 22380 46716 22432
rect 47952 22423 48004 22432
rect 47952 22389 47961 22423
rect 47961 22389 47995 22423
rect 47995 22389 48004 22423
rect 47952 22380 48004 22389
rect 49608 22380 49660 22432
rect 53932 22380 53984 22432
rect 54116 22380 54168 22432
rect 54484 22559 54536 22568
rect 54484 22525 54493 22559
rect 54493 22525 54527 22559
rect 54527 22525 54536 22559
rect 54484 22516 54536 22525
rect 54576 22516 54628 22568
rect 55128 22559 55180 22568
rect 55128 22525 55137 22559
rect 55137 22525 55171 22559
rect 55171 22525 55180 22559
rect 55128 22516 55180 22525
rect 57244 22559 57296 22568
rect 57244 22525 57253 22559
rect 57253 22525 57287 22559
rect 57287 22525 57296 22559
rect 57244 22516 57296 22525
rect 8172 22278 8224 22330
rect 8236 22278 8288 22330
rect 8300 22278 8352 22330
rect 8364 22278 8416 22330
rect 8428 22278 8480 22330
rect 22616 22278 22668 22330
rect 22680 22278 22732 22330
rect 22744 22278 22796 22330
rect 22808 22278 22860 22330
rect 22872 22278 22924 22330
rect 37060 22278 37112 22330
rect 37124 22278 37176 22330
rect 37188 22278 37240 22330
rect 37252 22278 37304 22330
rect 37316 22278 37368 22330
rect 51504 22278 51556 22330
rect 51568 22278 51620 22330
rect 51632 22278 51684 22330
rect 51696 22278 51748 22330
rect 51760 22278 51812 22330
rect 3700 22176 3752 22228
rect 4896 22176 4948 22228
rect 7104 22219 7156 22228
rect 7104 22185 7113 22219
rect 7113 22185 7147 22219
rect 7147 22185 7156 22219
rect 7104 22176 7156 22185
rect 9772 22176 9824 22228
rect 11152 22176 11204 22228
rect 12072 22176 12124 22228
rect 13820 22219 13872 22228
rect 13820 22185 13829 22219
rect 13829 22185 13863 22219
rect 13863 22185 13872 22219
rect 13820 22176 13872 22185
rect 10140 22083 10192 22092
rect 10140 22049 10149 22083
rect 10149 22049 10183 22083
rect 10183 22049 10192 22083
rect 10140 22040 10192 22049
rect 12164 22083 12216 22092
rect 12164 22049 12173 22083
rect 12173 22049 12207 22083
rect 12207 22049 12216 22083
rect 12164 22040 12216 22049
rect 2964 22015 3016 22024
rect 2964 21981 2973 22015
rect 2973 21981 3007 22015
rect 3007 21981 3016 22015
rect 2964 21972 3016 21981
rect 4712 22015 4764 22024
rect 4712 21981 4721 22015
rect 4721 21981 4755 22015
rect 4755 21981 4764 22015
rect 4712 21972 4764 21981
rect 6460 21972 6512 22024
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 9036 21972 9088 22024
rect 16396 22176 16448 22228
rect 20720 22219 20772 22228
rect 20720 22185 20729 22219
rect 20729 22185 20763 22219
rect 20763 22185 20772 22219
rect 20720 22176 20772 22185
rect 23388 22219 23440 22228
rect 23388 22185 23397 22219
rect 23397 22185 23431 22219
rect 23431 22185 23440 22219
rect 23388 22176 23440 22185
rect 26332 22176 26384 22228
rect 26792 22176 26844 22228
rect 29184 22176 29236 22228
rect 31576 22176 31628 22228
rect 17132 22108 17184 22160
rect 4252 21879 4304 21888
rect 4252 21845 4261 21879
rect 4261 21845 4295 21879
rect 4295 21845 4304 21879
rect 4252 21836 4304 21845
rect 4620 21836 4672 21888
rect 4988 21836 5040 21888
rect 5264 21879 5316 21888
rect 5264 21845 5273 21879
rect 5273 21845 5307 21879
rect 5307 21845 5316 21879
rect 5264 21836 5316 21845
rect 6092 21904 6144 21956
rect 10140 21904 10192 21956
rect 11336 21904 11388 21956
rect 15108 21972 15160 22024
rect 15384 22040 15436 22092
rect 16304 22040 16356 22092
rect 16488 22083 16540 22092
rect 16488 22049 16497 22083
rect 16497 22049 16531 22083
rect 16531 22049 16540 22083
rect 16488 22040 16540 22049
rect 16672 22040 16724 22092
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 17684 22083 17736 22092
rect 17684 22049 17693 22083
rect 17693 22049 17727 22083
rect 17727 22049 17736 22083
rect 17684 22040 17736 22049
rect 17868 22108 17920 22160
rect 21732 22040 21784 22092
rect 22376 22083 22428 22092
rect 22376 22049 22385 22083
rect 22385 22049 22419 22083
rect 22419 22049 22428 22083
rect 22376 22040 22428 22049
rect 22560 22040 22612 22092
rect 30564 22108 30616 22160
rect 34336 22176 34388 22228
rect 35072 22176 35124 22228
rect 35808 22176 35860 22228
rect 24032 22083 24084 22092
rect 24032 22049 24041 22083
rect 24041 22049 24075 22083
rect 24075 22049 24084 22083
rect 24032 22040 24084 22049
rect 18880 21972 18932 22024
rect 19248 21972 19300 22024
rect 20812 21972 20864 22024
rect 22192 21972 22244 22024
rect 7196 21879 7248 21888
rect 7196 21845 7205 21879
rect 7205 21845 7239 21879
rect 7239 21845 7248 21879
rect 7196 21836 7248 21845
rect 9864 21836 9916 21888
rect 10876 21836 10928 21888
rect 10968 21836 11020 21888
rect 12440 21836 12492 21888
rect 17960 21904 18012 21956
rect 12808 21879 12860 21888
rect 12808 21845 12817 21879
rect 12817 21845 12851 21879
rect 12851 21845 12860 21879
rect 12808 21836 12860 21845
rect 14280 21836 14332 21888
rect 14556 21879 14608 21888
rect 14556 21845 14565 21879
rect 14565 21845 14599 21879
rect 14599 21845 14608 21879
rect 14556 21836 14608 21845
rect 14924 21879 14976 21888
rect 14924 21845 14933 21879
rect 14933 21845 14967 21879
rect 14967 21845 14976 21879
rect 14924 21836 14976 21845
rect 16856 21836 16908 21888
rect 19800 21904 19852 21956
rect 23204 21972 23256 22024
rect 24860 22040 24912 22092
rect 24952 22015 25004 22024
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 32036 22083 32088 22092
rect 26700 21972 26752 22024
rect 26976 21972 27028 22024
rect 29368 21972 29420 22024
rect 31576 21972 31628 22024
rect 32036 22049 32045 22083
rect 32045 22049 32079 22083
rect 32079 22049 32088 22083
rect 32036 22040 32088 22049
rect 35440 22083 35492 22092
rect 32588 21972 32640 22024
rect 35440 22049 35449 22083
rect 35449 22049 35483 22083
rect 35483 22049 35492 22083
rect 35440 22040 35492 22049
rect 39120 22108 39172 22160
rect 40592 22176 40644 22228
rect 42064 22176 42116 22228
rect 42616 22219 42668 22228
rect 42616 22185 42625 22219
rect 42625 22185 42659 22219
rect 42659 22185 42668 22219
rect 42616 22176 42668 22185
rect 41144 22108 41196 22160
rect 48872 22176 48924 22228
rect 49424 22176 49476 22228
rect 35256 22015 35308 22024
rect 35256 21981 35265 22015
rect 35265 21981 35299 22015
rect 35299 21981 35308 22015
rect 35256 21972 35308 21981
rect 37832 22040 37884 22092
rect 38660 22083 38712 22092
rect 38660 22049 38669 22083
rect 38669 22049 38703 22083
rect 38703 22049 38712 22083
rect 38660 22040 38712 22049
rect 38936 22083 38988 22092
rect 38936 22049 38945 22083
rect 38945 22049 38979 22083
rect 38979 22049 38988 22083
rect 38936 22040 38988 22049
rect 40040 22040 40092 22092
rect 40500 22083 40552 22092
rect 40500 22049 40509 22083
rect 40509 22049 40543 22083
rect 40543 22049 40552 22083
rect 40500 22040 40552 22049
rect 38384 22015 38436 22024
rect 38384 21981 38393 22015
rect 38393 21981 38427 22015
rect 38427 21981 38436 22015
rect 38384 21972 38436 21981
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 19064 21836 19116 21888
rect 19432 21836 19484 21888
rect 22468 21836 22520 21888
rect 23112 21836 23164 21888
rect 27436 21879 27488 21888
rect 27436 21845 27445 21879
rect 27445 21845 27479 21879
rect 27479 21845 27488 21879
rect 27436 21836 27488 21845
rect 27804 21947 27856 21956
rect 27804 21913 27838 21947
rect 27838 21913 27856 21947
rect 27804 21904 27856 21913
rect 27988 21904 28040 21956
rect 32220 21904 32272 21956
rect 33416 21904 33468 21956
rect 36360 21904 36412 21956
rect 41420 21972 41472 22024
rect 42524 22040 42576 22092
rect 42708 22040 42760 22092
rect 46572 22108 46624 22160
rect 47952 22108 48004 22160
rect 48596 22083 48648 22092
rect 48596 22049 48605 22083
rect 48605 22049 48639 22083
rect 48639 22049 48648 22083
rect 48596 22040 48648 22049
rect 50068 22176 50120 22228
rect 51080 22176 51132 22228
rect 43444 22015 43496 22024
rect 43444 21981 43453 22015
rect 43453 21981 43487 22015
rect 43487 21981 43496 22015
rect 43444 21972 43496 21981
rect 29460 21836 29512 21888
rect 29552 21879 29604 21888
rect 29552 21845 29561 21879
rect 29561 21845 29595 21879
rect 29595 21845 29604 21879
rect 29552 21836 29604 21845
rect 30656 21879 30708 21888
rect 30656 21845 30665 21879
rect 30665 21845 30699 21879
rect 30699 21845 30708 21879
rect 30656 21836 30708 21845
rect 31484 21836 31536 21888
rect 33048 21836 33100 21888
rect 34152 21879 34204 21888
rect 34152 21845 34161 21879
rect 34161 21845 34195 21879
rect 34195 21845 34204 21879
rect 34152 21836 34204 21845
rect 34704 21879 34756 21888
rect 34704 21845 34713 21879
rect 34713 21845 34747 21879
rect 34747 21845 34756 21879
rect 34704 21836 34756 21845
rect 36820 21879 36872 21888
rect 36820 21845 36829 21879
rect 36829 21845 36863 21879
rect 36863 21845 36872 21879
rect 36820 21836 36872 21845
rect 36912 21879 36964 21888
rect 36912 21845 36921 21879
rect 36921 21845 36955 21879
rect 36955 21845 36964 21879
rect 36912 21836 36964 21845
rect 37556 21836 37608 21888
rect 39028 21836 39080 21888
rect 39580 21836 39632 21888
rect 43628 21904 43680 21956
rect 46664 21972 46716 22024
rect 40132 21836 40184 21888
rect 42524 21836 42576 21888
rect 43812 21836 43864 21888
rect 45284 21879 45336 21888
rect 45284 21845 45293 21879
rect 45293 21845 45327 21879
rect 45327 21845 45336 21879
rect 45284 21836 45336 21845
rect 45376 21879 45428 21888
rect 45376 21845 45385 21879
rect 45385 21845 45419 21879
rect 45419 21845 45428 21879
rect 45376 21836 45428 21845
rect 45468 21836 45520 21888
rect 48136 21904 48188 21956
rect 49516 21904 49568 21956
rect 50160 22040 50212 22092
rect 51908 22176 51960 22228
rect 52552 22108 52604 22160
rect 54576 22083 54628 22092
rect 54576 22049 54585 22083
rect 54585 22049 54619 22083
rect 54619 22049 54628 22083
rect 54576 22040 54628 22049
rect 54668 22083 54720 22092
rect 54668 22049 54677 22083
rect 54677 22049 54711 22083
rect 54711 22049 54720 22083
rect 54668 22040 54720 22049
rect 55220 22040 55272 22092
rect 54024 21972 54076 22024
rect 56048 21972 56100 22024
rect 50252 21904 50304 21956
rect 52736 21904 52788 21956
rect 53472 21947 53524 21956
rect 53472 21913 53481 21947
rect 53481 21913 53515 21947
rect 53515 21913 53524 21947
rect 53472 21904 53524 21913
rect 47952 21879 48004 21888
rect 47952 21845 47961 21879
rect 47961 21845 47995 21879
rect 47995 21845 48004 21879
rect 47952 21836 48004 21845
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 49424 21836 49476 21888
rect 50896 21879 50948 21888
rect 50896 21845 50905 21879
rect 50905 21845 50939 21879
rect 50939 21845 50948 21879
rect 50896 21836 50948 21845
rect 52920 21879 52972 21888
rect 52920 21845 52929 21879
rect 52929 21845 52963 21879
rect 52963 21845 52972 21879
rect 52920 21836 52972 21845
rect 53288 21836 53340 21888
rect 54116 21879 54168 21888
rect 54116 21845 54125 21879
rect 54125 21845 54159 21879
rect 54159 21845 54168 21879
rect 54116 21836 54168 21845
rect 54576 21836 54628 21888
rect 57244 21836 57296 21888
rect 15394 21734 15446 21786
rect 15458 21734 15510 21786
rect 15522 21734 15574 21786
rect 15586 21734 15638 21786
rect 15650 21734 15702 21786
rect 29838 21734 29890 21786
rect 29902 21734 29954 21786
rect 29966 21734 30018 21786
rect 30030 21734 30082 21786
rect 30094 21734 30146 21786
rect 44282 21734 44334 21786
rect 44346 21734 44398 21786
rect 44410 21734 44462 21786
rect 44474 21734 44526 21786
rect 44538 21734 44590 21786
rect 58726 21734 58778 21786
rect 58790 21734 58842 21786
rect 58854 21734 58906 21786
rect 58918 21734 58970 21786
rect 58982 21734 59034 21786
rect 2964 21632 3016 21684
rect 4712 21632 4764 21684
rect 5724 21675 5776 21684
rect 5724 21641 5733 21675
rect 5733 21641 5767 21675
rect 5767 21641 5776 21675
rect 5724 21632 5776 21641
rect 6644 21632 6696 21684
rect 7196 21632 7248 21684
rect 10048 21632 10100 21684
rect 10692 21632 10744 21684
rect 11060 21675 11112 21684
rect 11060 21641 11069 21675
rect 11069 21641 11103 21675
rect 11103 21641 11112 21675
rect 11060 21632 11112 21641
rect 11980 21632 12032 21684
rect 12808 21632 12860 21684
rect 14372 21632 14424 21684
rect 16120 21632 16172 21684
rect 21088 21632 21140 21684
rect 22376 21632 22428 21684
rect 24952 21632 25004 21684
rect 3056 21607 3108 21616
rect 3056 21573 3074 21607
rect 3074 21573 3108 21607
rect 3056 21564 3108 21573
rect 3700 21539 3752 21548
rect 3700 21505 3734 21539
rect 3734 21505 3752 21539
rect 3700 21496 3752 21505
rect 4252 21496 4304 21548
rect 6184 21496 6236 21548
rect 9220 21564 9272 21616
rect 9864 21564 9916 21616
rect 20812 21564 20864 21616
rect 27988 21632 28040 21684
rect 25596 21607 25648 21616
rect 6460 21471 6512 21480
rect 6460 21437 6469 21471
rect 6469 21437 6503 21471
rect 6503 21437 6512 21471
rect 6460 21428 6512 21437
rect 10140 21496 10192 21548
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 13636 21496 13688 21548
rect 14556 21496 14608 21548
rect 18788 21496 18840 21548
rect 25596 21573 25630 21607
rect 25630 21573 25648 21607
rect 25596 21564 25648 21573
rect 23296 21496 23348 21548
rect 25320 21539 25372 21548
rect 25320 21505 25329 21539
rect 25329 21505 25363 21539
rect 25363 21505 25372 21539
rect 25320 21496 25372 21505
rect 7932 21335 7984 21344
rect 7932 21301 7941 21335
rect 7941 21301 7975 21335
rect 7975 21301 7984 21335
rect 7932 21292 7984 21301
rect 9036 21292 9088 21344
rect 22100 21360 22152 21412
rect 13544 21292 13596 21344
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 16212 21292 16264 21344
rect 16580 21292 16632 21344
rect 17684 21292 17736 21344
rect 18420 21292 18472 21344
rect 19064 21292 19116 21344
rect 19248 21292 19300 21344
rect 27436 21428 27488 21480
rect 27804 21428 27856 21480
rect 28448 21496 28500 21548
rect 28080 21428 28132 21480
rect 29552 21632 29604 21684
rect 31668 21632 31720 21684
rect 29460 21564 29512 21616
rect 31024 21564 31076 21616
rect 31484 21564 31536 21616
rect 33324 21632 33376 21684
rect 34060 21675 34112 21684
rect 34060 21641 34069 21675
rect 34069 21641 34103 21675
rect 34103 21641 34112 21675
rect 34060 21632 34112 21641
rect 34428 21632 34480 21684
rect 37464 21632 37516 21684
rect 37832 21632 37884 21684
rect 39580 21675 39632 21684
rect 39580 21641 39589 21675
rect 39589 21641 39623 21675
rect 39623 21641 39632 21675
rect 39580 21632 39632 21641
rect 40408 21632 40460 21684
rect 32956 21539 33008 21548
rect 26700 21403 26752 21412
rect 26700 21369 26709 21403
rect 26709 21369 26743 21403
rect 26743 21369 26752 21403
rect 26700 21360 26752 21369
rect 28356 21360 28408 21412
rect 30104 21428 30156 21480
rect 32956 21505 32974 21539
rect 32974 21505 33008 21539
rect 32956 21496 33008 21505
rect 33048 21539 33100 21548
rect 33048 21505 33057 21539
rect 33057 21505 33091 21539
rect 33091 21505 33100 21539
rect 33048 21496 33100 21505
rect 33784 21539 33836 21548
rect 33784 21505 33793 21539
rect 33793 21505 33827 21539
rect 33827 21505 33836 21539
rect 33784 21496 33836 21505
rect 24032 21292 24084 21344
rect 27620 21292 27672 21344
rect 28264 21292 28316 21344
rect 33324 21403 33376 21412
rect 33324 21369 33333 21403
rect 33333 21369 33367 21403
rect 33367 21369 33376 21403
rect 33324 21360 33376 21369
rect 33600 21428 33652 21480
rect 35440 21539 35492 21548
rect 35440 21505 35449 21539
rect 35449 21505 35483 21539
rect 35483 21505 35492 21539
rect 35440 21496 35492 21505
rect 35992 21496 36044 21548
rect 36820 21496 36872 21548
rect 38568 21564 38620 21616
rect 43444 21632 43496 21684
rect 45192 21675 45244 21684
rect 39212 21496 39264 21548
rect 40040 21539 40092 21548
rect 40040 21505 40049 21539
rect 40049 21505 40083 21539
rect 40083 21505 40092 21539
rect 40040 21496 40092 21505
rect 40776 21496 40828 21548
rect 42708 21607 42760 21616
rect 42708 21573 42717 21607
rect 42717 21573 42751 21607
rect 42751 21573 42760 21607
rect 42708 21564 42760 21573
rect 41512 21496 41564 21548
rect 43628 21496 43680 21548
rect 43812 21539 43864 21548
rect 43812 21505 43821 21539
rect 43821 21505 43855 21539
rect 43855 21505 43864 21539
rect 43812 21496 43864 21505
rect 45192 21641 45201 21675
rect 45201 21641 45235 21675
rect 45235 21641 45244 21675
rect 45192 21632 45244 21641
rect 45560 21675 45612 21684
rect 45560 21641 45569 21675
rect 45569 21641 45603 21675
rect 45603 21641 45612 21675
rect 45560 21632 45612 21641
rect 49056 21675 49108 21684
rect 49056 21641 49065 21675
rect 49065 21641 49099 21675
rect 49099 21641 49108 21675
rect 49056 21632 49108 21641
rect 49148 21632 49200 21684
rect 51172 21675 51224 21684
rect 51172 21641 51181 21675
rect 51181 21641 51215 21675
rect 51215 21641 51224 21675
rect 51172 21632 51224 21641
rect 52552 21675 52604 21684
rect 52552 21641 52561 21675
rect 52561 21641 52595 21675
rect 52595 21641 52604 21675
rect 52552 21632 52604 21641
rect 52736 21675 52788 21684
rect 52736 21641 52745 21675
rect 52745 21641 52779 21675
rect 52779 21641 52788 21675
rect 52736 21632 52788 21641
rect 54024 21632 54076 21684
rect 54208 21675 54260 21684
rect 54208 21641 54217 21675
rect 54217 21641 54251 21675
rect 54251 21641 54260 21675
rect 54208 21632 54260 21641
rect 45284 21564 45336 21616
rect 52920 21564 52972 21616
rect 40132 21471 40184 21480
rect 40132 21437 40141 21471
rect 40141 21437 40175 21471
rect 40175 21437 40184 21471
rect 40132 21428 40184 21437
rect 29276 21292 29328 21344
rect 31852 21335 31904 21344
rect 31852 21301 31861 21335
rect 31861 21301 31895 21335
rect 31895 21301 31904 21335
rect 31852 21292 31904 21301
rect 33508 21292 33560 21344
rect 33784 21292 33836 21344
rect 34060 21292 34112 21344
rect 44824 21428 44876 21480
rect 44916 21471 44968 21480
rect 44916 21437 44925 21471
rect 44925 21437 44959 21471
rect 44959 21437 44968 21471
rect 44916 21428 44968 21437
rect 45008 21428 45060 21480
rect 45376 21428 45428 21480
rect 45560 21496 45612 21548
rect 47952 21496 48004 21548
rect 49240 21496 49292 21548
rect 50896 21496 50948 21548
rect 53288 21539 53340 21548
rect 53288 21505 53297 21539
rect 53297 21505 53331 21539
rect 53331 21505 53340 21539
rect 53288 21496 53340 21505
rect 54116 21496 54168 21548
rect 42432 21360 42484 21412
rect 45560 21360 45612 21412
rect 48964 21360 49016 21412
rect 49332 21360 49384 21412
rect 40408 21292 40460 21344
rect 40776 21335 40828 21344
rect 40776 21301 40785 21335
rect 40785 21301 40819 21335
rect 40819 21301 40828 21335
rect 40776 21292 40828 21301
rect 44732 21292 44784 21344
rect 46572 21292 46624 21344
rect 48596 21292 48648 21344
rect 55220 21403 55272 21412
rect 50160 21292 50212 21344
rect 55220 21369 55229 21403
rect 55229 21369 55263 21403
rect 55263 21369 55272 21403
rect 55220 21360 55272 21369
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 22616 21190 22668 21242
rect 22680 21190 22732 21242
rect 22744 21190 22796 21242
rect 22808 21190 22860 21242
rect 22872 21190 22924 21242
rect 37060 21190 37112 21242
rect 37124 21190 37176 21242
rect 37188 21190 37240 21242
rect 37252 21190 37304 21242
rect 37316 21190 37368 21242
rect 51504 21190 51556 21242
rect 51568 21190 51620 21242
rect 51632 21190 51684 21242
rect 51696 21190 51748 21242
rect 51760 21190 51812 21242
rect 4436 21088 4488 21140
rect 5264 21020 5316 21072
rect 4620 20952 4672 21004
rect 7748 21088 7800 21140
rect 7932 21088 7984 21140
rect 7012 20952 7064 21004
rect 7104 20995 7156 21004
rect 7104 20961 7113 20995
rect 7113 20961 7147 20995
rect 7147 20961 7156 20995
rect 7104 20952 7156 20961
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 5908 20927 5960 20936
rect 5908 20893 5917 20927
rect 5917 20893 5951 20927
rect 5951 20893 5960 20927
rect 5908 20884 5960 20893
rect 12440 21088 12492 21140
rect 16856 21088 16908 21140
rect 22192 21131 22244 21140
rect 10876 21020 10928 21072
rect 9036 20884 9088 20936
rect 9312 20816 9364 20868
rect 4252 20748 4304 20800
rect 6092 20748 6144 20800
rect 6184 20748 6236 20800
rect 8760 20748 8812 20800
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 11152 20952 11204 21004
rect 11244 20995 11296 21004
rect 11244 20961 11253 20995
rect 11253 20961 11287 20995
rect 11287 20961 11296 20995
rect 11244 20952 11296 20961
rect 14280 21020 14332 21072
rect 16672 21020 16724 21072
rect 11796 20995 11848 21004
rect 11796 20961 11805 20995
rect 11805 20961 11839 20995
rect 11839 20961 11848 20995
rect 11796 20952 11848 20961
rect 15384 20952 15436 21004
rect 16396 20995 16448 21004
rect 16396 20961 16405 20995
rect 16405 20961 16439 20995
rect 16439 20961 16448 20995
rect 16396 20952 16448 20961
rect 11612 20927 11664 20936
rect 11612 20893 11646 20927
rect 11646 20893 11664 20927
rect 11612 20884 11664 20893
rect 15016 20927 15068 20936
rect 15016 20893 15025 20927
rect 15025 20893 15059 20927
rect 15059 20893 15068 20927
rect 15016 20884 15068 20893
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 20720 20952 20772 21004
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 18880 20884 18932 20936
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 20168 20816 20220 20868
rect 12072 20748 12124 20800
rect 13912 20748 13964 20800
rect 14372 20748 14424 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16488 20748 16540 20757
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17408 20791 17460 20800
rect 17408 20757 17417 20791
rect 17417 20757 17451 20791
rect 17451 20757 17460 20791
rect 17408 20748 17460 20757
rect 20720 20791 20772 20800
rect 20720 20757 20729 20791
rect 20729 20757 20763 20791
rect 20763 20757 20772 20791
rect 20720 20748 20772 20757
rect 21272 20995 21324 21004
rect 21272 20961 21281 20995
rect 21281 20961 21315 20995
rect 21315 20961 21324 20995
rect 21272 20952 21324 20961
rect 22192 21097 22201 21131
rect 22201 21097 22235 21131
rect 22235 21097 22244 21131
rect 22192 21088 22244 21097
rect 22284 21131 22336 21140
rect 22284 21097 22293 21131
rect 22293 21097 22327 21131
rect 22327 21097 22336 21131
rect 22284 21088 22336 21097
rect 24032 21088 24084 21140
rect 23388 20952 23440 21004
rect 25320 21088 25372 21140
rect 29368 21131 29420 21140
rect 29368 21097 29377 21131
rect 29377 21097 29411 21131
rect 29411 21097 29420 21131
rect 29368 21088 29420 21097
rect 31852 21088 31904 21140
rect 32220 21131 32272 21140
rect 32220 21097 32229 21131
rect 32229 21097 32263 21131
rect 32263 21097 32272 21131
rect 32220 21088 32272 21097
rect 33324 21088 33376 21140
rect 33968 21131 34020 21140
rect 33968 21097 33977 21131
rect 33977 21097 34011 21131
rect 34011 21097 34020 21131
rect 33968 21088 34020 21097
rect 34704 21088 34756 21140
rect 36360 21131 36412 21140
rect 36360 21097 36369 21131
rect 36369 21097 36403 21131
rect 36403 21097 36412 21131
rect 36360 21088 36412 21097
rect 38568 21088 38620 21140
rect 23204 20884 23256 20936
rect 27988 20995 28040 21004
rect 27988 20961 27997 20995
rect 27997 20961 28031 20995
rect 28031 20961 28040 20995
rect 27988 20952 28040 20961
rect 32588 20995 32640 21004
rect 21272 20816 21324 20868
rect 29644 20884 29696 20936
rect 30104 20927 30156 20936
rect 30104 20893 30113 20927
rect 30113 20893 30147 20927
rect 30147 20893 30156 20927
rect 32588 20961 32597 20995
rect 32597 20961 32631 20995
rect 32631 20961 32640 20995
rect 32588 20952 32640 20961
rect 30104 20884 30156 20893
rect 25964 20816 26016 20868
rect 27804 20816 27856 20868
rect 28724 20816 28776 20868
rect 30564 20816 30616 20868
rect 23112 20748 23164 20800
rect 26424 20791 26476 20800
rect 26424 20757 26433 20791
rect 26433 20757 26467 20791
rect 26467 20757 26476 20791
rect 26424 20748 26476 20757
rect 26516 20791 26568 20800
rect 26516 20757 26525 20791
rect 26525 20757 26559 20791
rect 26559 20757 26568 20791
rect 26516 20748 26568 20757
rect 26976 20791 27028 20800
rect 26976 20757 26985 20791
rect 26985 20757 27019 20791
rect 27019 20757 27028 20791
rect 26976 20748 27028 20757
rect 37648 21063 37700 21072
rect 37648 21029 37657 21063
rect 37657 21029 37691 21063
rect 37691 21029 37700 21063
rect 37648 21020 37700 21029
rect 38384 21020 38436 21072
rect 36912 20995 36964 21004
rect 36912 20961 36921 20995
rect 36921 20961 36955 20995
rect 36955 20961 36964 20995
rect 36912 20952 36964 20961
rect 40408 21131 40460 21140
rect 40408 21097 40417 21131
rect 40417 21097 40451 21131
rect 40451 21097 40460 21131
rect 40408 21088 40460 21097
rect 43812 21088 43864 21140
rect 44824 21088 44876 21140
rect 45192 21131 45244 21140
rect 45192 21097 45201 21131
rect 45201 21097 45235 21131
rect 45235 21097 45244 21131
rect 45192 21088 45244 21097
rect 45560 21131 45612 21140
rect 45560 21097 45569 21131
rect 45569 21097 45603 21131
rect 45603 21097 45612 21131
rect 45560 21088 45612 21097
rect 49056 21088 49108 21140
rect 49516 21088 49568 21140
rect 54668 21088 54720 21140
rect 42616 20952 42668 21004
rect 40776 20884 40828 20936
rect 44916 21020 44968 21072
rect 54484 21020 54536 21072
rect 56508 21020 56560 21072
rect 48136 20995 48188 21004
rect 48136 20961 48145 20995
rect 48145 20961 48179 20995
rect 48179 20961 48188 20995
rect 48136 20952 48188 20961
rect 48780 20952 48832 21004
rect 55220 20952 55272 21004
rect 55864 20927 55916 20936
rect 55864 20893 55873 20927
rect 55873 20893 55907 20927
rect 55907 20893 55916 20927
rect 55864 20884 55916 20893
rect 56048 20927 56100 20936
rect 56048 20893 56057 20927
rect 56057 20893 56091 20927
rect 56091 20893 56100 20927
rect 56048 20884 56100 20893
rect 57336 20927 57388 20936
rect 57336 20893 57345 20927
rect 57345 20893 57379 20927
rect 57379 20893 57388 20927
rect 57336 20884 57388 20893
rect 55404 20816 55456 20868
rect 33784 20748 33836 20800
rect 37832 20748 37884 20800
rect 48596 20748 48648 20800
rect 49056 20791 49108 20800
rect 49056 20757 49065 20791
rect 49065 20757 49099 20791
rect 49099 20757 49108 20791
rect 49056 20748 49108 20757
rect 52460 20748 52512 20800
rect 53840 20748 53892 20800
rect 55312 20791 55364 20800
rect 55312 20757 55321 20791
rect 55321 20757 55355 20791
rect 55355 20757 55364 20791
rect 55312 20748 55364 20757
rect 56692 20791 56744 20800
rect 56692 20757 56701 20791
rect 56701 20757 56735 20791
rect 56735 20757 56744 20791
rect 56692 20748 56744 20757
rect 56784 20791 56836 20800
rect 56784 20757 56793 20791
rect 56793 20757 56827 20791
rect 56827 20757 56836 20791
rect 56784 20748 56836 20757
rect 15394 20646 15446 20698
rect 15458 20646 15510 20698
rect 15522 20646 15574 20698
rect 15586 20646 15638 20698
rect 15650 20646 15702 20698
rect 29838 20646 29890 20698
rect 29902 20646 29954 20698
rect 29966 20646 30018 20698
rect 30030 20646 30082 20698
rect 30094 20646 30146 20698
rect 44282 20646 44334 20698
rect 44346 20646 44398 20698
rect 44410 20646 44462 20698
rect 44474 20646 44526 20698
rect 44538 20646 44590 20698
rect 58726 20646 58778 20698
rect 58790 20646 58842 20698
rect 58854 20646 58906 20698
rect 58918 20646 58970 20698
rect 58982 20646 59034 20698
rect 6092 20544 6144 20596
rect 7012 20544 7064 20596
rect 11612 20544 11664 20596
rect 11796 20544 11848 20596
rect 15016 20544 15068 20596
rect 17408 20544 17460 20596
rect 20168 20587 20220 20596
rect 20168 20553 20177 20587
rect 20177 20553 20211 20587
rect 20211 20553 20220 20587
rect 20168 20544 20220 20553
rect 21088 20587 21140 20596
rect 21088 20553 21097 20587
rect 21097 20553 21131 20587
rect 21131 20553 21140 20587
rect 21088 20544 21140 20553
rect 22468 20544 22520 20596
rect 23296 20544 23348 20596
rect 25964 20587 26016 20596
rect 25964 20553 25973 20587
rect 25973 20553 26007 20587
rect 26007 20553 26016 20587
rect 25964 20544 26016 20553
rect 27804 20544 27856 20596
rect 27896 20587 27948 20596
rect 27896 20553 27905 20587
rect 27905 20553 27939 20587
rect 27939 20553 27948 20587
rect 27896 20544 27948 20553
rect 28448 20544 28500 20596
rect 28724 20587 28776 20596
rect 28724 20553 28733 20587
rect 28733 20553 28767 20587
rect 28767 20553 28776 20587
rect 28724 20544 28776 20553
rect 30564 20587 30616 20596
rect 30564 20553 30573 20587
rect 30573 20553 30607 20587
rect 30607 20553 30616 20587
rect 30564 20544 30616 20553
rect 37648 20587 37700 20596
rect 37648 20553 37657 20587
rect 37657 20553 37691 20587
rect 37691 20553 37700 20587
rect 37648 20544 37700 20553
rect 54668 20544 54720 20596
rect 55864 20544 55916 20596
rect 22100 20476 22152 20528
rect 23388 20476 23440 20528
rect 26976 20476 27028 20528
rect 28264 20519 28316 20528
rect 28264 20485 28273 20519
rect 28273 20485 28307 20519
rect 28307 20485 28316 20519
rect 28264 20476 28316 20485
rect 44640 20476 44692 20528
rect 50252 20476 50304 20528
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 15844 20408 15896 20460
rect 4528 20383 4580 20392
rect 4528 20349 4537 20383
rect 4537 20349 4571 20383
rect 4571 20349 4580 20383
rect 4528 20340 4580 20349
rect 5908 20340 5960 20392
rect 10048 20383 10100 20392
rect 10048 20349 10057 20383
rect 10057 20349 10091 20383
rect 10091 20349 10100 20383
rect 10048 20340 10100 20349
rect 10140 20340 10192 20392
rect 14924 20383 14976 20392
rect 14924 20349 14933 20383
rect 14933 20349 14967 20383
rect 14967 20349 14976 20383
rect 14924 20340 14976 20349
rect 15200 20340 15252 20392
rect 16028 20340 16080 20392
rect 17132 20340 17184 20392
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 26424 20408 26476 20460
rect 26516 20451 26568 20460
rect 26516 20417 26525 20451
rect 26525 20417 26559 20451
rect 26559 20417 26568 20451
rect 26516 20408 26568 20417
rect 29276 20451 29328 20460
rect 29276 20417 29285 20451
rect 29285 20417 29319 20451
rect 29319 20417 29328 20451
rect 29276 20408 29328 20417
rect 30656 20408 30708 20460
rect 54576 20451 54628 20460
rect 22468 20340 22520 20392
rect 23480 20383 23532 20392
rect 23480 20349 23489 20383
rect 23489 20349 23523 20383
rect 23523 20349 23532 20383
rect 23480 20340 23532 20349
rect 28448 20383 28500 20392
rect 28448 20349 28457 20383
rect 28457 20349 28491 20383
rect 28491 20349 28500 20383
rect 28448 20340 28500 20349
rect 45560 20383 45612 20392
rect 45560 20349 45569 20383
rect 45569 20349 45603 20383
rect 45603 20349 45612 20383
rect 45560 20340 45612 20349
rect 48228 20383 48280 20392
rect 48228 20349 48237 20383
rect 48237 20349 48271 20383
rect 48271 20349 48280 20383
rect 48228 20340 48280 20349
rect 48412 20383 48464 20392
rect 48412 20349 48421 20383
rect 48421 20349 48455 20383
rect 48455 20349 48464 20383
rect 48412 20340 48464 20349
rect 54576 20417 54585 20451
rect 54585 20417 54619 20451
rect 54619 20417 54628 20451
rect 54576 20408 54628 20417
rect 54208 20383 54260 20392
rect 54208 20349 54217 20383
rect 54217 20349 54251 20383
rect 54251 20349 54260 20383
rect 54208 20340 54260 20349
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 6552 20247 6604 20256
rect 6552 20213 6561 20247
rect 6561 20213 6595 20247
rect 6595 20213 6604 20247
rect 6552 20204 6604 20213
rect 7288 20204 7340 20256
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 14096 20204 14148 20256
rect 49332 20315 49384 20324
rect 49332 20281 49341 20315
rect 49341 20281 49375 20315
rect 49375 20281 49384 20315
rect 49332 20272 49384 20281
rect 50252 20272 50304 20324
rect 55128 20408 55180 20460
rect 55404 20408 55456 20460
rect 56784 20476 56836 20528
rect 56876 20408 56928 20460
rect 16488 20204 16540 20256
rect 18604 20204 18656 20256
rect 23020 20204 23072 20256
rect 38108 20204 38160 20256
rect 39764 20247 39816 20256
rect 39764 20213 39773 20247
rect 39773 20213 39807 20247
rect 39807 20213 39816 20247
rect 39764 20204 39816 20213
rect 44548 20204 44600 20256
rect 44824 20247 44876 20256
rect 44824 20213 44833 20247
rect 44833 20213 44867 20247
rect 44867 20213 44876 20247
rect 44824 20204 44876 20213
rect 45376 20204 45428 20256
rect 47308 20204 47360 20256
rect 48688 20204 48740 20256
rect 53656 20247 53708 20256
rect 53656 20213 53665 20247
rect 53665 20213 53699 20247
rect 53699 20213 53708 20247
rect 53656 20204 53708 20213
rect 56324 20383 56376 20392
rect 56324 20349 56333 20383
rect 56333 20349 56367 20383
rect 56367 20349 56376 20383
rect 56324 20340 56376 20349
rect 56692 20204 56744 20256
rect 57244 20204 57296 20256
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 22616 20102 22668 20154
rect 22680 20102 22732 20154
rect 22744 20102 22796 20154
rect 22808 20102 22860 20154
rect 22872 20102 22924 20154
rect 37060 20102 37112 20154
rect 37124 20102 37176 20154
rect 37188 20102 37240 20154
rect 37252 20102 37304 20154
rect 37316 20102 37368 20154
rect 51504 20102 51556 20154
rect 51568 20102 51620 20154
rect 51632 20102 51684 20154
rect 51696 20102 51748 20154
rect 51760 20102 51812 20154
rect 4528 20043 4580 20052
rect 4528 20009 4537 20043
rect 4537 20009 4571 20043
rect 4571 20009 4580 20043
rect 4528 20000 4580 20009
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 6092 19728 6144 19780
rect 18696 20000 18748 20052
rect 21732 20043 21784 20052
rect 21732 20009 21741 20043
rect 21741 20009 21775 20043
rect 21775 20009 21784 20043
rect 21732 20000 21784 20009
rect 23480 20000 23532 20052
rect 9312 19975 9364 19984
rect 9312 19941 9321 19975
rect 9321 19941 9355 19975
rect 9355 19941 9364 19975
rect 9312 19932 9364 19941
rect 9404 19932 9456 19984
rect 11244 19932 11296 19984
rect 15292 19932 15344 19984
rect 16672 19932 16724 19984
rect 17408 19932 17460 19984
rect 13820 19864 13872 19916
rect 15844 19864 15896 19916
rect 14372 19839 14424 19848
rect 14372 19805 14406 19839
rect 14406 19805 14424 19839
rect 14372 19796 14424 19805
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 18052 19796 18104 19848
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 22468 19864 22520 19916
rect 23112 19907 23164 19916
rect 23112 19873 23121 19907
rect 23121 19873 23155 19907
rect 23155 19873 23164 19907
rect 23112 19864 23164 19873
rect 23204 19864 23256 19916
rect 23388 19932 23440 19984
rect 28448 20000 28500 20052
rect 38844 19932 38896 19984
rect 24952 19839 25004 19848
rect 24952 19805 24961 19839
rect 24961 19805 24995 19839
rect 24995 19805 25004 19839
rect 24952 19796 25004 19805
rect 26240 19839 26292 19848
rect 26240 19805 26249 19839
rect 26249 19805 26283 19839
rect 26283 19805 26292 19839
rect 26240 19796 26292 19805
rect 26516 19839 26568 19848
rect 26516 19805 26525 19839
rect 26525 19805 26559 19839
rect 26559 19805 26568 19839
rect 26516 19796 26568 19805
rect 9680 19728 9732 19780
rect 10048 19728 10100 19780
rect 17868 19728 17920 19780
rect 17960 19728 18012 19780
rect 18604 19771 18656 19780
rect 18604 19737 18622 19771
rect 18622 19737 18656 19771
rect 18604 19728 18656 19737
rect 21088 19771 21140 19780
rect 21088 19737 21097 19771
rect 21097 19737 21131 19771
rect 21131 19737 21140 19771
rect 21088 19728 21140 19737
rect 4252 19660 4304 19712
rect 6460 19660 6512 19712
rect 9128 19660 9180 19712
rect 10784 19660 10836 19712
rect 11244 19660 11296 19712
rect 12256 19660 12308 19712
rect 14280 19660 14332 19712
rect 16948 19660 17000 19712
rect 22928 19728 22980 19780
rect 36912 19864 36964 19916
rect 38108 19864 38160 19916
rect 48228 20043 48280 20052
rect 48228 20009 48237 20043
rect 48237 20009 48271 20043
rect 48271 20009 48280 20043
rect 48228 20000 48280 20009
rect 48412 20000 48464 20052
rect 49332 20000 49384 20052
rect 50252 20000 50304 20052
rect 54576 20000 54628 20052
rect 56692 20000 56744 20052
rect 56876 20000 56928 20052
rect 44916 19932 44968 19984
rect 39764 19864 39816 19916
rect 44548 19864 44600 19916
rect 44640 19907 44692 19916
rect 44640 19873 44649 19907
rect 44649 19873 44683 19907
rect 44683 19873 44692 19907
rect 44640 19864 44692 19873
rect 44824 19864 44876 19916
rect 46664 19864 46716 19916
rect 30656 19839 30708 19848
rect 30656 19805 30665 19839
rect 30665 19805 30699 19839
rect 30699 19805 30708 19839
rect 30656 19796 30708 19805
rect 31392 19839 31444 19848
rect 31392 19805 31401 19839
rect 31401 19805 31435 19839
rect 31435 19805 31444 19839
rect 31392 19796 31444 19805
rect 33784 19771 33836 19780
rect 33784 19737 33793 19771
rect 33793 19737 33827 19771
rect 33827 19737 33836 19771
rect 33784 19728 33836 19737
rect 37648 19839 37700 19848
rect 37648 19805 37657 19839
rect 37657 19805 37691 19839
rect 37691 19805 37700 19839
rect 37648 19796 37700 19805
rect 39028 19796 39080 19848
rect 41972 19839 42024 19848
rect 41972 19805 41981 19839
rect 41981 19805 42015 19839
rect 42015 19805 42024 19839
rect 41972 19796 42024 19805
rect 42708 19796 42760 19848
rect 45008 19796 45060 19848
rect 47308 19796 47360 19848
rect 47860 19796 47912 19848
rect 48688 19907 48740 19916
rect 48688 19873 48697 19907
rect 48697 19873 48731 19907
rect 48731 19873 48740 19907
rect 48688 19864 48740 19873
rect 48780 19907 48832 19916
rect 48780 19873 48789 19907
rect 48789 19873 48823 19907
rect 48823 19873 48832 19907
rect 48780 19864 48832 19873
rect 49240 19864 49292 19916
rect 56508 19975 56560 19984
rect 56508 19941 56517 19975
rect 56517 19941 56551 19975
rect 56551 19941 56560 19975
rect 56508 19932 56560 19941
rect 55404 19864 55456 19916
rect 49332 19796 49384 19848
rect 49608 19839 49660 19848
rect 49608 19805 49617 19839
rect 49617 19805 49651 19839
rect 49651 19805 49660 19839
rect 49608 19796 49660 19805
rect 50344 19796 50396 19848
rect 51908 19796 51960 19848
rect 39580 19771 39632 19780
rect 39580 19737 39589 19771
rect 39589 19737 39623 19771
rect 39623 19737 39632 19771
rect 39580 19728 39632 19737
rect 48412 19728 48464 19780
rect 53656 19796 53708 19848
rect 53932 19796 53984 19848
rect 56140 19839 56192 19848
rect 56140 19805 56158 19839
rect 56158 19805 56192 19839
rect 56140 19796 56192 19805
rect 57244 19864 57296 19916
rect 57428 19907 57480 19916
rect 57428 19873 57437 19907
rect 57437 19873 57471 19907
rect 57471 19873 57480 19907
rect 57428 19864 57480 19873
rect 19708 19703 19760 19712
rect 19708 19669 19717 19703
rect 19717 19669 19751 19703
rect 19751 19669 19760 19703
rect 19708 19660 19760 19669
rect 22284 19660 22336 19712
rect 22836 19660 22888 19712
rect 23848 19703 23900 19712
rect 23848 19669 23857 19703
rect 23857 19669 23891 19703
rect 23891 19669 23900 19703
rect 23848 19660 23900 19669
rect 25596 19703 25648 19712
rect 25596 19669 25605 19703
rect 25605 19669 25639 19703
rect 25639 19669 25648 19703
rect 25596 19660 25648 19669
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 27436 19703 27488 19712
rect 27436 19669 27445 19703
rect 27445 19669 27479 19703
rect 27479 19669 27488 19703
rect 27436 19660 27488 19669
rect 29736 19660 29788 19712
rect 30840 19703 30892 19712
rect 30840 19669 30849 19703
rect 30849 19669 30883 19703
rect 30883 19669 30892 19703
rect 30840 19660 30892 19669
rect 31760 19703 31812 19712
rect 31760 19669 31769 19703
rect 31769 19669 31803 19703
rect 31803 19669 31812 19703
rect 31760 19660 31812 19669
rect 32312 19660 32364 19712
rect 33692 19660 33744 19712
rect 35348 19703 35400 19712
rect 35348 19669 35357 19703
rect 35357 19669 35391 19703
rect 35391 19669 35400 19703
rect 35348 19660 35400 19669
rect 37556 19660 37608 19712
rect 37740 19660 37792 19712
rect 38476 19660 38528 19712
rect 38660 19660 38712 19712
rect 38936 19703 38988 19712
rect 38936 19669 38945 19703
rect 38945 19669 38979 19703
rect 38979 19669 38988 19703
rect 38936 19660 38988 19669
rect 39028 19703 39080 19712
rect 39028 19669 39037 19703
rect 39037 19669 39071 19703
rect 39071 19669 39080 19703
rect 39028 19660 39080 19669
rect 39120 19660 39172 19712
rect 40592 19703 40644 19712
rect 40592 19669 40601 19703
rect 40601 19669 40635 19703
rect 40635 19669 40644 19703
rect 40592 19660 40644 19669
rect 41420 19703 41472 19712
rect 41420 19669 41429 19703
rect 41429 19669 41463 19703
rect 41463 19669 41472 19703
rect 41420 19660 41472 19669
rect 44180 19660 44232 19712
rect 44640 19660 44692 19712
rect 45376 19703 45428 19712
rect 45376 19669 45385 19703
rect 45385 19669 45419 19703
rect 45419 19669 45428 19703
rect 45376 19660 45428 19669
rect 45836 19703 45888 19712
rect 45836 19669 45845 19703
rect 45845 19669 45879 19703
rect 45879 19669 45888 19703
rect 45836 19660 45888 19669
rect 48780 19660 48832 19712
rect 49424 19660 49476 19712
rect 49884 19660 49936 19712
rect 51724 19703 51776 19712
rect 51724 19669 51733 19703
rect 51733 19669 51767 19703
rect 51767 19669 51776 19703
rect 51724 19660 51776 19669
rect 55220 19728 55272 19780
rect 54392 19703 54444 19712
rect 54392 19669 54401 19703
rect 54401 19669 54435 19703
rect 54435 19669 54444 19703
rect 54392 19660 54444 19669
rect 57520 19703 57572 19712
rect 57520 19669 57529 19703
rect 57529 19669 57563 19703
rect 57563 19669 57572 19703
rect 57520 19660 57572 19669
rect 57612 19703 57664 19712
rect 57612 19669 57621 19703
rect 57621 19669 57655 19703
rect 57655 19669 57664 19703
rect 57612 19660 57664 19669
rect 57980 19703 58032 19712
rect 57980 19669 57989 19703
rect 57989 19669 58023 19703
rect 58023 19669 58032 19703
rect 57980 19660 58032 19669
rect 15394 19558 15446 19610
rect 15458 19558 15510 19610
rect 15522 19558 15574 19610
rect 15586 19558 15638 19610
rect 15650 19558 15702 19610
rect 29838 19558 29890 19610
rect 29902 19558 29954 19610
rect 29966 19558 30018 19610
rect 30030 19558 30082 19610
rect 30094 19558 30146 19610
rect 44282 19558 44334 19610
rect 44346 19558 44398 19610
rect 44410 19558 44462 19610
rect 44474 19558 44526 19610
rect 44538 19558 44590 19610
rect 58726 19558 58778 19610
rect 58790 19558 58842 19610
rect 58854 19558 58906 19610
rect 58918 19558 58970 19610
rect 58982 19558 59034 19610
rect 4804 19456 4856 19508
rect 11244 19456 11296 19508
rect 15200 19499 15252 19508
rect 15200 19465 15209 19499
rect 15209 19465 15243 19499
rect 15243 19465 15252 19499
rect 15200 19456 15252 19465
rect 16488 19456 16540 19508
rect 17960 19456 18012 19508
rect 2412 19320 2464 19372
rect 2780 19363 2832 19372
rect 2780 19329 2814 19363
rect 2814 19329 2832 19363
rect 2780 19320 2832 19329
rect 5080 19363 5132 19372
rect 5080 19329 5098 19363
rect 5098 19329 5132 19363
rect 5080 19320 5132 19329
rect 6460 19320 6512 19372
rect 7932 19252 7984 19304
rect 14924 19388 14976 19440
rect 17132 19388 17184 19440
rect 11060 19320 11112 19372
rect 13820 19363 13872 19372
rect 13820 19329 13829 19363
rect 13829 19329 13863 19363
rect 13863 19329 13872 19363
rect 13820 19320 13872 19329
rect 14372 19320 14424 19372
rect 16028 19320 16080 19372
rect 17960 19320 18012 19372
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 20260 19456 20312 19508
rect 21088 19456 21140 19508
rect 20628 19320 20680 19372
rect 21916 19320 21968 19372
rect 22928 19456 22980 19508
rect 23296 19456 23348 19508
rect 25596 19456 25648 19508
rect 26516 19499 26568 19508
rect 26516 19465 26525 19499
rect 26525 19465 26559 19499
rect 26559 19465 26568 19499
rect 26516 19456 26568 19465
rect 30656 19456 30708 19508
rect 30840 19456 30892 19508
rect 35256 19456 35308 19508
rect 37648 19456 37700 19508
rect 39120 19456 39172 19508
rect 35992 19388 36044 19440
rect 10232 19295 10284 19304
rect 10232 19261 10241 19295
rect 10241 19261 10275 19295
rect 10275 19261 10284 19295
rect 10232 19252 10284 19261
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 12072 19252 12124 19304
rect 12624 19295 12676 19304
rect 12624 19261 12633 19295
rect 12633 19261 12667 19295
rect 12667 19261 12676 19295
rect 12624 19252 12676 19261
rect 15844 19295 15896 19304
rect 15844 19261 15853 19295
rect 15853 19261 15887 19295
rect 15887 19261 15896 19295
rect 15844 19252 15896 19261
rect 19340 19252 19392 19304
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 6000 19116 6052 19168
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 9772 19116 9824 19168
rect 11888 19116 11940 19168
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 16212 19116 16264 19168
rect 21180 19184 21232 19236
rect 22836 19295 22888 19346
rect 27528 19320 27580 19372
rect 31484 19320 31536 19372
rect 35440 19320 35492 19372
rect 38476 19320 38528 19372
rect 40224 19456 40276 19508
rect 45560 19456 45612 19508
rect 45836 19456 45888 19508
rect 49148 19456 49200 19508
rect 50344 19499 50396 19508
rect 50344 19465 50353 19499
rect 50353 19465 50387 19499
rect 50387 19465 50396 19499
rect 50344 19456 50396 19465
rect 51724 19456 51776 19508
rect 39580 19388 39632 19440
rect 47860 19431 47912 19440
rect 47860 19397 47869 19431
rect 47869 19397 47903 19431
rect 47903 19397 47912 19431
rect 47860 19388 47912 19397
rect 48412 19431 48464 19440
rect 48412 19397 48421 19431
rect 48421 19397 48455 19431
rect 48455 19397 48464 19431
rect 48412 19388 48464 19397
rect 22836 19294 22870 19295
rect 22870 19294 22888 19295
rect 23204 19252 23256 19304
rect 23848 19295 23900 19304
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 19340 19116 19392 19168
rect 21088 19116 21140 19168
rect 22284 19184 22336 19236
rect 22468 19227 22520 19236
rect 22468 19193 22477 19227
rect 22477 19193 22511 19227
rect 22511 19193 22520 19227
rect 22468 19184 22520 19193
rect 21548 19116 21600 19168
rect 23848 19261 23857 19295
rect 23857 19261 23891 19295
rect 23891 19261 23900 19295
rect 23848 19252 23900 19261
rect 24860 19252 24912 19304
rect 27160 19295 27212 19304
rect 27160 19261 27169 19295
rect 27169 19261 27203 19295
rect 27203 19261 27212 19295
rect 27160 19252 27212 19261
rect 30196 19295 30248 19304
rect 30196 19261 30205 19295
rect 30205 19261 30239 19295
rect 30239 19261 30248 19295
rect 30196 19252 30248 19261
rect 29276 19184 29328 19236
rect 31300 19295 31352 19304
rect 31300 19261 31309 19295
rect 31309 19261 31343 19295
rect 31343 19261 31352 19295
rect 31300 19252 31352 19261
rect 32128 19252 32180 19304
rect 32588 19252 32640 19304
rect 34704 19295 34756 19304
rect 34704 19261 34713 19295
rect 34713 19261 34747 19295
rect 34747 19261 34756 19295
rect 34704 19252 34756 19261
rect 38384 19295 38436 19304
rect 38384 19261 38393 19295
rect 38393 19261 38427 19295
rect 38427 19261 38436 19295
rect 38384 19252 38436 19261
rect 31760 19184 31812 19236
rect 24492 19159 24544 19168
rect 24492 19125 24501 19159
rect 24501 19125 24535 19159
rect 24535 19125 24544 19159
rect 24492 19116 24544 19125
rect 27896 19116 27948 19168
rect 29552 19159 29604 19168
rect 29552 19125 29561 19159
rect 29561 19125 29595 19159
rect 29595 19125 29604 19159
rect 29552 19116 29604 19125
rect 31944 19159 31996 19168
rect 31944 19125 31953 19159
rect 31953 19125 31987 19159
rect 31987 19125 31996 19159
rect 31944 19116 31996 19125
rect 32404 19159 32456 19168
rect 32404 19125 32413 19159
rect 32413 19125 32447 19159
rect 32447 19125 32456 19159
rect 32404 19116 32456 19125
rect 36728 19116 36780 19168
rect 37648 19116 37700 19168
rect 37924 19116 37976 19168
rect 39212 19252 39264 19304
rect 40960 19252 41012 19304
rect 42432 19295 42484 19304
rect 42432 19261 42441 19295
rect 42441 19261 42475 19295
rect 42475 19261 42484 19295
rect 42432 19252 42484 19261
rect 43444 19252 43496 19304
rect 49148 19320 49200 19372
rect 49332 19363 49384 19372
rect 49332 19329 49341 19363
rect 49341 19329 49375 19363
rect 49375 19329 49384 19363
rect 49332 19320 49384 19329
rect 51908 19320 51960 19372
rect 44180 19295 44232 19304
rect 44180 19261 44189 19295
rect 44189 19261 44223 19295
rect 44223 19261 44232 19295
rect 44180 19252 44232 19261
rect 46296 19295 46348 19304
rect 46296 19261 46305 19295
rect 46305 19261 46339 19295
rect 46339 19261 46348 19295
rect 46296 19252 46348 19261
rect 46756 19295 46808 19304
rect 46756 19261 46765 19295
rect 46765 19261 46799 19295
rect 46799 19261 46808 19295
rect 46756 19252 46808 19261
rect 47768 19295 47820 19304
rect 47768 19261 47777 19295
rect 47777 19261 47811 19295
rect 47811 19261 47820 19295
rect 47768 19252 47820 19261
rect 49056 19295 49108 19304
rect 49056 19261 49065 19295
rect 49065 19261 49099 19295
rect 49099 19261 49108 19295
rect 49056 19252 49108 19261
rect 39856 19116 39908 19168
rect 41052 19159 41104 19168
rect 41052 19125 41061 19159
rect 41061 19125 41095 19159
rect 41095 19125 41104 19159
rect 41052 19116 41104 19125
rect 41880 19116 41932 19168
rect 42892 19116 42944 19168
rect 43260 19116 43312 19168
rect 44088 19184 44140 19236
rect 43536 19159 43588 19168
rect 43536 19125 43545 19159
rect 43545 19125 43579 19159
rect 43579 19125 43588 19159
rect 43536 19116 43588 19125
rect 44640 19116 44692 19168
rect 45836 19116 45888 19168
rect 46940 19116 46992 19168
rect 48136 19116 48188 19168
rect 48320 19159 48372 19168
rect 48320 19125 48329 19159
rect 48329 19125 48363 19159
rect 48363 19125 48372 19159
rect 48320 19116 48372 19125
rect 50068 19295 50120 19304
rect 50068 19261 50077 19295
rect 50077 19261 50111 19295
rect 50111 19261 50120 19295
rect 50068 19252 50120 19261
rect 49608 19227 49660 19236
rect 49608 19193 49617 19227
rect 49617 19193 49651 19227
rect 49651 19193 49660 19227
rect 49608 19184 49660 19193
rect 56048 19456 56100 19508
rect 58256 19456 58308 19508
rect 54576 19363 54628 19372
rect 54576 19329 54585 19363
rect 54585 19329 54619 19363
rect 54619 19329 54628 19363
rect 54576 19320 54628 19329
rect 55312 19320 55364 19372
rect 56324 19363 56376 19372
rect 56324 19329 56333 19363
rect 56333 19329 56367 19363
rect 56367 19329 56376 19363
rect 56324 19320 56376 19329
rect 57980 19320 58032 19372
rect 52368 19116 52420 19168
rect 52460 19159 52512 19168
rect 52460 19125 52469 19159
rect 52469 19125 52503 19159
rect 52503 19125 52512 19159
rect 52460 19116 52512 19125
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 22616 19014 22668 19066
rect 22680 19014 22732 19066
rect 22744 19014 22796 19066
rect 22808 19014 22860 19066
rect 22872 19014 22924 19066
rect 37060 19014 37112 19066
rect 37124 19014 37176 19066
rect 37188 19014 37240 19066
rect 37252 19014 37304 19066
rect 37316 19014 37368 19066
rect 51504 19014 51556 19066
rect 51568 19014 51620 19066
rect 51632 19014 51684 19066
rect 51696 19014 51748 19066
rect 51760 19014 51812 19066
rect 2780 18912 2832 18964
rect 5908 18912 5960 18964
rect 7932 18955 7984 18964
rect 7932 18921 7941 18955
rect 7941 18921 7975 18955
rect 7975 18921 7984 18955
rect 7932 18912 7984 18921
rect 9680 18955 9732 18964
rect 9680 18921 9689 18955
rect 9689 18921 9723 18955
rect 9723 18921 9732 18955
rect 9680 18912 9732 18921
rect 10232 18912 10284 18964
rect 12624 18912 12676 18964
rect 13084 18912 13136 18964
rect 14372 18912 14424 18964
rect 16396 18912 16448 18964
rect 6828 18844 6880 18896
rect 4804 18819 4856 18828
rect 4804 18785 4813 18819
rect 4813 18785 4847 18819
rect 4847 18785 4856 18819
rect 4804 18776 4856 18785
rect 6000 18776 6052 18828
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 7748 18776 7800 18828
rect 8576 18776 8628 18828
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 10416 18819 10468 18828
rect 10416 18785 10425 18819
rect 10425 18785 10459 18819
rect 10459 18785 10468 18819
rect 10416 18776 10468 18785
rect 17960 18912 18012 18964
rect 20536 18912 20588 18964
rect 21456 18912 21508 18964
rect 24952 18912 25004 18964
rect 26240 18912 26292 18964
rect 27160 18912 27212 18964
rect 27436 18912 27488 18964
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 16764 18819 16816 18828
rect 16764 18785 16773 18819
rect 16773 18785 16807 18819
rect 16807 18785 16816 18819
rect 16764 18776 16816 18785
rect 18144 18776 18196 18828
rect 4252 18683 4304 18692
rect 4252 18649 4261 18683
rect 4261 18649 4295 18683
rect 4295 18649 4304 18683
rect 7472 18683 7524 18692
rect 4252 18640 4304 18649
rect 7472 18649 7481 18683
rect 7481 18649 7515 18683
rect 7515 18649 7524 18683
rect 7472 18640 7524 18649
rect 5816 18572 5868 18624
rect 10876 18640 10928 18692
rect 12164 18708 12216 18760
rect 13820 18751 13872 18760
rect 13820 18717 13829 18751
rect 13829 18717 13863 18751
rect 13863 18717 13872 18751
rect 13820 18708 13872 18717
rect 19156 18708 19208 18760
rect 22468 18751 22520 18760
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 11060 18640 11112 18692
rect 11336 18640 11388 18692
rect 14096 18640 14148 18692
rect 19340 18640 19392 18692
rect 19708 18640 19760 18692
rect 21916 18640 21968 18692
rect 22192 18683 22244 18692
rect 22192 18649 22210 18683
rect 22210 18649 22244 18683
rect 22192 18640 22244 18649
rect 23020 18640 23072 18692
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 10232 18615 10284 18624
rect 10232 18581 10241 18615
rect 10241 18581 10275 18615
rect 10275 18581 10284 18615
rect 10232 18572 10284 18581
rect 10968 18572 11020 18624
rect 11704 18572 11756 18624
rect 12992 18572 13044 18624
rect 15200 18572 15252 18624
rect 15844 18572 15896 18624
rect 17132 18572 17184 18624
rect 22008 18572 22060 18624
rect 25596 18751 25648 18760
rect 25596 18717 25605 18751
rect 25605 18717 25639 18751
rect 25639 18717 25648 18751
rect 25596 18708 25648 18717
rect 26976 18708 27028 18760
rect 27160 18640 27212 18692
rect 25044 18615 25096 18624
rect 25044 18581 25053 18615
rect 25053 18581 25087 18615
rect 25087 18581 25096 18615
rect 25044 18572 25096 18581
rect 26240 18615 26292 18624
rect 26240 18581 26249 18615
rect 26249 18581 26283 18615
rect 26283 18581 26292 18615
rect 26240 18572 26292 18581
rect 26424 18572 26476 18624
rect 26516 18572 26568 18624
rect 27712 18708 27764 18760
rect 29644 18819 29696 18828
rect 29644 18785 29653 18819
rect 29653 18785 29687 18819
rect 29687 18785 29696 18819
rect 29644 18776 29696 18785
rect 29552 18708 29604 18760
rect 31300 18912 31352 18964
rect 32404 18912 32456 18964
rect 31852 18844 31904 18896
rect 34704 18912 34756 18964
rect 36912 18955 36964 18964
rect 36912 18921 36921 18955
rect 36921 18921 36955 18955
rect 36955 18921 36964 18955
rect 36912 18912 36964 18921
rect 37648 18912 37700 18964
rect 39212 18912 39264 18964
rect 40960 18912 41012 18964
rect 41972 18912 42024 18964
rect 42524 18912 42576 18964
rect 45836 18912 45888 18964
rect 46756 18912 46808 18964
rect 31944 18776 31996 18828
rect 32312 18751 32364 18760
rect 32312 18717 32321 18751
rect 32321 18717 32355 18751
rect 32355 18717 32364 18751
rect 32312 18708 32364 18717
rect 32772 18776 32824 18828
rect 32588 18751 32640 18760
rect 32588 18717 32597 18751
rect 32597 18717 32631 18751
rect 32631 18717 32640 18751
rect 32588 18708 32640 18717
rect 29644 18640 29696 18692
rect 31760 18640 31812 18692
rect 33416 18708 33468 18760
rect 33692 18819 33744 18828
rect 33692 18785 33701 18819
rect 33701 18785 33735 18819
rect 33735 18785 33744 18819
rect 33692 18776 33744 18785
rect 35256 18819 35308 18828
rect 35256 18785 35265 18819
rect 35265 18785 35299 18819
rect 35299 18785 35308 18819
rect 35256 18776 35308 18785
rect 35440 18776 35492 18828
rect 36728 18776 36780 18828
rect 37924 18776 37976 18828
rect 37740 18640 37792 18692
rect 27804 18615 27856 18624
rect 27804 18581 27813 18615
rect 27813 18581 27847 18615
rect 27847 18581 27856 18615
rect 27804 18572 27856 18581
rect 28816 18572 28868 18624
rect 30380 18572 30432 18624
rect 32864 18572 32916 18624
rect 36084 18615 36136 18624
rect 36084 18581 36093 18615
rect 36093 18581 36127 18615
rect 36127 18581 36136 18615
rect 36084 18572 36136 18581
rect 37280 18615 37332 18624
rect 37280 18581 37289 18615
rect 37289 18581 37323 18615
rect 37323 18581 37332 18615
rect 37280 18572 37332 18581
rect 37464 18572 37516 18624
rect 38660 18708 38712 18760
rect 39948 18708 40000 18760
rect 41052 18776 41104 18828
rect 41880 18776 41932 18828
rect 43352 18776 43404 18828
rect 40224 18751 40276 18760
rect 40224 18717 40233 18751
rect 40233 18717 40267 18751
rect 40267 18717 40276 18751
rect 40224 18708 40276 18717
rect 42892 18708 42944 18760
rect 44088 18819 44140 18828
rect 44088 18785 44097 18819
rect 44097 18785 44131 18819
rect 44131 18785 44140 18819
rect 44088 18776 44140 18785
rect 44640 18776 44692 18828
rect 43720 18751 43772 18760
rect 43720 18717 43738 18751
rect 43738 18717 43772 18751
rect 43720 18708 43772 18717
rect 43812 18751 43864 18760
rect 43812 18717 43821 18751
rect 43821 18717 43855 18751
rect 43855 18717 43864 18751
rect 43812 18708 43864 18717
rect 45376 18708 45428 18760
rect 38476 18640 38528 18692
rect 38936 18640 38988 18692
rect 45008 18683 45060 18692
rect 45008 18649 45017 18683
rect 45017 18649 45051 18683
rect 45051 18649 45060 18683
rect 48228 18912 48280 18964
rect 48872 18912 48924 18964
rect 49700 18912 49752 18964
rect 50068 18912 50120 18964
rect 48136 18776 48188 18828
rect 48320 18708 48372 18760
rect 45008 18640 45060 18649
rect 39856 18572 39908 18624
rect 40132 18615 40184 18624
rect 40132 18581 40141 18615
rect 40141 18581 40175 18615
rect 40175 18581 40184 18615
rect 40132 18572 40184 18581
rect 42616 18572 42668 18624
rect 44180 18572 44232 18624
rect 45284 18572 45336 18624
rect 49056 18683 49108 18692
rect 49056 18649 49065 18683
rect 49065 18649 49099 18683
rect 49099 18649 49108 18683
rect 49056 18640 49108 18649
rect 51908 18708 51960 18760
rect 47400 18572 47452 18624
rect 51172 18640 51224 18692
rect 51632 18640 51684 18692
rect 52736 18640 52788 18692
rect 54208 18912 54260 18964
rect 53656 18844 53708 18896
rect 54484 18844 54536 18896
rect 55220 18776 55272 18828
rect 54392 18708 54444 18760
rect 56140 18912 56192 18964
rect 57336 18912 57388 18964
rect 57520 18912 57572 18964
rect 58256 18819 58308 18828
rect 58256 18785 58265 18819
rect 58265 18785 58299 18819
rect 58299 18785 58308 18819
rect 58256 18776 58308 18785
rect 57244 18708 57296 18760
rect 53196 18615 53248 18624
rect 53196 18581 53205 18615
rect 53205 18581 53239 18615
rect 53239 18581 53248 18615
rect 53196 18572 53248 18581
rect 53288 18615 53340 18624
rect 53288 18581 53297 18615
rect 53297 18581 53331 18615
rect 53331 18581 53340 18615
rect 53288 18572 53340 18581
rect 53748 18615 53800 18624
rect 53748 18581 53757 18615
rect 53757 18581 53791 18615
rect 53791 18581 53800 18615
rect 53748 18572 53800 18581
rect 54668 18572 54720 18624
rect 57612 18572 57664 18624
rect 15394 18470 15446 18522
rect 15458 18470 15510 18522
rect 15522 18470 15574 18522
rect 15586 18470 15638 18522
rect 15650 18470 15702 18522
rect 29838 18470 29890 18522
rect 29902 18470 29954 18522
rect 29966 18470 30018 18522
rect 30030 18470 30082 18522
rect 30094 18470 30146 18522
rect 44282 18470 44334 18522
rect 44346 18470 44398 18522
rect 44410 18470 44462 18522
rect 44474 18470 44526 18522
rect 44538 18470 44590 18522
rect 58726 18470 58778 18522
rect 58790 18470 58842 18522
rect 58854 18470 58906 18522
rect 58918 18470 58970 18522
rect 58982 18470 59034 18522
rect 4804 18368 4856 18420
rect 7472 18368 7524 18420
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 11060 18368 11112 18420
rect 13912 18368 13964 18420
rect 19156 18368 19208 18420
rect 20812 18368 20864 18420
rect 21088 18411 21140 18420
rect 21088 18377 21097 18411
rect 21097 18377 21131 18411
rect 21131 18377 21140 18411
rect 21088 18368 21140 18377
rect 21180 18368 21232 18420
rect 6460 18232 6512 18284
rect 6920 18232 6972 18284
rect 7748 18232 7800 18284
rect 9128 18232 9180 18284
rect 9772 18232 9824 18284
rect 10968 18232 11020 18284
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 11888 18232 11940 18284
rect 20720 18300 20772 18352
rect 22100 18300 22152 18352
rect 19708 18232 19760 18284
rect 21732 18232 21784 18284
rect 11244 18207 11296 18216
rect 11244 18173 11253 18207
rect 11253 18173 11287 18207
rect 11287 18173 11296 18207
rect 11244 18164 11296 18173
rect 12072 18164 12124 18216
rect 12532 18207 12584 18216
rect 12532 18173 12566 18207
rect 12566 18173 12584 18207
rect 12532 18164 12584 18173
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 16396 18164 16448 18216
rect 20996 18164 21048 18216
rect 22008 18164 22060 18216
rect 22560 18164 22612 18216
rect 23020 18164 23072 18216
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 11060 18096 11112 18148
rect 12256 18096 12308 18148
rect 13728 18096 13780 18148
rect 21916 18096 21968 18148
rect 9864 18028 9916 18080
rect 14096 18028 14148 18080
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 20720 18028 20772 18080
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 22468 18028 22520 18080
rect 23388 18028 23440 18080
rect 24860 18232 24912 18284
rect 25044 18343 25096 18352
rect 25044 18309 25078 18343
rect 25078 18309 25096 18343
rect 27988 18368 28040 18420
rect 28172 18368 28224 18420
rect 25044 18300 25096 18309
rect 28816 18343 28868 18352
rect 28816 18309 28825 18343
rect 28825 18309 28859 18343
rect 28859 18309 28868 18343
rect 28816 18300 28868 18309
rect 29644 18368 29696 18420
rect 26240 18232 26292 18284
rect 27068 18232 27120 18284
rect 26884 18164 26936 18216
rect 27160 18207 27212 18216
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 29828 18343 29880 18352
rect 29828 18309 29862 18343
rect 29862 18309 29880 18343
rect 29828 18300 29880 18309
rect 30196 18368 30248 18420
rect 31944 18368 31996 18420
rect 32864 18368 32916 18420
rect 35992 18411 36044 18420
rect 35992 18377 36001 18411
rect 36001 18377 36035 18411
rect 36035 18377 36044 18411
rect 35992 18368 36044 18377
rect 36084 18368 36136 18420
rect 37924 18411 37976 18420
rect 37924 18377 37933 18411
rect 37933 18377 37967 18411
rect 37967 18377 37976 18411
rect 37924 18368 37976 18377
rect 38476 18411 38528 18420
rect 38476 18377 38485 18411
rect 38485 18377 38519 18411
rect 38519 18377 38528 18411
rect 38476 18368 38528 18377
rect 38936 18368 38988 18420
rect 39028 18368 39080 18420
rect 39580 18368 39632 18420
rect 32036 18300 32088 18352
rect 27988 18207 28040 18216
rect 27988 18173 28022 18207
rect 28022 18173 28040 18207
rect 27988 18164 28040 18173
rect 28356 18164 28408 18216
rect 26148 18071 26200 18080
rect 26148 18037 26157 18071
rect 26157 18037 26191 18071
rect 26191 18037 26200 18071
rect 26148 18028 26200 18037
rect 27620 18139 27672 18148
rect 27620 18105 27629 18139
rect 27629 18105 27663 18139
rect 27663 18105 27672 18139
rect 27620 18096 27672 18105
rect 29000 18096 29052 18148
rect 31484 18207 31536 18216
rect 31484 18173 31493 18207
rect 31493 18173 31527 18207
rect 31527 18173 31536 18207
rect 31484 18164 31536 18173
rect 31576 18207 31628 18216
rect 31576 18173 31585 18207
rect 31585 18173 31619 18207
rect 31619 18173 31628 18207
rect 31576 18164 31628 18173
rect 31392 18096 31444 18148
rect 31944 18232 31996 18284
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32128 18232 32180 18241
rect 33140 18232 33192 18284
rect 33416 18232 33468 18284
rect 33508 18232 33560 18284
rect 37280 18300 37332 18352
rect 34520 18164 34572 18216
rect 36728 18232 36780 18284
rect 37556 18232 37608 18284
rect 38844 18232 38896 18284
rect 39856 18275 39908 18284
rect 39856 18241 39865 18275
rect 39865 18241 39899 18275
rect 39899 18241 39908 18275
rect 39856 18232 39908 18241
rect 42432 18368 42484 18420
rect 41420 18300 41472 18352
rect 42708 18300 42760 18352
rect 40868 18275 40920 18284
rect 40868 18241 40877 18275
rect 40877 18241 40911 18275
rect 40911 18241 40920 18275
rect 40868 18232 40920 18241
rect 45008 18368 45060 18420
rect 46296 18368 46348 18420
rect 47768 18411 47820 18420
rect 47768 18377 47777 18411
rect 47777 18377 47811 18411
rect 47811 18377 47820 18411
rect 47768 18368 47820 18377
rect 50068 18368 50120 18420
rect 51632 18411 51684 18420
rect 51632 18377 51641 18411
rect 51641 18377 51675 18411
rect 51675 18377 51684 18411
rect 51632 18368 51684 18377
rect 52736 18411 52788 18420
rect 52736 18377 52745 18411
rect 52745 18377 52779 18411
rect 52779 18377 52788 18411
rect 52736 18368 52788 18377
rect 53288 18368 53340 18420
rect 53748 18368 53800 18420
rect 43536 18300 43588 18352
rect 45284 18300 45336 18352
rect 43628 18232 43680 18284
rect 28172 18028 28224 18080
rect 32036 18096 32088 18148
rect 42524 18207 42576 18216
rect 42524 18173 42533 18207
rect 42533 18173 42567 18207
rect 42567 18173 42576 18207
rect 42524 18164 42576 18173
rect 44824 18232 44876 18284
rect 35716 18096 35768 18148
rect 39764 18096 39816 18148
rect 42800 18096 42852 18148
rect 32772 18028 32824 18080
rect 33600 18071 33652 18080
rect 33600 18037 33609 18071
rect 33609 18037 33643 18071
rect 33643 18037 33652 18071
rect 33600 18028 33652 18037
rect 33692 18028 33744 18080
rect 39948 18028 40000 18080
rect 43168 18071 43220 18080
rect 43168 18037 43177 18071
rect 43177 18037 43211 18071
rect 43211 18037 43220 18071
rect 43168 18028 43220 18037
rect 44088 18028 44140 18080
rect 47308 18028 47360 18080
rect 47952 18028 48004 18080
rect 49608 18028 49660 18080
rect 49700 18071 49752 18080
rect 49700 18037 49709 18071
rect 49709 18037 49743 18071
rect 49743 18037 49752 18071
rect 49700 18028 49752 18037
rect 49884 18028 49936 18080
rect 52828 18164 52880 18216
rect 53196 18164 53248 18216
rect 58072 18164 58124 18216
rect 52644 18028 52696 18080
rect 53656 18028 53708 18080
rect 54484 18071 54536 18080
rect 54484 18037 54493 18071
rect 54493 18037 54527 18071
rect 54527 18037 54536 18071
rect 54484 18028 54536 18037
rect 57888 18071 57940 18080
rect 57888 18037 57897 18071
rect 57897 18037 57931 18071
rect 57931 18037 57940 18071
rect 57888 18028 57940 18037
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 22616 17926 22668 17978
rect 22680 17926 22732 17978
rect 22744 17926 22796 17978
rect 22808 17926 22860 17978
rect 22872 17926 22924 17978
rect 37060 17926 37112 17978
rect 37124 17926 37176 17978
rect 37188 17926 37240 17978
rect 37252 17926 37304 17978
rect 37316 17926 37368 17978
rect 51504 17926 51556 17978
rect 51568 17926 51620 17978
rect 51632 17926 51684 17978
rect 51696 17926 51748 17978
rect 51760 17926 51812 17978
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 6828 17756 6880 17808
rect 7380 17756 7432 17808
rect 11060 17824 11112 17876
rect 11244 17867 11296 17876
rect 11244 17833 11253 17867
rect 11253 17833 11287 17867
rect 11287 17833 11296 17867
rect 11244 17824 11296 17833
rect 13820 17824 13872 17876
rect 16764 17824 16816 17876
rect 19708 17824 19760 17876
rect 22192 17824 22244 17876
rect 22468 17824 22520 17876
rect 24860 17824 24912 17876
rect 25320 17867 25372 17876
rect 25320 17833 25329 17867
rect 25329 17833 25363 17867
rect 25363 17833 25372 17867
rect 25320 17824 25372 17833
rect 25596 17824 25648 17876
rect 10968 17756 11020 17808
rect 27896 17824 27948 17876
rect 28080 17824 28132 17876
rect 28172 17824 28224 17876
rect 33140 17824 33192 17876
rect 33508 17824 33560 17876
rect 7840 17688 7892 17740
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 11336 17688 11388 17740
rect 11888 17688 11940 17740
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 20720 17731 20772 17740
rect 20720 17697 20729 17731
rect 20729 17697 20763 17731
rect 20763 17697 20772 17731
rect 20720 17688 20772 17697
rect 3516 17663 3568 17672
rect 3516 17629 3525 17663
rect 3525 17629 3559 17663
rect 3559 17629 3568 17663
rect 3516 17620 3568 17629
rect 3792 17663 3844 17672
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 9588 17552 9640 17604
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 4252 17484 4304 17536
rect 8392 17484 8444 17536
rect 12440 17552 12492 17604
rect 15292 17620 15344 17672
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 16212 17620 16264 17672
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 12164 17484 12216 17536
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 17224 17484 17276 17536
rect 17776 17484 17828 17536
rect 18052 17484 18104 17536
rect 20720 17484 20772 17536
rect 20996 17527 21048 17536
rect 20996 17493 21005 17527
rect 21005 17493 21039 17527
rect 21039 17493 21048 17527
rect 20996 17484 21048 17493
rect 21824 17688 21876 17740
rect 34520 17867 34572 17876
rect 34520 17833 34529 17867
rect 34529 17833 34563 17867
rect 34563 17833 34572 17867
rect 34520 17824 34572 17833
rect 35716 17824 35768 17876
rect 40868 17824 40920 17876
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 26056 17620 26108 17672
rect 32680 17731 32732 17740
rect 32680 17697 32689 17731
rect 32689 17697 32723 17731
rect 32723 17697 32732 17731
rect 32680 17688 32732 17697
rect 33416 17688 33468 17740
rect 27528 17620 27580 17672
rect 31944 17620 31996 17672
rect 34244 17688 34296 17740
rect 36084 17620 36136 17672
rect 38108 17688 38160 17740
rect 53656 17824 53708 17876
rect 57060 17824 57112 17876
rect 43812 17756 43864 17808
rect 53472 17756 53524 17808
rect 43168 17688 43220 17740
rect 44180 17688 44232 17740
rect 54576 17688 54628 17740
rect 44732 17620 44784 17672
rect 53012 17663 53064 17672
rect 53012 17629 53021 17663
rect 53021 17629 53055 17663
rect 53055 17629 53064 17663
rect 53012 17620 53064 17629
rect 53104 17663 53156 17672
rect 53104 17629 53113 17663
rect 53113 17629 53147 17663
rect 53147 17629 53156 17663
rect 53104 17620 53156 17629
rect 53840 17620 53892 17672
rect 55864 17663 55916 17672
rect 55864 17629 55873 17663
rect 55873 17629 55907 17663
rect 55907 17629 55916 17663
rect 55864 17620 55916 17629
rect 56048 17663 56100 17672
rect 56048 17629 56057 17663
rect 56057 17629 56091 17663
rect 56091 17629 56100 17663
rect 56048 17620 56100 17629
rect 27896 17552 27948 17604
rect 21732 17484 21784 17536
rect 24400 17527 24452 17536
rect 24400 17493 24409 17527
rect 24409 17493 24443 17527
rect 24443 17493 24452 17527
rect 24400 17484 24452 17493
rect 24584 17484 24636 17536
rect 25872 17527 25924 17536
rect 25872 17493 25881 17527
rect 25881 17493 25915 17527
rect 25915 17493 25924 17527
rect 25872 17484 25924 17493
rect 26424 17484 26476 17536
rect 29000 17484 29052 17536
rect 37832 17552 37884 17604
rect 41144 17552 41196 17604
rect 57520 17552 57572 17604
rect 30380 17484 30432 17536
rect 32772 17484 32824 17536
rect 35808 17527 35860 17536
rect 35808 17493 35817 17527
rect 35817 17493 35851 17527
rect 35851 17493 35860 17527
rect 35808 17484 35860 17493
rect 37464 17527 37516 17536
rect 37464 17493 37473 17527
rect 37473 17493 37507 17527
rect 37507 17493 37516 17527
rect 37464 17484 37516 17493
rect 43996 17527 44048 17536
rect 43996 17493 44005 17527
rect 44005 17493 44039 17527
rect 44039 17493 44048 17527
rect 43996 17484 44048 17493
rect 52184 17527 52236 17536
rect 52184 17493 52193 17527
rect 52193 17493 52227 17527
rect 52227 17493 52236 17527
rect 52184 17484 52236 17493
rect 52368 17527 52420 17536
rect 52368 17493 52377 17527
rect 52377 17493 52411 17527
rect 52411 17493 52420 17527
rect 52368 17484 52420 17493
rect 53656 17484 53708 17536
rect 55312 17527 55364 17536
rect 55312 17493 55321 17527
rect 55321 17493 55355 17527
rect 55355 17493 55364 17527
rect 55312 17484 55364 17493
rect 56600 17484 56652 17536
rect 58256 17527 58308 17536
rect 58256 17493 58265 17527
rect 58265 17493 58299 17527
rect 58299 17493 58308 17527
rect 58256 17484 58308 17493
rect 15394 17382 15446 17434
rect 15458 17382 15510 17434
rect 15522 17382 15574 17434
rect 15586 17382 15638 17434
rect 15650 17382 15702 17434
rect 29838 17382 29890 17434
rect 29902 17382 29954 17434
rect 29966 17382 30018 17434
rect 30030 17382 30082 17434
rect 30094 17382 30146 17434
rect 44282 17382 44334 17434
rect 44346 17382 44398 17434
rect 44410 17382 44462 17434
rect 44474 17382 44526 17434
rect 44538 17382 44590 17434
rect 58726 17382 58778 17434
rect 58790 17382 58842 17434
rect 58854 17382 58906 17434
rect 58918 17382 58970 17434
rect 58982 17382 59034 17434
rect 2964 17280 3016 17332
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 9864 17280 9916 17332
rect 10324 17280 10376 17332
rect 10508 17280 10560 17332
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 15292 17323 15344 17332
rect 15292 17289 15301 17323
rect 15301 17289 15335 17323
rect 15335 17289 15344 17323
rect 15292 17280 15344 17289
rect 16948 17280 17000 17332
rect 19340 17280 19392 17332
rect 20536 17280 20588 17332
rect 22376 17280 22428 17332
rect 24400 17280 24452 17332
rect 25872 17280 25924 17332
rect 27988 17280 28040 17332
rect 31576 17280 31628 17332
rect 31760 17280 31812 17332
rect 32680 17280 32732 17332
rect 33508 17280 33560 17332
rect 35808 17280 35860 17332
rect 42800 17323 42852 17332
rect 42800 17289 42809 17323
rect 42809 17289 42843 17323
rect 42843 17289 42852 17323
rect 42800 17280 42852 17289
rect 52368 17280 52420 17332
rect 53104 17280 53156 17332
rect 53472 17280 53524 17332
rect 55312 17280 55364 17332
rect 56048 17280 56100 17332
rect 8392 17255 8444 17264
rect 8392 17221 8401 17255
rect 8401 17221 8435 17255
rect 8435 17221 8444 17255
rect 8392 17212 8444 17221
rect 6460 17144 6512 17196
rect 6920 17187 6972 17196
rect 6920 17153 6954 17187
rect 6954 17153 6972 17187
rect 6920 17144 6972 17153
rect 1584 17076 1636 17128
rect 2412 17119 2464 17128
rect 2412 17085 2421 17119
rect 2421 17085 2455 17119
rect 2455 17085 2464 17119
rect 2412 17076 2464 17085
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 12532 17212 12584 17264
rect 15844 17212 15896 17264
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 17224 17144 17276 17196
rect 19248 17144 19300 17196
rect 23388 17187 23440 17196
rect 23388 17153 23397 17187
rect 23397 17153 23431 17187
rect 23431 17153 23440 17187
rect 23388 17144 23440 17153
rect 28080 17212 28132 17264
rect 29000 17255 29052 17264
rect 29000 17221 29009 17255
rect 29009 17221 29043 17255
rect 29043 17221 29052 17255
rect 29000 17212 29052 17221
rect 26056 17144 26108 17196
rect 26148 17187 26200 17196
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 15016 17076 15068 17128
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 20904 17119 20956 17128
rect 20904 17085 20913 17119
rect 20913 17085 20947 17119
rect 20947 17085 20956 17119
rect 20904 17076 20956 17085
rect 22376 17119 22428 17128
rect 22376 17085 22385 17119
rect 22385 17085 22419 17119
rect 22419 17085 22428 17119
rect 22376 17076 22428 17085
rect 12164 17008 12216 17060
rect 16304 17051 16356 17060
rect 16304 17017 16313 17051
rect 16313 17017 16347 17051
rect 16347 17017 16356 17051
rect 16304 17008 16356 17017
rect 4528 16983 4580 16992
rect 4528 16949 4537 16983
rect 4537 16949 4571 16983
rect 4571 16949 4580 16983
rect 4528 16940 4580 16949
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11796 16940 11848 16992
rect 12716 16940 12768 16992
rect 15016 16940 15068 16992
rect 15200 16983 15252 16992
rect 15200 16949 15209 16983
rect 15209 16949 15243 16983
rect 15243 16949 15252 16983
rect 15200 16940 15252 16949
rect 21088 17008 21140 17060
rect 21732 17008 21784 17060
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 27620 17076 27672 17128
rect 28172 17076 28224 17128
rect 27896 17008 27948 17060
rect 31668 17144 31720 17196
rect 31944 17076 31996 17128
rect 33784 17144 33836 17196
rect 35256 17144 35308 17196
rect 44088 17212 44140 17264
rect 37924 17119 37976 17128
rect 37924 17085 37933 17119
rect 37933 17085 37967 17119
rect 37967 17085 37976 17119
rect 37924 17076 37976 17085
rect 38660 17119 38712 17128
rect 38660 17085 38669 17119
rect 38669 17085 38703 17119
rect 38703 17085 38712 17119
rect 38660 17076 38712 17085
rect 22192 16940 22244 16992
rect 24400 16940 24452 16992
rect 24860 16983 24912 16992
rect 24860 16949 24869 16983
rect 24869 16949 24903 16983
rect 24903 16949 24912 16983
rect 24860 16940 24912 16949
rect 25044 16940 25096 16992
rect 27252 16983 27304 16992
rect 27252 16949 27261 16983
rect 27261 16949 27295 16983
rect 27295 16949 27304 16983
rect 27252 16940 27304 16949
rect 27712 16940 27764 16992
rect 32956 16983 33008 16992
rect 32956 16949 32965 16983
rect 32965 16949 32999 16983
rect 32999 16949 33008 16983
rect 32956 16940 33008 16949
rect 33784 16983 33836 16992
rect 33784 16949 33793 16983
rect 33793 16949 33827 16983
rect 33827 16949 33836 16983
rect 34520 16983 34572 16992
rect 33784 16940 33836 16949
rect 34520 16949 34529 16983
rect 34529 16949 34563 16983
rect 34563 16949 34572 16983
rect 34520 16940 34572 16949
rect 35808 16983 35860 16992
rect 35808 16949 35817 16983
rect 35817 16949 35851 16983
rect 35851 16949 35860 16983
rect 35808 16940 35860 16949
rect 36176 16940 36228 16992
rect 37464 17008 37516 17060
rect 43812 17144 43864 17196
rect 48136 17187 48188 17196
rect 48136 17153 48145 17187
rect 48145 17153 48179 17187
rect 48179 17153 48188 17187
rect 48136 17144 48188 17153
rect 51172 17187 51224 17196
rect 51172 17153 51181 17187
rect 51181 17153 51215 17187
rect 51215 17153 51224 17187
rect 51172 17144 51224 17153
rect 52644 17212 52696 17264
rect 54576 17187 54628 17196
rect 54576 17153 54585 17187
rect 54585 17153 54619 17187
rect 54619 17153 54628 17187
rect 54576 17144 54628 17153
rect 40040 17119 40092 17128
rect 40040 17085 40049 17119
rect 40049 17085 40083 17119
rect 40083 17085 40092 17119
rect 40040 17076 40092 17085
rect 40224 17076 40276 17128
rect 44180 17119 44232 17128
rect 44180 17085 44189 17119
rect 44189 17085 44223 17119
rect 44223 17085 44232 17119
rect 44180 17076 44232 17085
rect 40316 17008 40368 17060
rect 50896 17119 50948 17128
rect 50896 17085 50905 17119
rect 50905 17085 50939 17119
rect 50939 17085 50948 17119
rect 50896 17076 50948 17085
rect 52184 17076 52236 17128
rect 52920 17076 52972 17128
rect 57428 17280 57480 17332
rect 57888 17212 57940 17264
rect 56876 17187 56928 17196
rect 56876 17153 56885 17187
rect 56885 17153 56919 17187
rect 56919 17153 56928 17187
rect 56876 17144 56928 17153
rect 57336 17008 57388 17060
rect 37556 16940 37608 16992
rect 38016 16983 38068 16992
rect 38016 16949 38025 16983
rect 38025 16949 38059 16983
rect 38059 16949 38068 16983
rect 38016 16940 38068 16949
rect 40684 16983 40736 16992
rect 40684 16949 40693 16983
rect 40693 16949 40727 16983
rect 40727 16949 40736 16983
rect 40684 16940 40736 16949
rect 43536 16983 43588 16992
rect 43536 16949 43545 16983
rect 43545 16949 43579 16983
rect 43579 16949 43588 16983
rect 43536 16940 43588 16949
rect 50252 16983 50304 16992
rect 50252 16949 50261 16983
rect 50261 16949 50295 16983
rect 50295 16949 50304 16983
rect 50252 16940 50304 16949
rect 53564 16983 53616 16992
rect 53564 16949 53573 16983
rect 53573 16949 53607 16983
rect 53607 16949 53616 16983
rect 53564 16940 53616 16949
rect 56324 16983 56376 16992
rect 56324 16949 56333 16983
rect 56333 16949 56367 16983
rect 56367 16949 56376 16983
rect 56324 16940 56376 16949
rect 56508 16940 56560 16992
rect 56784 16940 56836 16992
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 22616 16838 22668 16890
rect 22680 16838 22732 16890
rect 22744 16838 22796 16890
rect 22808 16838 22860 16890
rect 22872 16838 22924 16890
rect 37060 16838 37112 16890
rect 37124 16838 37176 16890
rect 37188 16838 37240 16890
rect 37252 16838 37304 16890
rect 37316 16838 37368 16890
rect 51504 16838 51556 16890
rect 51568 16838 51620 16890
rect 51632 16838 51684 16890
rect 51696 16838 51748 16890
rect 51760 16838 51812 16890
rect 3884 16711 3936 16720
rect 3884 16677 3893 16711
rect 3893 16677 3927 16711
rect 3927 16677 3936 16711
rect 3884 16668 3936 16677
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 6920 16736 6972 16788
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 9588 16779 9640 16788
rect 9588 16745 9597 16779
rect 9597 16745 9631 16779
rect 9631 16745 9640 16779
rect 9588 16736 9640 16745
rect 11796 16736 11848 16788
rect 15936 16779 15988 16788
rect 15936 16745 15945 16779
rect 15945 16745 15979 16779
rect 15979 16745 15988 16779
rect 15936 16736 15988 16745
rect 18144 16736 18196 16788
rect 18880 16736 18932 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 22376 16736 22428 16788
rect 22468 16736 22520 16788
rect 22836 16736 22888 16788
rect 24860 16736 24912 16788
rect 27620 16736 27672 16788
rect 27712 16736 27764 16788
rect 27896 16736 27948 16788
rect 28080 16736 28132 16788
rect 30380 16736 30432 16788
rect 3332 16532 3384 16584
rect 2504 16464 2556 16516
rect 4896 16464 4948 16516
rect 2964 16439 3016 16448
rect 2964 16405 2973 16439
rect 2973 16405 3007 16439
rect 3007 16405 3016 16439
rect 2964 16396 3016 16405
rect 3056 16439 3108 16448
rect 3056 16405 3065 16439
rect 3065 16405 3099 16439
rect 3099 16405 3108 16439
rect 3056 16396 3108 16405
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 4620 16396 4672 16448
rect 5540 16396 5592 16448
rect 6828 16396 6880 16448
rect 7472 16532 7524 16584
rect 8208 16464 8260 16516
rect 17868 16668 17920 16720
rect 9772 16600 9824 16652
rect 16304 16600 16356 16652
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 17592 16600 17644 16652
rect 18236 16600 18288 16652
rect 14280 16532 14332 16584
rect 15108 16532 15160 16584
rect 17040 16532 17092 16584
rect 17776 16532 17828 16584
rect 18420 16532 18472 16584
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 22192 16600 22244 16652
rect 22560 16668 22612 16720
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 20812 16532 20864 16584
rect 22928 16532 22980 16584
rect 24492 16532 24544 16584
rect 25320 16600 25372 16652
rect 33140 16600 33192 16652
rect 33692 16600 33744 16652
rect 34520 16600 34572 16652
rect 35348 16736 35400 16788
rect 36176 16736 36228 16788
rect 37464 16736 37516 16788
rect 36084 16711 36136 16720
rect 36084 16677 36093 16711
rect 36093 16677 36127 16711
rect 36127 16677 36136 16711
rect 36084 16668 36136 16677
rect 40040 16643 40092 16652
rect 40040 16609 40049 16643
rect 40049 16609 40083 16643
rect 40083 16609 40092 16643
rect 40040 16600 40092 16609
rect 40684 16736 40736 16788
rect 41420 16643 41472 16652
rect 41420 16609 41429 16643
rect 41429 16609 41463 16643
rect 41463 16609 41472 16643
rect 41420 16600 41472 16609
rect 45192 16736 45244 16788
rect 48136 16736 48188 16788
rect 50896 16736 50948 16788
rect 53012 16736 53064 16788
rect 55864 16736 55916 16788
rect 56600 16736 56652 16788
rect 56784 16736 56836 16788
rect 56876 16736 56928 16788
rect 18604 16507 18656 16516
rect 18604 16473 18613 16507
rect 18613 16473 18647 16507
rect 18647 16473 18656 16507
rect 18604 16464 18656 16473
rect 21180 16464 21232 16516
rect 24584 16464 24636 16516
rect 26056 16532 26108 16584
rect 24952 16464 25004 16516
rect 25964 16464 26016 16516
rect 27804 16464 27856 16516
rect 28724 16575 28776 16584
rect 28724 16541 28733 16575
rect 28733 16541 28767 16575
rect 28767 16541 28776 16575
rect 28724 16532 28776 16541
rect 30196 16575 30248 16584
rect 30196 16541 30205 16575
rect 30205 16541 30239 16575
rect 30239 16541 30248 16575
rect 30196 16532 30248 16541
rect 31760 16532 31812 16584
rect 32128 16575 32180 16584
rect 32128 16541 32137 16575
rect 32137 16541 32171 16575
rect 32171 16541 32180 16575
rect 32128 16532 32180 16541
rect 29460 16464 29512 16516
rect 29552 16507 29604 16516
rect 29552 16473 29561 16507
rect 29561 16473 29595 16507
rect 29595 16473 29604 16507
rect 34152 16575 34204 16584
rect 34152 16541 34161 16575
rect 34161 16541 34195 16575
rect 34195 16541 34204 16575
rect 34152 16532 34204 16541
rect 35808 16532 35860 16584
rect 37556 16532 37608 16584
rect 29552 16464 29604 16473
rect 19984 16439 20036 16448
rect 19984 16405 19993 16439
rect 19993 16405 20027 16439
rect 20027 16405 20036 16439
rect 19984 16396 20036 16405
rect 21272 16396 21324 16448
rect 22192 16439 22244 16448
rect 22192 16405 22201 16439
rect 22201 16405 22235 16439
rect 22235 16405 22244 16439
rect 22192 16396 22244 16405
rect 22560 16396 22612 16448
rect 22744 16396 22796 16448
rect 23112 16439 23164 16448
rect 23112 16405 23121 16439
rect 23121 16405 23155 16439
rect 23155 16405 23164 16439
rect 23112 16396 23164 16405
rect 23296 16396 23348 16448
rect 37464 16464 37516 16516
rect 26884 16439 26936 16448
rect 26884 16405 26893 16439
rect 26893 16405 26927 16439
rect 26927 16405 26936 16439
rect 26884 16396 26936 16405
rect 29368 16439 29420 16448
rect 29368 16405 29377 16439
rect 29377 16405 29411 16439
rect 29411 16405 29420 16439
rect 29368 16396 29420 16405
rect 31300 16439 31352 16448
rect 31300 16405 31309 16439
rect 31309 16405 31343 16439
rect 31343 16405 31352 16439
rect 31300 16396 31352 16405
rect 31392 16396 31444 16448
rect 31484 16439 31536 16448
rect 31484 16405 31493 16439
rect 31493 16405 31527 16439
rect 31527 16405 31536 16439
rect 31484 16396 31536 16405
rect 33600 16439 33652 16448
rect 33600 16405 33609 16439
rect 33609 16405 33643 16439
rect 33643 16405 33652 16439
rect 33600 16396 33652 16405
rect 38660 16464 38712 16516
rect 38936 16464 38988 16516
rect 40592 16532 40644 16584
rect 42156 16532 42208 16584
rect 49056 16600 49108 16652
rect 50160 16600 50212 16652
rect 51172 16600 51224 16652
rect 51724 16643 51776 16652
rect 51724 16609 51733 16643
rect 51733 16609 51767 16643
rect 51767 16609 51776 16643
rect 51724 16600 51776 16609
rect 53656 16643 53708 16652
rect 53656 16609 53665 16643
rect 53665 16609 53699 16643
rect 53699 16609 53708 16643
rect 53656 16600 53708 16609
rect 53748 16643 53800 16652
rect 53748 16609 53757 16643
rect 53757 16609 53791 16643
rect 53791 16609 53800 16643
rect 53748 16600 53800 16609
rect 53840 16600 53892 16652
rect 54208 16600 54260 16652
rect 43536 16532 43588 16584
rect 47676 16575 47728 16584
rect 47676 16541 47685 16575
rect 47685 16541 47719 16575
rect 47719 16541 47728 16575
rect 47676 16532 47728 16541
rect 37648 16439 37700 16448
rect 37648 16405 37657 16439
rect 37657 16405 37691 16439
rect 37691 16405 37700 16439
rect 37648 16396 37700 16405
rect 39028 16396 39080 16448
rect 40684 16439 40736 16448
rect 40684 16405 40693 16439
rect 40693 16405 40727 16439
rect 40727 16405 40736 16439
rect 40684 16396 40736 16405
rect 42340 16439 42392 16448
rect 42340 16405 42349 16439
rect 42349 16405 42383 16439
rect 42383 16405 42392 16439
rect 42340 16396 42392 16405
rect 43168 16396 43220 16448
rect 45008 16396 45060 16448
rect 47032 16439 47084 16448
rect 47032 16405 47041 16439
rect 47041 16405 47075 16439
rect 47075 16405 47084 16439
rect 47032 16396 47084 16405
rect 50988 16575 51040 16584
rect 50988 16541 50997 16575
rect 50997 16541 51031 16575
rect 51031 16541 51040 16575
rect 50988 16532 51040 16541
rect 53564 16532 53616 16584
rect 52368 16464 52420 16516
rect 56784 16600 56836 16652
rect 57888 16600 57940 16652
rect 58164 16643 58216 16652
rect 58164 16609 58173 16643
rect 58173 16609 58207 16643
rect 58207 16609 58216 16643
rect 58164 16600 58216 16609
rect 56324 16575 56376 16584
rect 56324 16541 56333 16575
rect 56333 16541 56367 16575
rect 56367 16541 56376 16575
rect 56324 16532 56376 16541
rect 56416 16532 56468 16584
rect 56600 16575 56652 16584
rect 56600 16541 56609 16575
rect 56609 16541 56643 16575
rect 56643 16541 56652 16575
rect 56600 16532 56652 16541
rect 48228 16396 48280 16448
rect 49240 16439 49292 16448
rect 49240 16405 49249 16439
rect 49249 16405 49283 16439
rect 49283 16405 49292 16439
rect 49240 16396 49292 16405
rect 49424 16396 49476 16448
rect 50252 16396 50304 16448
rect 50620 16439 50672 16448
rect 50620 16405 50629 16439
rect 50629 16405 50663 16439
rect 50663 16405 50672 16439
rect 50620 16396 50672 16405
rect 52552 16396 52604 16448
rect 53564 16439 53616 16448
rect 53564 16405 53573 16439
rect 53573 16405 53607 16439
rect 53607 16405 53616 16439
rect 53564 16396 53616 16405
rect 55220 16396 55272 16448
rect 56876 16396 56928 16448
rect 57612 16439 57664 16448
rect 57612 16405 57621 16439
rect 57621 16405 57655 16439
rect 57655 16405 57664 16439
rect 57612 16396 57664 16405
rect 57888 16396 57940 16448
rect 15394 16294 15446 16346
rect 15458 16294 15510 16346
rect 15522 16294 15574 16346
rect 15586 16294 15638 16346
rect 15650 16294 15702 16346
rect 29838 16294 29890 16346
rect 29902 16294 29954 16346
rect 29966 16294 30018 16346
rect 30030 16294 30082 16346
rect 30094 16294 30146 16346
rect 44282 16294 44334 16346
rect 44346 16294 44398 16346
rect 44410 16294 44462 16346
rect 44474 16294 44526 16346
rect 44538 16294 44590 16346
rect 58726 16294 58778 16346
rect 58790 16294 58842 16346
rect 58854 16294 58906 16346
rect 58918 16294 58970 16346
rect 58982 16294 59034 16346
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 2964 16192 3016 16244
rect 3424 16192 3476 16244
rect 4896 16235 4948 16244
rect 4896 16201 4905 16235
rect 4905 16201 4939 16235
rect 4939 16201 4948 16235
rect 4896 16192 4948 16201
rect 16580 16192 16632 16244
rect 17040 16192 17092 16244
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 20904 16235 20956 16244
rect 20904 16201 20913 16235
rect 20913 16201 20947 16235
rect 20947 16201 20956 16235
rect 20904 16192 20956 16201
rect 21272 16235 21324 16244
rect 21272 16201 21281 16235
rect 21281 16201 21315 16235
rect 21315 16201 21324 16235
rect 21272 16192 21324 16201
rect 22744 16192 22796 16244
rect 23112 16192 23164 16244
rect 3056 16099 3108 16108
rect 3056 16065 3065 16099
rect 3065 16065 3099 16099
rect 3099 16065 3108 16099
rect 3056 16056 3108 16065
rect 4528 16124 4580 16176
rect 4620 16056 4672 16108
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 5632 16056 5684 16108
rect 18328 16124 18380 16176
rect 20352 16124 20404 16176
rect 8208 16099 8260 16108
rect 8208 16065 8217 16099
rect 8217 16065 8251 16099
rect 8251 16065 8260 16099
rect 8208 16056 8260 16065
rect 6736 16031 6788 16040
rect 6736 15997 6745 16031
rect 6745 15997 6779 16031
rect 6779 15997 6788 16031
rect 6736 15988 6788 15997
rect 7288 15988 7340 16040
rect 7472 16031 7524 16040
rect 7472 15997 7481 16031
rect 7481 15997 7515 16031
rect 7515 15997 7524 16031
rect 8760 16056 8812 16108
rect 7472 15988 7524 15997
rect 6000 15852 6052 15904
rect 6552 15852 6604 15904
rect 14832 16056 14884 16108
rect 16120 16056 16172 16108
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 12440 15988 12492 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 15568 15988 15620 16040
rect 15844 15988 15896 16040
rect 9496 15920 9548 15972
rect 15936 15920 15988 15972
rect 9588 15852 9640 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11612 15852 11664 15904
rect 12072 15852 12124 15904
rect 12348 15852 12400 15904
rect 13176 15895 13228 15904
rect 13176 15861 13185 15895
rect 13185 15861 13219 15895
rect 13219 15861 13228 15895
rect 13176 15852 13228 15861
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 16396 15852 16448 15904
rect 19248 15988 19300 16040
rect 20720 15988 20772 16040
rect 21180 15988 21232 16040
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 22744 16099 22796 16108
rect 22744 16065 22753 16099
rect 22753 16065 22787 16099
rect 22787 16065 22796 16099
rect 22744 16056 22796 16065
rect 25320 16192 25372 16244
rect 26424 16235 26476 16244
rect 26424 16201 26433 16235
rect 26433 16201 26467 16235
rect 26467 16201 26476 16235
rect 26424 16192 26476 16201
rect 29368 16192 29420 16244
rect 30196 16192 30248 16244
rect 30380 16235 30432 16244
rect 30380 16201 30389 16235
rect 30389 16201 30423 16235
rect 30423 16201 30432 16235
rect 30380 16192 30432 16201
rect 31484 16192 31536 16244
rect 31944 16235 31996 16244
rect 31944 16201 31953 16235
rect 31953 16201 31987 16235
rect 31987 16201 31996 16235
rect 31944 16192 31996 16201
rect 32128 16235 32180 16244
rect 32128 16201 32137 16235
rect 32137 16201 32171 16235
rect 32171 16201 32180 16235
rect 32128 16192 32180 16201
rect 32496 16192 32548 16244
rect 32956 16192 33008 16244
rect 34152 16192 34204 16244
rect 37648 16192 37700 16244
rect 37924 16192 37976 16244
rect 40684 16192 40736 16244
rect 43996 16192 44048 16244
rect 45192 16235 45244 16244
rect 45192 16201 45201 16235
rect 45201 16201 45235 16235
rect 45235 16201 45244 16235
rect 45192 16192 45244 16201
rect 47032 16192 47084 16244
rect 27252 16167 27304 16176
rect 27252 16133 27286 16167
rect 27286 16133 27304 16167
rect 27252 16124 27304 16133
rect 26056 16056 26108 16108
rect 27068 16056 27120 16108
rect 22928 15988 22980 16040
rect 23112 15988 23164 16040
rect 24308 16031 24360 16040
rect 24308 15997 24317 16031
rect 24317 15997 24351 16031
rect 24351 15997 24360 16031
rect 24308 15988 24360 15997
rect 24400 15988 24452 16040
rect 23020 15963 23072 15972
rect 23020 15929 23029 15963
rect 23029 15929 23063 15963
rect 23063 15929 23072 15963
rect 23020 15920 23072 15929
rect 26332 16031 26384 16040
rect 26332 15997 26341 16031
rect 26341 15997 26375 16031
rect 26375 15997 26384 16031
rect 26332 15988 26384 15997
rect 21916 15852 21968 15904
rect 22468 15852 22520 15904
rect 23204 15852 23256 15904
rect 25504 15895 25556 15904
rect 25504 15861 25513 15895
rect 25513 15861 25547 15895
rect 25547 15861 25556 15895
rect 25504 15852 25556 15861
rect 26792 15895 26844 15904
rect 26792 15861 26801 15895
rect 26801 15861 26835 15895
rect 26835 15861 26844 15895
rect 26792 15852 26844 15861
rect 28080 15988 28132 16040
rect 28540 16031 28592 16040
rect 28540 15997 28549 16031
rect 28549 15997 28583 16031
rect 28583 15997 28592 16031
rect 28540 15988 28592 15997
rect 31300 16056 31352 16108
rect 33692 16056 33744 16108
rect 34428 16056 34480 16108
rect 36176 16099 36228 16108
rect 36176 16065 36185 16099
rect 36185 16065 36219 16099
rect 36219 16065 36228 16099
rect 36176 16056 36228 16065
rect 32956 15988 33008 16040
rect 33140 16031 33192 16040
rect 33140 15997 33149 16031
rect 33149 15997 33183 16031
rect 33183 15997 33192 16031
rect 33140 15988 33192 15997
rect 33784 16031 33836 16040
rect 33784 15997 33793 16031
rect 33793 15997 33827 16031
rect 33827 15997 33836 16031
rect 33784 15988 33836 15997
rect 35716 15988 35768 16040
rect 35992 15988 36044 16040
rect 36820 15988 36872 16040
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 38016 16056 38068 16108
rect 43168 16056 43220 16108
rect 47308 16167 47360 16176
rect 47308 16133 47317 16167
rect 47317 16133 47351 16167
rect 47351 16133 47360 16167
rect 47308 16124 47360 16133
rect 45468 16056 45520 16108
rect 45928 16099 45980 16108
rect 45928 16065 45962 16099
rect 45962 16065 45980 16099
rect 45928 16056 45980 16065
rect 48228 16099 48280 16108
rect 48228 16065 48237 16099
rect 48237 16065 48271 16099
rect 48271 16065 48280 16099
rect 48228 16056 48280 16065
rect 50988 16192 51040 16244
rect 52552 16192 52604 16244
rect 53564 16192 53616 16244
rect 54576 16192 54628 16244
rect 55312 16192 55364 16244
rect 56508 16192 56560 16244
rect 57520 16192 57572 16244
rect 57612 16192 57664 16244
rect 53012 16124 53064 16176
rect 51724 16056 51776 16108
rect 52736 16056 52788 16108
rect 54392 16099 54444 16108
rect 54392 16065 54426 16099
rect 54426 16065 54444 16099
rect 54392 16056 54444 16065
rect 57336 16124 57388 16176
rect 32588 15920 32640 15972
rect 28172 15852 28224 15904
rect 28908 15852 28960 15904
rect 30472 15852 30524 15904
rect 31576 15852 31628 15904
rect 35440 15920 35492 15972
rect 36360 15920 36412 15972
rect 35164 15895 35216 15904
rect 35164 15861 35173 15895
rect 35173 15861 35207 15895
rect 35207 15861 35216 15895
rect 35164 15852 35216 15861
rect 36544 15852 36596 15904
rect 37556 15852 37608 15904
rect 39028 15852 39080 15904
rect 39580 15852 39632 15904
rect 41604 15988 41656 16040
rect 41972 15988 42024 16040
rect 42800 15988 42852 16040
rect 42340 15920 42392 15972
rect 44088 15988 44140 16040
rect 44180 15988 44232 16040
rect 45008 15988 45060 16040
rect 48412 16031 48464 16040
rect 48412 15997 48430 16031
rect 48430 15997 48464 16031
rect 48412 15988 48464 15997
rect 49332 15988 49384 16040
rect 49424 16031 49476 16040
rect 49424 15997 49433 16031
rect 49433 15997 49467 16031
rect 49467 15997 49476 16031
rect 49424 15988 49476 15997
rect 48688 15920 48740 15972
rect 48872 15920 48924 15972
rect 58072 15988 58124 16040
rect 40224 15895 40276 15904
rect 40224 15861 40233 15895
rect 40233 15861 40267 15895
rect 40267 15861 40276 15895
rect 40224 15852 40276 15861
rect 41236 15895 41288 15904
rect 41236 15861 41245 15895
rect 41245 15861 41279 15895
rect 41279 15861 41288 15895
rect 41236 15852 41288 15861
rect 42156 15895 42208 15904
rect 42156 15861 42165 15895
rect 42165 15861 42199 15895
rect 42199 15861 42208 15895
rect 42156 15852 42208 15861
rect 47032 15895 47084 15904
rect 47032 15861 47041 15895
rect 47041 15861 47075 15895
rect 47075 15861 47084 15895
rect 47032 15852 47084 15861
rect 49792 15852 49844 15904
rect 52368 15852 52420 15904
rect 55496 15895 55548 15904
rect 55496 15861 55505 15895
rect 55505 15861 55539 15895
rect 55539 15861 55548 15895
rect 55496 15852 55548 15861
rect 56324 15852 56376 15904
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 22616 15750 22668 15802
rect 22680 15750 22732 15802
rect 22744 15750 22796 15802
rect 22808 15750 22860 15802
rect 22872 15750 22924 15802
rect 37060 15750 37112 15802
rect 37124 15750 37176 15802
rect 37188 15750 37240 15802
rect 37252 15750 37304 15802
rect 37316 15750 37368 15802
rect 51504 15750 51556 15802
rect 51568 15750 51620 15802
rect 51632 15750 51684 15802
rect 51696 15750 51748 15802
rect 51760 15750 51812 15802
rect 3516 15648 3568 15700
rect 3424 15580 3476 15632
rect 4528 15580 4580 15632
rect 5356 15648 5408 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 6552 15691 6604 15700
rect 6552 15657 6561 15691
rect 6561 15657 6595 15691
rect 6595 15657 6604 15691
rect 6552 15648 6604 15657
rect 7472 15648 7524 15700
rect 10876 15648 10928 15700
rect 13728 15648 13780 15700
rect 14832 15648 14884 15700
rect 15752 15648 15804 15700
rect 15936 15648 15988 15700
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 17868 15648 17920 15700
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21272 15648 21324 15700
rect 24308 15648 24360 15700
rect 25964 15691 26016 15700
rect 25964 15657 25973 15691
rect 25973 15657 26007 15691
rect 26007 15657 26016 15691
rect 25964 15648 26016 15657
rect 26332 15648 26384 15700
rect 26792 15648 26844 15700
rect 28724 15648 28776 15700
rect 28908 15648 28960 15700
rect 2596 15444 2648 15496
rect 2872 15419 2924 15428
rect 2872 15385 2881 15419
rect 2881 15385 2915 15419
rect 2915 15385 2924 15419
rect 2872 15376 2924 15385
rect 4252 15444 4304 15496
rect 4344 15444 4396 15496
rect 4436 15487 4488 15496
rect 4436 15453 4445 15487
rect 4445 15453 4479 15487
rect 4479 15453 4488 15487
rect 4436 15444 4488 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 5172 15376 5224 15428
rect 5540 15419 5592 15428
rect 5540 15385 5549 15419
rect 5549 15385 5583 15419
rect 5583 15385 5592 15419
rect 5540 15376 5592 15385
rect 4620 15308 4672 15360
rect 5724 15351 5776 15360
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 6460 15580 6512 15632
rect 7380 15580 7432 15632
rect 9220 15623 9272 15632
rect 9220 15589 9229 15623
rect 9229 15589 9263 15623
rect 9263 15589 9272 15623
rect 9220 15580 9272 15589
rect 6828 15512 6880 15564
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6736 15444 6788 15496
rect 6552 15419 6604 15428
rect 6552 15385 6593 15419
rect 6593 15385 6604 15419
rect 7012 15444 7064 15496
rect 7196 15444 7248 15496
rect 10416 15512 10468 15564
rect 16764 15512 16816 15564
rect 17776 15512 17828 15564
rect 26884 15512 26936 15564
rect 29276 15648 29328 15700
rect 30380 15648 30432 15700
rect 9496 15444 9548 15496
rect 11704 15444 11756 15496
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 12348 15487 12400 15496
rect 12348 15453 12382 15487
rect 12382 15453 12400 15487
rect 12348 15444 12400 15453
rect 18052 15444 18104 15496
rect 19248 15487 19300 15496
rect 19248 15453 19257 15487
rect 19257 15453 19291 15487
rect 19291 15453 19300 15487
rect 19248 15444 19300 15453
rect 21364 15444 21416 15496
rect 23480 15444 23532 15496
rect 29552 15580 29604 15632
rect 31852 15555 31904 15564
rect 31852 15521 31861 15555
rect 31861 15521 31895 15555
rect 31895 15521 31904 15555
rect 31852 15512 31904 15521
rect 32496 15555 32548 15564
rect 32496 15521 32505 15555
rect 32505 15521 32539 15555
rect 32539 15521 32548 15555
rect 32496 15512 32548 15521
rect 33600 15648 33652 15700
rect 35164 15648 35216 15700
rect 37556 15648 37608 15700
rect 38936 15648 38988 15700
rect 42524 15691 42576 15700
rect 42524 15657 42533 15691
rect 42533 15657 42567 15691
rect 42567 15657 42576 15691
rect 42524 15648 42576 15657
rect 45468 15648 45520 15700
rect 47676 15648 47728 15700
rect 48136 15691 48188 15700
rect 48136 15657 48145 15691
rect 48145 15657 48179 15691
rect 48179 15657 48188 15691
rect 48136 15648 48188 15657
rect 48872 15648 48924 15700
rect 49056 15691 49108 15700
rect 49056 15657 49065 15691
rect 49065 15657 49099 15691
rect 49099 15657 49108 15691
rect 49056 15648 49108 15657
rect 49240 15648 49292 15700
rect 6552 15376 6604 15385
rect 7380 15419 7432 15428
rect 7380 15385 7389 15419
rect 7389 15385 7423 15419
rect 7423 15385 7432 15419
rect 7380 15376 7432 15385
rect 8668 15376 8720 15428
rect 9128 15376 9180 15428
rect 14280 15376 14332 15428
rect 18236 15376 18288 15428
rect 19800 15376 19852 15428
rect 21824 15376 21876 15428
rect 23296 15376 23348 15428
rect 29460 15376 29512 15428
rect 30472 15444 30524 15496
rect 31300 15487 31352 15496
rect 31300 15453 31309 15487
rect 31309 15453 31343 15487
rect 31343 15453 31352 15487
rect 31300 15444 31352 15453
rect 31392 15444 31444 15496
rect 31576 15487 31628 15496
rect 31576 15453 31585 15487
rect 31585 15453 31619 15487
rect 31619 15453 31628 15487
rect 31576 15444 31628 15453
rect 32588 15487 32640 15496
rect 32588 15453 32597 15487
rect 32597 15453 32631 15487
rect 32631 15453 32640 15487
rect 32588 15444 32640 15453
rect 35072 15580 35124 15632
rect 36084 15580 36136 15632
rect 36820 15580 36872 15632
rect 35808 15512 35860 15564
rect 36360 15512 36412 15564
rect 36636 15512 36688 15564
rect 33692 15444 33744 15496
rect 34336 15444 34388 15496
rect 35992 15444 36044 15496
rect 41972 15512 42024 15564
rect 42156 15512 42208 15564
rect 44916 15512 44968 15564
rect 46848 15555 46900 15564
rect 46848 15521 46857 15555
rect 46857 15521 46891 15555
rect 46891 15521 46900 15555
rect 46848 15512 46900 15521
rect 47584 15555 47636 15564
rect 47584 15521 47593 15555
rect 47593 15521 47627 15555
rect 47627 15521 47636 15555
rect 47584 15512 47636 15521
rect 48504 15555 48556 15564
rect 48504 15521 48513 15555
rect 48513 15521 48547 15555
rect 48547 15521 48556 15555
rect 48504 15512 48556 15521
rect 55496 15648 55548 15700
rect 55312 15580 55364 15632
rect 52368 15555 52420 15564
rect 52368 15521 52377 15555
rect 52377 15521 52411 15555
rect 52411 15521 52420 15555
rect 52368 15512 52420 15521
rect 52644 15555 52696 15564
rect 52644 15521 52653 15555
rect 52653 15521 52687 15555
rect 52687 15521 52696 15555
rect 52644 15512 52696 15521
rect 53472 15512 53524 15564
rect 53656 15512 53708 15564
rect 39856 15444 39908 15496
rect 41604 15444 41656 15496
rect 42064 15444 42116 15496
rect 43720 15444 43772 15496
rect 46664 15487 46716 15496
rect 46664 15453 46673 15487
rect 46673 15453 46707 15487
rect 46707 15453 46716 15487
rect 46664 15444 46716 15453
rect 7840 15308 7892 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10692 15308 10744 15360
rect 14556 15308 14608 15360
rect 15568 15308 15620 15360
rect 15844 15308 15896 15360
rect 17960 15308 18012 15360
rect 18328 15308 18380 15360
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 21272 15308 21324 15360
rect 21732 15308 21784 15360
rect 22468 15308 22520 15360
rect 22652 15351 22704 15360
rect 22652 15317 22661 15351
rect 22661 15317 22695 15351
rect 22695 15317 22704 15351
rect 22652 15308 22704 15317
rect 23756 15308 23808 15360
rect 24584 15351 24636 15360
rect 24584 15317 24593 15351
rect 24593 15317 24627 15351
rect 24627 15317 24636 15351
rect 24584 15308 24636 15317
rect 28264 15308 28316 15360
rect 29092 15351 29144 15360
rect 29092 15317 29101 15351
rect 29101 15317 29135 15351
rect 29135 15317 29144 15351
rect 29092 15308 29144 15317
rect 29276 15308 29328 15360
rect 31760 15308 31812 15360
rect 33968 15351 34020 15360
rect 33968 15317 33977 15351
rect 33977 15317 34011 15351
rect 34011 15317 34020 15351
rect 33968 15308 34020 15317
rect 34612 15308 34664 15360
rect 34704 15351 34756 15360
rect 34704 15317 34713 15351
rect 34713 15317 34747 15351
rect 34747 15317 34756 15351
rect 34704 15308 34756 15317
rect 35256 15376 35308 15428
rect 37648 15376 37700 15428
rect 40776 15376 40828 15428
rect 36636 15351 36688 15360
rect 36636 15317 36645 15351
rect 36645 15317 36679 15351
rect 36679 15317 36688 15351
rect 36636 15308 36688 15317
rect 38476 15308 38528 15360
rect 39580 15351 39632 15360
rect 39580 15317 39589 15351
rect 39589 15317 39623 15351
rect 39623 15317 39632 15351
rect 39580 15308 39632 15317
rect 44732 15376 44784 15428
rect 48228 15376 48280 15428
rect 49424 15444 49476 15496
rect 50620 15444 50672 15496
rect 52552 15487 52604 15496
rect 52552 15453 52570 15487
rect 52570 15453 52604 15487
rect 52552 15444 52604 15453
rect 54484 15512 54536 15564
rect 49240 15376 49292 15428
rect 56416 15648 56468 15700
rect 56784 15648 56836 15700
rect 56784 15512 56836 15564
rect 57888 15691 57940 15700
rect 57888 15657 57897 15691
rect 57897 15657 57931 15691
rect 57931 15657 57940 15691
rect 57888 15648 57940 15657
rect 58256 15512 58308 15564
rect 53932 15376 53984 15428
rect 41972 15308 42024 15360
rect 42800 15308 42852 15360
rect 43352 15308 43404 15360
rect 44180 15308 44232 15360
rect 44640 15308 44692 15360
rect 46204 15351 46256 15360
rect 46204 15317 46213 15351
rect 46213 15317 46247 15351
rect 46247 15317 46256 15351
rect 46204 15308 46256 15317
rect 47308 15308 47360 15360
rect 48596 15308 48648 15360
rect 50160 15308 50212 15360
rect 54668 15308 54720 15360
rect 55220 15308 55272 15360
rect 55772 15308 55824 15360
rect 56784 15308 56836 15360
rect 57520 15351 57572 15360
rect 57520 15317 57529 15351
rect 57529 15317 57563 15351
rect 57563 15317 57572 15351
rect 57520 15308 57572 15317
rect 15394 15206 15446 15258
rect 15458 15206 15510 15258
rect 15522 15206 15574 15258
rect 15586 15206 15638 15258
rect 15650 15206 15702 15258
rect 29838 15206 29890 15258
rect 29902 15206 29954 15258
rect 29966 15206 30018 15258
rect 30030 15206 30082 15258
rect 30094 15206 30146 15258
rect 44282 15206 44334 15258
rect 44346 15206 44398 15258
rect 44410 15206 44462 15258
rect 44474 15206 44526 15258
rect 44538 15206 44590 15258
rect 58726 15206 58778 15258
rect 58790 15206 58842 15258
rect 58854 15206 58906 15258
rect 58918 15206 58970 15258
rect 58982 15206 59034 15258
rect 2596 15147 2648 15156
rect 2596 15113 2605 15147
rect 2605 15113 2639 15147
rect 2639 15113 2648 15147
rect 2596 15104 2648 15113
rect 2872 15104 2924 15156
rect 3056 15104 3108 15156
rect 3516 15104 3568 15156
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 3148 15011 3200 15020
rect 3148 14977 3157 15011
rect 3157 14977 3191 15011
rect 3191 14977 3200 15011
rect 3148 14968 3200 14977
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 4344 15104 4396 15156
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 4712 15104 4764 15156
rect 5724 15104 5776 15156
rect 6000 15104 6052 15156
rect 6092 15104 6144 15156
rect 2780 14832 2832 14884
rect 3884 14900 3936 14952
rect 5540 14968 5592 15020
rect 5632 14900 5684 14952
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 9220 15104 9272 15156
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 12624 15104 12676 15156
rect 14280 15104 14332 15156
rect 16396 15104 16448 15156
rect 18052 15104 18104 15156
rect 18880 15104 18932 15156
rect 19800 15147 19852 15156
rect 19800 15113 19809 15147
rect 19809 15113 19843 15147
rect 19843 15113 19852 15147
rect 19800 15104 19852 15113
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 23112 15147 23164 15156
rect 23112 15113 23121 15147
rect 23121 15113 23155 15147
rect 23155 15113 23164 15147
rect 23112 15104 23164 15113
rect 29092 15104 29144 15156
rect 32036 15104 32088 15156
rect 33692 15147 33744 15156
rect 33692 15113 33701 15147
rect 33701 15113 33735 15147
rect 33735 15113 33744 15147
rect 33692 15104 33744 15113
rect 34428 15147 34480 15156
rect 34428 15113 34437 15147
rect 34437 15113 34471 15147
rect 34471 15113 34480 15147
rect 34428 15104 34480 15113
rect 40776 15104 40828 15156
rect 10324 15036 10376 15088
rect 13176 15036 13228 15088
rect 17868 15036 17920 15088
rect 18788 15079 18840 15088
rect 18788 15045 18797 15079
rect 18797 15045 18831 15079
rect 18831 15045 18840 15079
rect 18788 15036 18840 15045
rect 29184 15036 29236 15088
rect 29460 15036 29512 15088
rect 41236 15036 41288 15088
rect 7012 14900 7064 14952
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 11612 14900 11664 14952
rect 12256 14900 12308 14952
rect 3976 14764 4028 14816
rect 4068 14764 4120 14816
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 11704 14764 11756 14816
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 14096 14943 14148 14952
rect 14096 14909 14105 14943
rect 14105 14909 14139 14943
rect 14139 14909 14148 14943
rect 19984 14968 20036 15020
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 22652 14968 22704 15020
rect 28264 14968 28316 15020
rect 28540 14968 28592 15020
rect 14096 14900 14148 14909
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 15016 14900 15068 14952
rect 12716 14875 12768 14884
rect 12716 14841 12725 14875
rect 12725 14841 12759 14875
rect 12759 14841 12768 14875
rect 12716 14832 12768 14841
rect 15200 14832 15252 14884
rect 16028 14900 16080 14952
rect 20076 14832 20128 14884
rect 31576 14968 31628 15020
rect 33968 14968 34020 15020
rect 34704 14968 34756 15020
rect 43260 15104 43312 15156
rect 44732 15104 44784 15156
rect 45928 15104 45980 15156
rect 47216 15104 47268 15156
rect 47584 15104 47636 15156
rect 48228 15147 48280 15156
rect 48228 15113 48237 15147
rect 48237 15113 48271 15147
rect 48271 15113 48280 15147
rect 48228 15104 48280 15113
rect 52368 15104 52420 15156
rect 54392 15147 54444 15156
rect 54392 15113 54401 15147
rect 54401 15113 54435 15147
rect 54435 15113 54444 15147
rect 54392 15104 54444 15113
rect 41972 15011 42024 15020
rect 41972 14977 41981 15011
rect 41981 14977 42015 15011
rect 42015 14977 42024 15011
rect 41972 14968 42024 14977
rect 43168 14968 43220 15020
rect 43352 15011 43404 15020
rect 43352 14977 43361 15011
rect 43361 14977 43395 15011
rect 43395 14977 43404 15011
rect 43352 14968 43404 14977
rect 44180 14968 44232 15020
rect 44640 14968 44692 15020
rect 46204 14968 46256 15020
rect 47032 14968 47084 15020
rect 48504 14968 48556 15020
rect 54116 14968 54168 15020
rect 54668 14968 54720 15020
rect 31300 14900 31352 14952
rect 32312 14900 32364 14952
rect 35716 14943 35768 14952
rect 35716 14909 35725 14943
rect 35725 14909 35759 14943
rect 35759 14909 35768 14943
rect 35716 14900 35768 14909
rect 39028 14900 39080 14952
rect 39856 14943 39908 14952
rect 39856 14909 39865 14943
rect 39865 14909 39899 14943
rect 39899 14909 39908 14943
rect 39856 14900 39908 14909
rect 41512 14900 41564 14952
rect 41696 14900 41748 14952
rect 41420 14832 41472 14884
rect 42248 14832 42300 14884
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 13636 14764 13688 14816
rect 16764 14764 16816 14816
rect 21272 14764 21324 14816
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 24216 14764 24268 14816
rect 34612 14764 34664 14816
rect 35808 14764 35860 14816
rect 42432 14807 42484 14816
rect 42432 14773 42441 14807
rect 42441 14773 42475 14807
rect 42475 14773 42484 14807
rect 42432 14764 42484 14773
rect 49608 14943 49660 14952
rect 49608 14909 49617 14943
rect 49617 14909 49651 14943
rect 49651 14909 49660 14943
rect 49608 14900 49660 14909
rect 50252 14943 50304 14952
rect 50252 14909 50261 14943
rect 50261 14909 50295 14943
rect 50295 14909 50304 14943
rect 50252 14900 50304 14909
rect 51908 14875 51960 14884
rect 51908 14841 51917 14875
rect 51917 14841 51951 14875
rect 51951 14841 51960 14875
rect 51908 14832 51960 14841
rect 43812 14764 43864 14816
rect 46848 14764 46900 14816
rect 48872 14764 48924 14816
rect 49332 14764 49384 14816
rect 51080 14764 51132 14816
rect 57428 14807 57480 14816
rect 57428 14773 57437 14807
rect 57437 14773 57471 14807
rect 57471 14773 57480 14807
rect 57428 14764 57480 14773
rect 58164 14764 58216 14816
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 22616 14662 22668 14714
rect 22680 14662 22732 14714
rect 22744 14662 22796 14714
rect 22808 14662 22860 14714
rect 22872 14662 22924 14714
rect 37060 14662 37112 14714
rect 37124 14662 37176 14714
rect 37188 14662 37240 14714
rect 37252 14662 37304 14714
rect 37316 14662 37368 14714
rect 51504 14662 51556 14714
rect 51568 14662 51620 14714
rect 51632 14662 51684 14714
rect 51696 14662 51748 14714
rect 51760 14662 51812 14714
rect 3148 14560 3200 14612
rect 3332 14560 3384 14612
rect 4068 14560 4120 14612
rect 4712 14560 4764 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 6552 14560 6604 14612
rect 6736 14560 6788 14612
rect 3516 14492 3568 14544
rect 3884 14356 3936 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 9864 14560 9916 14612
rect 11520 14560 11572 14612
rect 14280 14603 14332 14612
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 14832 14560 14884 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 21180 14603 21232 14612
rect 21180 14569 21189 14603
rect 21189 14569 21223 14603
rect 21223 14569 21232 14603
rect 21180 14560 21232 14569
rect 21364 14560 21416 14612
rect 3608 14331 3660 14340
rect 3608 14297 3617 14331
rect 3617 14297 3651 14331
rect 3651 14297 3660 14331
rect 7012 14356 7064 14408
rect 16120 14492 16172 14544
rect 28540 14560 28592 14612
rect 28908 14560 28960 14612
rect 32588 14560 32640 14612
rect 35072 14560 35124 14612
rect 35440 14560 35492 14612
rect 37464 14560 37516 14612
rect 38200 14560 38252 14612
rect 39856 14560 39908 14612
rect 42156 14560 42208 14612
rect 42432 14560 42484 14612
rect 42616 14560 42668 14612
rect 47216 14560 47268 14612
rect 48596 14560 48648 14612
rect 12072 14424 12124 14476
rect 14096 14424 14148 14476
rect 8668 14356 8720 14408
rect 16764 14424 16816 14476
rect 19064 14424 19116 14476
rect 22100 14424 22152 14476
rect 26056 14467 26108 14476
rect 26056 14433 26065 14467
rect 26065 14433 26099 14467
rect 26099 14433 26108 14467
rect 26056 14424 26108 14433
rect 31024 14492 31076 14544
rect 31116 14424 31168 14476
rect 41512 14424 41564 14476
rect 42248 14424 42300 14476
rect 16028 14356 16080 14408
rect 16672 14356 16724 14408
rect 17316 14356 17368 14408
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 22376 14399 22428 14408
rect 22376 14365 22385 14399
rect 22385 14365 22419 14399
rect 22419 14365 22428 14399
rect 22376 14356 22428 14365
rect 24676 14356 24728 14408
rect 25320 14399 25372 14408
rect 25320 14365 25329 14399
rect 25329 14365 25363 14399
rect 25363 14365 25372 14399
rect 25320 14356 25372 14365
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 3608 14288 3660 14297
rect 3332 14220 3384 14272
rect 4528 14288 4580 14340
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 9956 14331 10008 14340
rect 9956 14297 9990 14331
rect 9990 14297 10008 14331
rect 9956 14288 10008 14297
rect 10876 14288 10928 14340
rect 13268 14288 13320 14340
rect 15292 14288 15344 14340
rect 20720 14331 20772 14340
rect 20720 14297 20729 14331
rect 20729 14297 20763 14331
rect 20763 14297 20772 14331
rect 20720 14288 20772 14297
rect 21548 14288 21600 14340
rect 26148 14288 26200 14340
rect 27252 14288 27304 14340
rect 32404 14356 32456 14408
rect 36084 14399 36136 14408
rect 36084 14365 36093 14399
rect 36093 14365 36127 14399
rect 36127 14365 36136 14399
rect 36084 14356 36136 14365
rect 36176 14356 36228 14408
rect 37832 14356 37884 14408
rect 38660 14356 38712 14408
rect 42524 14492 42576 14544
rect 49148 14492 49200 14544
rect 49608 14560 49660 14612
rect 54116 14603 54168 14612
rect 54116 14569 54125 14603
rect 54125 14569 54159 14603
rect 54159 14569 54168 14603
rect 54116 14560 54168 14569
rect 56600 14560 56652 14612
rect 43720 14467 43772 14476
rect 43720 14433 43729 14467
rect 43729 14433 43763 14467
rect 43763 14433 43772 14467
rect 43720 14424 43772 14433
rect 44824 14424 44876 14476
rect 44916 14356 44968 14408
rect 46664 14399 46716 14408
rect 46664 14365 46673 14399
rect 46673 14365 46707 14399
rect 46707 14365 46716 14399
rect 46664 14356 46716 14365
rect 30380 14288 30432 14340
rect 34428 14288 34480 14340
rect 38384 14288 38436 14340
rect 41696 14331 41748 14340
rect 41696 14297 41705 14331
rect 41705 14297 41739 14331
rect 41739 14297 41748 14331
rect 41696 14288 41748 14297
rect 41788 14288 41840 14340
rect 10600 14220 10652 14272
rect 12256 14220 12308 14272
rect 14924 14220 14976 14272
rect 15936 14263 15988 14272
rect 15936 14229 15945 14263
rect 15945 14229 15979 14263
rect 15979 14229 15988 14263
rect 15936 14220 15988 14229
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 24216 14220 24268 14272
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 26056 14220 26108 14272
rect 27436 14263 27488 14272
rect 27436 14229 27445 14263
rect 27445 14229 27479 14263
rect 27479 14229 27488 14263
rect 27436 14220 27488 14229
rect 29644 14220 29696 14272
rect 31024 14220 31076 14272
rect 31576 14220 31628 14272
rect 36820 14220 36872 14272
rect 36912 14220 36964 14272
rect 37004 14220 37056 14272
rect 37924 14263 37976 14272
rect 37924 14229 37933 14263
rect 37933 14229 37967 14263
rect 37967 14229 37976 14263
rect 37924 14220 37976 14229
rect 42340 14263 42392 14272
rect 42340 14229 42349 14263
rect 42349 14229 42383 14263
rect 42383 14229 42392 14263
rect 42340 14220 42392 14229
rect 43812 14263 43864 14272
rect 43812 14229 43821 14263
rect 43821 14229 43855 14263
rect 43855 14229 43864 14263
rect 43812 14220 43864 14229
rect 44180 14263 44232 14272
rect 44180 14229 44189 14263
rect 44189 14229 44223 14263
rect 44223 14229 44232 14263
rect 44180 14220 44232 14229
rect 45928 14220 45980 14272
rect 46204 14220 46256 14272
rect 48596 14220 48648 14272
rect 49240 14399 49292 14408
rect 49240 14365 49249 14399
rect 49249 14365 49283 14399
rect 49283 14365 49292 14399
rect 49240 14356 49292 14365
rect 49332 14399 49384 14408
rect 49332 14365 49341 14399
rect 49341 14365 49375 14399
rect 49375 14365 49384 14399
rect 49332 14356 49384 14365
rect 52552 14492 52604 14544
rect 51908 14424 51960 14476
rect 49700 14220 49752 14272
rect 54852 14399 54904 14408
rect 54852 14365 54861 14399
rect 54861 14365 54895 14399
rect 54895 14365 54904 14399
rect 54852 14356 54904 14365
rect 58440 14399 58492 14408
rect 58440 14365 58449 14399
rect 58449 14365 58483 14399
rect 58483 14365 58492 14399
rect 58440 14356 58492 14365
rect 51540 14288 51592 14340
rect 53012 14288 53064 14340
rect 51908 14220 51960 14272
rect 52092 14263 52144 14272
rect 52092 14229 52101 14263
rect 52101 14229 52135 14263
rect 52135 14229 52144 14263
rect 52092 14220 52144 14229
rect 54300 14263 54352 14272
rect 54300 14229 54309 14263
rect 54309 14229 54343 14263
rect 54343 14229 54352 14263
rect 54300 14220 54352 14229
rect 56876 14220 56928 14272
rect 57244 14220 57296 14272
rect 15394 14118 15446 14170
rect 15458 14118 15510 14170
rect 15522 14118 15574 14170
rect 15586 14118 15638 14170
rect 15650 14118 15702 14170
rect 29838 14118 29890 14170
rect 29902 14118 29954 14170
rect 29966 14118 30018 14170
rect 30030 14118 30082 14170
rect 30094 14118 30146 14170
rect 44282 14118 44334 14170
rect 44346 14118 44398 14170
rect 44410 14118 44462 14170
rect 44474 14118 44526 14170
rect 44538 14118 44590 14170
rect 58726 14118 58778 14170
rect 58790 14118 58842 14170
rect 58854 14118 58906 14170
rect 58918 14118 58970 14170
rect 58982 14118 59034 14170
rect 3332 14059 3384 14068
rect 3332 14025 3341 14059
rect 3341 14025 3375 14059
rect 3375 14025 3384 14059
rect 3332 14016 3384 14025
rect 4344 14016 4396 14068
rect 7196 14016 7248 14068
rect 7288 14016 7340 14068
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 3976 13948 4028 14000
rect 3884 13880 3936 13932
rect 4068 13812 4120 13864
rect 6368 13880 6420 13932
rect 9864 14016 9916 14068
rect 9956 14016 10008 14068
rect 9680 13880 9732 13932
rect 10600 14059 10652 14068
rect 10600 14025 10609 14059
rect 10609 14025 10643 14059
rect 10643 14025 10652 14059
rect 10600 14016 10652 14025
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 10876 14016 10928 14068
rect 11336 14016 11388 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 12716 14016 12768 14068
rect 13176 14016 13228 14068
rect 13268 14059 13320 14068
rect 13268 14025 13277 14059
rect 13277 14025 13311 14059
rect 13311 14025 13320 14059
rect 13268 14016 13320 14025
rect 13452 14016 13504 14068
rect 15936 14016 15988 14068
rect 16028 14059 16080 14068
rect 16028 14025 16037 14059
rect 16037 14025 16071 14059
rect 16071 14025 16080 14059
rect 16028 14016 16080 14025
rect 16212 14016 16264 14068
rect 15200 13991 15252 14000
rect 15200 13957 15209 13991
rect 15209 13957 15243 13991
rect 15243 13957 15252 13991
rect 15200 13948 15252 13957
rect 16580 13948 16632 14000
rect 16948 13991 17000 14000
rect 16948 13957 16971 13991
rect 16971 13957 17000 13991
rect 16948 13948 17000 13957
rect 18604 14016 18656 14068
rect 5908 13812 5960 13864
rect 9128 13812 9180 13864
rect 10508 13812 10560 13864
rect 2596 13676 2648 13728
rect 6828 13676 6880 13728
rect 9680 13744 9732 13796
rect 13912 13880 13964 13932
rect 15752 13880 15804 13932
rect 18052 13880 18104 13932
rect 12256 13744 12308 13796
rect 14372 13812 14424 13864
rect 15292 13812 15344 13864
rect 16212 13812 16264 13864
rect 16396 13812 16448 13864
rect 11336 13676 11388 13728
rect 11612 13676 11664 13728
rect 15292 13676 15344 13728
rect 16028 13676 16080 13728
rect 20904 13880 20956 13932
rect 21824 13880 21876 13932
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 25320 14016 25372 14068
rect 26148 14059 26200 14068
rect 26148 14025 26157 14059
rect 26157 14025 26191 14059
rect 26191 14025 26200 14059
rect 26148 14016 26200 14025
rect 27252 14059 27304 14068
rect 27252 14025 27261 14059
rect 27261 14025 27295 14059
rect 27295 14025 27304 14059
rect 27252 14016 27304 14025
rect 27436 14016 27488 14068
rect 24216 13948 24268 14000
rect 19800 13812 19852 13864
rect 19984 13812 20036 13864
rect 20352 13812 20404 13864
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 18052 13744 18104 13796
rect 18328 13744 18380 13796
rect 21272 13744 21324 13796
rect 18972 13719 19024 13728
rect 18972 13685 18981 13719
rect 18981 13685 19015 13719
rect 19015 13685 19024 13719
rect 18972 13676 19024 13685
rect 20076 13719 20128 13728
rect 20076 13685 20085 13719
rect 20085 13685 20119 13719
rect 20119 13685 20128 13719
rect 20076 13676 20128 13685
rect 20720 13676 20772 13728
rect 20812 13676 20864 13728
rect 22100 13744 22152 13796
rect 22468 13744 22520 13796
rect 23480 13855 23532 13864
rect 23480 13821 23489 13855
rect 23489 13821 23523 13855
rect 23523 13821 23532 13855
rect 23480 13812 23532 13821
rect 24400 13923 24452 13932
rect 24400 13889 24434 13923
rect 24434 13889 24452 13923
rect 24400 13880 24452 13889
rect 30380 14016 30432 14068
rect 32404 14016 32456 14068
rect 36084 14016 36136 14068
rect 36544 14016 36596 14068
rect 38384 14016 38436 14068
rect 29276 13880 29328 13932
rect 30932 13948 30984 14000
rect 31668 13948 31720 14000
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 31116 13923 31168 13932
rect 31116 13889 31125 13923
rect 31125 13889 31159 13923
rect 31159 13889 31168 13923
rect 31116 13880 31168 13889
rect 34060 13948 34112 14000
rect 34336 13948 34388 14000
rect 34428 13923 34480 13932
rect 34428 13889 34437 13923
rect 34437 13889 34471 13923
rect 34471 13889 34480 13923
rect 34428 13880 34480 13889
rect 25872 13855 25924 13864
rect 25872 13821 25881 13855
rect 25881 13821 25915 13855
rect 25915 13821 25924 13855
rect 25872 13812 25924 13821
rect 26700 13812 26752 13864
rect 26792 13855 26844 13864
rect 26792 13821 26801 13855
rect 26801 13821 26835 13855
rect 26835 13821 26844 13855
rect 26792 13812 26844 13821
rect 27528 13812 27580 13864
rect 29460 13855 29512 13864
rect 29460 13821 29469 13855
rect 29469 13821 29503 13855
rect 29503 13821 29512 13855
rect 29460 13812 29512 13821
rect 23020 13676 23072 13728
rect 23296 13676 23348 13728
rect 24032 13719 24084 13728
rect 24032 13685 24041 13719
rect 24041 13685 24075 13719
rect 24075 13685 24084 13719
rect 24032 13676 24084 13685
rect 25136 13744 25188 13796
rect 37924 13880 37976 13932
rect 31852 13812 31904 13864
rect 32864 13812 32916 13864
rect 33508 13855 33560 13864
rect 33508 13821 33517 13855
rect 33517 13821 33551 13855
rect 33551 13821 33560 13855
rect 33508 13812 33560 13821
rect 34152 13855 34204 13864
rect 34152 13821 34161 13855
rect 34161 13821 34195 13855
rect 34195 13821 34204 13855
rect 34152 13812 34204 13821
rect 36084 13812 36136 13864
rect 36636 13812 36688 13864
rect 37832 13855 37884 13864
rect 37832 13821 37841 13855
rect 37841 13821 37875 13855
rect 37875 13821 37884 13855
rect 37832 13812 37884 13821
rect 38016 13812 38068 13864
rect 38200 13855 38252 13864
rect 38200 13821 38209 13855
rect 38209 13821 38243 13855
rect 38243 13821 38252 13855
rect 38200 13812 38252 13821
rect 39764 14016 39816 14068
rect 40316 14016 40368 14068
rect 42156 14016 42208 14068
rect 42524 14016 42576 14068
rect 43812 14016 43864 14068
rect 46204 14016 46256 14068
rect 46664 14016 46716 14068
rect 46756 14059 46808 14068
rect 46756 14025 46765 14059
rect 46765 14025 46799 14059
rect 46799 14025 46808 14059
rect 46756 14016 46808 14025
rect 50252 14016 50304 14068
rect 51540 14059 51592 14068
rect 51540 14025 51549 14059
rect 51549 14025 51583 14059
rect 51583 14025 51592 14059
rect 51540 14016 51592 14025
rect 54852 14016 54904 14068
rect 56600 14016 56652 14068
rect 57244 14059 57296 14068
rect 57244 14025 57253 14059
rect 57253 14025 57287 14059
rect 57287 14025 57296 14059
rect 57244 14016 57296 14025
rect 57520 14016 57572 14068
rect 42708 13948 42760 14000
rect 52460 13948 52512 14000
rect 33968 13744 34020 13796
rect 34336 13744 34388 13796
rect 37004 13744 37056 13796
rect 37648 13744 37700 13796
rect 41052 13855 41104 13864
rect 41052 13821 41061 13855
rect 41061 13821 41095 13855
rect 41095 13821 41104 13855
rect 41052 13812 41104 13821
rect 44088 13923 44140 13932
rect 44088 13889 44097 13923
rect 44097 13889 44131 13923
rect 44131 13889 44140 13923
rect 44088 13880 44140 13889
rect 44180 13880 44232 13932
rect 48320 13880 48372 13932
rect 48596 13923 48648 13932
rect 48596 13889 48605 13923
rect 48605 13889 48639 13923
rect 48639 13889 48648 13923
rect 48596 13880 48648 13889
rect 48872 13923 48924 13932
rect 48872 13889 48906 13923
rect 48906 13889 48924 13923
rect 48872 13880 48924 13889
rect 49148 13880 49200 13932
rect 41604 13855 41656 13864
rect 41604 13821 41613 13855
rect 41613 13821 41647 13855
rect 41647 13821 41656 13855
rect 41604 13812 41656 13821
rect 42248 13812 42300 13864
rect 42524 13812 42576 13864
rect 45560 13855 45612 13864
rect 45560 13821 45569 13855
rect 45569 13821 45603 13855
rect 45603 13821 45612 13855
rect 45560 13812 45612 13821
rect 26424 13676 26476 13728
rect 28816 13676 28868 13728
rect 35716 13676 35768 13728
rect 35808 13676 35860 13728
rect 36728 13676 36780 13728
rect 38752 13676 38804 13728
rect 44272 13719 44324 13728
rect 44272 13685 44281 13719
rect 44281 13685 44315 13719
rect 44315 13685 44324 13719
rect 44272 13676 44324 13685
rect 46480 13676 46532 13728
rect 47584 13855 47636 13864
rect 47584 13821 47593 13855
rect 47593 13821 47627 13855
rect 47627 13821 47636 13855
rect 47584 13812 47636 13821
rect 47768 13812 47820 13864
rect 50068 13855 50120 13864
rect 50068 13821 50077 13855
rect 50077 13821 50111 13855
rect 50111 13821 50120 13855
rect 50068 13812 50120 13821
rect 52092 13923 52144 13932
rect 52092 13889 52101 13923
rect 52101 13889 52135 13923
rect 52135 13889 52144 13923
rect 52092 13880 52144 13889
rect 55128 13948 55180 14000
rect 55864 13880 55916 13932
rect 52368 13812 52420 13864
rect 53288 13855 53340 13864
rect 53288 13821 53297 13855
rect 53297 13821 53331 13855
rect 53331 13821 53340 13855
rect 53288 13812 53340 13821
rect 53472 13855 53524 13864
rect 53472 13821 53481 13855
rect 53481 13821 53515 13855
rect 53515 13821 53524 13855
rect 53472 13812 53524 13821
rect 54116 13812 54168 13864
rect 55312 13855 55364 13864
rect 55312 13821 55321 13855
rect 55321 13821 55355 13855
rect 55355 13821 55364 13855
rect 55312 13812 55364 13821
rect 56600 13855 56652 13864
rect 56600 13821 56609 13855
rect 56609 13821 56643 13855
rect 56643 13821 56652 13855
rect 56600 13812 56652 13821
rect 53104 13744 53156 13796
rect 50712 13719 50764 13728
rect 50712 13685 50721 13719
rect 50721 13685 50755 13719
rect 50755 13685 50764 13719
rect 50712 13676 50764 13685
rect 54024 13676 54076 13728
rect 56048 13719 56100 13728
rect 56048 13685 56057 13719
rect 56057 13685 56091 13719
rect 56091 13685 56100 13719
rect 56048 13676 56100 13685
rect 57888 13719 57940 13728
rect 57888 13685 57897 13719
rect 57897 13685 57931 13719
rect 57931 13685 57940 13719
rect 57888 13676 57940 13685
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 22616 13574 22668 13626
rect 22680 13574 22732 13626
rect 22744 13574 22796 13626
rect 22808 13574 22860 13626
rect 22872 13574 22924 13626
rect 37060 13574 37112 13626
rect 37124 13574 37176 13626
rect 37188 13574 37240 13626
rect 37252 13574 37304 13626
rect 37316 13574 37368 13626
rect 51504 13574 51556 13626
rect 51568 13574 51620 13626
rect 51632 13574 51684 13626
rect 51696 13574 51748 13626
rect 51760 13574 51812 13626
rect 2780 13472 2832 13524
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 4068 13515 4120 13524
rect 4068 13481 4077 13515
rect 4077 13481 4111 13515
rect 4111 13481 4120 13515
rect 4068 13472 4120 13481
rect 4436 13472 4488 13524
rect 6368 13472 6420 13524
rect 6828 13472 6880 13524
rect 7380 13515 7432 13524
rect 7380 13481 7389 13515
rect 7389 13481 7423 13515
rect 7423 13481 7432 13515
rect 7380 13472 7432 13481
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 2964 13268 3016 13320
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 5908 13447 5960 13456
rect 5908 13413 5917 13447
rect 5917 13413 5951 13447
rect 5951 13413 5960 13447
rect 5908 13404 5960 13413
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 10692 13472 10744 13524
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 15016 13472 15068 13524
rect 16580 13472 16632 13524
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 8760 13243 8812 13252
rect 8760 13209 8769 13243
rect 8769 13209 8803 13243
rect 8803 13209 8812 13243
rect 8760 13200 8812 13209
rect 6644 13132 6696 13184
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 10416 13132 10468 13184
rect 11060 13132 11112 13184
rect 12900 13336 12952 13388
rect 13728 13336 13780 13388
rect 14280 13336 14332 13388
rect 16304 13404 16356 13456
rect 18328 13515 18380 13524
rect 18328 13481 18337 13515
rect 18337 13481 18371 13515
rect 18371 13481 18380 13515
rect 18328 13472 18380 13481
rect 18880 13472 18932 13524
rect 21180 13472 21232 13524
rect 22376 13472 22428 13524
rect 23296 13515 23348 13524
rect 23296 13481 23305 13515
rect 23305 13481 23339 13515
rect 23339 13481 23348 13515
rect 23296 13472 23348 13481
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 24676 13472 24728 13524
rect 17592 13447 17644 13456
rect 16488 13336 16540 13388
rect 17592 13413 17601 13447
rect 17601 13413 17635 13447
rect 17635 13413 17644 13447
rect 17592 13404 17644 13413
rect 14924 13311 14976 13320
rect 11520 13200 11572 13252
rect 12072 13243 12124 13252
rect 12072 13209 12081 13243
rect 12081 13209 12115 13243
rect 12115 13209 12124 13243
rect 12072 13200 12124 13209
rect 14924 13277 14958 13311
rect 14958 13277 14976 13311
rect 14924 13268 14976 13277
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 18604 13336 18656 13388
rect 18880 13379 18932 13388
rect 18880 13345 18889 13379
rect 18889 13345 18923 13379
rect 18923 13345 18932 13379
rect 18880 13336 18932 13345
rect 17132 13268 17184 13320
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 12992 13243 13044 13252
rect 12992 13209 13001 13243
rect 13001 13209 13035 13243
rect 13035 13209 13044 13243
rect 12992 13200 13044 13209
rect 11612 13132 11664 13184
rect 20352 13447 20404 13456
rect 20352 13413 20361 13447
rect 20361 13413 20395 13447
rect 20395 13413 20404 13447
rect 20352 13404 20404 13413
rect 20720 13404 20772 13456
rect 19800 13379 19852 13388
rect 19800 13345 19809 13379
rect 19809 13345 19843 13379
rect 19843 13345 19852 13379
rect 19800 13336 19852 13345
rect 20812 13379 20864 13388
rect 20812 13345 20821 13379
rect 20821 13345 20855 13379
rect 20855 13345 20864 13379
rect 20812 13336 20864 13345
rect 21640 13268 21692 13320
rect 19800 13200 19852 13252
rect 18144 13132 18196 13184
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 22192 13132 22244 13184
rect 22468 13311 22520 13320
rect 22468 13277 22486 13311
rect 22486 13277 22520 13311
rect 24216 13336 24268 13388
rect 26056 13472 26108 13524
rect 26792 13472 26844 13524
rect 29460 13472 29512 13524
rect 34244 13472 34296 13524
rect 36636 13472 36688 13524
rect 25136 13404 25188 13456
rect 26332 13404 26384 13456
rect 24952 13379 25004 13388
rect 24952 13345 24961 13379
rect 24961 13345 24995 13379
rect 24995 13345 25004 13379
rect 24952 13336 25004 13345
rect 22468 13268 22520 13277
rect 24492 13268 24544 13320
rect 26148 13379 26200 13388
rect 26148 13345 26157 13379
rect 26157 13345 26191 13379
rect 26191 13345 26200 13379
rect 26148 13336 26200 13345
rect 27252 13336 27304 13388
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 23296 13200 23348 13252
rect 27436 13268 27488 13320
rect 28540 13311 28592 13320
rect 28540 13277 28549 13311
rect 28549 13277 28583 13311
rect 28583 13277 28592 13311
rect 28540 13268 28592 13277
rect 28632 13268 28684 13320
rect 33048 13404 33100 13456
rect 32588 13379 32640 13388
rect 32588 13345 32597 13379
rect 32597 13345 32631 13379
rect 32631 13345 32640 13379
rect 32588 13336 32640 13345
rect 37740 13472 37792 13524
rect 39120 13472 39172 13524
rect 41144 13515 41196 13524
rect 41144 13481 41153 13515
rect 41153 13481 41187 13515
rect 41187 13481 41196 13515
rect 41144 13472 41196 13481
rect 41696 13472 41748 13524
rect 42064 13472 42116 13524
rect 45560 13472 45612 13524
rect 47584 13472 47636 13524
rect 51908 13472 51960 13524
rect 35992 13404 36044 13456
rect 37004 13447 37056 13456
rect 37004 13413 37013 13447
rect 37013 13413 37047 13447
rect 37047 13413 37056 13447
rect 37004 13404 37056 13413
rect 47400 13447 47452 13456
rect 47400 13413 47409 13447
rect 47409 13413 47443 13447
rect 47443 13413 47452 13447
rect 47400 13404 47452 13413
rect 48964 13404 49016 13456
rect 34336 13336 34388 13388
rect 35256 13379 35308 13388
rect 35256 13345 35265 13379
rect 35265 13345 35299 13379
rect 35299 13345 35308 13379
rect 35256 13336 35308 13345
rect 35440 13379 35492 13388
rect 35440 13345 35449 13379
rect 35449 13345 35483 13379
rect 35483 13345 35492 13379
rect 35440 13336 35492 13345
rect 35716 13336 35768 13388
rect 36728 13379 36780 13388
rect 36728 13345 36737 13379
rect 36737 13345 36771 13379
rect 36771 13345 36780 13379
rect 36728 13336 36780 13345
rect 37924 13336 37976 13388
rect 42156 13336 42208 13388
rect 42616 13336 42668 13388
rect 48228 13379 48280 13388
rect 48228 13345 48237 13379
rect 48237 13345 48271 13379
rect 48271 13345 48280 13379
rect 48228 13336 48280 13345
rect 48320 13336 48372 13388
rect 49332 13336 49384 13388
rect 51356 13404 51408 13456
rect 53288 13404 53340 13456
rect 36636 13311 36688 13320
rect 36636 13277 36654 13311
rect 36654 13277 36688 13311
rect 36636 13268 36688 13277
rect 37648 13311 37700 13320
rect 37648 13277 37657 13311
rect 37657 13277 37691 13311
rect 37691 13277 37700 13311
rect 37648 13268 37700 13277
rect 39028 13268 39080 13320
rect 43260 13311 43312 13320
rect 43260 13277 43269 13311
rect 43269 13277 43303 13311
rect 43303 13277 43312 13311
rect 43260 13268 43312 13277
rect 44088 13268 44140 13320
rect 45560 13268 45612 13320
rect 45928 13311 45980 13320
rect 45928 13277 45962 13311
rect 45962 13277 45980 13311
rect 27528 13243 27580 13252
rect 27528 13209 27537 13243
rect 27537 13209 27571 13243
rect 27571 13209 27580 13243
rect 27528 13200 27580 13209
rect 29552 13243 29604 13252
rect 29552 13209 29561 13243
rect 29561 13209 29595 13243
rect 29595 13209 29604 13243
rect 29552 13200 29604 13209
rect 22928 13132 22980 13184
rect 25136 13132 25188 13184
rect 26608 13132 26660 13184
rect 27344 13132 27396 13184
rect 30748 13132 30800 13184
rect 33140 13200 33192 13252
rect 34796 13175 34848 13184
rect 34796 13141 34805 13175
rect 34805 13141 34839 13175
rect 34839 13141 34848 13175
rect 34796 13132 34848 13141
rect 35164 13175 35216 13184
rect 35164 13141 35173 13175
rect 35173 13141 35207 13175
rect 35207 13141 35216 13175
rect 35164 13132 35216 13141
rect 38568 13132 38620 13184
rect 38844 13243 38896 13252
rect 38844 13209 38862 13243
rect 38862 13209 38896 13243
rect 38844 13200 38896 13209
rect 39672 13200 39724 13252
rect 41328 13200 41380 13252
rect 41972 13200 42024 13252
rect 42616 13200 42668 13252
rect 44272 13200 44324 13252
rect 45928 13268 45980 13277
rect 46204 13268 46256 13320
rect 48504 13311 48556 13320
rect 48504 13277 48513 13311
rect 48513 13277 48547 13311
rect 48547 13277 48556 13311
rect 48504 13268 48556 13277
rect 50712 13336 50764 13388
rect 53104 13379 53156 13388
rect 53104 13345 53113 13379
rect 53113 13345 53147 13379
rect 53147 13345 53156 13379
rect 53104 13336 53156 13345
rect 55312 13472 55364 13524
rect 58440 13472 58492 13524
rect 49240 13200 49292 13252
rect 41696 13175 41748 13184
rect 41696 13141 41705 13175
rect 41705 13141 41739 13175
rect 41739 13141 41748 13175
rect 41696 13132 41748 13141
rect 42340 13132 42392 13184
rect 47584 13175 47636 13184
rect 47584 13141 47593 13175
rect 47593 13141 47627 13175
rect 47627 13141 47636 13175
rect 47584 13132 47636 13141
rect 48412 13132 48464 13184
rect 52460 13311 52512 13320
rect 52460 13277 52469 13311
rect 52469 13277 52503 13311
rect 52503 13277 52512 13311
rect 52460 13268 52512 13277
rect 55312 13311 55364 13320
rect 55312 13277 55321 13311
rect 55321 13277 55355 13311
rect 55355 13277 55364 13311
rect 56876 13311 56928 13320
rect 55312 13268 55364 13277
rect 56876 13277 56885 13311
rect 56885 13277 56919 13311
rect 56919 13277 56928 13311
rect 56876 13268 56928 13277
rect 57888 13268 57940 13320
rect 53196 13200 53248 13252
rect 50988 13175 51040 13184
rect 50988 13141 50997 13175
rect 50997 13141 51031 13175
rect 51031 13141 51040 13175
rect 50988 13132 51040 13141
rect 51816 13175 51868 13184
rect 51816 13141 51825 13175
rect 51825 13141 51859 13175
rect 51859 13141 51868 13175
rect 51816 13132 51868 13141
rect 53748 13132 53800 13184
rect 54300 13200 54352 13252
rect 56048 13200 56100 13252
rect 55128 13132 55180 13184
rect 56692 13175 56744 13184
rect 56692 13141 56701 13175
rect 56701 13141 56735 13175
rect 56735 13141 56744 13175
rect 56692 13132 56744 13141
rect 15394 13030 15446 13082
rect 15458 13030 15510 13082
rect 15522 13030 15574 13082
rect 15586 13030 15638 13082
rect 15650 13030 15702 13082
rect 29838 13030 29890 13082
rect 29902 13030 29954 13082
rect 29966 13030 30018 13082
rect 30030 13030 30082 13082
rect 30094 13030 30146 13082
rect 44282 13030 44334 13082
rect 44346 13030 44398 13082
rect 44410 13030 44462 13082
rect 44474 13030 44526 13082
rect 44538 13030 44590 13082
rect 58726 13030 58778 13082
rect 58790 13030 58842 13082
rect 58854 13030 58906 13082
rect 58918 13030 58970 13082
rect 58982 13030 59034 13082
rect 4068 12928 4120 12980
rect 6460 12860 6512 12912
rect 6644 12792 6696 12844
rect 16304 12971 16356 12980
rect 16304 12937 16313 12971
rect 16313 12937 16347 12971
rect 16347 12937 16356 12971
rect 16304 12928 16356 12937
rect 16396 12928 16448 12980
rect 17960 12928 18012 12980
rect 20996 12928 21048 12980
rect 21916 12928 21968 12980
rect 22928 12928 22980 12980
rect 24952 12928 25004 12980
rect 25136 12928 25188 12980
rect 9220 12860 9272 12912
rect 10140 12860 10192 12912
rect 11060 12903 11112 12912
rect 11060 12869 11069 12903
rect 11069 12869 11103 12903
rect 11103 12869 11112 12903
rect 11060 12860 11112 12869
rect 13360 12860 13412 12912
rect 18972 12860 19024 12912
rect 9772 12835 9824 12844
rect 9772 12801 9790 12835
rect 9790 12801 9824 12835
rect 9772 12792 9824 12801
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 3424 12699 3476 12708
rect 3424 12665 3433 12699
rect 3433 12665 3467 12699
rect 3467 12665 3476 12699
rect 3424 12656 3476 12665
rect 10968 12724 11020 12776
rect 12164 12724 12216 12776
rect 13636 12792 13688 12844
rect 15016 12792 15068 12844
rect 15108 12792 15160 12844
rect 13820 12724 13872 12776
rect 14464 12767 14516 12776
rect 14464 12733 14473 12767
rect 14473 12733 14507 12767
rect 14507 12733 14516 12767
rect 14464 12724 14516 12733
rect 15568 12724 15620 12776
rect 17132 12724 17184 12776
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 19984 12835 20036 12844
rect 19984 12801 20018 12835
rect 20018 12801 20036 12835
rect 19984 12792 20036 12801
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 24032 12835 24084 12844
rect 24032 12801 24066 12835
rect 24066 12801 24084 12835
rect 24032 12792 24084 12801
rect 26148 12792 26200 12844
rect 28540 12928 28592 12980
rect 28632 12928 28684 12980
rect 29736 12928 29788 12980
rect 33508 12971 33560 12980
rect 33508 12937 33517 12971
rect 33517 12937 33551 12971
rect 33551 12937 33560 12971
rect 33508 12928 33560 12937
rect 35256 12928 35308 12980
rect 36084 12928 36136 12980
rect 36728 12928 36780 12980
rect 36820 12928 36872 12980
rect 37004 12928 37056 12980
rect 38660 12971 38712 12980
rect 38660 12937 38669 12971
rect 38669 12937 38703 12971
rect 38703 12937 38712 12971
rect 38660 12928 38712 12937
rect 38844 12928 38896 12980
rect 39672 12971 39724 12980
rect 39672 12937 39681 12971
rect 39681 12937 39715 12971
rect 39715 12937 39724 12971
rect 39672 12928 39724 12937
rect 41052 12928 41104 12980
rect 42708 12971 42760 12980
rect 42708 12937 42717 12971
rect 42717 12937 42751 12971
rect 42751 12937 42760 12971
rect 42708 12928 42760 12937
rect 43260 12928 43312 12980
rect 45560 12971 45612 12980
rect 45560 12937 45569 12971
rect 45569 12937 45603 12971
rect 45603 12937 45612 12971
rect 45560 12928 45612 12937
rect 47584 12928 47636 12980
rect 26700 12860 26752 12912
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27344 12792 27396 12801
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 18880 12724 18932 12776
rect 5724 12588 5776 12640
rect 8944 12588 8996 12640
rect 10508 12588 10560 12640
rect 11704 12588 11756 12640
rect 16212 12588 16264 12640
rect 24860 12724 24912 12776
rect 25136 12724 25188 12776
rect 26424 12724 26476 12776
rect 27528 12767 27580 12776
rect 27528 12733 27537 12767
rect 27537 12733 27571 12767
rect 27571 12733 27580 12767
rect 28816 12903 28868 12912
rect 28816 12869 28850 12903
rect 28850 12869 28868 12903
rect 28816 12860 28868 12869
rect 31852 12792 31904 12844
rect 33232 12792 33284 12844
rect 36544 12860 36596 12912
rect 34428 12792 34480 12844
rect 34612 12835 34664 12844
rect 34612 12801 34646 12835
rect 34646 12801 34664 12835
rect 34612 12792 34664 12801
rect 38752 12792 38804 12844
rect 38936 12792 38988 12844
rect 40684 12792 40736 12844
rect 41144 12792 41196 12844
rect 42892 12792 42944 12844
rect 46020 12835 46072 12844
rect 46020 12801 46054 12835
rect 46054 12801 46072 12835
rect 46020 12792 46072 12801
rect 48320 12860 48372 12912
rect 50068 12928 50120 12980
rect 50988 12928 51040 12980
rect 51816 12928 51868 12980
rect 52460 12928 52512 12980
rect 54024 12928 54076 12980
rect 54760 12928 54812 12980
rect 56600 12928 56652 12980
rect 56692 12928 56744 12980
rect 27528 12724 27580 12733
rect 21456 12588 21508 12640
rect 22100 12631 22152 12640
rect 22100 12597 22109 12631
rect 22109 12597 22143 12631
rect 22143 12597 22152 12631
rect 22100 12588 22152 12597
rect 23296 12631 23348 12640
rect 23296 12597 23305 12631
rect 23305 12597 23339 12631
rect 23339 12597 23348 12631
rect 23296 12588 23348 12597
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 27804 12656 27856 12708
rect 26976 12631 27028 12640
rect 26976 12597 26985 12631
rect 26985 12597 27019 12631
rect 27019 12597 27028 12631
rect 26976 12588 27028 12597
rect 35808 12724 35860 12776
rect 36452 12767 36504 12776
rect 36452 12733 36461 12767
rect 36461 12733 36495 12767
rect 36495 12733 36504 12767
rect 36452 12724 36504 12733
rect 36912 12724 36964 12776
rect 39304 12767 39356 12776
rect 39304 12733 39313 12767
rect 39313 12733 39347 12767
rect 39347 12733 39356 12767
rect 39304 12724 39356 12733
rect 41420 12724 41472 12776
rect 45100 12767 45152 12776
rect 45100 12733 45109 12767
rect 45109 12733 45143 12767
rect 45143 12733 45152 12767
rect 45100 12724 45152 12733
rect 45744 12767 45796 12776
rect 45744 12733 45753 12767
rect 45753 12733 45787 12767
rect 45787 12733 45796 12767
rect 45744 12724 45796 12733
rect 47492 12724 47544 12776
rect 49792 12792 49844 12844
rect 50344 12767 50396 12776
rect 50344 12733 50353 12767
rect 50353 12733 50387 12767
rect 50387 12733 50396 12767
rect 50344 12724 50396 12733
rect 53196 12835 53248 12844
rect 53196 12801 53205 12835
rect 53205 12801 53239 12835
rect 53239 12801 53248 12835
rect 53196 12792 53248 12801
rect 51172 12767 51224 12776
rect 51172 12733 51181 12767
rect 51181 12733 51215 12767
rect 51215 12733 51224 12767
rect 51172 12724 51224 12733
rect 53748 12860 53800 12912
rect 53932 12860 53984 12912
rect 54760 12792 54812 12844
rect 54668 12767 54720 12776
rect 54668 12733 54677 12767
rect 54677 12733 54711 12767
rect 54711 12733 54720 12767
rect 54668 12724 54720 12733
rect 54944 12767 54996 12776
rect 54944 12733 54953 12767
rect 54953 12733 54987 12767
rect 54987 12733 54996 12767
rect 54944 12724 54996 12733
rect 55128 12724 55180 12776
rect 33600 12631 33652 12640
rect 33600 12597 33609 12631
rect 33609 12597 33643 12631
rect 33643 12597 33652 12631
rect 33600 12588 33652 12597
rect 35716 12631 35768 12640
rect 35716 12597 35725 12631
rect 35725 12597 35759 12631
rect 35759 12597 35768 12631
rect 35716 12588 35768 12597
rect 42432 12588 42484 12640
rect 42708 12588 42760 12640
rect 44456 12631 44508 12640
rect 44456 12597 44465 12631
rect 44465 12597 44499 12631
rect 44499 12597 44508 12631
rect 44456 12588 44508 12597
rect 46756 12588 46808 12640
rect 53472 12656 53524 12708
rect 55220 12699 55272 12708
rect 55220 12665 55229 12699
rect 55229 12665 55263 12699
rect 55263 12665 55272 12699
rect 55220 12656 55272 12665
rect 55864 12767 55916 12776
rect 55864 12733 55873 12767
rect 55873 12733 55907 12767
rect 55907 12733 55916 12767
rect 55864 12724 55916 12733
rect 56508 12767 56560 12776
rect 56508 12733 56517 12767
rect 56517 12733 56551 12767
rect 56551 12733 56560 12767
rect 56508 12724 56560 12733
rect 57152 12724 57204 12776
rect 49700 12631 49752 12640
rect 49700 12597 49709 12631
rect 49709 12597 49743 12631
rect 49743 12597 49752 12631
rect 49700 12588 49752 12597
rect 51356 12588 51408 12640
rect 56140 12588 56192 12640
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 22616 12486 22668 12538
rect 22680 12486 22732 12538
rect 22744 12486 22796 12538
rect 22808 12486 22860 12538
rect 22872 12486 22924 12538
rect 37060 12486 37112 12538
rect 37124 12486 37176 12538
rect 37188 12486 37240 12538
rect 37252 12486 37304 12538
rect 37316 12486 37368 12538
rect 51504 12486 51556 12538
rect 51568 12486 51620 12538
rect 51632 12486 51684 12538
rect 51696 12486 51748 12538
rect 51760 12486 51812 12538
rect 4252 12384 4304 12436
rect 5172 12384 5224 12436
rect 9772 12384 9824 12436
rect 10600 12384 10652 12436
rect 11796 12384 11848 12436
rect 12256 12384 12308 12436
rect 14556 12384 14608 12436
rect 17500 12384 17552 12436
rect 3516 12316 3568 12368
rect 2596 12291 2648 12300
rect 2596 12257 2605 12291
rect 2605 12257 2639 12291
rect 2639 12257 2648 12291
rect 2596 12248 2648 12257
rect 6460 12316 6512 12368
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 3792 12180 3844 12232
rect 3884 12180 3936 12232
rect 5724 12180 5776 12232
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 5172 12112 5224 12164
rect 6828 12112 6880 12164
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 8944 12180 8996 12232
rect 10968 12248 11020 12300
rect 11152 12248 11204 12300
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 11796 12248 11848 12300
rect 12624 12248 12676 12300
rect 15108 12316 15160 12368
rect 17132 12316 17184 12368
rect 13912 12248 13964 12300
rect 11428 12180 11480 12232
rect 12164 12180 12216 12232
rect 9128 12112 9180 12164
rect 4160 12044 4212 12096
rect 4620 12044 4672 12096
rect 13912 12112 13964 12164
rect 15844 12248 15896 12300
rect 16212 12248 16264 12300
rect 16488 12248 16540 12300
rect 18236 12248 18288 12300
rect 19340 12248 19392 12300
rect 19708 12384 19760 12436
rect 22468 12384 22520 12436
rect 24492 12427 24544 12436
rect 24492 12393 24501 12427
rect 24501 12393 24535 12427
rect 24535 12393 24544 12427
rect 24492 12384 24544 12393
rect 26240 12384 26292 12436
rect 27528 12384 27580 12436
rect 29736 12384 29788 12436
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 19892 12112 19944 12164
rect 21272 12248 21324 12300
rect 21640 12248 21692 12300
rect 25136 12291 25188 12300
rect 25136 12257 25145 12291
rect 25145 12257 25179 12291
rect 25179 12257 25188 12291
rect 25136 12248 25188 12257
rect 26976 12291 27028 12300
rect 26976 12257 26985 12291
rect 26985 12257 27019 12291
rect 27019 12257 27028 12291
rect 26976 12248 27028 12257
rect 30380 12316 30432 12368
rect 32680 12316 32732 12368
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21916 12223 21968 12232
rect 21916 12189 21950 12223
rect 21950 12189 21968 12223
rect 21916 12180 21968 12189
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 22100 12180 22152 12189
rect 27804 12223 27856 12232
rect 27804 12189 27813 12223
rect 27813 12189 27847 12223
rect 27847 12189 27856 12223
rect 29736 12223 29788 12232
rect 27804 12180 27856 12189
rect 29736 12189 29745 12223
rect 29745 12189 29779 12223
rect 29779 12189 29788 12223
rect 29736 12180 29788 12189
rect 31576 12291 31628 12300
rect 31576 12257 31585 12291
rect 31585 12257 31619 12291
rect 31619 12257 31628 12291
rect 31576 12248 31628 12257
rect 31944 12248 31996 12300
rect 34336 12316 34388 12368
rect 34612 12316 34664 12368
rect 35164 12316 35216 12368
rect 36636 12316 36688 12368
rect 39304 12316 39356 12368
rect 41328 12359 41380 12368
rect 41328 12325 41337 12359
rect 41337 12325 41371 12359
rect 41371 12325 41380 12359
rect 41328 12316 41380 12325
rect 41604 12316 41656 12368
rect 42708 12316 42760 12368
rect 45100 12384 45152 12436
rect 47032 12427 47084 12436
rect 47032 12393 47041 12427
rect 47041 12393 47075 12427
rect 47075 12393 47084 12427
rect 47032 12384 47084 12393
rect 47308 12384 47360 12436
rect 30380 12223 30432 12232
rect 30380 12189 30389 12223
rect 30389 12189 30423 12223
rect 30423 12189 30432 12223
rect 30380 12180 30432 12189
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 33600 12248 33652 12300
rect 34060 12291 34112 12300
rect 34060 12257 34069 12291
rect 34069 12257 34103 12291
rect 34103 12257 34112 12291
rect 34060 12248 34112 12257
rect 34796 12248 34848 12300
rect 35716 12248 35768 12300
rect 35900 12248 35952 12300
rect 36728 12248 36780 12300
rect 36820 12248 36872 12300
rect 38108 12248 38160 12300
rect 38660 12291 38712 12300
rect 38660 12257 38669 12291
rect 38669 12257 38703 12291
rect 38703 12257 38712 12291
rect 38660 12248 38712 12257
rect 41512 12248 41564 12300
rect 42340 12291 42392 12300
rect 42340 12257 42349 12291
rect 42349 12257 42383 12291
rect 42383 12257 42392 12291
rect 42340 12248 42392 12257
rect 32956 12223 33008 12232
rect 32956 12189 32965 12223
rect 32965 12189 32999 12223
rect 32999 12189 33008 12223
rect 32956 12180 33008 12189
rect 37648 12180 37700 12232
rect 39948 12223 40000 12232
rect 12716 12044 12768 12096
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 14004 12044 14056 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 15200 12087 15252 12096
rect 15200 12053 15209 12087
rect 15209 12053 15243 12087
rect 15243 12053 15252 12087
rect 15200 12044 15252 12053
rect 15752 12044 15804 12096
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 19800 12044 19852 12096
rect 20812 12087 20864 12096
rect 20812 12053 20821 12087
rect 20821 12053 20855 12087
rect 20855 12053 20864 12087
rect 20812 12044 20864 12053
rect 28540 12087 28592 12096
rect 28540 12053 28549 12087
rect 28549 12053 28583 12087
rect 28583 12053 28592 12087
rect 28540 12044 28592 12053
rect 29000 12087 29052 12096
rect 29000 12053 29009 12087
rect 29009 12053 29043 12087
rect 29043 12053 29052 12087
rect 29000 12044 29052 12053
rect 29276 12044 29328 12096
rect 34152 12112 34204 12164
rect 39948 12189 39957 12223
rect 39957 12189 39991 12223
rect 39991 12189 40000 12223
rect 39948 12180 40000 12189
rect 42064 12223 42116 12232
rect 42064 12189 42073 12223
rect 42073 12189 42107 12223
rect 42107 12189 42116 12223
rect 42064 12180 42116 12189
rect 40960 12112 41012 12164
rect 43168 12180 43220 12232
rect 44456 12248 44508 12300
rect 43536 12180 43588 12232
rect 30656 12087 30708 12096
rect 30656 12053 30665 12087
rect 30665 12053 30699 12087
rect 30699 12053 30708 12087
rect 30656 12044 30708 12053
rect 30840 12044 30892 12096
rect 32956 12044 33008 12096
rect 33324 12087 33376 12096
rect 33324 12053 33333 12087
rect 33333 12053 33367 12087
rect 33367 12053 33376 12087
rect 33324 12044 33376 12053
rect 33416 12087 33468 12096
rect 33416 12053 33425 12087
rect 33425 12053 33459 12087
rect 33459 12053 33468 12087
rect 33416 12044 33468 12053
rect 35900 12044 35952 12096
rect 36452 12087 36504 12096
rect 36452 12053 36461 12087
rect 36461 12053 36495 12087
rect 36495 12053 36504 12087
rect 36452 12044 36504 12053
rect 36544 12044 36596 12096
rect 38936 12087 38988 12096
rect 38936 12053 38945 12087
rect 38945 12053 38979 12087
rect 38979 12053 38988 12087
rect 38936 12044 38988 12053
rect 39120 12044 39172 12096
rect 42432 12044 42484 12096
rect 42524 12044 42576 12096
rect 45560 12044 45612 12096
rect 46756 12248 46808 12300
rect 47676 12291 47728 12300
rect 47676 12257 47685 12291
rect 47685 12257 47719 12291
rect 47719 12257 47728 12291
rect 47676 12248 47728 12257
rect 50344 12384 50396 12436
rect 53932 12427 53984 12436
rect 53932 12393 53941 12427
rect 53941 12393 53975 12427
rect 53975 12393 53984 12427
rect 53932 12384 53984 12393
rect 54944 12384 54996 12436
rect 55496 12427 55548 12436
rect 55496 12393 55505 12427
rect 55505 12393 55539 12427
rect 55539 12393 55548 12427
rect 55496 12384 55548 12393
rect 48504 12248 48556 12300
rect 48964 12248 49016 12300
rect 51080 12180 51132 12232
rect 48412 12044 48464 12096
rect 49884 12087 49936 12096
rect 49884 12053 49893 12087
rect 49893 12053 49927 12087
rect 49927 12053 49936 12087
rect 49884 12044 49936 12053
rect 50896 12044 50948 12096
rect 51264 12044 51316 12096
rect 52368 12180 52420 12232
rect 56048 12223 56100 12232
rect 56048 12189 56057 12223
rect 56057 12189 56091 12223
rect 56091 12189 56100 12223
rect 56048 12180 56100 12189
rect 56692 12223 56744 12232
rect 56692 12189 56701 12223
rect 56701 12189 56735 12223
rect 56735 12189 56744 12223
rect 56692 12180 56744 12189
rect 55220 12112 55272 12164
rect 54392 12044 54444 12096
rect 54668 12087 54720 12096
rect 54668 12053 54677 12087
rect 54677 12053 54711 12087
rect 54711 12053 54720 12087
rect 54668 12044 54720 12053
rect 56232 12044 56284 12096
rect 57520 12044 57572 12096
rect 15394 11942 15446 11994
rect 15458 11942 15510 11994
rect 15522 11942 15574 11994
rect 15586 11942 15638 11994
rect 15650 11942 15702 11994
rect 29838 11942 29890 11994
rect 29902 11942 29954 11994
rect 29966 11942 30018 11994
rect 30030 11942 30082 11994
rect 30094 11942 30146 11994
rect 44282 11942 44334 11994
rect 44346 11942 44398 11994
rect 44410 11942 44462 11994
rect 44474 11942 44526 11994
rect 44538 11942 44590 11994
rect 58726 11942 58778 11994
rect 58790 11942 58842 11994
rect 58854 11942 58906 11994
rect 58918 11942 58970 11994
rect 58982 11942 59034 11994
rect 2964 11883 3016 11892
rect 2964 11849 2973 11883
rect 2973 11849 3007 11883
rect 3007 11849 3016 11883
rect 2964 11840 3016 11849
rect 3792 11883 3844 11892
rect 3792 11849 3801 11883
rect 3801 11849 3835 11883
rect 3835 11849 3844 11883
rect 3792 11840 3844 11849
rect 5540 11840 5592 11892
rect 5816 11840 5868 11892
rect 8208 11840 8260 11892
rect 9128 11840 9180 11892
rect 11428 11840 11480 11892
rect 11704 11840 11756 11892
rect 6460 11772 6512 11824
rect 6644 11772 6696 11824
rect 6828 11772 6880 11824
rect 10692 11772 10744 11824
rect 10784 11772 10836 11824
rect 12256 11840 12308 11892
rect 15016 11883 15068 11892
rect 15016 11849 15025 11883
rect 15025 11849 15059 11883
rect 15059 11849 15068 11883
rect 15016 11840 15068 11849
rect 15200 11840 15252 11892
rect 21916 11840 21968 11892
rect 28540 11840 28592 11892
rect 29000 11840 29052 11892
rect 30656 11840 30708 11892
rect 33324 11840 33376 11892
rect 33416 11840 33468 11892
rect 36912 11840 36964 11892
rect 38108 11840 38160 11892
rect 39120 11840 39172 11892
rect 39948 11840 40000 11892
rect 42248 11840 42300 11892
rect 42892 11840 42944 11892
rect 46020 11840 46072 11892
rect 47032 11840 47084 11892
rect 49792 11840 49844 11892
rect 50160 11840 50212 11892
rect 50896 11883 50948 11892
rect 50896 11849 50905 11883
rect 50905 11849 50939 11883
rect 50939 11849 50948 11883
rect 50896 11840 50948 11849
rect 54576 11840 54628 11892
rect 56048 11840 56100 11892
rect 56692 11840 56744 11892
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 3884 11704 3936 11756
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 10508 11704 10560 11756
rect 10968 11704 11020 11756
rect 14464 11772 14516 11824
rect 14096 11704 14148 11756
rect 20812 11772 20864 11824
rect 9588 11636 9640 11688
rect 8944 11568 8996 11620
rect 14556 11636 14608 11688
rect 31760 11772 31812 11824
rect 31852 11704 31904 11756
rect 40960 11815 41012 11824
rect 40960 11781 40969 11815
rect 40969 11781 41003 11815
rect 41003 11781 41012 11815
rect 40960 11772 41012 11781
rect 42064 11772 42116 11824
rect 34336 11704 34388 11756
rect 36176 11704 36228 11756
rect 41512 11704 41564 11756
rect 41696 11704 41748 11756
rect 49240 11704 49292 11756
rect 11796 11568 11848 11620
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 6368 11500 6420 11552
rect 7380 11500 7432 11552
rect 10600 11500 10652 11552
rect 11336 11500 11388 11552
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 13544 11500 13596 11552
rect 15844 11568 15896 11620
rect 16396 11568 16448 11620
rect 23296 11636 23348 11688
rect 23572 11679 23624 11688
rect 23572 11645 23581 11679
rect 23581 11645 23615 11679
rect 23615 11645 23624 11679
rect 23572 11636 23624 11645
rect 25412 11679 25464 11688
rect 25412 11645 25421 11679
rect 25421 11645 25455 11679
rect 25455 11645 25464 11679
rect 25412 11636 25464 11645
rect 20720 11568 20772 11620
rect 22100 11568 22152 11620
rect 25504 11568 25556 11620
rect 16028 11500 16080 11552
rect 16488 11500 16540 11552
rect 19800 11500 19852 11552
rect 20076 11543 20128 11552
rect 20076 11509 20085 11543
rect 20085 11509 20119 11543
rect 20119 11509 20128 11543
rect 20076 11500 20128 11509
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 26056 11500 26108 11552
rect 26148 11500 26200 11552
rect 28172 11500 28224 11552
rect 32588 11636 32640 11688
rect 33140 11636 33192 11688
rect 33232 11636 33284 11688
rect 31852 11568 31904 11620
rect 32864 11568 32916 11620
rect 36268 11636 36320 11688
rect 34060 11568 34112 11620
rect 38936 11611 38988 11620
rect 38936 11577 38945 11611
rect 38945 11577 38979 11611
rect 38979 11577 38988 11611
rect 38936 11568 38988 11577
rect 42524 11636 42576 11688
rect 43536 11636 43588 11688
rect 53104 11704 53156 11756
rect 56508 11704 56560 11756
rect 56968 11704 57020 11756
rect 57152 11747 57204 11756
rect 57152 11713 57161 11747
rect 57161 11713 57195 11747
rect 57195 11713 57204 11747
rect 57152 11704 57204 11713
rect 51448 11679 51500 11688
rect 51448 11645 51457 11679
rect 51457 11645 51491 11679
rect 51491 11645 51500 11679
rect 51448 11636 51500 11645
rect 52368 11636 52420 11688
rect 57428 11679 57480 11688
rect 57428 11645 57437 11679
rect 57437 11645 57471 11679
rect 57471 11645 57480 11679
rect 57428 11636 57480 11645
rect 57520 11636 57572 11688
rect 41420 11568 41472 11620
rect 46848 11568 46900 11620
rect 31300 11500 31352 11552
rect 32036 11500 32088 11552
rect 32496 11500 32548 11552
rect 35348 11543 35400 11552
rect 35348 11509 35357 11543
rect 35357 11509 35391 11543
rect 35391 11509 35400 11543
rect 35348 11500 35400 11509
rect 35716 11500 35768 11552
rect 40040 11543 40092 11552
rect 40040 11509 40049 11543
rect 40049 11509 40083 11543
rect 40083 11509 40092 11543
rect 40040 11500 40092 11509
rect 45652 11543 45704 11552
rect 45652 11509 45661 11543
rect 45661 11509 45695 11543
rect 45695 11509 45704 11543
rect 45652 11500 45704 11509
rect 51356 11500 51408 11552
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 22616 11398 22668 11450
rect 22680 11398 22732 11450
rect 22744 11398 22796 11450
rect 22808 11398 22860 11450
rect 22872 11398 22924 11450
rect 37060 11398 37112 11450
rect 37124 11398 37176 11450
rect 37188 11398 37240 11450
rect 37252 11398 37304 11450
rect 37316 11398 37368 11450
rect 51504 11398 51556 11450
rect 51568 11398 51620 11450
rect 51632 11398 51684 11450
rect 51696 11398 51748 11450
rect 51760 11398 51812 11450
rect 4620 11296 4672 11348
rect 4160 11271 4212 11280
rect 4160 11237 4169 11271
rect 4169 11237 4203 11271
rect 4203 11237 4212 11271
rect 4160 11228 4212 11237
rect 6460 11228 6512 11280
rect 3792 11067 3844 11076
rect 3792 11033 3801 11067
rect 3801 11033 3835 11067
rect 3835 11033 3844 11067
rect 3792 11024 3844 11033
rect 4712 11160 4764 11212
rect 5724 11160 5776 11212
rect 6828 11160 6880 11212
rect 11152 11296 11204 11348
rect 13360 11296 13412 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16028 11296 16080 11348
rect 19892 11339 19944 11348
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 20076 11296 20128 11348
rect 22284 11296 22336 11348
rect 25412 11339 25464 11348
rect 25412 11305 25421 11339
rect 25421 11305 25455 11339
rect 25455 11305 25464 11339
rect 25412 11296 25464 11305
rect 30380 11296 30432 11348
rect 32588 11339 32640 11348
rect 32588 11305 32597 11339
rect 32597 11305 32631 11339
rect 32631 11305 32640 11339
rect 32588 11296 32640 11305
rect 32772 11339 32824 11348
rect 32772 11305 32781 11339
rect 32781 11305 32815 11339
rect 32815 11305 32824 11339
rect 32772 11296 32824 11305
rect 2596 10956 2648 11008
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 6644 11092 6696 11144
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 4252 10956 4304 11008
rect 4436 10956 4488 11008
rect 5816 11024 5868 11076
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 9588 11024 9640 11076
rect 10784 11160 10836 11212
rect 12072 11228 12124 11280
rect 12164 11160 12216 11212
rect 14188 11228 14240 11280
rect 14372 11228 14424 11280
rect 21916 11228 21968 11280
rect 27252 11228 27304 11280
rect 35716 11228 35768 11280
rect 40132 11296 40184 11348
rect 42248 11339 42300 11348
rect 42248 11305 42257 11339
rect 42257 11305 42291 11339
rect 42291 11305 42300 11339
rect 42248 11296 42300 11305
rect 42616 11339 42668 11348
rect 42616 11305 42625 11339
rect 42625 11305 42659 11339
rect 42659 11305 42668 11339
rect 42616 11296 42668 11305
rect 43536 11296 43588 11348
rect 57060 11296 57112 11348
rect 45652 11228 45704 11280
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 15200 11092 15252 11144
rect 17868 11092 17920 11144
rect 18236 11092 18288 11144
rect 22008 11160 22060 11212
rect 24124 11160 24176 11212
rect 26148 11160 26200 11212
rect 36084 11160 36136 11212
rect 36820 11160 36872 11212
rect 21916 11092 21968 11144
rect 22560 11135 22612 11144
rect 22560 11101 22569 11135
rect 22569 11101 22603 11135
rect 22603 11101 22612 11135
rect 22560 11092 22612 11101
rect 24216 11092 24268 11144
rect 24860 11092 24912 11144
rect 25596 11092 25648 11144
rect 26424 11092 26476 11144
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 33600 11135 33652 11144
rect 33600 11101 33609 11135
rect 33609 11101 33643 11135
rect 33643 11101 33652 11135
rect 33600 11092 33652 11101
rect 34336 11135 34388 11144
rect 34336 11101 34345 11135
rect 34345 11101 34379 11135
rect 34379 11101 34388 11135
rect 34336 11092 34388 11101
rect 35348 11135 35400 11144
rect 35348 11101 35357 11135
rect 35357 11101 35391 11135
rect 35391 11101 35400 11135
rect 35348 11092 35400 11101
rect 36452 11092 36504 11144
rect 36728 11092 36780 11144
rect 37280 11092 37332 11144
rect 38752 11135 38804 11144
rect 38752 11101 38761 11135
rect 38761 11101 38795 11135
rect 38795 11101 38804 11135
rect 38752 11092 38804 11101
rect 39580 11135 39632 11144
rect 39580 11101 39589 11135
rect 39589 11101 39623 11135
rect 39623 11101 39632 11135
rect 39580 11092 39632 11101
rect 40132 11092 40184 11144
rect 41236 11092 41288 11144
rect 43812 11135 43864 11144
rect 43812 11101 43821 11135
rect 43821 11101 43855 11135
rect 43855 11101 43864 11135
rect 43812 11092 43864 11101
rect 44180 11092 44232 11144
rect 44824 11092 44876 11144
rect 45836 11135 45888 11144
rect 45836 11101 45845 11135
rect 45845 11101 45879 11135
rect 45879 11101 45888 11135
rect 45836 11092 45888 11101
rect 47032 11135 47084 11144
rect 47032 11101 47041 11135
rect 47041 11101 47075 11135
rect 47075 11101 47084 11135
rect 47032 11092 47084 11101
rect 10876 11024 10928 11076
rect 11612 11024 11664 11076
rect 12256 11024 12308 11076
rect 13176 11067 13228 11076
rect 13176 11033 13185 11067
rect 13185 11033 13219 11067
rect 13219 11033 13228 11067
rect 13176 11024 13228 11033
rect 14004 11024 14056 11076
rect 16488 11024 16540 11076
rect 18052 11024 18104 11076
rect 20812 11067 20864 11076
rect 20812 11033 20821 11067
rect 20821 11033 20855 11067
rect 20855 11033 20864 11067
rect 20812 11024 20864 11033
rect 23112 11024 23164 11076
rect 5172 10956 5224 11008
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 7840 10999 7892 11008
rect 7840 10965 7849 10999
rect 7849 10965 7883 10999
rect 7883 10965 7892 10999
rect 7840 10956 7892 10965
rect 11060 10999 11112 11008
rect 11060 10965 11069 10999
rect 11069 10965 11103 10999
rect 11103 10965 11112 10999
rect 11060 10956 11112 10965
rect 15016 10956 15068 11008
rect 17684 10956 17736 11008
rect 22008 10999 22060 11008
rect 22008 10965 22017 10999
rect 22017 10965 22051 10999
rect 22051 10965 22060 10999
rect 22008 10956 22060 10965
rect 25504 10956 25556 11008
rect 28540 11067 28592 11076
rect 28540 11033 28549 11067
rect 28549 11033 28583 11067
rect 28583 11033 28592 11067
rect 28540 11024 28592 11033
rect 33324 11024 33376 11076
rect 26332 10956 26384 11008
rect 32680 10956 32732 11008
rect 33232 10956 33284 11008
rect 33784 10999 33836 11008
rect 33784 10965 33793 10999
rect 33793 10965 33827 10999
rect 33827 10965 33836 10999
rect 33784 10956 33836 10965
rect 34888 10999 34940 11008
rect 34888 10965 34897 10999
rect 34897 10965 34931 10999
rect 34931 10965 34940 10999
rect 34888 10956 34940 10965
rect 36820 11024 36872 11076
rect 40408 11067 40460 11076
rect 40408 11033 40417 11067
rect 40417 11033 40451 11067
rect 40451 11033 40460 11067
rect 40408 11024 40460 11033
rect 42064 11024 42116 11076
rect 35440 10956 35492 11008
rect 35808 10956 35860 11008
rect 36452 10999 36504 11008
rect 36452 10965 36461 10999
rect 36461 10965 36495 10999
rect 36495 10965 36504 10999
rect 36452 10956 36504 10965
rect 36636 10956 36688 11008
rect 38200 10999 38252 11008
rect 38200 10965 38209 10999
rect 38209 10965 38243 10999
rect 38243 10965 38252 10999
rect 38200 10956 38252 10965
rect 39028 10956 39080 11008
rect 41144 10956 41196 11008
rect 41328 10999 41380 11008
rect 41328 10965 41337 10999
rect 41337 10965 41371 10999
rect 41371 10965 41380 10999
rect 41328 10956 41380 10965
rect 43168 10999 43220 11008
rect 43168 10965 43177 10999
rect 43177 10965 43211 10999
rect 43211 10965 43220 10999
rect 43168 10956 43220 10965
rect 43904 10999 43956 11008
rect 43904 10965 43913 10999
rect 43913 10965 43947 10999
rect 43947 10965 43956 10999
rect 43904 10956 43956 10965
rect 44640 10956 44692 11008
rect 46204 10956 46256 11008
rect 46480 10999 46532 11008
rect 46480 10965 46489 10999
rect 46489 10965 46523 10999
rect 46523 10965 46532 10999
rect 46480 10956 46532 10965
rect 50344 11160 50396 11212
rect 50620 11160 50672 11212
rect 52092 11160 52144 11212
rect 56784 11203 56836 11212
rect 56784 11169 56793 11203
rect 56793 11169 56827 11203
rect 56827 11169 56836 11203
rect 56784 11160 56836 11169
rect 50712 11135 50764 11144
rect 50712 11101 50721 11135
rect 50721 11101 50755 11135
rect 50755 11101 50764 11135
rect 50712 11092 50764 11101
rect 52184 11135 52236 11144
rect 52184 11101 52193 11135
rect 52193 11101 52227 11135
rect 52227 11101 52236 11135
rect 52184 11092 52236 11101
rect 56140 11092 56192 11144
rect 49608 11024 49660 11076
rect 51080 11024 51132 11076
rect 54392 11024 54444 11076
rect 56784 11024 56836 11076
rect 48320 10956 48372 11008
rect 48504 10956 48556 11008
rect 50160 10999 50212 11008
rect 50160 10965 50169 10999
rect 50169 10965 50203 10999
rect 50203 10965 50212 10999
rect 50160 10956 50212 10965
rect 51172 10956 51224 11008
rect 56232 10956 56284 11008
rect 56876 10999 56928 11008
rect 56876 10965 56885 10999
rect 56885 10965 56919 10999
rect 56919 10965 56928 10999
rect 56876 10956 56928 10965
rect 57336 10999 57388 11008
rect 57336 10965 57345 10999
rect 57345 10965 57379 10999
rect 57379 10965 57388 10999
rect 57336 10956 57388 10965
rect 15394 10854 15446 10906
rect 15458 10854 15510 10906
rect 15522 10854 15574 10906
rect 15586 10854 15638 10906
rect 15650 10854 15702 10906
rect 29838 10854 29890 10906
rect 29902 10854 29954 10906
rect 29966 10854 30018 10906
rect 30030 10854 30082 10906
rect 30094 10854 30146 10906
rect 44282 10854 44334 10906
rect 44346 10854 44398 10906
rect 44410 10854 44462 10906
rect 44474 10854 44526 10906
rect 44538 10854 44590 10906
rect 58726 10854 58778 10906
rect 58790 10854 58842 10906
rect 58854 10854 58906 10906
rect 58918 10854 58970 10906
rect 58982 10854 59034 10906
rect 5356 10795 5408 10804
rect 5356 10761 5365 10795
rect 5365 10761 5399 10795
rect 5399 10761 5408 10795
rect 5356 10752 5408 10761
rect 5172 10684 5224 10736
rect 3516 10548 3568 10600
rect 3700 10591 3752 10600
rect 3700 10557 3709 10591
rect 3709 10557 3743 10591
rect 3743 10557 3752 10591
rect 3700 10548 3752 10557
rect 1584 10480 1636 10532
rect 2688 10480 2740 10532
rect 4896 10616 4948 10668
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 6000 10548 6052 10600
rect 6644 10752 6696 10804
rect 7840 10752 7892 10804
rect 10140 10752 10192 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 12624 10752 12676 10804
rect 15016 10752 15068 10804
rect 17040 10752 17092 10804
rect 18236 10752 18288 10804
rect 9036 10684 9088 10736
rect 20536 10684 20588 10736
rect 30748 10684 30800 10736
rect 33784 10684 33836 10736
rect 34244 10684 34296 10736
rect 8944 10616 8996 10668
rect 11060 10659 11112 10668
rect 11060 10625 11069 10659
rect 11069 10625 11103 10659
rect 11103 10625 11112 10659
rect 11060 10616 11112 10625
rect 10600 10548 10652 10600
rect 11520 10548 11572 10600
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 12624 10548 12676 10600
rect 14556 10616 14608 10668
rect 5724 10523 5776 10532
rect 5724 10489 5733 10523
rect 5733 10489 5767 10523
rect 5767 10489 5776 10523
rect 5724 10480 5776 10489
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 4988 10412 5040 10464
rect 5264 10412 5316 10464
rect 5908 10412 5960 10464
rect 13544 10548 13596 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 23480 10616 23532 10668
rect 24676 10659 24728 10668
rect 24676 10625 24685 10659
rect 24685 10625 24719 10659
rect 24719 10625 24728 10659
rect 24676 10616 24728 10625
rect 16856 10548 16908 10600
rect 19984 10548 20036 10600
rect 21916 10591 21968 10600
rect 21916 10557 21925 10591
rect 21925 10557 21959 10591
rect 21959 10557 21968 10591
rect 21916 10548 21968 10557
rect 22100 10591 22152 10600
rect 22100 10557 22109 10591
rect 22109 10557 22143 10591
rect 22143 10557 22152 10591
rect 22100 10548 22152 10557
rect 24032 10591 24084 10600
rect 24032 10557 24041 10591
rect 24041 10557 24075 10591
rect 24075 10557 24084 10591
rect 24032 10548 24084 10557
rect 24124 10548 24176 10600
rect 25688 10616 25740 10668
rect 26056 10659 26108 10668
rect 26056 10625 26074 10659
rect 26074 10625 26108 10659
rect 26056 10616 26108 10625
rect 30564 10616 30616 10668
rect 31208 10616 31260 10668
rect 26332 10591 26384 10600
rect 26332 10557 26341 10591
rect 26341 10557 26375 10591
rect 26375 10557 26384 10591
rect 26332 10548 26384 10557
rect 19616 10480 19668 10532
rect 21824 10480 21876 10532
rect 23296 10480 23348 10532
rect 23572 10480 23624 10532
rect 26424 10480 26476 10532
rect 10508 10412 10560 10464
rect 14188 10412 14240 10464
rect 15292 10412 15344 10464
rect 15384 10412 15436 10464
rect 15844 10412 15896 10464
rect 16028 10412 16080 10464
rect 19432 10412 19484 10464
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 24584 10412 24636 10464
rect 29000 10548 29052 10600
rect 29276 10591 29328 10600
rect 29276 10557 29285 10591
rect 29285 10557 29319 10591
rect 29319 10557 29328 10591
rect 29276 10548 29328 10557
rect 29460 10548 29512 10600
rect 34888 10616 34940 10668
rect 36452 10684 36504 10736
rect 36544 10727 36596 10736
rect 36544 10693 36553 10727
rect 36553 10693 36587 10727
rect 36587 10693 36596 10727
rect 36544 10684 36596 10693
rect 36912 10684 36964 10736
rect 33968 10548 34020 10600
rect 36360 10659 36412 10668
rect 36360 10625 36369 10659
rect 36369 10625 36403 10659
rect 36403 10625 36412 10659
rect 36360 10616 36412 10625
rect 38200 10684 38252 10736
rect 40500 10752 40552 10804
rect 42248 10795 42300 10804
rect 42248 10761 42257 10795
rect 42257 10761 42291 10795
rect 42291 10761 42300 10795
rect 42248 10752 42300 10761
rect 43812 10795 43864 10804
rect 43812 10761 43821 10795
rect 43821 10761 43855 10795
rect 43855 10761 43864 10795
rect 43812 10752 43864 10761
rect 45836 10752 45888 10804
rect 49608 10752 49660 10804
rect 36820 10548 36872 10600
rect 38936 10616 38988 10668
rect 39120 10591 39172 10600
rect 39120 10557 39129 10591
rect 39129 10557 39163 10591
rect 39163 10557 39172 10591
rect 39120 10548 39172 10557
rect 39304 10659 39356 10668
rect 39304 10625 39313 10659
rect 39313 10625 39347 10659
rect 39347 10625 39356 10659
rect 39304 10616 39356 10625
rect 41328 10616 41380 10668
rect 33232 10480 33284 10532
rect 33600 10480 33652 10532
rect 37280 10480 37332 10532
rect 43904 10616 43956 10668
rect 45652 10684 45704 10736
rect 44640 10616 44692 10668
rect 46480 10684 46532 10736
rect 46664 10684 46716 10736
rect 48228 10684 48280 10736
rect 49056 10727 49108 10736
rect 49056 10693 49065 10727
rect 49065 10693 49099 10727
rect 49099 10693 49108 10727
rect 49056 10684 49108 10693
rect 46112 10616 46164 10668
rect 41604 10548 41656 10600
rect 41788 10591 41840 10600
rect 41788 10557 41797 10591
rect 41797 10557 41831 10591
rect 41831 10557 41840 10591
rect 41788 10548 41840 10557
rect 26700 10455 26752 10464
rect 26700 10421 26709 10455
rect 26709 10421 26743 10455
rect 26743 10421 26752 10455
rect 26700 10412 26752 10421
rect 29092 10412 29144 10464
rect 30840 10412 30892 10464
rect 31852 10455 31904 10464
rect 31852 10421 31861 10455
rect 31861 10421 31895 10455
rect 31895 10421 31904 10455
rect 31852 10412 31904 10421
rect 33048 10412 33100 10464
rect 37648 10412 37700 10464
rect 39580 10412 39632 10464
rect 40132 10412 40184 10464
rect 41880 10412 41932 10464
rect 48320 10548 48372 10600
rect 49884 10684 49936 10736
rect 50160 10684 50212 10736
rect 50620 10795 50672 10804
rect 50620 10761 50629 10795
rect 50629 10761 50663 10795
rect 50663 10761 50672 10795
rect 50620 10752 50672 10761
rect 50712 10795 50764 10804
rect 50712 10761 50721 10795
rect 50721 10761 50755 10795
rect 50755 10761 50764 10795
rect 50712 10752 50764 10761
rect 51172 10795 51224 10804
rect 51172 10761 51181 10795
rect 51181 10761 51215 10795
rect 51215 10761 51224 10795
rect 51172 10752 51224 10761
rect 52184 10752 52236 10804
rect 54208 10752 54260 10804
rect 56876 10752 56928 10804
rect 51816 10684 51868 10736
rect 51908 10659 51960 10668
rect 51908 10625 51917 10659
rect 51917 10625 51951 10659
rect 51951 10625 51960 10659
rect 51908 10616 51960 10625
rect 52644 10616 52696 10668
rect 57520 10659 57572 10668
rect 57520 10625 57529 10659
rect 57529 10625 57563 10659
rect 57563 10625 57572 10659
rect 57520 10616 57572 10625
rect 51356 10591 51408 10600
rect 51356 10557 51365 10591
rect 51365 10557 51399 10591
rect 51399 10557 51408 10591
rect 51356 10548 51408 10557
rect 52368 10548 52420 10600
rect 52552 10548 52604 10600
rect 54116 10591 54168 10600
rect 54116 10557 54125 10591
rect 54125 10557 54159 10591
rect 54159 10557 54168 10591
rect 54116 10548 54168 10557
rect 54760 10591 54812 10600
rect 54760 10557 54769 10591
rect 54769 10557 54803 10591
rect 54803 10557 54812 10591
rect 54760 10548 54812 10557
rect 55496 10591 55548 10600
rect 55496 10557 55505 10591
rect 55505 10557 55539 10591
rect 55539 10557 55548 10591
rect 55496 10548 55548 10557
rect 56324 10591 56376 10600
rect 56324 10557 56333 10591
rect 56333 10557 56367 10591
rect 56367 10557 56376 10591
rect 56324 10548 56376 10557
rect 56416 10548 56468 10600
rect 56600 10591 56652 10600
rect 56600 10557 56609 10591
rect 56609 10557 56643 10591
rect 56643 10557 56652 10591
rect 56600 10548 56652 10557
rect 56784 10548 56836 10600
rect 57336 10591 57388 10600
rect 57336 10557 57345 10591
rect 57345 10557 57379 10591
rect 57379 10557 57388 10591
rect 57336 10548 57388 10557
rect 58440 10591 58492 10600
rect 58440 10557 58449 10591
rect 58449 10557 58483 10591
rect 58483 10557 58492 10591
rect 58440 10548 58492 10557
rect 48228 10455 48280 10464
rect 48228 10421 48237 10455
rect 48237 10421 48271 10455
rect 48271 10421 48280 10455
rect 48228 10412 48280 10421
rect 48504 10455 48556 10464
rect 48504 10421 48513 10455
rect 48513 10421 48547 10455
rect 48547 10421 48556 10455
rect 48504 10412 48556 10421
rect 51816 10412 51868 10464
rect 54668 10480 54720 10532
rect 52000 10412 52052 10464
rect 53472 10455 53524 10464
rect 53472 10421 53481 10455
rect 53481 10421 53515 10455
rect 53515 10421 53524 10455
rect 53472 10412 53524 10421
rect 54208 10455 54260 10464
rect 54208 10421 54217 10455
rect 54217 10421 54251 10455
rect 54251 10421 54260 10455
rect 54208 10412 54260 10421
rect 54944 10455 54996 10464
rect 54944 10421 54953 10455
rect 54953 10421 54987 10455
rect 54987 10421 54996 10455
rect 54944 10412 54996 10421
rect 57888 10455 57940 10464
rect 57888 10421 57897 10455
rect 57897 10421 57931 10455
rect 57931 10421 57940 10455
rect 57888 10412 57940 10421
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 22616 10310 22668 10362
rect 22680 10310 22732 10362
rect 22744 10310 22796 10362
rect 22808 10310 22860 10362
rect 22872 10310 22924 10362
rect 37060 10310 37112 10362
rect 37124 10310 37176 10362
rect 37188 10310 37240 10362
rect 37252 10310 37304 10362
rect 37316 10310 37368 10362
rect 51504 10310 51556 10362
rect 51568 10310 51620 10362
rect 51632 10310 51684 10362
rect 51696 10310 51748 10362
rect 51760 10310 51812 10362
rect 2688 10208 2740 10260
rect 2136 10072 2188 10124
rect 2412 10072 2464 10124
rect 3516 10251 3568 10260
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 3700 10208 3752 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 4528 10140 4580 10192
rect 5448 10140 5500 10192
rect 5816 10251 5868 10260
rect 5816 10217 5825 10251
rect 5825 10217 5859 10251
rect 5859 10217 5868 10251
rect 5816 10208 5868 10217
rect 5908 10208 5960 10260
rect 6460 10183 6512 10192
rect 6460 10149 6469 10183
rect 6469 10149 6503 10183
rect 6503 10149 6512 10183
rect 6460 10140 6512 10149
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 4252 10004 4304 10056
rect 4712 10004 4764 10056
rect 6828 10208 6880 10260
rect 9036 10208 9088 10260
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 9772 10208 9824 10260
rect 12072 10208 12124 10260
rect 12164 10208 12216 10260
rect 8668 10140 8720 10192
rect 9496 10140 9548 10192
rect 13544 10208 13596 10260
rect 15016 10208 15068 10260
rect 5724 10072 5776 10124
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 14464 10072 14516 10124
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 14096 10004 14148 10056
rect 15936 10208 15988 10260
rect 15844 10072 15896 10124
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 21088 10208 21140 10260
rect 24032 10208 24084 10260
rect 24124 10251 24176 10260
rect 24124 10217 24133 10251
rect 24133 10217 24167 10251
rect 24167 10217 24176 10251
rect 24124 10208 24176 10217
rect 19984 10072 20036 10124
rect 24584 10208 24636 10260
rect 24676 10208 24728 10260
rect 25136 10115 25188 10124
rect 25136 10081 25145 10115
rect 25145 10081 25179 10115
rect 25179 10081 25188 10115
rect 25136 10072 25188 10081
rect 25688 10115 25740 10124
rect 25688 10081 25697 10115
rect 25697 10081 25731 10115
rect 25731 10081 25740 10115
rect 25688 10072 25740 10081
rect 26516 10072 26568 10124
rect 27436 10115 27488 10124
rect 27436 10081 27445 10115
rect 27445 10081 27479 10115
rect 27479 10081 27488 10115
rect 27436 10072 27488 10081
rect 31116 10115 31168 10124
rect 31116 10081 31125 10115
rect 31125 10081 31159 10115
rect 31159 10081 31168 10115
rect 34888 10208 34940 10260
rect 35624 10208 35676 10260
rect 34336 10140 34388 10192
rect 36176 10208 36228 10260
rect 36452 10208 36504 10260
rect 38752 10208 38804 10260
rect 41788 10208 41840 10260
rect 44180 10208 44232 10260
rect 31116 10072 31168 10081
rect 34244 10115 34296 10124
rect 34244 10081 34253 10115
rect 34253 10081 34287 10115
rect 34287 10081 34296 10115
rect 34244 10072 34296 10081
rect 35900 10115 35952 10124
rect 35900 10081 35909 10115
rect 35909 10081 35943 10115
rect 35943 10081 35952 10115
rect 35900 10072 35952 10081
rect 15384 10047 15436 10056
rect 15384 10013 15402 10047
rect 15402 10013 15436 10047
rect 15384 10004 15436 10013
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 16580 10004 16632 10056
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 20076 10047 20128 10056
rect 20076 10013 20085 10047
rect 20085 10013 20119 10047
rect 20119 10013 20128 10047
rect 20076 10004 20128 10013
rect 22008 10047 22060 10056
rect 22008 10013 22026 10047
rect 22026 10013 22060 10047
rect 22008 10004 22060 10013
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 23204 10004 23256 10056
rect 24860 10004 24912 10056
rect 25504 10047 25556 10056
rect 25504 10013 25538 10047
rect 25538 10013 25556 10047
rect 25504 10004 25556 10013
rect 26608 10004 26660 10056
rect 5264 9936 5316 9988
rect 12992 9936 13044 9988
rect 18052 9936 18104 9988
rect 23020 9936 23072 9988
rect 10324 9911 10376 9920
rect 10324 9877 10333 9911
rect 10333 9877 10367 9911
rect 10367 9877 10376 9911
rect 10324 9868 10376 9877
rect 15752 9868 15804 9920
rect 19524 9911 19576 9920
rect 19524 9877 19533 9911
rect 19533 9877 19567 9911
rect 19567 9877 19576 9911
rect 19524 9868 19576 9877
rect 19616 9868 19668 9920
rect 26148 9868 26200 9920
rect 26240 9868 26292 9920
rect 32680 10004 32732 10056
rect 33968 10047 34020 10056
rect 33968 10013 33977 10047
rect 33977 10013 34011 10047
rect 34011 10013 34020 10047
rect 33968 10004 34020 10013
rect 34428 10004 34480 10056
rect 35348 10047 35400 10056
rect 35348 10013 35357 10047
rect 35357 10013 35391 10047
rect 35391 10013 35400 10047
rect 35348 10004 35400 10013
rect 35624 10047 35676 10056
rect 35624 10013 35633 10047
rect 35633 10013 35667 10047
rect 35667 10013 35676 10047
rect 35624 10004 35676 10013
rect 36636 10072 36688 10124
rect 39028 10115 39080 10124
rect 39028 10081 39037 10115
rect 39037 10081 39071 10115
rect 39071 10081 39080 10115
rect 39028 10072 39080 10081
rect 39212 10115 39264 10124
rect 39212 10081 39221 10115
rect 39221 10081 39255 10115
rect 39255 10081 39264 10115
rect 39212 10072 39264 10081
rect 41328 10115 41380 10124
rect 41328 10081 41337 10115
rect 41337 10081 41371 10115
rect 41371 10081 41380 10115
rect 41328 10072 41380 10081
rect 41512 10072 41564 10124
rect 41880 10115 41932 10124
rect 41880 10081 41889 10115
rect 41889 10081 41923 10115
rect 41923 10081 41932 10115
rect 41880 10072 41932 10081
rect 45652 10140 45704 10192
rect 43168 10072 43220 10124
rect 45192 10072 45244 10124
rect 46388 10208 46440 10260
rect 46480 10208 46532 10260
rect 46112 10140 46164 10192
rect 48504 10208 48556 10260
rect 49056 10208 49108 10260
rect 50436 10208 50488 10260
rect 52460 10208 52512 10260
rect 52644 10208 52696 10260
rect 54116 10251 54168 10260
rect 54116 10217 54125 10251
rect 54125 10217 54159 10251
rect 54159 10217 54168 10251
rect 54116 10208 54168 10217
rect 54208 10208 54260 10260
rect 55496 10208 55548 10260
rect 52000 10183 52052 10192
rect 52000 10149 52009 10183
rect 52009 10149 52043 10183
rect 52043 10149 52052 10183
rect 52000 10140 52052 10149
rect 47768 10115 47820 10124
rect 47768 10081 47777 10115
rect 47777 10081 47811 10115
rect 47811 10081 47820 10115
rect 47768 10072 47820 10081
rect 48228 10072 48280 10124
rect 51264 10072 51316 10124
rect 28448 9936 28500 9988
rect 30748 9936 30800 9988
rect 34520 9936 34572 9988
rect 36544 10047 36596 10056
rect 36544 10013 36553 10047
rect 36553 10013 36587 10047
rect 36587 10013 36596 10047
rect 36544 10004 36596 10013
rect 36820 10004 36872 10056
rect 41144 10004 41196 10056
rect 41604 10004 41656 10056
rect 42524 10004 42576 10056
rect 28172 9868 28224 9920
rect 29368 9911 29420 9920
rect 29368 9877 29377 9911
rect 29377 9877 29411 9911
rect 29411 9877 29420 9911
rect 29368 9868 29420 9877
rect 29644 9868 29696 9920
rect 33600 9911 33652 9920
rect 33600 9877 33609 9911
rect 33609 9877 33643 9911
rect 33643 9877 33652 9911
rect 33600 9868 33652 9877
rect 34704 9911 34756 9920
rect 34704 9877 34713 9911
rect 34713 9877 34747 9911
rect 34747 9877 34756 9911
rect 34704 9868 34756 9877
rect 37004 9936 37056 9988
rect 37556 9936 37608 9988
rect 37648 9936 37700 9988
rect 41512 9936 41564 9988
rect 46848 10047 46900 10056
rect 46848 10013 46857 10047
rect 46857 10013 46891 10047
rect 46891 10013 46900 10047
rect 46848 10004 46900 10013
rect 47584 10047 47636 10056
rect 47584 10013 47593 10047
rect 47593 10013 47627 10047
rect 47627 10013 47636 10047
rect 47584 10004 47636 10013
rect 44088 9936 44140 9988
rect 46020 9936 46072 9988
rect 35624 9868 35676 9920
rect 35808 9868 35860 9920
rect 37464 9868 37516 9920
rect 38476 9911 38528 9920
rect 38476 9877 38485 9911
rect 38485 9877 38519 9911
rect 38519 9877 38528 9911
rect 38476 9868 38528 9877
rect 38660 9868 38712 9920
rect 39120 9868 39172 9920
rect 42800 9868 42852 9920
rect 45008 9911 45060 9920
rect 45008 9877 45017 9911
rect 45017 9877 45051 9911
rect 45051 9877 45060 9911
rect 45008 9868 45060 9877
rect 45468 9911 45520 9920
rect 45468 9877 45477 9911
rect 45477 9877 45511 9911
rect 45511 9877 45520 9911
rect 45468 9868 45520 9877
rect 47860 9911 47912 9920
rect 47860 9877 47869 9911
rect 47869 9877 47903 9911
rect 47903 9877 47912 9911
rect 47860 9868 47912 9877
rect 48320 9936 48372 9988
rect 49148 9936 49200 9988
rect 49976 10047 50028 10056
rect 49976 10013 49985 10047
rect 49985 10013 50019 10047
rect 50019 10013 50028 10047
rect 49976 10004 50028 10013
rect 51448 10047 51500 10056
rect 51448 10013 51457 10047
rect 51457 10013 51491 10047
rect 51491 10013 51500 10047
rect 51448 10004 51500 10013
rect 51632 10047 51684 10056
rect 51632 10013 51650 10047
rect 51650 10013 51684 10047
rect 51632 10004 51684 10013
rect 50344 9979 50396 9988
rect 50344 9945 50353 9979
rect 50353 9945 50387 9979
rect 50387 9945 50396 9979
rect 50344 9936 50396 9945
rect 52736 10047 52788 10056
rect 52736 10013 52745 10047
rect 52745 10013 52779 10047
rect 52779 10013 52788 10047
rect 52736 10004 52788 10013
rect 53472 9936 53524 9988
rect 53840 9936 53892 9988
rect 56692 10072 56744 10124
rect 55128 10004 55180 10056
rect 55404 9936 55456 9988
rect 56048 9936 56100 9988
rect 57612 9936 57664 9988
rect 48412 9868 48464 9920
rect 49332 9911 49384 9920
rect 49332 9877 49341 9911
rect 49341 9877 49375 9911
rect 49375 9877 49384 9911
rect 49332 9868 49384 9877
rect 50436 9868 50488 9920
rect 51448 9868 51500 9920
rect 56416 9868 56468 9920
rect 56692 9911 56744 9920
rect 56692 9877 56701 9911
rect 56701 9877 56735 9911
rect 56735 9877 56744 9911
rect 56692 9868 56744 9877
rect 58164 9911 58216 9920
rect 58164 9877 58173 9911
rect 58173 9877 58207 9911
rect 58207 9877 58216 9911
rect 58164 9868 58216 9877
rect 15394 9766 15446 9818
rect 15458 9766 15510 9818
rect 15522 9766 15574 9818
rect 15586 9766 15638 9818
rect 15650 9766 15702 9818
rect 29838 9766 29890 9818
rect 29902 9766 29954 9818
rect 29966 9766 30018 9818
rect 30030 9766 30082 9818
rect 30094 9766 30146 9818
rect 44282 9766 44334 9818
rect 44346 9766 44398 9818
rect 44410 9766 44462 9818
rect 44474 9766 44526 9818
rect 44538 9766 44590 9818
rect 58726 9766 58778 9818
rect 58790 9766 58842 9818
rect 58854 9766 58906 9818
rect 58918 9766 58970 9818
rect 58982 9766 59034 9818
rect 4252 9707 4304 9716
rect 4252 9673 4261 9707
rect 4261 9673 4295 9707
rect 4295 9673 4304 9707
rect 4252 9664 4304 9673
rect 4804 9664 4856 9716
rect 5448 9664 5500 9716
rect 12992 9707 13044 9716
rect 12992 9673 13001 9707
rect 13001 9673 13035 9707
rect 13035 9673 13044 9707
rect 12992 9664 13044 9673
rect 18236 9664 18288 9716
rect 25228 9664 25280 9716
rect 29460 9707 29512 9716
rect 29460 9673 29469 9707
rect 29469 9673 29503 9707
rect 29503 9673 29512 9707
rect 29460 9664 29512 9673
rect 34704 9664 34756 9716
rect 36176 9664 36228 9716
rect 36636 9664 36688 9716
rect 37004 9664 37056 9716
rect 37832 9664 37884 9716
rect 3056 9596 3108 9648
rect 4160 9596 4212 9648
rect 2044 9528 2096 9580
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 4988 9639 5040 9648
rect 4988 9605 4997 9639
rect 4997 9605 5031 9639
rect 5031 9605 5040 9639
rect 4988 9596 5040 9605
rect 5172 9639 5224 9648
rect 5172 9605 5181 9639
rect 5181 9605 5215 9639
rect 5215 9605 5224 9639
rect 5172 9596 5224 9605
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 39304 9664 39356 9716
rect 5816 9596 5868 9648
rect 8760 9596 8812 9648
rect 10324 9596 10376 9648
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 10048 9528 10100 9580
rect 12624 9528 12676 9580
rect 15292 9596 15344 9648
rect 17684 9596 17736 9648
rect 13176 9528 13228 9580
rect 14464 9528 14516 9580
rect 17960 9528 18012 9580
rect 19248 9596 19300 9648
rect 19524 9596 19576 9648
rect 22284 9639 22336 9648
rect 22284 9605 22293 9639
rect 22293 9605 22327 9639
rect 22327 9605 22336 9639
rect 22284 9596 22336 9605
rect 25504 9596 25556 9648
rect 27068 9596 27120 9648
rect 28540 9596 28592 9648
rect 18328 9528 18380 9580
rect 35440 9596 35492 9648
rect 23020 9528 23072 9580
rect 23480 9528 23532 9580
rect 26516 9528 26568 9580
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 29644 9528 29696 9580
rect 3332 9435 3384 9444
rect 3332 9401 3341 9435
rect 3341 9401 3375 9435
rect 3375 9401 3384 9435
rect 3332 9392 3384 9401
rect 3792 9392 3844 9444
rect 7564 9460 7616 9512
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 9680 9460 9732 9512
rect 4436 9324 4488 9376
rect 5448 9324 5500 9376
rect 6644 9324 6696 9376
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 8576 9324 8628 9376
rect 10600 9324 10652 9376
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 14372 9324 14424 9376
rect 15844 9324 15896 9376
rect 16580 9324 16632 9376
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 24216 9460 24268 9512
rect 24400 9503 24452 9512
rect 24400 9469 24409 9503
rect 24409 9469 24443 9503
rect 24443 9469 24452 9503
rect 24400 9460 24452 9469
rect 25504 9460 25556 9512
rect 26700 9460 26752 9512
rect 28080 9503 28132 9512
rect 28080 9469 28089 9503
rect 28089 9469 28123 9503
rect 28123 9469 28132 9503
rect 28080 9460 28132 9469
rect 30564 9571 30616 9580
rect 30564 9537 30598 9571
rect 30598 9537 30616 9571
rect 30564 9528 30616 9537
rect 33140 9528 33192 9580
rect 34612 9528 34664 9580
rect 34796 9571 34848 9580
rect 34796 9537 34830 9571
rect 34830 9537 34848 9571
rect 34796 9528 34848 9537
rect 35164 9528 35216 9580
rect 25136 9392 25188 9444
rect 19432 9324 19484 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 23848 9367 23900 9376
rect 23848 9333 23857 9367
rect 23857 9333 23891 9367
rect 23891 9333 23900 9367
rect 23848 9324 23900 9333
rect 25044 9324 25096 9376
rect 30288 9460 30340 9512
rect 30472 9503 30524 9512
rect 30472 9469 30481 9503
rect 30481 9469 30515 9503
rect 30515 9469 30524 9503
rect 30472 9460 30524 9469
rect 30196 9435 30248 9444
rect 30196 9401 30205 9435
rect 30205 9401 30239 9435
rect 30239 9401 30248 9435
rect 30196 9392 30248 9401
rect 31944 9460 31996 9512
rect 32128 9460 32180 9512
rect 37924 9596 37976 9648
rect 38660 9596 38712 9648
rect 37464 9571 37516 9580
rect 37464 9537 37473 9571
rect 37473 9537 37507 9571
rect 37507 9537 37516 9571
rect 37464 9528 37516 9537
rect 38016 9571 38068 9580
rect 38016 9537 38025 9571
rect 38025 9537 38059 9571
rect 38059 9537 38068 9571
rect 38016 9528 38068 9537
rect 38568 9460 38620 9512
rect 39304 9571 39356 9580
rect 39304 9537 39313 9571
rect 39313 9537 39347 9571
rect 39347 9537 39356 9571
rect 39304 9528 39356 9537
rect 39580 9571 39632 9580
rect 39580 9537 39589 9571
rect 39589 9537 39623 9571
rect 39623 9537 39632 9571
rect 39580 9528 39632 9537
rect 41328 9664 41380 9716
rect 41512 9664 41564 9716
rect 41604 9707 41656 9716
rect 41604 9673 41613 9707
rect 41613 9673 41647 9707
rect 41647 9673 41656 9707
rect 41604 9664 41656 9673
rect 42524 9664 42576 9716
rect 43996 9664 44048 9716
rect 44088 9707 44140 9716
rect 44088 9673 44097 9707
rect 44097 9673 44131 9707
rect 44131 9673 44140 9707
rect 44088 9664 44140 9673
rect 45008 9528 45060 9580
rect 45468 9664 45520 9716
rect 46020 9664 46072 9716
rect 46388 9664 46440 9716
rect 46480 9664 46532 9716
rect 46664 9664 46716 9716
rect 47768 9664 47820 9716
rect 53472 9664 53524 9716
rect 54668 9664 54720 9716
rect 46204 9596 46256 9648
rect 46848 9596 46900 9648
rect 49332 9596 49384 9648
rect 54944 9596 54996 9648
rect 40500 9503 40552 9512
rect 40500 9469 40509 9503
rect 40509 9469 40543 9503
rect 40543 9469 40552 9503
rect 40500 9460 40552 9469
rect 40684 9503 40736 9512
rect 40684 9469 40693 9503
rect 40693 9469 40727 9503
rect 40727 9469 40736 9503
rect 40684 9460 40736 9469
rect 45652 9571 45704 9580
rect 45652 9537 45661 9571
rect 45661 9537 45695 9571
rect 45695 9537 45704 9571
rect 45652 9528 45704 9537
rect 47768 9528 47820 9580
rect 47860 9528 47912 9580
rect 48320 9571 48372 9580
rect 48320 9537 48329 9571
rect 48329 9537 48363 9571
rect 48363 9537 48372 9571
rect 48320 9528 48372 9537
rect 49700 9528 49752 9580
rect 52000 9528 52052 9580
rect 30840 9324 30892 9376
rect 32036 9324 32088 9376
rect 32404 9324 32456 9376
rect 33784 9367 33836 9376
rect 33784 9333 33793 9367
rect 33793 9333 33827 9367
rect 33827 9333 33836 9367
rect 33784 9324 33836 9333
rect 35900 9367 35952 9376
rect 35900 9333 35909 9367
rect 35909 9333 35943 9367
rect 35943 9333 35952 9367
rect 35900 9324 35952 9333
rect 36728 9367 36780 9376
rect 36728 9333 36737 9367
rect 36737 9333 36771 9367
rect 36771 9333 36780 9367
rect 36728 9324 36780 9333
rect 37648 9367 37700 9376
rect 37648 9333 37657 9367
rect 37657 9333 37691 9367
rect 37691 9333 37700 9367
rect 37648 9324 37700 9333
rect 39304 9324 39356 9376
rect 39488 9324 39540 9376
rect 44824 9435 44876 9444
rect 44824 9401 44833 9435
rect 44833 9401 44867 9435
rect 44867 9401 44876 9435
rect 44824 9392 44876 9401
rect 45560 9392 45612 9444
rect 53748 9503 53800 9512
rect 53748 9469 53757 9503
rect 53757 9469 53791 9503
rect 53791 9469 53800 9503
rect 53748 9460 53800 9469
rect 56048 9707 56100 9716
rect 56048 9673 56057 9707
rect 56057 9673 56091 9707
rect 56091 9673 56100 9707
rect 56048 9664 56100 9673
rect 57336 9664 57388 9716
rect 56600 9596 56652 9648
rect 55404 9528 55456 9580
rect 56968 9528 57020 9580
rect 58164 9528 58216 9580
rect 55588 9392 55640 9444
rect 57336 9503 57388 9512
rect 57336 9469 57345 9503
rect 57345 9469 57379 9503
rect 57379 9469 57388 9503
rect 57336 9460 57388 9469
rect 57428 9503 57480 9512
rect 57428 9469 57437 9503
rect 57437 9469 57471 9503
rect 57471 9469 57480 9503
rect 57428 9460 57480 9469
rect 41328 9367 41380 9376
rect 41328 9333 41337 9367
rect 41337 9333 41371 9367
rect 41371 9333 41380 9367
rect 41328 9324 41380 9333
rect 46388 9324 46440 9376
rect 46572 9367 46624 9376
rect 46572 9333 46581 9367
rect 46581 9333 46615 9367
rect 46615 9333 46624 9367
rect 46572 9324 46624 9333
rect 47584 9367 47636 9376
rect 47584 9333 47593 9367
rect 47593 9333 47627 9367
rect 47627 9333 47636 9367
rect 47584 9324 47636 9333
rect 47952 9324 48004 9376
rect 50344 9324 50396 9376
rect 51356 9324 51408 9376
rect 51632 9367 51684 9376
rect 51632 9333 51641 9367
rect 51641 9333 51675 9367
rect 51675 9333 51684 9367
rect 51632 9324 51684 9333
rect 52920 9324 52972 9376
rect 54760 9324 54812 9376
rect 55312 9324 55364 9376
rect 56876 9367 56928 9376
rect 56876 9333 56885 9367
rect 56885 9333 56919 9367
rect 56919 9333 56928 9367
rect 56876 9324 56928 9333
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 22616 9222 22668 9274
rect 22680 9222 22732 9274
rect 22744 9222 22796 9274
rect 22808 9222 22860 9274
rect 22872 9222 22924 9274
rect 37060 9222 37112 9274
rect 37124 9222 37176 9274
rect 37188 9222 37240 9274
rect 37252 9222 37304 9274
rect 37316 9222 37368 9274
rect 51504 9222 51556 9274
rect 51568 9222 51620 9274
rect 51632 9222 51684 9274
rect 51696 9222 51748 9274
rect 51760 9222 51812 9274
rect 6092 9120 6144 9172
rect 6368 9120 6420 9172
rect 7012 9120 7064 9172
rect 7104 9120 7156 9172
rect 8944 9120 8996 9172
rect 10876 9120 10928 9172
rect 11520 9120 11572 9172
rect 16212 9120 16264 9172
rect 16672 9120 16724 9172
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 18144 9120 18196 9172
rect 20076 9120 20128 9172
rect 23020 9120 23072 9172
rect 23848 9120 23900 9172
rect 25044 9120 25096 9172
rect 26516 9163 26568 9172
rect 26516 9129 26525 9163
rect 26525 9129 26559 9163
rect 26559 9129 26568 9163
rect 26516 9120 26568 9129
rect 28080 9120 28132 9172
rect 31116 9120 31168 9172
rect 31760 9120 31812 9172
rect 33140 9163 33192 9172
rect 33140 9129 33149 9163
rect 33149 9129 33183 9163
rect 33183 9129 33192 9163
rect 33140 9120 33192 9129
rect 33784 9120 33836 9172
rect 34520 9163 34572 9172
rect 34520 9129 34529 9163
rect 34529 9129 34563 9163
rect 34563 9129 34572 9163
rect 34520 9120 34572 9129
rect 8852 9052 8904 9104
rect 10508 9052 10560 9104
rect 4528 8984 4580 9036
rect 11612 9095 11664 9104
rect 11612 9061 11621 9095
rect 11621 9061 11655 9095
rect 11655 9061 11664 9095
rect 11612 9052 11664 9061
rect 3792 8916 3844 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7656 8959 7708 8968
rect 7656 8925 7690 8959
rect 7690 8925 7708 8959
rect 7656 8916 7708 8925
rect 6828 8848 6880 8900
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 11152 8984 11204 9036
rect 16856 8984 16908 9036
rect 19616 8984 19668 9036
rect 21272 8984 21324 9036
rect 4620 8780 4672 8832
rect 6460 8780 6512 8832
rect 8024 8780 8076 8832
rect 9220 8848 9272 8900
rect 9496 8780 9548 8832
rect 10140 8780 10192 8832
rect 10692 8780 10744 8832
rect 11336 8848 11388 8900
rect 11612 8848 11664 8900
rect 16028 8848 16080 8900
rect 23664 8916 23716 8968
rect 24400 8916 24452 8968
rect 24860 8916 24912 8968
rect 11796 8780 11848 8832
rect 12348 8823 12400 8832
rect 12348 8789 12357 8823
rect 12357 8789 12391 8823
rect 12391 8789 12400 8823
rect 12348 8780 12400 8789
rect 16212 8780 16264 8832
rect 17408 8823 17460 8832
rect 17408 8789 17417 8823
rect 17417 8789 17451 8823
rect 17451 8789 17460 8823
rect 17408 8780 17460 8789
rect 18788 8780 18840 8832
rect 19800 8848 19852 8900
rect 20352 8848 20404 8900
rect 30196 9052 30248 9104
rect 28908 8984 28960 9036
rect 26148 8916 26200 8968
rect 33600 8984 33652 9036
rect 36544 9120 36596 9172
rect 37556 9163 37608 9172
rect 37556 9129 37565 9163
rect 37565 9129 37599 9163
rect 37599 9129 37608 9163
rect 37556 9120 37608 9129
rect 37648 9120 37700 9172
rect 37924 9120 37976 9172
rect 38016 9120 38068 9172
rect 39212 9120 39264 9172
rect 41972 9120 42024 9172
rect 42432 9120 42484 9172
rect 43996 9163 44048 9172
rect 43996 9129 44005 9163
rect 44005 9129 44039 9163
rect 44039 9129 44048 9163
rect 43996 9120 44048 9129
rect 45836 9163 45888 9172
rect 45836 9129 45845 9163
rect 45845 9129 45879 9163
rect 45879 9129 45888 9163
rect 45836 9120 45888 9129
rect 46480 9120 46532 9172
rect 49148 9120 49200 9172
rect 49700 9163 49752 9172
rect 49700 9129 49709 9163
rect 49709 9129 49743 9163
rect 49743 9129 49752 9163
rect 49700 9120 49752 9129
rect 50344 9163 50396 9172
rect 50344 9129 50353 9163
rect 50353 9129 50387 9163
rect 50387 9129 50396 9163
rect 50344 9120 50396 9129
rect 52552 9120 52604 9172
rect 52736 9120 52788 9172
rect 53748 9120 53800 9172
rect 55128 9163 55180 9172
rect 55128 9129 55137 9163
rect 55137 9129 55171 9163
rect 55171 9129 55180 9163
rect 55128 9120 55180 9129
rect 55312 9120 55364 9172
rect 56600 9120 56652 9172
rect 56876 9120 56928 9172
rect 57612 9163 57664 9172
rect 57612 9129 57621 9163
rect 57621 9129 57655 9163
rect 57655 9129 57664 9163
rect 57612 9120 57664 9129
rect 30288 8916 30340 8968
rect 29000 8891 29052 8900
rect 29000 8857 29009 8891
rect 29009 8857 29043 8891
rect 29043 8857 29052 8891
rect 29000 8848 29052 8857
rect 19432 8780 19484 8832
rect 19524 8780 19576 8832
rect 22468 8780 22520 8832
rect 23204 8780 23256 8832
rect 24860 8823 24912 8832
rect 24860 8789 24869 8823
rect 24869 8789 24903 8823
rect 24903 8789 24912 8823
rect 24860 8780 24912 8789
rect 25504 8780 25556 8832
rect 26700 8780 26752 8832
rect 28632 8823 28684 8832
rect 28632 8789 28641 8823
rect 28641 8789 28675 8823
rect 28675 8789 28684 8823
rect 28632 8780 28684 8789
rect 29092 8823 29144 8832
rect 29092 8789 29101 8823
rect 29101 8789 29135 8823
rect 29135 8789 29144 8823
rect 29092 8780 29144 8789
rect 30196 8780 30248 8832
rect 34520 8848 34572 8900
rect 35164 8848 35216 8900
rect 35900 9027 35952 9036
rect 35900 8993 35909 9027
rect 35909 8993 35943 9027
rect 35943 8993 35952 9027
rect 35900 8984 35952 8993
rect 40684 9052 40736 9104
rect 42800 9052 42852 9104
rect 46388 9095 46440 9104
rect 46388 9061 46397 9095
rect 46397 9061 46431 9095
rect 46431 9061 46440 9095
rect 46388 9052 46440 9061
rect 38476 8984 38528 9036
rect 38568 8984 38620 9036
rect 40592 8984 40644 9036
rect 44916 8984 44968 9036
rect 37832 8916 37884 8968
rect 39488 8916 39540 8968
rect 43444 8959 43496 8968
rect 43444 8925 43453 8959
rect 43453 8925 43487 8959
rect 43487 8925 43496 8959
rect 43444 8916 43496 8925
rect 45284 8959 45336 8968
rect 45284 8925 45293 8959
rect 45293 8925 45327 8959
rect 45327 8925 45336 8959
rect 45284 8916 45336 8925
rect 36084 8848 36136 8900
rect 38384 8848 38436 8900
rect 41972 8848 42024 8900
rect 42156 8891 42208 8900
rect 42156 8857 42165 8891
rect 42165 8857 42199 8891
rect 42199 8857 42208 8891
rect 42156 8848 42208 8857
rect 47768 8984 47820 9036
rect 53840 9052 53892 9104
rect 54024 9095 54076 9104
rect 54024 9061 54033 9095
rect 54033 9061 54067 9095
rect 54067 9061 54076 9095
rect 54024 9052 54076 9061
rect 54668 9095 54720 9104
rect 54668 9061 54677 9095
rect 54677 9061 54711 9095
rect 54711 9061 54720 9095
rect 54668 9052 54720 9061
rect 56416 9052 56468 9104
rect 56692 8984 56744 9036
rect 47952 8959 48004 8968
rect 47952 8925 47961 8959
rect 47961 8925 47995 8959
rect 47995 8925 48004 8959
rect 47952 8916 48004 8925
rect 51080 8959 51132 8968
rect 51080 8925 51114 8959
rect 51114 8925 51132 8959
rect 51080 8916 51132 8925
rect 58256 8959 58308 8968
rect 58256 8925 58265 8959
rect 58265 8925 58299 8959
rect 58299 8925 58308 8959
rect 58256 8916 58308 8925
rect 52920 8891 52972 8900
rect 30472 8823 30524 8832
rect 30472 8789 30481 8823
rect 30481 8789 30515 8823
rect 30515 8789 30524 8823
rect 30472 8780 30524 8789
rect 31760 8780 31812 8832
rect 32404 8780 32456 8832
rect 35716 8823 35768 8832
rect 35716 8789 35725 8823
rect 35725 8789 35759 8823
rect 35759 8789 35768 8823
rect 35716 8780 35768 8789
rect 42892 8823 42944 8832
rect 42892 8789 42901 8823
rect 42901 8789 42935 8823
rect 42935 8789 42944 8823
rect 42892 8780 42944 8789
rect 52920 8857 52929 8891
rect 52929 8857 52963 8891
rect 52963 8857 52972 8891
rect 52920 8848 52972 8857
rect 56600 8848 56652 8900
rect 45560 8780 45612 8832
rect 57704 8823 57756 8832
rect 57704 8789 57713 8823
rect 57713 8789 57747 8823
rect 57747 8789 57756 8823
rect 57704 8780 57756 8789
rect 15394 8678 15446 8730
rect 15458 8678 15510 8730
rect 15522 8678 15574 8730
rect 15586 8678 15638 8730
rect 15650 8678 15702 8730
rect 29838 8678 29890 8730
rect 29902 8678 29954 8730
rect 29966 8678 30018 8730
rect 30030 8678 30082 8730
rect 30094 8678 30146 8730
rect 44282 8678 44334 8730
rect 44346 8678 44398 8730
rect 44410 8678 44462 8730
rect 44474 8678 44526 8730
rect 44538 8678 44590 8730
rect 58726 8678 58778 8730
rect 58790 8678 58842 8730
rect 58854 8678 58906 8730
rect 58918 8678 58970 8730
rect 58982 8678 59034 8730
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 7564 8619 7616 8628
rect 7564 8585 7573 8619
rect 7573 8585 7607 8619
rect 7607 8585 7616 8619
rect 7564 8576 7616 8585
rect 9220 8576 9272 8628
rect 11152 8576 11204 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 17960 8576 18012 8628
rect 18788 8576 18840 8628
rect 6368 8508 6420 8560
rect 6828 8508 6880 8560
rect 8576 8508 8628 8560
rect 7104 8440 7156 8492
rect 4528 8304 4580 8356
rect 8024 8440 8076 8492
rect 7748 8372 7800 8424
rect 8668 8440 8720 8492
rect 8576 8372 8628 8424
rect 8852 8372 8904 8424
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 16396 8508 16448 8560
rect 17408 8440 17460 8492
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 11520 8372 11572 8424
rect 11612 8415 11664 8424
rect 11612 8381 11621 8415
rect 11621 8381 11655 8415
rect 11655 8381 11664 8415
rect 11612 8372 11664 8381
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 19524 8508 19576 8560
rect 20076 8440 20128 8492
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 4988 8236 5040 8288
rect 5540 8236 5592 8288
rect 5908 8236 5960 8288
rect 10600 8304 10652 8356
rect 12532 8304 12584 8356
rect 17960 8304 18012 8356
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 19340 8372 19392 8424
rect 25228 8619 25280 8628
rect 25228 8585 25237 8619
rect 25237 8585 25271 8619
rect 25271 8585 25280 8619
rect 25228 8576 25280 8585
rect 28448 8619 28500 8628
rect 28448 8585 28457 8619
rect 28457 8585 28491 8619
rect 28491 8585 28500 8619
rect 28448 8576 28500 8585
rect 28632 8576 28684 8628
rect 29092 8576 29144 8628
rect 30380 8576 30432 8628
rect 30748 8619 30800 8628
rect 30748 8585 30757 8619
rect 30757 8585 30791 8619
rect 30791 8585 30800 8619
rect 30748 8576 30800 8585
rect 30840 8619 30892 8628
rect 30840 8585 30849 8619
rect 30849 8585 30883 8619
rect 30883 8585 30892 8619
rect 30840 8576 30892 8585
rect 34796 8576 34848 8628
rect 35716 8576 35768 8628
rect 36084 8576 36136 8628
rect 42892 8576 42944 8628
rect 48320 8576 48372 8628
rect 49976 8576 50028 8628
rect 50344 8576 50396 8628
rect 52736 8576 52788 8628
rect 55772 8576 55824 8628
rect 20352 8508 20404 8560
rect 25136 8508 25188 8560
rect 26700 8440 26752 8492
rect 29368 8483 29420 8492
rect 29368 8449 29377 8483
rect 29377 8449 29411 8483
rect 29411 8449 29420 8483
rect 29368 8440 29420 8449
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 45284 8508 45336 8560
rect 23756 8372 23808 8424
rect 24032 8415 24084 8424
rect 24032 8381 24041 8415
rect 24041 8381 24075 8415
rect 24075 8381 24084 8415
rect 24032 8372 24084 8381
rect 26884 8372 26936 8424
rect 31392 8415 31444 8424
rect 31392 8381 31401 8415
rect 31401 8381 31435 8415
rect 31435 8381 31444 8415
rect 31392 8372 31444 8381
rect 22376 8304 22428 8356
rect 10324 8236 10376 8288
rect 15108 8236 15160 8288
rect 20168 8236 20220 8288
rect 23572 8236 23624 8288
rect 24676 8236 24728 8288
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 28908 8304 28960 8356
rect 31852 8304 31904 8356
rect 35992 8304 36044 8356
rect 32036 8236 32088 8288
rect 34428 8236 34480 8288
rect 35348 8236 35400 8288
rect 39396 8440 39448 8492
rect 42524 8483 42576 8492
rect 42524 8449 42533 8483
rect 42533 8449 42567 8483
rect 42567 8449 42576 8483
rect 42524 8440 42576 8449
rect 42616 8440 42668 8492
rect 36636 8415 36688 8424
rect 36636 8381 36645 8415
rect 36645 8381 36679 8415
rect 36679 8381 36688 8415
rect 36636 8372 36688 8381
rect 41420 8415 41472 8424
rect 41420 8381 41429 8415
rect 41429 8381 41463 8415
rect 41463 8381 41472 8415
rect 41420 8372 41472 8381
rect 41604 8415 41656 8424
rect 41604 8381 41613 8415
rect 41613 8381 41647 8415
rect 41647 8381 41656 8415
rect 41604 8372 41656 8381
rect 44180 8304 44232 8356
rect 47584 8415 47636 8424
rect 47584 8381 47593 8415
rect 47593 8381 47627 8415
rect 47627 8381 47636 8415
rect 47584 8372 47636 8381
rect 51356 8508 51408 8560
rect 57060 8508 57112 8560
rect 52000 8440 52052 8492
rect 52184 8440 52236 8492
rect 54024 8372 54076 8424
rect 52092 8304 52144 8356
rect 52920 8347 52972 8356
rect 52920 8313 52929 8347
rect 52929 8313 52963 8347
rect 52963 8313 52972 8347
rect 52920 8304 52972 8313
rect 56692 8440 56744 8492
rect 57244 8483 57296 8492
rect 57244 8449 57253 8483
rect 57253 8449 57287 8483
rect 57287 8449 57296 8483
rect 57244 8440 57296 8449
rect 54576 8415 54628 8424
rect 54576 8381 54585 8415
rect 54585 8381 54619 8415
rect 54619 8381 54628 8415
rect 54576 8372 54628 8381
rect 55772 8372 55824 8424
rect 37464 8236 37516 8288
rect 38384 8279 38436 8288
rect 38384 8245 38393 8279
rect 38393 8245 38427 8279
rect 38427 8245 38436 8279
rect 38384 8236 38436 8245
rect 40776 8279 40828 8288
rect 40776 8245 40785 8279
rect 40785 8245 40819 8279
rect 40819 8245 40828 8279
rect 40776 8236 40828 8245
rect 41236 8236 41288 8288
rect 43168 8236 43220 8288
rect 43996 8279 44048 8288
rect 43996 8245 44005 8279
rect 44005 8245 44039 8279
rect 44039 8245 44048 8279
rect 43996 8236 44048 8245
rect 48228 8279 48280 8288
rect 48228 8245 48237 8279
rect 48237 8245 48271 8279
rect 48271 8245 48280 8279
rect 48228 8236 48280 8245
rect 51172 8236 51224 8288
rect 53932 8279 53984 8288
rect 53932 8245 53941 8279
rect 53941 8245 53975 8279
rect 53975 8245 53984 8279
rect 53932 8236 53984 8245
rect 54392 8236 54444 8288
rect 54760 8236 54812 8288
rect 55680 8304 55732 8356
rect 56600 8372 56652 8424
rect 57428 8415 57480 8424
rect 57428 8381 57437 8415
rect 57437 8381 57471 8415
rect 57471 8381 57480 8415
rect 57428 8372 57480 8381
rect 58440 8415 58492 8424
rect 58440 8381 58449 8415
rect 58449 8381 58483 8415
rect 58483 8381 58492 8415
rect 58440 8372 58492 8381
rect 56232 8236 56284 8288
rect 56784 8279 56836 8288
rect 56784 8245 56793 8279
rect 56793 8245 56827 8279
rect 56827 8245 56836 8279
rect 56784 8236 56836 8245
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 22616 8134 22668 8186
rect 22680 8134 22732 8186
rect 22744 8134 22796 8186
rect 22808 8134 22860 8186
rect 22872 8134 22924 8186
rect 37060 8134 37112 8186
rect 37124 8134 37176 8186
rect 37188 8134 37240 8186
rect 37252 8134 37304 8186
rect 37316 8134 37368 8186
rect 51504 8134 51556 8186
rect 51568 8134 51620 8186
rect 51632 8134 51684 8186
rect 51696 8134 51748 8186
rect 51760 8134 51812 8186
rect 7748 8032 7800 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 10324 8032 10376 8084
rect 11612 8032 11664 8084
rect 12900 8032 12952 8084
rect 6368 7939 6420 7948
rect 6368 7905 6377 7939
rect 6377 7905 6411 7939
rect 6411 7905 6420 7939
rect 6368 7896 6420 7905
rect 7104 7964 7156 8016
rect 14096 8032 14148 8084
rect 14832 8032 14884 8084
rect 19248 8032 19300 8084
rect 19892 8032 19944 8084
rect 20812 8032 20864 8084
rect 24124 8075 24176 8084
rect 24124 8041 24133 8075
rect 24133 8041 24167 8075
rect 24167 8041 24176 8075
rect 24124 8032 24176 8041
rect 31392 8032 31444 8084
rect 34152 8032 34204 8084
rect 34888 8032 34940 8084
rect 35164 8032 35216 8084
rect 41420 8032 41472 8084
rect 42800 8075 42852 8084
rect 42800 8041 42809 8075
rect 42809 8041 42843 8075
rect 42843 8041 42852 8075
rect 42800 8032 42852 8041
rect 43444 8032 43496 8084
rect 7012 7828 7064 7880
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8300 7828 8352 7880
rect 9680 7828 9732 7880
rect 11060 7828 11112 7880
rect 17316 8007 17368 8016
rect 17316 7973 17325 8007
rect 17325 7973 17359 8007
rect 17359 7973 17368 8007
rect 17316 7964 17368 7973
rect 20352 7964 20404 8016
rect 22468 7964 22520 8016
rect 23480 7964 23532 8016
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 19708 7896 19760 7948
rect 20076 7939 20128 7948
rect 20076 7905 20094 7939
rect 20094 7905 20128 7939
rect 20076 7896 20128 7905
rect 20168 7939 20220 7948
rect 20168 7905 20177 7939
rect 20177 7905 20211 7939
rect 20211 7905 20220 7939
rect 20168 7896 20220 7905
rect 21272 7896 21324 7948
rect 22376 7896 22428 7948
rect 23664 7939 23716 7948
rect 23664 7905 23673 7939
rect 23673 7905 23707 7939
rect 23707 7905 23716 7939
rect 23664 7896 23716 7905
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 17592 7828 17644 7880
rect 8576 7760 8628 7812
rect 10232 7760 10284 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 5080 7692 5132 7744
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 10600 7692 10652 7744
rect 12992 7760 13044 7812
rect 17500 7803 17552 7812
rect 17500 7769 17509 7803
rect 17509 7769 17543 7803
rect 17543 7769 17552 7803
rect 17500 7760 17552 7769
rect 17960 7803 18012 7812
rect 17960 7769 17994 7803
rect 17994 7769 18012 7803
rect 17960 7760 18012 7769
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 14096 7735 14148 7744
rect 14096 7701 14105 7735
rect 14105 7701 14139 7735
rect 14139 7701 14148 7735
rect 14096 7692 14148 7701
rect 15108 7735 15160 7744
rect 15108 7701 15117 7735
rect 15117 7701 15151 7735
rect 15151 7701 15160 7735
rect 15108 7692 15160 7701
rect 16212 7692 16264 7744
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 20720 7828 20772 7880
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 23296 7828 23348 7880
rect 24676 7964 24728 8016
rect 27528 7964 27580 8016
rect 40592 7964 40644 8016
rect 24860 7896 24912 7948
rect 25412 7896 25464 7948
rect 26424 7896 26476 7948
rect 32128 7896 32180 7948
rect 41972 7896 42024 7948
rect 42616 7896 42668 7948
rect 43076 7964 43128 8016
rect 45836 8032 45888 8084
rect 46940 8075 46992 8084
rect 46940 8041 46949 8075
rect 46949 8041 46983 8075
rect 46983 8041 46992 8075
rect 46940 8032 46992 8041
rect 47584 8032 47636 8084
rect 50436 8075 50488 8084
rect 50436 8041 50445 8075
rect 50445 8041 50479 8075
rect 50479 8041 50488 8075
rect 50436 8032 50488 8041
rect 52736 8075 52788 8084
rect 52736 8041 52745 8075
rect 52745 8041 52779 8075
rect 52779 8041 52788 8075
rect 52736 8032 52788 8041
rect 52184 7964 52236 8016
rect 43996 7896 44048 7948
rect 48320 7939 48372 7948
rect 48320 7905 48329 7939
rect 48329 7905 48363 7939
rect 48363 7905 48372 7939
rect 48320 7896 48372 7905
rect 49332 7896 49384 7948
rect 50804 7939 50856 7948
rect 50804 7905 50813 7939
rect 50813 7905 50847 7939
rect 50847 7905 50856 7939
rect 50804 7896 50856 7905
rect 56600 8075 56652 8084
rect 56600 8041 56609 8075
rect 56609 8041 56643 8075
rect 56643 8041 56652 8075
rect 56600 8032 56652 8041
rect 58440 8032 58492 8084
rect 23940 7828 23992 7880
rect 25228 7828 25280 7880
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 31760 7828 31812 7837
rect 33140 7871 33192 7880
rect 33140 7837 33149 7871
rect 33149 7837 33183 7871
rect 33183 7837 33192 7871
rect 33140 7828 33192 7837
rect 36084 7871 36136 7880
rect 36084 7837 36093 7871
rect 36093 7837 36127 7871
rect 36127 7837 36136 7871
rect 36084 7828 36136 7837
rect 36820 7871 36872 7880
rect 36820 7837 36829 7871
rect 36829 7837 36863 7871
rect 36863 7837 36872 7871
rect 36820 7828 36872 7837
rect 37556 7871 37608 7880
rect 37556 7837 37565 7871
rect 37565 7837 37599 7871
rect 37599 7837 37608 7871
rect 37556 7828 37608 7837
rect 38108 7871 38160 7880
rect 38108 7837 38117 7871
rect 38117 7837 38151 7871
rect 38151 7837 38160 7871
rect 38108 7828 38160 7837
rect 39396 7871 39448 7880
rect 39396 7837 39405 7871
rect 39405 7837 39439 7871
rect 39439 7837 39448 7871
rect 39396 7828 39448 7837
rect 41236 7871 41288 7880
rect 41236 7837 41245 7871
rect 41245 7837 41279 7871
rect 41279 7837 41288 7871
rect 41236 7828 41288 7837
rect 41420 7828 41472 7880
rect 24860 7760 24912 7812
rect 35900 7760 35952 7812
rect 19800 7692 19852 7744
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 24400 7692 24452 7744
rect 25872 7692 25924 7744
rect 26700 7692 26752 7744
rect 32588 7735 32640 7744
rect 32588 7701 32597 7735
rect 32597 7701 32631 7735
rect 32631 7701 32640 7735
rect 32588 7692 32640 7701
rect 35532 7735 35584 7744
rect 35532 7701 35541 7735
rect 35541 7701 35575 7735
rect 35575 7701 35584 7735
rect 35532 7692 35584 7701
rect 36268 7735 36320 7744
rect 36268 7701 36277 7735
rect 36277 7701 36311 7735
rect 36311 7701 36320 7735
rect 36268 7692 36320 7701
rect 36728 7692 36780 7744
rect 38752 7735 38804 7744
rect 38752 7701 38761 7735
rect 38761 7701 38795 7735
rect 38795 7701 38804 7735
rect 38752 7692 38804 7701
rect 38844 7735 38896 7744
rect 38844 7701 38853 7735
rect 38853 7701 38887 7735
rect 38887 7701 38896 7735
rect 38844 7692 38896 7701
rect 41696 7735 41748 7744
rect 41696 7701 41705 7735
rect 41705 7701 41739 7735
rect 41739 7701 41748 7735
rect 41696 7692 41748 7701
rect 42892 7828 42944 7880
rect 43260 7828 43312 7880
rect 44640 7828 44692 7880
rect 48964 7871 49016 7880
rect 48964 7837 48973 7871
rect 48973 7837 49007 7871
rect 49007 7837 49016 7871
rect 48964 7828 49016 7837
rect 50620 7828 50672 7880
rect 52276 7871 52328 7880
rect 52276 7837 52285 7871
rect 52285 7837 52319 7871
rect 52319 7837 52328 7871
rect 52276 7828 52328 7837
rect 53840 7828 53892 7880
rect 55956 7871 56008 7880
rect 55956 7837 55965 7871
rect 55965 7837 55999 7871
rect 55999 7837 56008 7871
rect 55956 7828 56008 7837
rect 56416 7828 56468 7880
rect 56784 7828 56836 7880
rect 57428 7828 57480 7880
rect 51264 7760 51316 7812
rect 43352 7735 43404 7744
rect 43352 7701 43361 7735
rect 43361 7701 43395 7735
rect 43395 7701 43404 7735
rect 43352 7692 43404 7701
rect 43904 7735 43956 7744
rect 43904 7701 43913 7735
rect 43913 7701 43947 7735
rect 43947 7701 43956 7735
rect 43904 7692 43956 7701
rect 51632 7735 51684 7744
rect 51632 7701 51641 7735
rect 51641 7701 51675 7735
rect 51675 7701 51684 7735
rect 51632 7692 51684 7701
rect 55496 7692 55548 7744
rect 15394 7590 15446 7642
rect 15458 7590 15510 7642
rect 15522 7590 15574 7642
rect 15586 7590 15638 7642
rect 15650 7590 15702 7642
rect 29838 7590 29890 7642
rect 29902 7590 29954 7642
rect 29966 7590 30018 7642
rect 30030 7590 30082 7642
rect 30094 7590 30146 7642
rect 44282 7590 44334 7642
rect 44346 7590 44398 7642
rect 44410 7590 44462 7642
rect 44474 7590 44526 7642
rect 44538 7590 44590 7642
rect 58726 7590 58778 7642
rect 58790 7590 58842 7642
rect 58854 7590 58906 7642
rect 58918 7590 58970 7642
rect 58982 7590 59034 7642
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 5264 7488 5316 7540
rect 6368 7420 6420 7472
rect 8208 7488 8260 7540
rect 9220 7531 9272 7540
rect 9220 7497 9229 7531
rect 9229 7497 9263 7531
rect 9263 7497 9272 7531
rect 9220 7488 9272 7497
rect 10416 7488 10468 7540
rect 10692 7488 10744 7540
rect 12256 7488 12308 7540
rect 7380 7420 7432 7472
rect 8300 7420 8352 7472
rect 8668 7420 8720 7472
rect 11888 7420 11940 7472
rect 3148 7352 3200 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 7288 7352 7340 7404
rect 9036 7352 9088 7404
rect 9680 7352 9732 7404
rect 12900 7488 12952 7540
rect 14004 7488 14056 7540
rect 14556 7531 14608 7540
rect 14556 7497 14565 7531
rect 14565 7497 14599 7531
rect 14599 7497 14608 7531
rect 14556 7488 14608 7497
rect 14740 7488 14792 7540
rect 17592 7488 17644 7540
rect 19340 7488 19392 7540
rect 20168 7488 20220 7540
rect 15660 7463 15712 7472
rect 15660 7429 15669 7463
rect 15669 7429 15703 7463
rect 15703 7429 15712 7463
rect 15660 7420 15712 7429
rect 13820 7352 13872 7404
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 5172 7327 5224 7336
rect 5172 7293 5190 7327
rect 5190 7293 5224 7327
rect 5172 7284 5224 7293
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 6092 7284 6144 7336
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 8576 7284 8628 7336
rect 9128 7284 9180 7336
rect 10324 7284 10376 7336
rect 3884 7148 3936 7200
rect 5724 7148 5776 7200
rect 10692 7148 10744 7200
rect 11520 7148 11572 7200
rect 13820 7216 13872 7268
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 23020 7488 23072 7540
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 24032 7531 24084 7540
rect 24032 7497 24041 7531
rect 24041 7497 24075 7531
rect 24075 7497 24084 7531
rect 24032 7488 24084 7497
rect 25872 7488 25924 7540
rect 30472 7531 30524 7540
rect 30472 7497 30481 7531
rect 30481 7497 30515 7531
rect 30515 7497 30524 7531
rect 30472 7488 30524 7497
rect 30840 7488 30892 7540
rect 31760 7488 31812 7540
rect 33140 7488 33192 7540
rect 18052 7352 18104 7404
rect 19524 7352 19576 7404
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 18788 7284 18840 7336
rect 19248 7284 19300 7336
rect 23572 7420 23624 7472
rect 24676 7420 24728 7472
rect 20996 7352 21048 7404
rect 21456 7352 21508 7404
rect 22468 7352 22520 7404
rect 24400 7395 24452 7404
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 19800 7284 19852 7336
rect 25596 7395 25648 7404
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 25872 7395 25924 7404
rect 25872 7361 25881 7395
rect 25881 7361 25915 7395
rect 25915 7361 25924 7395
rect 25872 7352 25924 7361
rect 26424 7352 26476 7404
rect 33968 7420 34020 7472
rect 35164 7488 35216 7540
rect 35532 7488 35584 7540
rect 36636 7488 36688 7540
rect 39396 7488 39448 7540
rect 41604 7488 41656 7540
rect 41972 7531 42024 7540
rect 41972 7497 41981 7531
rect 41981 7497 42015 7531
rect 42015 7497 42024 7531
rect 41972 7488 42024 7497
rect 43352 7488 43404 7540
rect 36176 7420 36228 7472
rect 15936 7216 15988 7268
rect 13912 7148 13964 7200
rect 16212 7148 16264 7200
rect 17040 7148 17092 7200
rect 25688 7284 25740 7336
rect 27068 7284 27120 7336
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 28356 7327 28408 7336
rect 28356 7293 28365 7327
rect 28365 7293 28399 7327
rect 28399 7293 28408 7327
rect 28356 7284 28408 7293
rect 29368 7327 29420 7336
rect 29368 7293 29377 7327
rect 29377 7293 29411 7327
rect 29411 7293 29420 7327
rect 29368 7284 29420 7293
rect 30196 7284 30248 7336
rect 26056 7216 26108 7268
rect 18972 7191 19024 7200
rect 18972 7157 18981 7191
rect 18981 7157 19015 7191
rect 19015 7157 19024 7191
rect 18972 7148 19024 7157
rect 20720 7148 20772 7200
rect 27252 7216 27304 7268
rect 30932 7284 30984 7336
rect 33600 7327 33652 7336
rect 33600 7293 33609 7327
rect 33609 7293 33643 7327
rect 33643 7293 33652 7327
rect 33600 7284 33652 7293
rect 27620 7148 27672 7200
rect 29276 7148 29328 7200
rect 29460 7191 29512 7200
rect 29460 7157 29469 7191
rect 29469 7157 29503 7191
rect 29503 7157 29512 7191
rect 29460 7148 29512 7157
rect 35072 7352 35124 7404
rect 37648 7352 37700 7404
rect 40776 7420 40828 7472
rect 44640 7488 44692 7540
rect 47768 7488 47820 7540
rect 48228 7488 48280 7540
rect 48964 7488 49016 7540
rect 50804 7488 50856 7540
rect 47952 7463 48004 7472
rect 47952 7429 47961 7463
rect 47961 7429 47995 7463
rect 47995 7429 48004 7463
rect 47952 7420 48004 7429
rect 48504 7420 48556 7472
rect 51632 7488 51684 7540
rect 52276 7488 52328 7540
rect 53840 7488 53892 7540
rect 55312 7488 55364 7540
rect 56324 7488 56376 7540
rect 43076 7395 43128 7404
rect 43076 7361 43085 7395
rect 43085 7361 43119 7395
rect 43119 7361 43128 7395
rect 43076 7352 43128 7361
rect 43168 7352 43220 7404
rect 43352 7395 43404 7404
rect 43352 7361 43361 7395
rect 43361 7361 43395 7395
rect 43395 7361 43404 7395
rect 43352 7352 43404 7361
rect 48964 7395 49016 7404
rect 48964 7361 48973 7395
rect 48973 7361 49007 7395
rect 49007 7361 49016 7395
rect 48964 7352 49016 7361
rect 34520 7327 34572 7336
rect 34520 7293 34529 7327
rect 34529 7293 34563 7327
rect 34563 7293 34572 7327
rect 34520 7284 34572 7293
rect 36360 7216 36412 7268
rect 34704 7148 34756 7200
rect 35624 7148 35676 7200
rect 39120 7284 39172 7336
rect 44180 7284 44232 7336
rect 44916 7327 44968 7336
rect 44916 7293 44925 7327
rect 44925 7293 44959 7327
rect 44959 7293 44968 7327
rect 44916 7284 44968 7293
rect 45744 7327 45796 7336
rect 45744 7293 45753 7327
rect 45753 7293 45787 7327
rect 45787 7293 45796 7327
rect 45744 7284 45796 7293
rect 46480 7327 46532 7336
rect 46480 7293 46489 7327
rect 46489 7293 46523 7327
rect 46523 7293 46532 7327
rect 46480 7284 46532 7293
rect 46664 7327 46716 7336
rect 46664 7293 46673 7327
rect 46673 7293 46707 7327
rect 46707 7293 46716 7327
rect 46664 7284 46716 7293
rect 47400 7284 47452 7336
rect 50712 7352 50764 7404
rect 51264 7352 51316 7404
rect 52000 7352 52052 7404
rect 53932 7420 53984 7472
rect 57336 7420 57388 7472
rect 56232 7395 56284 7404
rect 56232 7361 56241 7395
rect 56241 7361 56275 7395
rect 56275 7361 56284 7395
rect 56232 7352 56284 7361
rect 56324 7352 56376 7404
rect 56508 7395 56560 7404
rect 56508 7361 56517 7395
rect 56517 7361 56551 7395
rect 56551 7361 56560 7395
rect 56508 7352 56560 7361
rect 57244 7395 57296 7404
rect 57244 7361 57253 7395
rect 57253 7361 57287 7395
rect 57287 7361 57296 7395
rect 57244 7352 57296 7361
rect 58440 7395 58492 7404
rect 58440 7361 58449 7395
rect 58449 7361 58483 7395
rect 58483 7361 58492 7395
rect 58440 7352 58492 7361
rect 43996 7216 44048 7268
rect 45652 7216 45704 7268
rect 38936 7148 38988 7200
rect 45192 7148 45244 7200
rect 45560 7148 45612 7200
rect 47584 7148 47636 7200
rect 49884 7148 49936 7200
rect 50620 7148 50672 7200
rect 50712 7148 50764 7200
rect 53288 7327 53340 7336
rect 53288 7293 53297 7327
rect 53297 7293 53331 7327
rect 53331 7293 53340 7327
rect 53288 7284 53340 7293
rect 52736 7191 52788 7200
rect 52736 7157 52745 7191
rect 52745 7157 52779 7191
rect 52779 7157 52788 7191
rect 52736 7148 52788 7157
rect 54208 7148 54260 7200
rect 54760 7148 54812 7200
rect 57336 7284 57388 7336
rect 56324 7148 56376 7200
rect 56876 7148 56928 7200
rect 57520 7148 57572 7200
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 22616 7046 22668 7098
rect 22680 7046 22732 7098
rect 22744 7046 22796 7098
rect 22808 7046 22860 7098
rect 22872 7046 22924 7098
rect 37060 7046 37112 7098
rect 37124 7046 37176 7098
rect 37188 7046 37240 7098
rect 37252 7046 37304 7098
rect 37316 7046 37368 7098
rect 51504 7046 51556 7098
rect 51568 7046 51620 7098
rect 51632 7046 51684 7098
rect 51696 7046 51748 7098
rect 51760 7046 51812 7098
rect 3608 6944 3660 6996
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 4620 6876 4672 6928
rect 11520 6808 11572 6860
rect 17316 6944 17368 6996
rect 18052 6944 18104 6996
rect 19800 6944 19852 6996
rect 20996 6987 21048 6996
rect 20996 6953 21005 6987
rect 21005 6953 21039 6987
rect 21039 6953 21048 6987
rect 20996 6944 21048 6953
rect 15384 6919 15436 6928
rect 15384 6885 15393 6919
rect 15393 6885 15427 6919
rect 15427 6885 15436 6919
rect 15384 6876 15436 6885
rect 15844 6876 15896 6928
rect 24860 6944 24912 6996
rect 25688 6944 25740 6996
rect 24952 6876 25004 6928
rect 26700 6944 26752 6996
rect 15660 6808 15712 6860
rect 18972 6851 19024 6860
rect 18972 6817 18981 6851
rect 18981 6817 19015 6851
rect 19015 6817 19024 6851
rect 18972 6808 19024 6817
rect 19432 6808 19484 6860
rect 20260 6851 20312 6860
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 22100 6808 22152 6860
rect 22468 6851 22520 6860
rect 22468 6817 22477 6851
rect 22477 6817 22511 6851
rect 22511 6817 22520 6851
rect 22468 6808 22520 6817
rect 24124 6808 24176 6860
rect 25504 6851 25556 6860
rect 25504 6817 25513 6851
rect 25513 6817 25547 6851
rect 25547 6817 25556 6851
rect 25504 6808 25556 6817
rect 29368 6987 29420 6996
rect 29368 6953 29377 6987
rect 29377 6953 29411 6987
rect 29411 6953 29420 6987
rect 29368 6944 29420 6953
rect 33600 6944 33652 6996
rect 36820 6944 36872 6996
rect 38108 6944 38160 6996
rect 38200 6944 38252 6996
rect 33692 6876 33744 6928
rect 27896 6808 27948 6860
rect 2136 6740 2188 6792
rect 2964 6672 3016 6724
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 5080 6672 5132 6724
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 7656 6740 7708 6792
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 12348 6740 12400 6792
rect 9036 6672 9088 6724
rect 12808 6715 12860 6724
rect 12808 6681 12842 6715
rect 12842 6681 12860 6715
rect 12808 6672 12860 6681
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 13176 6604 13228 6656
rect 14188 6647 14240 6656
rect 14188 6613 14197 6647
rect 14197 6613 14231 6647
rect 14231 6613 14240 6647
rect 14188 6604 14240 6613
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 14924 6740 14976 6792
rect 15200 6604 15252 6656
rect 16212 6740 16264 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 20720 6740 20772 6792
rect 19616 6672 19668 6724
rect 17040 6604 17092 6656
rect 19524 6604 19576 6656
rect 19892 6604 19944 6656
rect 22468 6672 22520 6724
rect 22928 6672 22980 6724
rect 23940 6604 23992 6656
rect 25136 6672 25188 6724
rect 26056 6740 26108 6792
rect 33968 6851 34020 6860
rect 33968 6817 33977 6851
rect 33977 6817 34011 6851
rect 34011 6817 34020 6851
rect 33968 6808 34020 6817
rect 34152 6851 34204 6860
rect 34152 6817 34161 6851
rect 34161 6817 34195 6851
rect 34195 6817 34204 6851
rect 34152 6808 34204 6817
rect 36452 6808 36504 6860
rect 36820 6851 36872 6860
rect 36820 6817 36829 6851
rect 36829 6817 36863 6851
rect 36863 6817 36872 6851
rect 36820 6808 36872 6817
rect 46664 6944 46716 6996
rect 53288 6944 53340 6996
rect 55956 6944 56008 6996
rect 41788 6876 41840 6928
rect 51172 6876 51224 6928
rect 25320 6715 25372 6724
rect 25320 6681 25329 6715
rect 25329 6681 25363 6715
rect 25363 6681 25372 6715
rect 25320 6672 25372 6681
rect 26976 6672 27028 6724
rect 28264 6715 28316 6724
rect 28264 6681 28298 6715
rect 28298 6681 28316 6715
rect 28264 6672 28316 6681
rect 28356 6672 28408 6724
rect 29460 6672 29512 6724
rect 24400 6604 24452 6656
rect 26332 6604 26384 6656
rect 32128 6740 32180 6792
rect 34520 6740 34572 6792
rect 37648 6740 37700 6792
rect 32588 6672 32640 6724
rect 36268 6672 36320 6724
rect 31024 6647 31076 6656
rect 31024 6613 31033 6647
rect 31033 6613 31067 6647
rect 31067 6613 31076 6647
rect 31024 6604 31076 6613
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 33876 6647 33928 6656
rect 33876 6613 33885 6647
rect 33885 6613 33919 6647
rect 33919 6613 33928 6647
rect 33876 6604 33928 6613
rect 37556 6672 37608 6724
rect 38016 6672 38068 6724
rect 38568 6672 38620 6724
rect 38752 6808 38804 6860
rect 38936 6740 38988 6792
rect 39856 6740 39908 6792
rect 40960 6740 41012 6792
rect 41696 6740 41748 6792
rect 46940 6808 46992 6860
rect 47124 6808 47176 6860
rect 47492 6851 47544 6860
rect 47492 6817 47501 6851
rect 47501 6817 47535 6851
rect 47535 6817 47544 6851
rect 47492 6808 47544 6817
rect 47609 6851 47661 6860
rect 47609 6817 47618 6851
rect 47618 6817 47652 6851
rect 47652 6817 47661 6851
rect 47609 6808 47661 6817
rect 48412 6808 48464 6860
rect 49056 6851 49108 6860
rect 49056 6817 49065 6851
rect 49065 6817 49099 6851
rect 49099 6817 49108 6851
rect 49056 6808 49108 6817
rect 50620 6808 50672 6860
rect 51356 6808 51408 6860
rect 52184 6808 52236 6860
rect 54024 6808 54076 6860
rect 55588 6808 55640 6860
rect 45008 6783 45060 6792
rect 45008 6749 45017 6783
rect 45017 6749 45051 6783
rect 45051 6749 45060 6783
rect 45008 6740 45060 6749
rect 45560 6740 45612 6792
rect 46756 6783 46808 6792
rect 46756 6749 46765 6783
rect 46765 6749 46799 6783
rect 46799 6749 46808 6783
rect 46756 6740 46808 6749
rect 47768 6783 47820 6792
rect 47768 6749 47777 6783
rect 47777 6749 47811 6783
rect 47811 6749 47820 6783
rect 47768 6740 47820 6749
rect 36544 6647 36596 6656
rect 36544 6613 36553 6647
rect 36553 6613 36587 6647
rect 36587 6613 36596 6647
rect 36544 6604 36596 6613
rect 36728 6604 36780 6656
rect 36820 6604 36872 6656
rect 38108 6604 38160 6656
rect 38660 6604 38712 6656
rect 39396 6604 39448 6656
rect 43904 6672 43956 6724
rect 43996 6672 44048 6724
rect 43260 6604 43312 6656
rect 45744 6604 45796 6656
rect 47124 6604 47176 6656
rect 49976 6783 50028 6792
rect 49976 6749 49985 6783
rect 49985 6749 50019 6783
rect 50019 6749 50028 6783
rect 49976 6740 50028 6749
rect 50804 6783 50856 6792
rect 50804 6749 50813 6783
rect 50813 6749 50847 6783
rect 50847 6749 50856 6783
rect 50804 6740 50856 6749
rect 51724 6740 51776 6792
rect 53840 6740 53892 6792
rect 54208 6672 54260 6724
rect 48320 6604 48372 6656
rect 49424 6604 49476 6656
rect 49884 6604 49936 6656
rect 51172 6604 51224 6656
rect 52460 6647 52512 6656
rect 52460 6613 52469 6647
rect 52469 6613 52503 6647
rect 52503 6613 52512 6647
rect 52460 6604 52512 6613
rect 54392 6647 54444 6656
rect 54392 6613 54401 6647
rect 54401 6613 54435 6647
rect 54435 6613 54444 6647
rect 54392 6604 54444 6613
rect 54576 6604 54628 6656
rect 56140 6740 56192 6792
rect 56416 6783 56468 6792
rect 56416 6749 56425 6783
rect 56425 6749 56459 6783
rect 56459 6749 56468 6783
rect 56416 6740 56468 6749
rect 57428 6740 57480 6792
rect 56508 6672 56560 6724
rect 55220 6604 55272 6656
rect 57060 6604 57112 6656
rect 57796 6647 57848 6656
rect 57796 6613 57805 6647
rect 57805 6613 57839 6647
rect 57839 6613 57848 6647
rect 57796 6604 57848 6613
rect 15394 6502 15446 6554
rect 15458 6502 15510 6554
rect 15522 6502 15574 6554
rect 15586 6502 15638 6554
rect 15650 6502 15702 6554
rect 29838 6502 29890 6554
rect 29902 6502 29954 6554
rect 29966 6502 30018 6554
rect 30030 6502 30082 6554
rect 30094 6502 30146 6554
rect 44282 6502 44334 6554
rect 44346 6502 44398 6554
rect 44410 6502 44462 6554
rect 44474 6502 44526 6554
rect 44538 6502 44590 6554
rect 58726 6502 58778 6554
rect 58790 6502 58842 6554
rect 58854 6502 58906 6554
rect 58918 6502 58970 6554
rect 58982 6502 59034 6554
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 4160 6400 4212 6452
rect 5172 6400 5224 6452
rect 7104 6400 7156 6452
rect 7288 6443 7340 6452
rect 7288 6409 7297 6443
rect 7297 6409 7331 6443
rect 7331 6409 7340 6443
rect 7288 6400 7340 6409
rect 7656 6443 7708 6452
rect 7656 6409 7665 6443
rect 7665 6409 7699 6443
rect 7699 6409 7708 6443
rect 7656 6400 7708 6409
rect 7748 6400 7800 6452
rect 10140 6400 10192 6452
rect 11428 6400 11480 6452
rect 12808 6400 12860 6452
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 4344 6332 4396 6384
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 2320 6239 2372 6248
rect 2320 6205 2329 6239
rect 2329 6205 2363 6239
rect 2363 6205 2372 6239
rect 2320 6196 2372 6205
rect 4068 6196 4120 6248
rect 6552 6196 6604 6248
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 14004 6400 14056 6452
rect 14188 6400 14240 6452
rect 16856 6400 16908 6452
rect 17040 6443 17092 6452
rect 17040 6409 17049 6443
rect 17049 6409 17083 6443
rect 17083 6409 17092 6443
rect 17040 6400 17092 6409
rect 18144 6400 18196 6452
rect 19248 6400 19300 6452
rect 20260 6400 20312 6452
rect 22928 6443 22980 6452
rect 22928 6409 22937 6443
rect 22937 6409 22971 6443
rect 22971 6409 22980 6443
rect 22928 6400 22980 6409
rect 25596 6400 25648 6452
rect 14096 6332 14148 6384
rect 15752 6332 15804 6384
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 11888 6264 11940 6316
rect 12532 6264 12584 6316
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 20720 6264 20772 6316
rect 23480 6307 23532 6316
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 1860 6060 1912 6112
rect 6368 6128 6420 6180
rect 15016 6128 15068 6180
rect 3332 6060 3384 6112
rect 4620 6060 4672 6112
rect 5908 6060 5960 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9496 6060 9548 6112
rect 11796 6060 11848 6112
rect 12348 6060 12400 6112
rect 12532 6060 12584 6112
rect 12808 6060 12860 6112
rect 13360 6060 13412 6112
rect 16488 6128 16540 6180
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 18144 6196 18196 6248
rect 19248 6196 19300 6248
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 18788 6060 18840 6112
rect 19340 6060 19392 6112
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 19800 6060 19852 6112
rect 21916 6196 21968 6248
rect 23940 6196 23992 6248
rect 26148 6400 26200 6452
rect 26424 6400 26476 6452
rect 26884 6400 26936 6452
rect 26976 6443 27028 6452
rect 26976 6409 26985 6443
rect 26985 6409 27019 6443
rect 27019 6409 27028 6443
rect 26976 6400 27028 6409
rect 27896 6443 27948 6452
rect 27896 6409 27905 6443
rect 27905 6409 27939 6443
rect 27939 6409 27948 6443
rect 27896 6400 27948 6409
rect 28264 6400 28316 6452
rect 30196 6400 30248 6452
rect 26332 6307 26384 6316
rect 26332 6273 26341 6307
rect 26341 6273 26375 6307
rect 26375 6273 26384 6307
rect 26332 6264 26384 6273
rect 27068 6264 27120 6316
rect 27620 6307 27672 6316
rect 27620 6273 27629 6307
rect 27629 6273 27663 6307
rect 27663 6273 27672 6307
rect 27620 6264 27672 6273
rect 29276 6307 29328 6316
rect 29276 6273 29285 6307
rect 29285 6273 29319 6307
rect 29319 6273 29328 6307
rect 29276 6264 29328 6273
rect 29644 6264 29696 6316
rect 30472 6332 30524 6384
rect 31024 6332 31076 6384
rect 26148 6128 26200 6180
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 22376 6060 22428 6112
rect 23664 6103 23716 6112
rect 23664 6069 23673 6103
rect 23673 6069 23707 6103
rect 23707 6069 23716 6103
rect 23664 6060 23716 6069
rect 30380 6196 30432 6248
rect 33692 6400 33744 6452
rect 35072 6400 35124 6452
rect 35164 6400 35216 6452
rect 36084 6400 36136 6452
rect 36820 6443 36872 6452
rect 36820 6409 36829 6443
rect 36829 6409 36863 6443
rect 36863 6409 36872 6443
rect 36820 6400 36872 6409
rect 36544 6332 36596 6384
rect 32128 6307 32180 6316
rect 32128 6273 32137 6307
rect 32137 6273 32171 6307
rect 32171 6273 32180 6307
rect 32128 6264 32180 6273
rect 32956 6264 33008 6316
rect 34704 6307 34756 6316
rect 34704 6273 34713 6307
rect 34713 6273 34747 6307
rect 34747 6273 34756 6307
rect 34704 6264 34756 6273
rect 35992 6264 36044 6316
rect 36728 6264 36780 6316
rect 38752 6400 38804 6452
rect 39304 6400 39356 6452
rect 41788 6400 41840 6452
rect 42892 6400 42944 6452
rect 44916 6400 44968 6452
rect 45468 6400 45520 6452
rect 46480 6400 46532 6452
rect 45008 6264 45060 6316
rect 45652 6264 45704 6316
rect 47676 6400 47728 6452
rect 49424 6400 49476 6452
rect 49976 6400 50028 6452
rect 50804 6400 50856 6452
rect 47952 6375 48004 6384
rect 47952 6341 47961 6375
rect 47961 6341 47995 6375
rect 47995 6341 48004 6375
rect 47952 6332 48004 6341
rect 46572 6264 46624 6316
rect 47584 6264 47636 6316
rect 49332 6307 49384 6316
rect 49332 6273 49341 6307
rect 49341 6273 49375 6307
rect 49375 6273 49384 6307
rect 49332 6264 49384 6273
rect 51172 6400 51224 6452
rect 52000 6400 52052 6452
rect 52460 6400 52512 6452
rect 54208 6443 54260 6452
rect 54208 6409 54217 6443
rect 54217 6409 54251 6443
rect 54251 6409 54260 6443
rect 54208 6400 54260 6409
rect 54392 6400 54444 6452
rect 55588 6400 55640 6452
rect 56416 6400 56468 6452
rect 57060 6443 57112 6452
rect 57060 6409 57069 6443
rect 57069 6409 57103 6443
rect 57103 6409 57112 6443
rect 57060 6400 57112 6409
rect 57428 6443 57480 6452
rect 57428 6409 57437 6443
rect 57437 6409 57471 6443
rect 57471 6409 57480 6443
rect 57428 6400 57480 6409
rect 57796 6400 57848 6452
rect 52736 6332 52788 6384
rect 33784 6196 33836 6248
rect 34428 6239 34480 6248
rect 34428 6205 34437 6239
rect 34437 6205 34471 6239
rect 34471 6205 34480 6239
rect 34428 6196 34480 6205
rect 34612 6239 34664 6248
rect 34612 6205 34630 6239
rect 34630 6205 34664 6239
rect 34612 6196 34664 6205
rect 34888 6128 34940 6180
rect 35808 6196 35860 6248
rect 37832 6239 37884 6248
rect 37832 6205 37841 6239
rect 37841 6205 37875 6239
rect 37875 6205 37884 6239
rect 37832 6196 37884 6205
rect 30380 6060 30432 6112
rect 33692 6060 33744 6112
rect 38016 6128 38068 6180
rect 38752 6196 38804 6248
rect 39028 6196 39080 6248
rect 39856 6196 39908 6248
rect 38200 6128 38252 6180
rect 42616 6128 42668 6180
rect 37464 6103 37516 6112
rect 37464 6069 37473 6103
rect 37473 6069 37507 6103
rect 37507 6069 37516 6103
rect 37464 6060 37516 6069
rect 38384 6060 38436 6112
rect 38844 6060 38896 6112
rect 39580 6103 39632 6112
rect 39580 6069 39589 6103
rect 39589 6069 39623 6103
rect 39623 6069 39632 6103
rect 39580 6060 39632 6069
rect 44088 6060 44140 6112
rect 47216 6196 47268 6248
rect 48136 6239 48188 6248
rect 48136 6205 48145 6239
rect 48145 6205 48179 6239
rect 48179 6205 48188 6239
rect 48136 6196 48188 6205
rect 51172 6307 51224 6316
rect 51172 6273 51181 6307
rect 51181 6273 51215 6307
rect 51215 6273 51224 6307
rect 51172 6264 51224 6273
rect 52552 6264 52604 6316
rect 46664 6060 46716 6112
rect 50252 6060 50304 6112
rect 50712 6103 50764 6112
rect 50712 6069 50721 6103
rect 50721 6069 50755 6103
rect 50755 6069 50764 6103
rect 50712 6060 50764 6069
rect 51264 6060 51316 6112
rect 52000 6196 52052 6248
rect 52092 6196 52144 6248
rect 52368 6060 52420 6112
rect 52736 6103 52788 6112
rect 52736 6069 52745 6103
rect 52745 6069 52779 6103
rect 52779 6069 52788 6103
rect 52736 6060 52788 6069
rect 55312 6307 55364 6316
rect 55312 6273 55321 6307
rect 55321 6273 55355 6307
rect 55355 6273 55364 6307
rect 55312 6264 55364 6273
rect 55496 6307 55548 6316
rect 55496 6273 55505 6307
rect 55505 6273 55539 6307
rect 55539 6273 55548 6307
rect 55496 6264 55548 6273
rect 56876 6239 56928 6248
rect 56876 6205 56885 6239
rect 56885 6205 56919 6239
rect 56919 6205 56928 6239
rect 56876 6196 56928 6205
rect 57336 6196 57388 6248
rect 55404 6060 55456 6112
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 22616 5958 22668 6010
rect 22680 5958 22732 6010
rect 22744 5958 22796 6010
rect 22808 5958 22860 6010
rect 22872 5958 22924 6010
rect 37060 5958 37112 6010
rect 37124 5958 37176 6010
rect 37188 5958 37240 6010
rect 37252 5958 37304 6010
rect 37316 5958 37368 6010
rect 51504 5958 51556 6010
rect 51568 5958 51620 6010
rect 51632 5958 51684 6010
rect 51696 5958 51748 6010
rect 51760 5958 51812 6010
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 2136 5856 2188 5908
rect 2320 5856 2372 5908
rect 3332 5831 3384 5840
rect 3332 5797 3341 5831
rect 3341 5797 3375 5831
rect 3375 5797 3384 5831
rect 3332 5788 3384 5797
rect 6092 5831 6144 5840
rect 6092 5797 6101 5831
rect 6101 5797 6135 5831
rect 6135 5797 6144 5831
rect 6092 5788 6144 5797
rect 6276 5788 6328 5840
rect 9220 5856 9272 5908
rect 9588 5856 9640 5908
rect 10784 5856 10836 5908
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13452 5856 13504 5908
rect 14924 5856 14976 5908
rect 15200 5899 15252 5908
rect 15200 5865 15209 5899
rect 15209 5865 15243 5899
rect 15243 5865 15252 5899
rect 15200 5856 15252 5865
rect 17040 5856 17092 5908
rect 19248 5899 19300 5908
rect 19248 5865 19257 5899
rect 19257 5865 19291 5899
rect 19291 5865 19300 5899
rect 19248 5856 19300 5865
rect 22008 5899 22060 5908
rect 22008 5865 22017 5899
rect 22017 5865 22051 5899
rect 22051 5865 22060 5899
rect 22008 5856 22060 5865
rect 24124 5856 24176 5908
rect 26148 5856 26200 5908
rect 27896 5856 27948 5908
rect 30380 5899 30432 5908
rect 30380 5865 30389 5899
rect 30389 5865 30423 5899
rect 30423 5865 30432 5899
rect 30380 5856 30432 5865
rect 30932 5856 30984 5908
rect 31116 5899 31168 5908
rect 31116 5865 31125 5899
rect 31125 5865 31159 5899
rect 31159 5865 31168 5899
rect 31116 5856 31168 5865
rect 32956 5899 33008 5908
rect 32956 5865 32965 5899
rect 32965 5865 32999 5899
rect 32999 5865 33008 5899
rect 32956 5856 33008 5865
rect 33508 5856 33560 5908
rect 33692 5856 33744 5908
rect 33876 5856 33928 5908
rect 34612 5856 34664 5908
rect 35808 5856 35860 5908
rect 37832 5856 37884 5908
rect 38384 5856 38436 5908
rect 38614 5856 38666 5908
rect 39120 5856 39172 5908
rect 45836 5856 45888 5908
rect 46572 5856 46624 5908
rect 47952 5856 48004 5908
rect 48136 5856 48188 5908
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 9312 5720 9364 5772
rect 4068 5652 4120 5704
rect 3056 5584 3108 5636
rect 4804 5584 4856 5636
rect 6184 5652 6236 5704
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 7748 5652 7800 5704
rect 10048 5720 10100 5772
rect 10876 5652 10928 5704
rect 10968 5652 11020 5704
rect 3700 5516 3752 5568
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4344 5516 4396 5568
rect 6092 5516 6144 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 7196 5516 7248 5568
rect 13912 5720 13964 5772
rect 14832 5652 14884 5704
rect 13360 5584 13412 5636
rect 18236 5720 18288 5772
rect 20628 5763 20680 5772
rect 20628 5729 20637 5763
rect 20637 5729 20671 5763
rect 20671 5729 20680 5763
rect 20628 5720 20680 5729
rect 22376 5720 22428 5772
rect 15292 5652 15344 5704
rect 16212 5652 16264 5704
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 26332 5763 26384 5772
rect 26332 5729 26341 5763
rect 26341 5729 26375 5763
rect 26375 5729 26384 5763
rect 26332 5720 26384 5729
rect 34428 5720 34480 5772
rect 37740 5720 37792 5772
rect 39856 5788 39908 5840
rect 45376 5788 45428 5840
rect 39028 5720 39080 5772
rect 24952 5695 25004 5704
rect 24952 5661 24961 5695
rect 24961 5661 24995 5695
rect 24995 5661 25004 5695
rect 24952 5652 25004 5661
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 40868 5720 40920 5772
rect 44088 5720 44140 5772
rect 39396 5695 39448 5704
rect 39396 5661 39405 5695
rect 39405 5661 39439 5695
rect 39439 5661 39448 5695
rect 39396 5652 39448 5661
rect 16488 5584 16540 5636
rect 19800 5584 19852 5636
rect 24216 5584 24268 5636
rect 24308 5584 24360 5636
rect 9496 5516 9548 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 10508 5516 10560 5568
rect 11796 5516 11848 5568
rect 13268 5516 13320 5568
rect 14004 5516 14056 5568
rect 16028 5516 16080 5568
rect 16672 5516 16724 5568
rect 17132 5516 17184 5568
rect 17684 5559 17736 5568
rect 17684 5525 17693 5559
rect 17693 5525 17727 5559
rect 17727 5525 17736 5559
rect 17684 5516 17736 5525
rect 19064 5559 19116 5568
rect 19064 5525 19073 5559
rect 19073 5525 19107 5559
rect 19107 5525 19116 5559
rect 19064 5516 19116 5525
rect 22192 5516 22244 5568
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 24860 5516 24912 5568
rect 29736 5584 29788 5636
rect 26884 5559 26936 5568
rect 26884 5525 26893 5559
rect 26893 5525 26927 5559
rect 26927 5525 26936 5559
rect 26884 5516 26936 5525
rect 30656 5516 30708 5568
rect 36820 5584 36872 5636
rect 38844 5584 38896 5636
rect 41420 5695 41472 5704
rect 41420 5661 41429 5695
rect 41429 5661 41463 5695
rect 41463 5661 41472 5695
rect 41420 5652 41472 5661
rect 41788 5695 41840 5704
rect 41788 5661 41797 5695
rect 41797 5661 41831 5695
rect 41831 5661 41840 5695
rect 41788 5652 41840 5661
rect 42340 5652 42392 5704
rect 42984 5695 43036 5704
rect 42984 5661 42993 5695
rect 42993 5661 43027 5695
rect 43027 5661 43036 5695
rect 42984 5652 43036 5661
rect 43076 5652 43128 5704
rect 44180 5652 44232 5704
rect 47584 5763 47636 5772
rect 47584 5729 47593 5763
rect 47593 5729 47627 5763
rect 47627 5729 47636 5763
rect 47584 5720 47636 5729
rect 48596 5856 48648 5908
rect 49056 5856 49108 5908
rect 50712 5856 50764 5908
rect 51264 5856 51316 5908
rect 52000 5899 52052 5908
rect 52000 5865 52009 5899
rect 52009 5865 52043 5899
rect 52043 5865 52052 5899
rect 52000 5856 52052 5865
rect 52920 5856 52972 5908
rect 34152 5516 34204 5568
rect 36912 5516 36964 5568
rect 37648 5516 37700 5568
rect 38108 5516 38160 5568
rect 39396 5516 39448 5568
rect 42708 5584 42760 5636
rect 40868 5559 40920 5568
rect 40868 5525 40877 5559
rect 40877 5525 40911 5559
rect 40911 5525 40920 5559
rect 40868 5516 40920 5525
rect 41696 5516 41748 5568
rect 43628 5516 43680 5568
rect 47032 5584 47084 5636
rect 47216 5516 47268 5568
rect 49884 5652 49936 5704
rect 50528 5652 50580 5704
rect 52828 5695 52880 5704
rect 52828 5661 52837 5695
rect 52837 5661 52871 5695
rect 52871 5661 52880 5695
rect 52828 5652 52880 5661
rect 53748 5652 53800 5704
rect 54852 5695 54904 5704
rect 54852 5661 54861 5695
rect 54861 5661 54895 5695
rect 54895 5661 54904 5695
rect 54852 5652 54904 5661
rect 55864 5695 55916 5704
rect 55864 5661 55873 5695
rect 55873 5661 55907 5695
rect 55907 5661 55916 5695
rect 55864 5652 55916 5661
rect 55956 5652 56008 5704
rect 57336 5695 57388 5704
rect 57336 5661 57345 5695
rect 57345 5661 57379 5695
rect 57379 5661 57388 5695
rect 57336 5652 57388 5661
rect 57796 5652 57848 5704
rect 52368 5584 52420 5636
rect 54484 5584 54536 5636
rect 48596 5516 48648 5568
rect 48688 5516 48740 5568
rect 49792 5516 49844 5568
rect 52000 5516 52052 5568
rect 53564 5559 53616 5568
rect 53564 5525 53573 5559
rect 53573 5525 53607 5559
rect 53607 5525 53616 5559
rect 53564 5516 53616 5525
rect 54208 5516 54260 5568
rect 54668 5516 54720 5568
rect 56048 5559 56100 5568
rect 56048 5525 56057 5559
rect 56057 5525 56091 5559
rect 56091 5525 56100 5559
rect 56048 5516 56100 5525
rect 56784 5559 56836 5568
rect 56784 5525 56793 5559
rect 56793 5525 56827 5559
rect 56827 5525 56836 5559
rect 56784 5516 56836 5525
rect 58164 5516 58216 5568
rect 15394 5414 15446 5466
rect 15458 5414 15510 5466
rect 15522 5414 15574 5466
rect 15586 5414 15638 5466
rect 15650 5414 15702 5466
rect 29838 5414 29890 5466
rect 29902 5414 29954 5466
rect 29966 5414 30018 5466
rect 30030 5414 30082 5466
rect 30094 5414 30146 5466
rect 44282 5414 44334 5466
rect 44346 5414 44398 5466
rect 44410 5414 44462 5466
rect 44474 5414 44526 5466
rect 44538 5414 44590 5466
rect 58726 5414 58778 5466
rect 58790 5414 58842 5466
rect 58854 5414 58906 5466
rect 58918 5414 58970 5466
rect 58982 5414 59034 5466
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3608 5312 3660 5364
rect 4436 5312 4488 5364
rect 5724 5355 5776 5364
rect 5724 5321 5733 5355
rect 5733 5321 5767 5355
rect 5767 5321 5776 5355
rect 5724 5312 5776 5321
rect 3884 5244 3936 5296
rect 4620 5244 4672 5296
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 6736 5312 6788 5364
rect 10968 5312 11020 5364
rect 11152 5312 11204 5364
rect 16120 5312 16172 5364
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 19708 5312 19760 5364
rect 21272 5312 21324 5364
rect 23848 5312 23900 5364
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 24308 5355 24360 5364
rect 24308 5321 24317 5355
rect 24317 5321 24351 5355
rect 24351 5321 24360 5355
rect 24308 5312 24360 5321
rect 24400 5355 24452 5364
rect 24400 5321 24409 5355
rect 24409 5321 24443 5355
rect 24443 5321 24452 5355
rect 24400 5312 24452 5321
rect 25872 5312 25924 5364
rect 8668 5244 8720 5296
rect 13820 5287 13872 5296
rect 13820 5253 13829 5287
rect 13829 5253 13863 5287
rect 13863 5253 13872 5287
rect 13820 5244 13872 5253
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 7012 5176 7064 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 5724 5040 5776 5092
rect 10508 5219 10560 5228
rect 10508 5185 10542 5219
rect 10542 5185 10560 5219
rect 10508 5176 10560 5185
rect 13268 5176 13320 5228
rect 16028 5176 16080 5228
rect 17684 5244 17736 5296
rect 19616 5287 19668 5296
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 9772 5108 9824 5160
rect 9312 5040 9364 5092
rect 11060 5108 11112 5160
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 14832 5108 14884 5160
rect 10232 5040 10284 5092
rect 11888 5040 11940 5092
rect 16212 5108 16264 5160
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 17960 5108 18012 5160
rect 19616 5253 19625 5287
rect 19625 5253 19659 5287
rect 19659 5253 19668 5287
rect 19616 5244 19668 5253
rect 23664 5244 23716 5296
rect 19064 5176 19116 5228
rect 19340 5176 19392 5228
rect 20168 5176 20220 5228
rect 4344 4972 4396 5024
rect 4712 4972 4764 5024
rect 6736 4972 6788 5024
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 9680 4972 9732 5024
rect 10876 4972 10928 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 12348 5015 12400 5024
rect 12348 4981 12357 5015
rect 12357 4981 12391 5015
rect 12391 4981 12400 5015
rect 12348 4972 12400 4981
rect 13452 5015 13504 5024
rect 13452 4981 13461 5015
rect 13461 4981 13495 5015
rect 13495 4981 13504 5015
rect 14096 5015 14148 5024
rect 13452 4972 13504 4981
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14556 4972 14608 5024
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 18696 5040 18748 5092
rect 19800 5108 19852 5160
rect 20720 5108 20772 5160
rect 21088 5151 21140 5160
rect 21088 5117 21097 5151
rect 21097 5117 21131 5151
rect 21131 5117 21140 5151
rect 21088 5108 21140 5117
rect 22100 5108 22152 5160
rect 26884 5312 26936 5364
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 27896 5312 27948 5364
rect 28448 5312 28500 5364
rect 35808 5312 35860 5364
rect 36912 5355 36964 5364
rect 36912 5321 36921 5355
rect 36921 5321 36955 5355
rect 36955 5321 36964 5355
rect 36912 5312 36964 5321
rect 22376 5040 22428 5092
rect 24952 5108 25004 5160
rect 27344 5219 27396 5228
rect 27344 5185 27353 5219
rect 27353 5185 27387 5219
rect 27387 5185 27396 5219
rect 27344 5176 27396 5185
rect 27528 5176 27580 5228
rect 37740 5244 37792 5296
rect 30564 5176 30616 5228
rect 30932 5176 30984 5228
rect 27436 5108 27488 5160
rect 30380 5151 30432 5160
rect 30380 5117 30389 5151
rect 30389 5117 30423 5151
rect 30423 5117 30432 5151
rect 30380 5108 30432 5117
rect 31300 5151 31352 5160
rect 31300 5117 31309 5151
rect 31309 5117 31343 5151
rect 31343 5117 31352 5151
rect 31300 5108 31352 5117
rect 35992 5108 36044 5160
rect 38292 5151 38344 5160
rect 38292 5117 38301 5151
rect 38301 5117 38335 5151
rect 38335 5117 38344 5151
rect 38292 5108 38344 5117
rect 33784 5083 33836 5092
rect 20904 5015 20956 5024
rect 20904 4981 20913 5015
rect 20913 4981 20947 5015
rect 20947 4981 20956 5015
rect 20904 4972 20956 4981
rect 21640 5015 21692 5024
rect 21640 4981 21649 5015
rect 21649 4981 21683 5015
rect 21683 4981 21692 5015
rect 21640 4972 21692 4981
rect 23756 4972 23808 5024
rect 27620 4972 27672 5024
rect 29460 4972 29512 5024
rect 31024 5015 31076 5024
rect 31024 4981 31033 5015
rect 31033 4981 31067 5015
rect 31067 4981 31076 5015
rect 31024 4972 31076 4981
rect 31576 4972 31628 5024
rect 33784 5049 33793 5083
rect 33793 5049 33827 5083
rect 33827 5049 33836 5083
rect 33784 5040 33836 5049
rect 35716 5083 35768 5092
rect 35716 5049 35725 5083
rect 35725 5049 35759 5083
rect 35759 5049 35768 5083
rect 39488 5108 39540 5160
rect 39672 5108 39724 5160
rect 41328 5312 41380 5364
rect 41512 5355 41564 5364
rect 41512 5321 41521 5355
rect 41521 5321 41555 5355
rect 41555 5321 41564 5355
rect 41512 5312 41564 5321
rect 41880 5244 41932 5296
rect 44180 5312 44232 5364
rect 46756 5355 46808 5364
rect 46756 5321 46765 5355
rect 46765 5321 46799 5355
rect 46799 5321 46808 5355
rect 46756 5312 46808 5321
rect 51172 5312 51224 5364
rect 54668 5355 54720 5364
rect 54668 5321 54677 5355
rect 54677 5321 54711 5355
rect 54711 5321 54720 5355
rect 54668 5312 54720 5321
rect 43260 5244 43312 5296
rect 43812 5176 43864 5228
rect 42432 5151 42484 5160
rect 42432 5117 42441 5151
rect 42441 5117 42475 5151
rect 42475 5117 42484 5151
rect 42432 5108 42484 5117
rect 42892 5108 42944 5160
rect 35716 5040 35768 5049
rect 32404 4972 32456 5024
rect 34888 4972 34940 5024
rect 35808 5015 35860 5024
rect 35808 4981 35817 5015
rect 35817 4981 35851 5015
rect 35851 4981 35860 5015
rect 35808 4972 35860 4981
rect 36636 4972 36688 5024
rect 37740 5015 37792 5024
rect 37740 4981 37749 5015
rect 37749 4981 37783 5015
rect 37783 4981 37792 5015
rect 37740 4972 37792 4981
rect 38568 5015 38620 5024
rect 38568 4981 38577 5015
rect 38577 4981 38611 5015
rect 38611 4981 38620 5015
rect 38568 4972 38620 4981
rect 38844 4972 38896 5024
rect 39304 5015 39356 5024
rect 39304 4981 39313 5015
rect 39313 4981 39347 5015
rect 39347 4981 39356 5015
rect 39304 4972 39356 4981
rect 40040 4972 40092 5024
rect 42616 5040 42668 5092
rect 49608 5244 49660 5296
rect 45284 5219 45336 5228
rect 45284 5185 45293 5219
rect 45293 5185 45327 5219
rect 45327 5185 45336 5219
rect 45284 5176 45336 5185
rect 48872 5176 48924 5228
rect 51264 5244 51316 5296
rect 55864 5312 55916 5364
rect 55956 5312 56008 5364
rect 56140 5312 56192 5364
rect 56048 5244 56100 5296
rect 56692 5312 56744 5364
rect 57888 5312 57940 5364
rect 51908 5176 51960 5228
rect 53288 5219 53340 5228
rect 53288 5185 53297 5219
rect 53297 5185 53331 5219
rect 53331 5185 53340 5219
rect 53288 5176 53340 5185
rect 54024 5176 54076 5228
rect 55220 5176 55272 5228
rect 56508 5219 56560 5228
rect 56508 5185 56517 5219
rect 56517 5185 56551 5219
rect 56551 5185 56560 5219
rect 56508 5176 56560 5185
rect 41420 4972 41472 5024
rect 42708 4972 42760 5024
rect 42800 4972 42852 5024
rect 43168 5015 43220 5024
rect 43168 4981 43177 5015
rect 43177 4981 43211 5015
rect 43211 4981 43220 5015
rect 43168 4972 43220 4981
rect 44732 5108 44784 5160
rect 51080 5108 51132 5160
rect 51356 5108 51408 5160
rect 52368 5151 52420 5160
rect 52368 5117 52377 5151
rect 52377 5117 52411 5151
rect 52411 5117 52420 5151
rect 52368 5108 52420 5117
rect 53196 5108 53248 5160
rect 54484 5151 54536 5160
rect 54484 5117 54493 5151
rect 54493 5117 54527 5151
rect 54527 5117 54536 5151
rect 54484 5108 54536 5117
rect 56692 5108 56744 5160
rect 57888 5108 57940 5160
rect 55128 5040 55180 5092
rect 46020 4972 46072 5024
rect 46572 5015 46624 5024
rect 46572 4981 46581 5015
rect 46581 4981 46615 5015
rect 46615 4981 46624 5015
rect 46572 4972 46624 4981
rect 50712 4972 50764 5024
rect 52920 5015 52972 5024
rect 52920 4981 52929 5015
rect 52929 4981 52963 5015
rect 52963 4981 52972 5015
rect 52920 4972 52972 4981
rect 55312 4972 55364 5024
rect 57704 4972 57756 5024
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 22616 4870 22668 4922
rect 22680 4870 22732 4922
rect 22744 4870 22796 4922
rect 22808 4870 22860 4922
rect 22872 4870 22924 4922
rect 37060 4870 37112 4922
rect 37124 4870 37176 4922
rect 37188 4870 37240 4922
rect 37252 4870 37304 4922
rect 37316 4870 37368 4922
rect 51504 4870 51556 4922
rect 51568 4870 51620 4922
rect 51632 4870 51684 4922
rect 51696 4870 51748 4922
rect 51760 4870 51812 4922
rect 1676 4632 1728 4684
rect 2136 4768 2188 4820
rect 3792 4768 3844 4820
rect 3884 4700 3936 4752
rect 4436 4743 4488 4752
rect 4436 4709 4445 4743
rect 4445 4709 4479 4743
rect 4479 4709 4488 4743
rect 4436 4700 4488 4709
rect 4804 4675 4856 4684
rect 4804 4641 4838 4675
rect 4838 4641 4856 4675
rect 4804 4632 4856 4641
rect 7564 4768 7616 4820
rect 10048 4700 10100 4752
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 2320 4496 2372 4548
rect 2688 4496 2740 4548
rect 8852 4632 8904 4684
rect 10232 4632 10284 4684
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 5816 4564 5868 4616
rect 6000 4564 6052 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7196 4564 7248 4616
rect 7932 4564 7984 4616
rect 5908 4496 5960 4548
rect 6092 4539 6144 4548
rect 6092 4505 6101 4539
rect 6101 4505 6135 4539
rect 6135 4505 6144 4539
rect 6092 4496 6144 4505
rect 9312 4496 9364 4548
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 11520 4768 11572 4820
rect 14096 4768 14148 4820
rect 15016 4768 15068 4820
rect 16212 4768 16264 4820
rect 17592 4811 17644 4820
rect 17592 4777 17601 4811
rect 17601 4777 17635 4811
rect 17635 4777 17644 4811
rect 17592 4768 17644 4777
rect 19708 4768 19760 4820
rect 20628 4768 20680 4820
rect 23848 4768 23900 4820
rect 24216 4811 24268 4820
rect 24216 4777 24225 4811
rect 24225 4777 24259 4811
rect 24259 4777 24268 4811
rect 24216 4768 24268 4777
rect 10968 4700 11020 4752
rect 16304 4700 16356 4752
rect 12440 4632 12492 4684
rect 16028 4632 16080 4684
rect 21548 4632 21600 4684
rect 13268 4564 13320 4616
rect 13912 4607 13964 4616
rect 13912 4573 13921 4607
rect 13921 4573 13955 4607
rect 13955 4573 13964 4607
rect 13912 4564 13964 4573
rect 14004 4564 14056 4616
rect 17040 4564 17092 4616
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 20444 4607 20496 4616
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 21180 4607 21232 4616
rect 21180 4573 21189 4607
rect 21189 4573 21223 4607
rect 21223 4573 21232 4607
rect 21180 4564 21232 4573
rect 21456 4607 21508 4616
rect 21456 4573 21465 4607
rect 21465 4573 21499 4607
rect 21499 4573 21508 4607
rect 21456 4564 21508 4573
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 22192 4564 22244 4616
rect 24400 4675 24452 4684
rect 24400 4641 24409 4675
rect 24409 4641 24443 4675
rect 24443 4641 24452 4675
rect 24400 4632 24452 4641
rect 24860 4700 24912 4752
rect 25136 4632 25188 4684
rect 27344 4768 27396 4820
rect 28448 4811 28500 4820
rect 28448 4777 28457 4811
rect 28457 4777 28491 4811
rect 28491 4777 28500 4811
rect 28448 4768 28500 4777
rect 27528 4632 27580 4684
rect 30472 4768 30524 4820
rect 31300 4768 31352 4820
rect 30196 4743 30248 4752
rect 30196 4709 30205 4743
rect 30205 4709 30239 4743
rect 30239 4709 30248 4743
rect 30196 4700 30248 4709
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 27712 4564 27764 4616
rect 28080 4607 28132 4616
rect 28080 4573 28089 4607
rect 28089 4573 28123 4607
rect 28123 4573 28132 4607
rect 28080 4564 28132 4573
rect 29368 4607 29420 4616
rect 29368 4573 29377 4607
rect 29377 4573 29411 4607
rect 29411 4573 29420 4607
rect 29368 4564 29420 4573
rect 16580 4496 16632 4548
rect 18696 4496 18748 4548
rect 23756 4496 23808 4548
rect 3608 4428 3660 4480
rect 8576 4428 8628 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 11244 4428 11296 4480
rect 12532 4428 12584 4480
rect 13084 4428 13136 4480
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 19248 4428 19300 4480
rect 19892 4471 19944 4480
rect 19892 4437 19901 4471
rect 19901 4437 19935 4471
rect 19935 4437 19944 4471
rect 19892 4428 19944 4437
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 22192 4428 22244 4480
rect 26792 4471 26844 4480
rect 26792 4437 26801 4471
rect 26801 4437 26835 4471
rect 26835 4437 26844 4471
rect 26792 4428 26844 4437
rect 27528 4471 27580 4480
rect 27528 4437 27537 4471
rect 27537 4437 27571 4471
rect 27571 4437 27580 4471
rect 27528 4428 27580 4437
rect 29000 4428 29052 4480
rect 29644 4564 29696 4616
rect 31576 4632 31628 4684
rect 33324 4768 33376 4820
rect 34428 4811 34480 4820
rect 34428 4777 34437 4811
rect 34437 4777 34471 4811
rect 34471 4777 34480 4811
rect 34428 4768 34480 4777
rect 35716 4768 35768 4820
rect 38292 4768 38344 4820
rect 38752 4811 38804 4820
rect 32404 4700 32456 4752
rect 33048 4743 33100 4752
rect 33048 4709 33057 4743
rect 33057 4709 33091 4743
rect 33091 4709 33100 4743
rect 33048 4700 33100 4709
rect 38752 4777 38761 4811
rect 38761 4777 38795 4811
rect 38795 4777 38804 4811
rect 38752 4768 38804 4777
rect 38844 4768 38896 4820
rect 36912 4632 36964 4684
rect 30472 4607 30524 4616
rect 30472 4573 30481 4607
rect 30481 4573 30515 4607
rect 30515 4573 30524 4607
rect 30472 4564 30524 4573
rect 31944 4607 31996 4616
rect 31944 4573 31953 4607
rect 31953 4573 31987 4607
rect 31987 4573 31996 4607
rect 31944 4564 31996 4573
rect 33876 4607 33928 4616
rect 33876 4573 33885 4607
rect 33885 4573 33919 4607
rect 33919 4573 33928 4607
rect 33876 4564 33928 4573
rect 35532 4607 35584 4616
rect 35532 4573 35541 4607
rect 35541 4573 35575 4607
rect 35575 4573 35584 4607
rect 35532 4564 35584 4573
rect 36268 4607 36320 4616
rect 36268 4573 36277 4607
rect 36277 4573 36311 4607
rect 36311 4573 36320 4607
rect 36268 4564 36320 4573
rect 40132 4700 40184 4752
rect 42432 4768 42484 4820
rect 43076 4700 43128 4752
rect 40040 4675 40092 4684
rect 40040 4641 40049 4675
rect 40049 4641 40083 4675
rect 40083 4641 40092 4675
rect 40040 4632 40092 4641
rect 43168 4632 43220 4684
rect 43720 4632 43772 4684
rect 45836 4700 45888 4752
rect 49608 4768 49660 4820
rect 45376 4632 45428 4684
rect 46020 4632 46072 4684
rect 48872 4700 48924 4752
rect 51264 4768 51316 4820
rect 52368 4768 52420 4820
rect 53288 4811 53340 4820
rect 53288 4777 53297 4811
rect 53297 4777 53331 4811
rect 53331 4777 53340 4811
rect 53288 4768 53340 4777
rect 36176 4496 36228 4548
rect 38016 4496 38068 4548
rect 38660 4564 38712 4616
rect 40960 4564 41012 4616
rect 42432 4607 42484 4616
rect 42432 4573 42441 4607
rect 42441 4573 42475 4607
rect 42475 4573 42484 4607
rect 42432 4564 42484 4573
rect 42800 4607 42852 4616
rect 42800 4573 42809 4607
rect 42809 4573 42843 4607
rect 42843 4573 42852 4607
rect 42800 4564 42852 4573
rect 43536 4607 43588 4616
rect 43536 4573 43545 4607
rect 43545 4573 43579 4607
rect 43579 4573 43588 4607
rect 43536 4564 43588 4573
rect 45468 4564 45520 4616
rect 46388 4607 46440 4616
rect 46388 4573 46397 4607
rect 46397 4573 46431 4607
rect 46431 4573 46440 4607
rect 46388 4564 46440 4573
rect 46756 4564 46808 4616
rect 40868 4496 40920 4548
rect 41696 4496 41748 4548
rect 30196 4428 30248 4480
rect 31484 4471 31536 4480
rect 31484 4437 31493 4471
rect 31493 4437 31527 4471
rect 31527 4437 31536 4471
rect 31484 4428 31536 4437
rect 34980 4471 35032 4480
rect 34980 4437 34989 4471
rect 34989 4437 35023 4471
rect 35023 4437 35032 4471
rect 34980 4428 35032 4437
rect 35716 4471 35768 4480
rect 35716 4437 35725 4471
rect 35725 4437 35759 4471
rect 35759 4437 35768 4471
rect 35716 4428 35768 4437
rect 36636 4471 36688 4480
rect 36636 4437 36645 4471
rect 36645 4437 36679 4471
rect 36679 4437 36688 4471
rect 36636 4428 36688 4437
rect 38108 4428 38160 4480
rect 41880 4471 41932 4480
rect 41880 4437 41889 4471
rect 41889 4437 41923 4471
rect 41923 4437 41932 4471
rect 41880 4428 41932 4437
rect 49056 4564 49108 4616
rect 50712 4564 50764 4616
rect 52276 4700 52328 4752
rect 52920 4700 52972 4752
rect 55036 4632 55088 4684
rect 55404 4700 55456 4752
rect 55220 4632 55272 4684
rect 55496 4632 55548 4684
rect 56324 4632 56376 4684
rect 51540 4564 51592 4616
rect 52276 4564 52328 4616
rect 53656 4564 53708 4616
rect 55128 4564 55180 4616
rect 58256 4607 58308 4616
rect 58256 4573 58265 4607
rect 58265 4573 58299 4607
rect 58299 4573 58308 4607
rect 58256 4564 58308 4573
rect 54944 4496 54996 4548
rect 56140 4496 56192 4548
rect 57152 4539 57204 4548
rect 57152 4505 57161 4539
rect 57161 4505 57195 4539
rect 57195 4505 57204 4539
rect 57152 4496 57204 4505
rect 43536 4428 43588 4480
rect 45008 4471 45060 4480
rect 45008 4437 45017 4471
rect 45017 4437 45051 4471
rect 45051 4437 45060 4471
rect 45008 4428 45060 4437
rect 45192 4428 45244 4480
rect 47952 4428 48004 4480
rect 49148 4471 49200 4480
rect 49148 4437 49157 4471
rect 49157 4437 49191 4471
rect 49191 4437 49200 4471
rect 49148 4428 49200 4437
rect 50436 4428 50488 4480
rect 52368 4471 52420 4480
rect 52368 4437 52377 4471
rect 52377 4437 52411 4471
rect 52411 4437 52420 4471
rect 52368 4428 52420 4437
rect 53472 4428 53524 4480
rect 53932 4428 53984 4480
rect 58072 4428 58124 4480
rect 15394 4326 15446 4378
rect 15458 4326 15510 4378
rect 15522 4326 15574 4378
rect 15586 4326 15638 4378
rect 15650 4326 15702 4378
rect 29838 4326 29890 4378
rect 29902 4326 29954 4378
rect 29966 4326 30018 4378
rect 30030 4326 30082 4378
rect 30094 4326 30146 4378
rect 44282 4326 44334 4378
rect 44346 4326 44398 4378
rect 44410 4326 44462 4378
rect 44474 4326 44526 4378
rect 44538 4326 44590 4378
rect 58726 4326 58778 4378
rect 58790 4326 58842 4378
rect 58854 4326 58906 4378
rect 58918 4326 58970 4378
rect 58982 4326 59034 4378
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 4252 4224 4304 4276
rect 4344 4224 4396 4276
rect 2780 4156 2832 4208
rect 6644 4156 6696 4208
rect 6920 4156 6972 4208
rect 4712 4088 4764 4140
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6460 4088 6512 4140
rect 3240 3952 3292 4004
rect 4068 4020 4120 4072
rect 4988 4020 5040 4072
rect 5448 4063 5500 4072
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 6092 4020 6144 4072
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 8852 4267 8904 4276
rect 8852 4233 8861 4267
rect 8861 4233 8895 4267
rect 8895 4233 8904 4267
rect 8852 4224 8904 4233
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 10416 4224 10468 4276
rect 12532 4224 12584 4276
rect 13452 4224 13504 4276
rect 15752 4224 15804 4276
rect 16120 4224 16172 4276
rect 18420 4224 18472 4276
rect 20168 4267 20220 4276
rect 20168 4233 20177 4267
rect 20177 4233 20211 4267
rect 20211 4233 20220 4267
rect 20168 4224 20220 4233
rect 20444 4224 20496 4276
rect 20628 4224 20680 4276
rect 20904 4224 20956 4276
rect 21548 4267 21600 4276
rect 21548 4233 21557 4267
rect 21557 4233 21591 4267
rect 21591 4233 21600 4267
rect 21548 4224 21600 4233
rect 7840 4088 7892 4140
rect 9220 4088 9272 4140
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 3884 3952 3936 4004
rect 4528 3952 4580 4004
rect 6644 3952 6696 4004
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 15936 4088 15988 4140
rect 1860 3884 1912 3936
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 10600 3952 10652 4004
rect 10968 3952 11020 4004
rect 12164 4020 12216 4072
rect 14924 4063 14976 4072
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 14924 4020 14976 4029
rect 16212 4088 16264 4140
rect 16948 4088 17000 4140
rect 17132 4131 17184 4140
rect 17132 4097 17166 4131
rect 17166 4097 17184 4131
rect 17132 4088 17184 4097
rect 10692 3884 10744 3936
rect 10876 3884 10928 3936
rect 11888 3884 11940 3936
rect 12072 3884 12124 3936
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 17868 4020 17920 4072
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 19524 4131 19576 4140
rect 19524 4097 19533 4131
rect 19533 4097 19567 4131
rect 19567 4097 19576 4131
rect 19524 4088 19576 4097
rect 24308 4224 24360 4276
rect 27528 4224 27580 4276
rect 27620 4224 27672 4276
rect 27712 4267 27764 4276
rect 27712 4233 27721 4267
rect 27721 4233 27755 4267
rect 27755 4233 27764 4267
rect 27712 4224 27764 4233
rect 28448 4224 28500 4276
rect 29368 4224 29420 4276
rect 30288 4224 30340 4276
rect 30472 4224 30524 4276
rect 31024 4267 31076 4276
rect 31024 4233 31033 4267
rect 31033 4233 31067 4267
rect 31067 4233 31076 4267
rect 31024 4224 31076 4233
rect 35532 4224 35584 4276
rect 35624 4224 35676 4276
rect 35808 4224 35860 4276
rect 36268 4224 36320 4276
rect 16396 3884 16448 3936
rect 17500 3884 17552 3936
rect 19064 4020 19116 4072
rect 23480 4020 23532 4072
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 26608 4063 26660 4072
rect 26608 4029 26617 4063
rect 26617 4029 26651 4063
rect 26651 4029 26660 4063
rect 26608 4020 26660 4029
rect 26700 4020 26752 4072
rect 27436 4020 27488 4072
rect 29460 4156 29512 4208
rect 19340 3884 19392 3936
rect 20812 3884 20864 3936
rect 22100 3927 22152 3936
rect 22100 3893 22109 3927
rect 22109 3893 22143 3927
rect 22143 3893 22152 3927
rect 22100 3884 22152 3893
rect 22468 3884 22520 3936
rect 23020 3884 23072 3936
rect 24860 3884 24912 3936
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 27160 3884 27212 3936
rect 30196 4131 30248 4140
rect 30196 4097 30205 4131
rect 30205 4097 30239 4131
rect 30239 4097 30248 4131
rect 30196 4088 30248 4097
rect 30196 3952 30248 4004
rect 30564 3995 30616 4004
rect 30564 3961 30573 3995
rect 30573 3961 30607 3995
rect 30607 3961 30616 3995
rect 30564 3952 30616 3961
rect 31668 4131 31720 4140
rect 31668 4097 31677 4131
rect 31677 4097 31711 4131
rect 31711 4097 31720 4131
rect 31668 4088 31720 4097
rect 38200 4224 38252 4276
rect 38660 4267 38712 4276
rect 38660 4233 38669 4267
rect 38669 4233 38703 4267
rect 38703 4233 38712 4267
rect 38660 4224 38712 4233
rect 39304 4224 39356 4276
rect 39488 4267 39540 4276
rect 39488 4233 39497 4267
rect 39497 4233 39531 4267
rect 39531 4233 39540 4267
rect 39488 4224 39540 4233
rect 39580 4224 39632 4276
rect 41696 4224 41748 4276
rect 42432 4224 42484 4276
rect 43168 4224 43220 4276
rect 37740 4156 37792 4208
rect 40960 4156 41012 4208
rect 44732 4267 44784 4276
rect 44732 4233 44741 4267
rect 44741 4233 44775 4267
rect 44775 4233 44784 4267
rect 44732 4224 44784 4233
rect 45008 4224 45060 4276
rect 46388 4224 46440 4276
rect 48780 4224 48832 4276
rect 49056 4267 49108 4276
rect 49056 4233 49065 4267
rect 49065 4233 49099 4267
rect 49099 4233 49108 4267
rect 49056 4224 49108 4233
rect 49700 4224 49752 4276
rect 50988 4224 51040 4276
rect 52276 4267 52328 4276
rect 52276 4233 52285 4267
rect 52285 4233 52319 4267
rect 52319 4233 52328 4267
rect 52276 4224 52328 4233
rect 52736 4224 52788 4276
rect 55036 4224 55088 4276
rect 55128 4224 55180 4276
rect 36912 4088 36964 4140
rect 31116 4063 31168 4072
rect 31116 4029 31125 4063
rect 31125 4029 31159 4063
rect 31159 4029 31168 4063
rect 31116 4020 31168 4029
rect 31576 4020 31628 4072
rect 33140 4020 33192 4072
rect 34152 4063 34204 4072
rect 34152 4029 34161 4063
rect 34161 4029 34195 4063
rect 34195 4029 34204 4063
rect 34152 4020 34204 4029
rect 34888 4063 34940 4072
rect 34888 4029 34897 4063
rect 34897 4029 34931 4063
rect 34931 4029 34940 4063
rect 34888 4020 34940 4029
rect 36360 4063 36412 4072
rect 36360 4029 36369 4063
rect 36369 4029 36403 4063
rect 36403 4029 36412 4063
rect 36360 4020 36412 4029
rect 36636 4020 36688 4072
rect 39764 4088 39816 4140
rect 40132 4131 40184 4140
rect 40132 4097 40141 4131
rect 40141 4097 40175 4131
rect 40175 4097 40184 4131
rect 40132 4088 40184 4097
rect 41512 4131 41564 4140
rect 41512 4097 41521 4131
rect 41521 4097 41555 4131
rect 41555 4097 41564 4131
rect 41512 4088 41564 4097
rect 42800 4088 42852 4140
rect 43628 4131 43680 4140
rect 43628 4097 43662 4131
rect 43662 4097 43680 4131
rect 30656 3884 30708 3936
rect 31208 3884 31260 3936
rect 32864 3927 32916 3936
rect 32864 3893 32873 3927
rect 32873 3893 32907 3927
rect 32907 3893 32916 3927
rect 32864 3884 32916 3893
rect 33232 3884 33284 3936
rect 34336 3927 34388 3936
rect 34336 3893 34345 3927
rect 34345 3893 34379 3927
rect 34379 3893 34388 3927
rect 34336 3884 34388 3893
rect 35900 3884 35952 3936
rect 39028 4020 39080 4072
rect 41420 4020 41472 4072
rect 37648 3884 37700 3936
rect 38016 3884 38068 3936
rect 43260 4020 43312 4072
rect 43168 3952 43220 4004
rect 39580 3927 39632 3936
rect 39580 3893 39589 3927
rect 39589 3893 39623 3927
rect 39623 3893 39632 3927
rect 39580 3884 39632 3893
rect 42064 3884 42116 3936
rect 43628 4088 43680 4097
rect 44916 4063 44968 4072
rect 44916 4029 44925 4063
rect 44925 4029 44959 4063
rect 44959 4029 44968 4063
rect 44916 4020 44968 4029
rect 48688 4088 48740 4140
rect 49792 4088 49844 4140
rect 51172 4088 51224 4140
rect 52000 4088 52052 4140
rect 53472 4156 53524 4208
rect 56140 4267 56192 4276
rect 56140 4233 56149 4267
rect 56149 4233 56183 4267
rect 56183 4233 56192 4267
rect 56140 4224 56192 4233
rect 46664 4020 46716 4072
rect 48136 4063 48188 4072
rect 48136 4029 48145 4063
rect 48145 4029 48179 4063
rect 48179 4029 48188 4063
rect 48136 4020 48188 4029
rect 46572 3952 46624 4004
rect 47308 3995 47360 4004
rect 47308 3961 47317 3995
rect 47317 3961 47351 3995
rect 47351 3961 47360 3995
rect 50252 4063 50304 4072
rect 50252 4029 50261 4063
rect 50261 4029 50295 4063
rect 50295 4029 50304 4063
rect 50252 4020 50304 4029
rect 47308 3952 47360 3961
rect 44272 3884 44324 3936
rect 44824 3884 44876 3936
rect 47584 3927 47636 3936
rect 47584 3893 47593 3927
rect 47593 3893 47627 3927
rect 47627 3893 47636 3927
rect 47584 3884 47636 3893
rect 47768 3884 47820 3936
rect 49240 3884 49292 3936
rect 51540 4020 51592 4072
rect 51356 3952 51408 4004
rect 52736 4020 52788 4072
rect 54208 4088 54260 4140
rect 53288 4020 53340 4072
rect 54024 4020 54076 4072
rect 54668 4088 54720 4140
rect 55312 4131 55364 4140
rect 55312 4097 55346 4131
rect 55346 4097 55364 4131
rect 55312 4088 55364 4097
rect 57980 4088 58032 4140
rect 53104 3884 53156 3936
rect 53380 3884 53432 3936
rect 56048 4020 56100 4072
rect 58348 4020 58400 4072
rect 54760 3952 54812 4004
rect 56140 3952 56192 4004
rect 58440 3952 58492 4004
rect 55588 3884 55640 3936
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 22616 3782 22668 3834
rect 22680 3782 22732 3834
rect 22744 3782 22796 3834
rect 22808 3782 22860 3834
rect 22872 3782 22924 3834
rect 37060 3782 37112 3834
rect 37124 3782 37176 3834
rect 37188 3782 37240 3834
rect 37252 3782 37304 3834
rect 37316 3782 37368 3834
rect 51504 3782 51556 3834
rect 51568 3782 51620 3834
rect 51632 3782 51684 3834
rect 51696 3782 51748 3834
rect 51760 3782 51812 3834
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 4804 3680 4856 3732
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 5448 3680 5500 3732
rect 3608 3587 3660 3596
rect 3608 3553 3617 3587
rect 3617 3553 3651 3587
rect 3651 3553 3660 3587
rect 3608 3544 3660 3553
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 4620 3544 4672 3596
rect 5816 3612 5868 3664
rect 1676 3476 1728 3528
rect 1860 3519 1912 3528
rect 1860 3485 1894 3519
rect 1894 3485 1912 3519
rect 1860 3476 1912 3485
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5724 3476 5776 3528
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 10784 3680 10836 3732
rect 10968 3680 11020 3732
rect 7380 3544 7432 3596
rect 11336 3680 11388 3732
rect 11888 3612 11940 3664
rect 12348 3612 12400 3664
rect 12440 3655 12492 3664
rect 12440 3621 12449 3655
rect 12449 3621 12483 3655
rect 12483 3621 12492 3655
rect 12440 3612 12492 3621
rect 13912 3680 13964 3732
rect 14740 3680 14792 3732
rect 14924 3680 14976 3732
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 5264 3408 5316 3460
rect 5908 3408 5960 3460
rect 6276 3408 6328 3460
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 5724 3340 5776 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 9680 3476 9732 3528
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 12532 3519 12584 3528
rect 12532 3485 12541 3519
rect 12541 3485 12575 3519
rect 12575 3485 12584 3519
rect 12532 3476 12584 3485
rect 13084 3476 13136 3528
rect 14280 3476 14332 3528
rect 14372 3476 14424 3528
rect 10968 3408 11020 3460
rect 11152 3340 11204 3392
rect 12256 3340 12308 3392
rect 14004 3340 14056 3392
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 15752 3476 15804 3528
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 16948 3680 17000 3732
rect 17500 3655 17552 3664
rect 16672 3544 16724 3596
rect 17500 3621 17509 3655
rect 17509 3621 17543 3655
rect 17543 3621 17552 3655
rect 17500 3612 17552 3621
rect 17868 3612 17920 3664
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 16672 3408 16724 3460
rect 19524 3680 19576 3732
rect 21180 3680 21232 3732
rect 23480 3680 23532 3732
rect 25136 3680 25188 3732
rect 28080 3680 28132 3732
rect 29736 3723 29788 3732
rect 29736 3689 29745 3723
rect 29745 3689 29779 3723
rect 29779 3689 29788 3723
rect 29736 3680 29788 3689
rect 33324 3680 33376 3732
rect 34152 3680 34204 3732
rect 34888 3680 34940 3732
rect 39028 3723 39080 3732
rect 39028 3689 39037 3723
rect 39037 3689 39071 3723
rect 39071 3689 39080 3723
rect 39028 3680 39080 3689
rect 39396 3680 39448 3732
rect 39580 3680 39632 3732
rect 40408 3680 40460 3732
rect 41788 3723 41840 3732
rect 41788 3689 41797 3723
rect 41797 3689 41831 3723
rect 41831 3689 41840 3723
rect 41788 3680 41840 3689
rect 41972 3680 42024 3732
rect 41696 3612 41748 3664
rect 18788 3519 18840 3528
rect 18788 3485 18806 3519
rect 18806 3485 18840 3519
rect 18788 3476 18840 3485
rect 19432 3476 19484 3528
rect 19708 3476 19760 3528
rect 19892 3519 19944 3528
rect 19892 3485 19926 3519
rect 19926 3485 19944 3519
rect 19892 3476 19944 3485
rect 22192 3519 22244 3528
rect 22192 3485 22210 3519
rect 22210 3485 22244 3519
rect 22192 3476 22244 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 20812 3408 20864 3460
rect 16396 3340 16448 3392
rect 21088 3383 21140 3392
rect 21088 3349 21097 3383
rect 21097 3349 21131 3383
rect 21131 3349 21140 3383
rect 21088 3340 21140 3349
rect 23020 3408 23072 3460
rect 25504 3476 25556 3528
rect 26792 3476 26844 3528
rect 27988 3476 28040 3528
rect 28816 3519 28868 3528
rect 28816 3485 28825 3519
rect 28825 3485 28859 3519
rect 28859 3485 28868 3519
rect 28816 3476 28868 3485
rect 29092 3476 29144 3528
rect 34704 3519 34756 3528
rect 34704 3485 34713 3519
rect 34713 3485 34747 3519
rect 34747 3485 34756 3519
rect 34704 3476 34756 3485
rect 24860 3408 24912 3460
rect 25596 3408 25648 3460
rect 32864 3408 32916 3460
rect 33600 3408 33652 3460
rect 35716 3408 35768 3460
rect 26608 3340 26660 3392
rect 27896 3383 27948 3392
rect 27896 3349 27905 3383
rect 27905 3349 27939 3383
rect 27939 3349 27948 3383
rect 27896 3340 27948 3349
rect 31944 3340 31996 3392
rect 37740 3476 37792 3528
rect 39764 3544 39816 3596
rect 39120 3519 39172 3528
rect 39120 3485 39129 3519
rect 39129 3485 39163 3519
rect 39163 3485 39172 3519
rect 39120 3476 39172 3485
rect 39856 3519 39908 3528
rect 39856 3485 39865 3519
rect 39865 3485 39899 3519
rect 39899 3485 39908 3519
rect 39856 3476 39908 3485
rect 37096 3451 37148 3460
rect 37096 3417 37105 3451
rect 37105 3417 37139 3451
rect 37139 3417 37148 3451
rect 37096 3408 37148 3417
rect 36820 3340 36872 3392
rect 40408 3340 40460 3392
rect 42340 3587 42392 3596
rect 42340 3553 42349 3587
rect 42349 3553 42383 3587
rect 42383 3553 42392 3587
rect 42340 3544 42392 3553
rect 42892 3723 42944 3732
rect 42892 3689 42901 3723
rect 42901 3689 42935 3723
rect 42935 3689 42944 3723
rect 42892 3680 42944 3689
rect 43168 3680 43220 3732
rect 43352 3680 43404 3732
rect 44548 3723 44600 3732
rect 44548 3689 44557 3723
rect 44557 3689 44591 3723
rect 44591 3689 44600 3723
rect 44548 3680 44600 3689
rect 46664 3680 46716 3732
rect 48964 3680 49016 3732
rect 49884 3680 49936 3732
rect 52736 3680 52788 3732
rect 52920 3680 52972 3732
rect 53196 3723 53248 3732
rect 53196 3689 53205 3723
rect 53205 3689 53239 3723
rect 53239 3689 53248 3723
rect 53196 3680 53248 3689
rect 41880 3476 41932 3528
rect 42248 3519 42300 3528
rect 42248 3485 42257 3519
rect 42257 3485 42291 3519
rect 42291 3485 42300 3519
rect 42248 3476 42300 3485
rect 44272 3587 44324 3596
rect 44272 3553 44281 3587
rect 44281 3553 44315 3587
rect 44315 3553 44324 3587
rect 44272 3544 44324 3553
rect 41144 3408 41196 3460
rect 43812 3408 43864 3460
rect 44824 3476 44876 3528
rect 48504 3476 48556 3528
rect 50252 3544 50304 3596
rect 53932 3680 53984 3732
rect 54852 3612 54904 3664
rect 54944 3655 54996 3664
rect 54944 3621 54953 3655
rect 54953 3621 54987 3655
rect 54987 3621 54996 3655
rect 54944 3612 54996 3621
rect 55588 3612 55640 3664
rect 49148 3476 49200 3528
rect 44916 3408 44968 3460
rect 45468 3408 45520 3460
rect 47584 3408 47636 3460
rect 41696 3340 41748 3392
rect 41880 3383 41932 3392
rect 41880 3349 41889 3383
rect 41889 3349 41923 3383
rect 41923 3349 41932 3383
rect 41880 3340 41932 3349
rect 46112 3340 46164 3392
rect 47676 3340 47728 3392
rect 48780 3340 48832 3392
rect 50528 3519 50580 3528
rect 50528 3485 50537 3519
rect 50537 3485 50571 3519
rect 50571 3485 50580 3519
rect 50528 3476 50580 3485
rect 51172 3476 51224 3528
rect 54300 3544 54352 3596
rect 53380 3476 53432 3528
rect 53564 3519 53616 3528
rect 53564 3485 53598 3519
rect 53598 3485 53616 3519
rect 53564 3476 53616 3485
rect 56508 3680 56560 3732
rect 57888 3680 57940 3732
rect 57796 3612 57848 3664
rect 58164 3587 58216 3596
rect 58164 3553 58173 3587
rect 58173 3553 58207 3587
rect 58207 3553 58216 3587
rect 58164 3544 58216 3553
rect 54208 3408 54260 3460
rect 57704 3476 57756 3528
rect 58072 3519 58124 3528
rect 58072 3485 58081 3519
rect 58081 3485 58115 3519
rect 58115 3485 58124 3519
rect 58072 3476 58124 3485
rect 56600 3408 56652 3460
rect 56692 3408 56744 3460
rect 57428 3408 57480 3460
rect 55496 3340 55548 3392
rect 57704 3340 57756 3392
rect 58532 3340 58584 3392
rect 15394 3238 15446 3290
rect 15458 3238 15510 3290
rect 15522 3238 15574 3290
rect 15586 3238 15638 3290
rect 15650 3238 15702 3290
rect 29838 3238 29890 3290
rect 29902 3238 29954 3290
rect 29966 3238 30018 3290
rect 30030 3238 30082 3290
rect 30094 3238 30146 3290
rect 44282 3238 44334 3290
rect 44346 3238 44398 3290
rect 44410 3238 44462 3290
rect 44474 3238 44526 3290
rect 44538 3238 44590 3290
rect 58726 3238 58778 3290
rect 58790 3238 58842 3290
rect 58854 3238 58906 3290
rect 58918 3238 58970 3290
rect 58982 3238 59034 3290
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 2780 3136 2832 3145
rect 2872 3136 2924 3188
rect 5080 3136 5132 3188
rect 1584 3111 1636 3120
rect 1584 3077 1593 3111
rect 1593 3077 1627 3111
rect 1627 3077 1636 3111
rect 1584 3068 1636 3077
rect 1676 3000 1728 3052
rect 2228 3000 2280 3052
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 5816 3111 5868 3120
rect 5816 3077 5825 3111
rect 5825 3077 5859 3111
rect 5859 3077 5868 3111
rect 5816 3068 5868 3077
rect 5724 3000 5776 3052
rect 6000 3000 6052 3052
rect 6644 3043 6696 3052
rect 6644 3009 6678 3043
rect 6678 3009 6696 3043
rect 5540 2932 5592 2984
rect 6000 2864 6052 2916
rect 5632 2796 5684 2848
rect 6644 3000 6696 3009
rect 7288 3136 7340 3188
rect 7932 3136 7984 3188
rect 11980 3179 12032 3188
rect 11980 3145 11989 3179
rect 11989 3145 12023 3179
rect 12023 3145 12032 3179
rect 11980 3136 12032 3145
rect 12072 3136 12124 3188
rect 15384 3136 15436 3188
rect 16396 3179 16448 3188
rect 16396 3145 16405 3179
rect 16405 3145 16439 3179
rect 16439 3145 16448 3179
rect 16396 3136 16448 3145
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 21456 3136 21508 3188
rect 22284 3136 22336 3188
rect 23112 3136 23164 3188
rect 25228 3136 25280 3188
rect 26056 3136 26108 3188
rect 26240 3136 26292 3188
rect 27068 3136 27120 3188
rect 27896 3136 27948 3188
rect 28816 3136 28868 3188
rect 31484 3136 31536 3188
rect 31576 3136 31628 3188
rect 32496 3179 32548 3188
rect 32496 3145 32505 3179
rect 32505 3145 32539 3179
rect 32539 3145 32548 3179
rect 32496 3136 32548 3145
rect 33140 3136 33192 3188
rect 33232 3136 33284 3188
rect 34336 3136 34388 3188
rect 35992 3179 36044 3188
rect 35992 3145 36001 3179
rect 36001 3145 36035 3179
rect 36035 3145 36044 3179
rect 35992 3136 36044 3145
rect 36360 3136 36412 3188
rect 36912 3136 36964 3188
rect 39672 3136 39724 3188
rect 39856 3136 39908 3188
rect 8024 3068 8076 3120
rect 8576 3000 8628 3052
rect 10968 3068 11020 3120
rect 11244 3000 11296 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 12532 3000 12584 3052
rect 13268 3043 13320 3052
rect 15844 3068 15896 3120
rect 13268 3009 13286 3043
rect 13286 3009 13320 3043
rect 13268 3000 13320 3009
rect 15200 3000 15252 3052
rect 15752 3043 15804 3052
rect 15752 3009 15754 3043
rect 15754 3009 15788 3043
rect 15788 3009 15804 3043
rect 15752 3000 15804 3009
rect 11336 2864 11388 2916
rect 11152 2796 11204 2848
rect 12900 2796 12952 2848
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17960 3068 18012 3120
rect 17868 3000 17920 3052
rect 19984 3000 20036 3052
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 18788 2932 18840 2984
rect 16304 2796 16356 2848
rect 18880 2796 18932 2848
rect 21456 3000 21508 3052
rect 21088 2975 21140 2984
rect 21088 2941 21097 2975
rect 21097 2941 21131 2975
rect 21131 2941 21140 2975
rect 21088 2932 21140 2941
rect 22192 2864 22244 2916
rect 24032 2975 24084 2984
rect 24032 2941 24041 2975
rect 24041 2941 24075 2975
rect 24075 2941 24084 2975
rect 24032 2932 24084 2941
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 25044 3000 25096 3009
rect 29000 3068 29052 3120
rect 28080 3000 28132 3052
rect 28448 3000 28500 3052
rect 26700 2932 26752 2984
rect 27068 2932 27120 2984
rect 30932 2975 30984 2984
rect 30932 2941 30941 2975
rect 30941 2941 30975 2975
rect 30975 2941 30984 2975
rect 30932 2932 30984 2941
rect 24584 2864 24636 2916
rect 33416 3111 33468 3120
rect 33416 3077 33425 3111
rect 33425 3077 33459 3111
rect 33459 3077 33468 3111
rect 33416 3068 33468 3077
rect 33600 3068 33652 3120
rect 34980 3068 35032 3120
rect 35348 3068 35400 3120
rect 37096 3068 37148 3120
rect 37740 3068 37792 3120
rect 42156 3136 42208 3188
rect 42800 3136 42852 3188
rect 47216 3136 47268 3188
rect 48136 3136 48188 3188
rect 34704 3000 34756 3052
rect 36820 3043 36872 3052
rect 36820 3009 36829 3043
rect 36829 3009 36863 3043
rect 36863 3009 36872 3043
rect 36820 3000 36872 3009
rect 38568 3000 38620 3052
rect 40408 3043 40460 3052
rect 40408 3009 40417 3043
rect 40417 3009 40451 3043
rect 40451 3009 40460 3043
rect 40408 3000 40460 3009
rect 40960 3000 41012 3052
rect 44640 3068 44692 3120
rect 31944 2932 31996 2984
rect 33048 2932 33100 2984
rect 36360 2932 36412 2984
rect 39488 2975 39540 2984
rect 39488 2941 39497 2975
rect 39497 2941 39531 2975
rect 39531 2941 39540 2975
rect 39488 2932 39540 2941
rect 42984 3000 43036 3052
rect 45100 3043 45152 3052
rect 45100 3009 45109 3043
rect 45109 3009 45143 3043
rect 45143 3009 45152 3043
rect 45100 3000 45152 3009
rect 46296 3043 46348 3052
rect 46296 3009 46305 3043
rect 46305 3009 46339 3043
rect 46339 3009 46348 3043
rect 46296 3000 46348 3009
rect 47584 3111 47636 3120
rect 47584 3077 47593 3111
rect 47593 3077 47627 3111
rect 47627 3077 47636 3111
rect 47584 3068 47636 3077
rect 47676 3068 47728 3120
rect 48320 3068 48372 3120
rect 42800 2932 42852 2984
rect 35992 2864 36044 2916
rect 36820 2864 36872 2916
rect 41972 2864 42024 2916
rect 43628 2932 43680 2984
rect 42984 2864 43036 2916
rect 46572 2932 46624 2984
rect 47216 3000 47268 3052
rect 48504 3043 48556 3052
rect 48504 3009 48520 3043
rect 48520 3009 48554 3043
rect 48554 3009 48556 3043
rect 48504 3000 48556 3009
rect 50528 3136 50580 3188
rect 50988 3179 51040 3188
rect 50988 3145 50997 3179
rect 50997 3145 51031 3179
rect 51031 3145 51040 3179
rect 50988 3136 51040 3145
rect 51172 3136 51224 3188
rect 50436 3068 50488 3120
rect 55680 3136 55732 3188
rect 56140 3179 56192 3188
rect 56140 3145 56149 3179
rect 56149 3145 56183 3179
rect 56183 3145 56192 3179
rect 56140 3136 56192 3145
rect 56508 3136 56560 3188
rect 56692 3136 56744 3188
rect 52368 3000 52420 3052
rect 48320 2864 48372 2916
rect 23756 2839 23808 2848
rect 23756 2805 23765 2839
rect 23765 2805 23799 2839
rect 23799 2805 23808 2839
rect 23756 2796 23808 2805
rect 47768 2796 47820 2848
rect 47860 2796 47912 2848
rect 51080 2864 51132 2916
rect 53104 3043 53156 3052
rect 53104 3009 53113 3043
rect 53113 3009 53147 3043
rect 53147 3009 53156 3043
rect 53104 3000 53156 3009
rect 53196 3043 53248 3052
rect 53196 3009 53205 3043
rect 53205 3009 53239 3043
rect 53239 3009 53248 3043
rect 53196 3000 53248 3009
rect 53012 2975 53064 2984
rect 53012 2941 53021 2975
rect 53021 2941 53055 2975
rect 53055 2941 53064 2975
rect 53012 2932 53064 2941
rect 53564 2932 53616 2984
rect 56784 3068 56836 3120
rect 58256 2932 58308 2984
rect 49976 2839 50028 2848
rect 49976 2805 49985 2839
rect 49985 2805 50019 2839
rect 50019 2805 50028 2839
rect 49976 2796 50028 2805
rect 51356 2796 51408 2848
rect 53748 2864 53800 2916
rect 54392 2864 54444 2916
rect 52828 2796 52880 2848
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 22616 2694 22668 2746
rect 22680 2694 22732 2746
rect 22744 2694 22796 2746
rect 22808 2694 22860 2746
rect 22872 2694 22924 2746
rect 37060 2694 37112 2746
rect 37124 2694 37176 2746
rect 37188 2694 37240 2746
rect 37252 2694 37304 2746
rect 37316 2694 37368 2746
rect 51504 2694 51556 2746
rect 51568 2694 51620 2746
rect 51632 2694 51684 2746
rect 51696 2694 51748 2746
rect 51760 2694 51812 2746
rect 2688 2592 2740 2644
rect 4436 2592 4488 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 9772 2592 9824 2644
rect 11796 2592 11848 2644
rect 16948 2592 17000 2644
rect 18880 2635 18932 2644
rect 18880 2601 18889 2635
rect 18889 2601 18923 2635
rect 18923 2601 18932 2635
rect 18880 2592 18932 2601
rect 21456 2592 21508 2644
rect 22376 2592 22428 2644
rect 25044 2592 25096 2644
rect 27160 2592 27212 2644
rect 29092 2592 29144 2644
rect 31668 2592 31720 2644
rect 34060 2592 34112 2644
rect 36176 2635 36228 2644
rect 36176 2601 36185 2635
rect 36185 2601 36219 2635
rect 36219 2601 36228 2635
rect 36176 2592 36228 2601
rect 39120 2592 39172 2644
rect 40960 2592 41012 2644
rect 42800 2592 42852 2644
rect 45284 2592 45336 2644
rect 47032 2635 47084 2644
rect 47032 2601 47041 2635
rect 47041 2601 47075 2635
rect 47075 2601 47084 2635
rect 47032 2592 47084 2601
rect 47400 2635 47452 2644
rect 47400 2601 47409 2635
rect 47409 2601 47443 2635
rect 47443 2601 47452 2635
rect 47400 2592 47452 2601
rect 48320 2592 48372 2644
rect 49976 2592 50028 2644
rect 51172 2592 51224 2644
rect 54208 2635 54260 2644
rect 54208 2601 54217 2635
rect 54217 2601 54251 2635
rect 54251 2601 54260 2635
rect 54208 2592 54260 2601
rect 57336 2592 57388 2644
rect 57796 2592 57848 2644
rect 16580 2524 16632 2576
rect 40500 2524 40552 2576
rect 3332 2456 3384 2508
rect 6460 2456 6512 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 3148 2388 3200 2440
rect 4896 2388 4948 2440
rect 3884 2320 3936 2372
rect 5908 2320 5960 2372
rect 6736 2363 6788 2372
rect 6736 2329 6745 2363
rect 6745 2329 6779 2363
rect 6779 2329 6788 2363
rect 6736 2320 6788 2329
rect 7196 2388 7248 2440
rect 12992 2456 13044 2508
rect 13820 2456 13872 2508
rect 15292 2456 15344 2508
rect 16672 2456 16724 2508
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 8852 2320 8904 2372
rect 10416 2363 10468 2372
rect 10416 2329 10425 2363
rect 10425 2329 10459 2363
rect 10459 2329 10468 2363
rect 10416 2320 10468 2329
rect 14004 2388 14056 2440
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 15384 2388 15436 2440
rect 17316 2456 17368 2508
rect 22100 2456 22152 2508
rect 28724 2499 28776 2508
rect 28724 2465 28733 2499
rect 28733 2465 28767 2499
rect 28767 2465 28776 2499
rect 28724 2456 28776 2465
rect 34060 2456 34112 2508
rect 37188 2456 37240 2508
rect 39028 2456 39080 2508
rect 42064 2456 42116 2508
rect 14280 2320 14332 2372
rect 20444 2363 20496 2372
rect 20444 2329 20453 2363
rect 20453 2329 20487 2363
rect 20487 2329 20496 2363
rect 20444 2320 20496 2329
rect 20996 2388 21048 2440
rect 21640 2388 21692 2440
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 23756 2388 23808 2440
rect 26056 2388 26108 2440
rect 26608 2431 26660 2440
rect 26608 2397 26617 2431
rect 26617 2397 26651 2431
rect 26651 2397 26660 2431
rect 26608 2388 26660 2397
rect 22652 2320 22704 2372
rect 25596 2363 25648 2372
rect 25596 2329 25605 2363
rect 25605 2329 25639 2363
rect 25639 2329 25648 2363
rect 25596 2320 25648 2329
rect 28172 2431 28224 2440
rect 28172 2397 28181 2431
rect 28181 2397 28215 2431
rect 28215 2397 28224 2431
rect 28172 2388 28224 2397
rect 31208 2388 31260 2440
rect 31944 2388 31996 2440
rect 33324 2431 33376 2440
rect 33324 2397 33333 2431
rect 33333 2397 33367 2431
rect 33367 2397 33376 2431
rect 33324 2388 33376 2397
rect 29368 2320 29420 2372
rect 30472 2320 30524 2372
rect 32036 2320 32088 2372
rect 32956 2320 33008 2372
rect 34796 2431 34848 2440
rect 34796 2397 34805 2431
rect 34805 2397 34839 2431
rect 34839 2397 34848 2431
rect 34796 2388 34848 2397
rect 34888 2388 34940 2440
rect 36820 2388 36872 2440
rect 37924 2388 37976 2440
rect 39672 2388 39724 2440
rect 40224 2388 40276 2440
rect 44180 2388 44232 2440
rect 9680 2252 9732 2304
rect 46664 2431 46716 2440
rect 46664 2397 46673 2431
rect 46673 2397 46707 2431
rect 46707 2397 46716 2431
rect 46664 2388 46716 2397
rect 48688 2456 48740 2508
rect 48780 2431 48832 2440
rect 48780 2397 48789 2431
rect 48789 2397 48823 2431
rect 48823 2397 48832 2431
rect 48780 2388 48832 2397
rect 50160 2431 50212 2440
rect 50160 2397 50169 2431
rect 50169 2397 50203 2431
rect 50203 2397 50212 2431
rect 50160 2388 50212 2397
rect 51080 2388 51132 2440
rect 52644 2388 52696 2440
rect 54760 2431 54812 2440
rect 54760 2397 54769 2431
rect 54769 2397 54803 2431
rect 54803 2397 54812 2431
rect 54760 2388 54812 2397
rect 57428 2499 57480 2508
rect 57428 2465 57437 2499
rect 57437 2465 57471 2499
rect 57471 2465 57480 2499
rect 57428 2456 57480 2465
rect 57612 2456 57664 2508
rect 58440 2499 58492 2508
rect 58440 2465 58449 2499
rect 58449 2465 58483 2499
rect 58483 2465 58492 2499
rect 58440 2456 58492 2465
rect 57244 2431 57296 2440
rect 57244 2397 57253 2431
rect 57253 2397 57287 2431
rect 57287 2397 57296 2431
rect 57244 2388 57296 2397
rect 45284 2320 45336 2372
rect 46940 2320 46992 2372
rect 52092 2320 52144 2372
rect 53656 2320 53708 2372
rect 55220 2320 55272 2372
rect 47584 2252 47636 2304
rect 15394 2150 15446 2202
rect 15458 2150 15510 2202
rect 15522 2150 15574 2202
rect 15586 2150 15638 2202
rect 15650 2150 15702 2202
rect 29838 2150 29890 2202
rect 29902 2150 29954 2202
rect 29966 2150 30018 2202
rect 30030 2150 30082 2202
rect 30094 2150 30146 2202
rect 44282 2150 44334 2202
rect 44346 2150 44398 2202
rect 44410 2150 44462 2202
rect 44474 2150 44526 2202
rect 44538 2150 44590 2202
rect 58726 2150 58778 2202
rect 58790 2150 58842 2202
rect 58854 2150 58906 2202
rect 58918 2150 58970 2202
rect 58982 2150 59034 2202
rect 2320 2048 2372 2100
rect 6368 2048 6420 2100
rect 14464 2048 14516 2100
rect 19616 2048 19668 2100
<< metal2 >>
rect 8172 27772 8480 27781
rect 8172 27770 8178 27772
rect 8234 27770 8258 27772
rect 8314 27770 8338 27772
rect 8394 27770 8418 27772
rect 8474 27770 8480 27772
rect 8234 27718 8236 27770
rect 8416 27718 8418 27770
rect 8172 27716 8178 27718
rect 8234 27716 8258 27718
rect 8314 27716 8338 27718
rect 8394 27716 8418 27718
rect 8474 27716 8480 27718
rect 8172 27707 8480 27716
rect 22616 27772 22924 27781
rect 22616 27770 22622 27772
rect 22678 27770 22702 27772
rect 22758 27770 22782 27772
rect 22838 27770 22862 27772
rect 22918 27770 22924 27772
rect 22678 27718 22680 27770
rect 22860 27718 22862 27770
rect 22616 27716 22622 27718
rect 22678 27716 22702 27718
rect 22758 27716 22782 27718
rect 22838 27716 22862 27718
rect 22918 27716 22924 27718
rect 22616 27707 22924 27716
rect 37060 27772 37368 27781
rect 37060 27770 37066 27772
rect 37122 27770 37146 27772
rect 37202 27770 37226 27772
rect 37282 27770 37306 27772
rect 37362 27770 37368 27772
rect 37122 27718 37124 27770
rect 37304 27718 37306 27770
rect 37060 27716 37066 27718
rect 37122 27716 37146 27718
rect 37202 27716 37226 27718
rect 37282 27716 37306 27718
rect 37362 27716 37368 27718
rect 37060 27707 37368 27716
rect 51504 27772 51812 27781
rect 51504 27770 51510 27772
rect 51566 27770 51590 27772
rect 51646 27770 51670 27772
rect 51726 27770 51750 27772
rect 51806 27770 51812 27772
rect 51566 27718 51568 27770
rect 51748 27718 51750 27770
rect 51504 27716 51510 27718
rect 51566 27716 51590 27718
rect 51646 27716 51670 27718
rect 51726 27716 51750 27718
rect 51806 27716 51812 27718
rect 51504 27707 51812 27716
rect 15394 27228 15702 27237
rect 15394 27226 15400 27228
rect 15456 27226 15480 27228
rect 15536 27226 15560 27228
rect 15616 27226 15640 27228
rect 15696 27226 15702 27228
rect 15456 27174 15458 27226
rect 15638 27174 15640 27226
rect 15394 27172 15400 27174
rect 15456 27172 15480 27174
rect 15536 27172 15560 27174
rect 15616 27172 15640 27174
rect 15696 27172 15702 27174
rect 15394 27163 15702 27172
rect 29838 27228 30146 27237
rect 29838 27226 29844 27228
rect 29900 27226 29924 27228
rect 29980 27226 30004 27228
rect 30060 27226 30084 27228
rect 30140 27226 30146 27228
rect 29900 27174 29902 27226
rect 30082 27174 30084 27226
rect 29838 27172 29844 27174
rect 29900 27172 29924 27174
rect 29980 27172 30004 27174
rect 30060 27172 30084 27174
rect 30140 27172 30146 27174
rect 29838 27163 30146 27172
rect 44282 27228 44590 27237
rect 44282 27226 44288 27228
rect 44344 27226 44368 27228
rect 44424 27226 44448 27228
rect 44504 27226 44528 27228
rect 44584 27226 44590 27228
rect 44344 27174 44346 27226
rect 44526 27174 44528 27226
rect 44282 27172 44288 27174
rect 44344 27172 44368 27174
rect 44424 27172 44448 27174
rect 44504 27172 44528 27174
rect 44584 27172 44590 27174
rect 44282 27163 44590 27172
rect 58726 27228 59034 27237
rect 58726 27226 58732 27228
rect 58788 27226 58812 27228
rect 58868 27226 58892 27228
rect 58948 27226 58972 27228
rect 59028 27226 59034 27228
rect 58788 27174 58790 27226
rect 58970 27174 58972 27226
rect 58726 27172 58732 27174
rect 58788 27172 58812 27174
rect 58868 27172 58892 27174
rect 58948 27172 58972 27174
rect 59028 27172 59034 27174
rect 58726 27163 59034 27172
rect 8172 26684 8480 26693
rect 8172 26682 8178 26684
rect 8234 26682 8258 26684
rect 8314 26682 8338 26684
rect 8394 26682 8418 26684
rect 8474 26682 8480 26684
rect 8234 26630 8236 26682
rect 8416 26630 8418 26682
rect 8172 26628 8178 26630
rect 8234 26628 8258 26630
rect 8314 26628 8338 26630
rect 8394 26628 8418 26630
rect 8474 26628 8480 26630
rect 8172 26619 8480 26628
rect 22616 26684 22924 26693
rect 22616 26682 22622 26684
rect 22678 26682 22702 26684
rect 22758 26682 22782 26684
rect 22838 26682 22862 26684
rect 22918 26682 22924 26684
rect 22678 26630 22680 26682
rect 22860 26630 22862 26682
rect 22616 26628 22622 26630
rect 22678 26628 22702 26630
rect 22758 26628 22782 26630
rect 22838 26628 22862 26630
rect 22918 26628 22924 26630
rect 22616 26619 22924 26628
rect 37060 26684 37368 26693
rect 37060 26682 37066 26684
rect 37122 26682 37146 26684
rect 37202 26682 37226 26684
rect 37282 26682 37306 26684
rect 37362 26682 37368 26684
rect 37122 26630 37124 26682
rect 37304 26630 37306 26682
rect 37060 26628 37066 26630
rect 37122 26628 37146 26630
rect 37202 26628 37226 26630
rect 37282 26628 37306 26630
rect 37362 26628 37368 26630
rect 37060 26619 37368 26628
rect 51504 26684 51812 26693
rect 51504 26682 51510 26684
rect 51566 26682 51590 26684
rect 51646 26682 51670 26684
rect 51726 26682 51750 26684
rect 51806 26682 51812 26684
rect 51566 26630 51568 26682
rect 51748 26630 51750 26682
rect 51504 26628 51510 26630
rect 51566 26628 51590 26630
rect 51646 26628 51670 26630
rect 51726 26628 51750 26630
rect 51806 26628 51812 26630
rect 51504 26619 51812 26628
rect 15394 26140 15702 26149
rect 15394 26138 15400 26140
rect 15456 26138 15480 26140
rect 15536 26138 15560 26140
rect 15616 26138 15640 26140
rect 15696 26138 15702 26140
rect 15456 26086 15458 26138
rect 15638 26086 15640 26138
rect 15394 26084 15400 26086
rect 15456 26084 15480 26086
rect 15536 26084 15560 26086
rect 15616 26084 15640 26086
rect 15696 26084 15702 26086
rect 15394 26075 15702 26084
rect 29838 26140 30146 26149
rect 29838 26138 29844 26140
rect 29900 26138 29924 26140
rect 29980 26138 30004 26140
rect 30060 26138 30084 26140
rect 30140 26138 30146 26140
rect 29900 26086 29902 26138
rect 30082 26086 30084 26138
rect 29838 26084 29844 26086
rect 29900 26084 29924 26086
rect 29980 26084 30004 26086
rect 30060 26084 30084 26086
rect 30140 26084 30146 26086
rect 29838 26075 30146 26084
rect 44282 26140 44590 26149
rect 44282 26138 44288 26140
rect 44344 26138 44368 26140
rect 44424 26138 44448 26140
rect 44504 26138 44528 26140
rect 44584 26138 44590 26140
rect 44344 26086 44346 26138
rect 44526 26086 44528 26138
rect 44282 26084 44288 26086
rect 44344 26084 44368 26086
rect 44424 26084 44448 26086
rect 44504 26084 44528 26086
rect 44584 26084 44590 26086
rect 44282 26075 44590 26084
rect 58726 26140 59034 26149
rect 58726 26138 58732 26140
rect 58788 26138 58812 26140
rect 58868 26138 58892 26140
rect 58948 26138 58972 26140
rect 59028 26138 59034 26140
rect 58788 26086 58790 26138
rect 58970 26086 58972 26138
rect 58726 26084 58732 26086
rect 58788 26084 58812 26086
rect 58868 26084 58892 26086
rect 58948 26084 58972 26086
rect 59028 26084 59034 26086
rect 58726 26075 59034 26084
rect 8172 25596 8480 25605
rect 8172 25594 8178 25596
rect 8234 25594 8258 25596
rect 8314 25594 8338 25596
rect 8394 25594 8418 25596
rect 8474 25594 8480 25596
rect 8234 25542 8236 25594
rect 8416 25542 8418 25594
rect 8172 25540 8178 25542
rect 8234 25540 8258 25542
rect 8314 25540 8338 25542
rect 8394 25540 8418 25542
rect 8474 25540 8480 25542
rect 8172 25531 8480 25540
rect 22616 25596 22924 25605
rect 22616 25594 22622 25596
rect 22678 25594 22702 25596
rect 22758 25594 22782 25596
rect 22838 25594 22862 25596
rect 22918 25594 22924 25596
rect 22678 25542 22680 25594
rect 22860 25542 22862 25594
rect 22616 25540 22622 25542
rect 22678 25540 22702 25542
rect 22758 25540 22782 25542
rect 22838 25540 22862 25542
rect 22918 25540 22924 25542
rect 22616 25531 22924 25540
rect 37060 25596 37368 25605
rect 37060 25594 37066 25596
rect 37122 25594 37146 25596
rect 37202 25594 37226 25596
rect 37282 25594 37306 25596
rect 37362 25594 37368 25596
rect 37122 25542 37124 25594
rect 37304 25542 37306 25594
rect 37060 25540 37066 25542
rect 37122 25540 37146 25542
rect 37202 25540 37226 25542
rect 37282 25540 37306 25542
rect 37362 25540 37368 25542
rect 37060 25531 37368 25540
rect 51504 25596 51812 25605
rect 51504 25594 51510 25596
rect 51566 25594 51590 25596
rect 51646 25594 51670 25596
rect 51726 25594 51750 25596
rect 51806 25594 51812 25596
rect 51566 25542 51568 25594
rect 51748 25542 51750 25594
rect 51504 25540 51510 25542
rect 51566 25540 51590 25542
rect 51646 25540 51670 25542
rect 51726 25540 51750 25542
rect 51806 25540 51812 25542
rect 51504 25531 51812 25540
rect 15394 25052 15702 25061
rect 15394 25050 15400 25052
rect 15456 25050 15480 25052
rect 15536 25050 15560 25052
rect 15616 25050 15640 25052
rect 15696 25050 15702 25052
rect 15456 24998 15458 25050
rect 15638 24998 15640 25050
rect 15394 24996 15400 24998
rect 15456 24996 15480 24998
rect 15536 24996 15560 24998
rect 15616 24996 15640 24998
rect 15696 24996 15702 24998
rect 15394 24987 15702 24996
rect 29838 25052 30146 25061
rect 29838 25050 29844 25052
rect 29900 25050 29924 25052
rect 29980 25050 30004 25052
rect 30060 25050 30084 25052
rect 30140 25050 30146 25052
rect 29900 24998 29902 25050
rect 30082 24998 30084 25050
rect 29838 24996 29844 24998
rect 29900 24996 29924 24998
rect 29980 24996 30004 24998
rect 30060 24996 30084 24998
rect 30140 24996 30146 24998
rect 29838 24987 30146 24996
rect 44282 25052 44590 25061
rect 44282 25050 44288 25052
rect 44344 25050 44368 25052
rect 44424 25050 44448 25052
rect 44504 25050 44528 25052
rect 44584 25050 44590 25052
rect 44344 24998 44346 25050
rect 44526 24998 44528 25050
rect 44282 24996 44288 24998
rect 44344 24996 44368 24998
rect 44424 24996 44448 24998
rect 44504 24996 44528 24998
rect 44584 24996 44590 24998
rect 44282 24987 44590 24996
rect 58726 25052 59034 25061
rect 58726 25050 58732 25052
rect 58788 25050 58812 25052
rect 58868 25050 58892 25052
rect 58948 25050 58972 25052
rect 59028 25050 59034 25052
rect 58788 24998 58790 25050
rect 58970 24998 58972 25050
rect 58726 24996 58732 24998
rect 58788 24996 58812 24998
rect 58868 24996 58892 24998
rect 58948 24996 58972 24998
rect 59028 24996 59034 24998
rect 58726 24987 59034 24996
rect 8172 24508 8480 24517
rect 8172 24506 8178 24508
rect 8234 24506 8258 24508
rect 8314 24506 8338 24508
rect 8394 24506 8418 24508
rect 8474 24506 8480 24508
rect 8234 24454 8236 24506
rect 8416 24454 8418 24506
rect 8172 24452 8178 24454
rect 8234 24452 8258 24454
rect 8314 24452 8338 24454
rect 8394 24452 8418 24454
rect 8474 24452 8480 24454
rect 8172 24443 8480 24452
rect 22616 24508 22924 24517
rect 22616 24506 22622 24508
rect 22678 24506 22702 24508
rect 22758 24506 22782 24508
rect 22838 24506 22862 24508
rect 22918 24506 22924 24508
rect 22678 24454 22680 24506
rect 22860 24454 22862 24506
rect 22616 24452 22622 24454
rect 22678 24452 22702 24454
rect 22758 24452 22782 24454
rect 22838 24452 22862 24454
rect 22918 24452 22924 24454
rect 22616 24443 22924 24452
rect 37060 24508 37368 24517
rect 37060 24506 37066 24508
rect 37122 24506 37146 24508
rect 37202 24506 37226 24508
rect 37282 24506 37306 24508
rect 37362 24506 37368 24508
rect 37122 24454 37124 24506
rect 37304 24454 37306 24506
rect 37060 24452 37066 24454
rect 37122 24452 37146 24454
rect 37202 24452 37226 24454
rect 37282 24452 37306 24454
rect 37362 24452 37368 24454
rect 37060 24443 37368 24452
rect 51504 24508 51812 24517
rect 51504 24506 51510 24508
rect 51566 24506 51590 24508
rect 51646 24506 51670 24508
rect 51726 24506 51750 24508
rect 51806 24506 51812 24508
rect 51566 24454 51568 24506
rect 51748 24454 51750 24506
rect 51504 24452 51510 24454
rect 51566 24452 51590 24454
rect 51646 24452 51670 24454
rect 51726 24452 51750 24454
rect 51806 24452 51812 24454
rect 51504 24443 51812 24452
rect 15394 23964 15702 23973
rect 15394 23962 15400 23964
rect 15456 23962 15480 23964
rect 15536 23962 15560 23964
rect 15616 23962 15640 23964
rect 15696 23962 15702 23964
rect 15456 23910 15458 23962
rect 15638 23910 15640 23962
rect 15394 23908 15400 23910
rect 15456 23908 15480 23910
rect 15536 23908 15560 23910
rect 15616 23908 15640 23910
rect 15696 23908 15702 23910
rect 15394 23899 15702 23908
rect 29838 23964 30146 23973
rect 29838 23962 29844 23964
rect 29900 23962 29924 23964
rect 29980 23962 30004 23964
rect 30060 23962 30084 23964
rect 30140 23962 30146 23964
rect 29900 23910 29902 23962
rect 30082 23910 30084 23962
rect 29838 23908 29844 23910
rect 29900 23908 29924 23910
rect 29980 23908 30004 23910
rect 30060 23908 30084 23910
rect 30140 23908 30146 23910
rect 29838 23899 30146 23908
rect 44282 23964 44590 23973
rect 44282 23962 44288 23964
rect 44344 23962 44368 23964
rect 44424 23962 44448 23964
rect 44504 23962 44528 23964
rect 44584 23962 44590 23964
rect 44344 23910 44346 23962
rect 44526 23910 44528 23962
rect 44282 23908 44288 23910
rect 44344 23908 44368 23910
rect 44424 23908 44448 23910
rect 44504 23908 44528 23910
rect 44584 23908 44590 23910
rect 44282 23899 44590 23908
rect 58726 23964 59034 23973
rect 58726 23962 58732 23964
rect 58788 23962 58812 23964
rect 58868 23962 58892 23964
rect 58948 23962 58972 23964
rect 59028 23962 59034 23964
rect 58788 23910 58790 23962
rect 58970 23910 58972 23962
rect 58726 23908 58732 23910
rect 58788 23908 58812 23910
rect 58868 23908 58892 23910
rect 58948 23908 58972 23910
rect 59028 23908 59034 23910
rect 58726 23899 59034 23908
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18236 23656 18288 23662
rect 18236 23598 18288 23604
rect 47584 23656 47636 23662
rect 47584 23598 47636 23604
rect 53288 23656 53340 23662
rect 53288 23598 53340 23604
rect 54024 23656 54076 23662
rect 54024 23598 54076 23604
rect 14556 23520 14608 23526
rect 14556 23462 14608 23468
rect 8172 23420 8480 23429
rect 8172 23418 8178 23420
rect 8234 23418 8258 23420
rect 8314 23418 8338 23420
rect 8394 23418 8418 23420
rect 8474 23418 8480 23420
rect 8234 23366 8236 23418
rect 8416 23366 8418 23418
rect 8172 23364 8178 23366
rect 8234 23364 8258 23366
rect 8314 23364 8338 23366
rect 8394 23364 8418 23366
rect 8474 23364 8480 23366
rect 8172 23355 8480 23364
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 4436 22568 4488 22574
rect 4436 22510 4488 22516
rect 3056 22432 3108 22438
rect 3056 22374 3108 22380
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 2976 21690 3004 21966
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 3068 21622 3096 22374
rect 3712 22234 3740 22510
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3056 21616 3108 21622
rect 3896 21570 3924 22374
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 3056 21558 3108 21564
rect 3712 21554 3924 21570
rect 4264 21554 4292 21830
rect 3700 21548 3924 21554
rect 3752 21542 3924 21548
rect 4252 21548 4304 21554
rect 3700 21490 3752 21496
rect 4252 21490 4304 21496
rect 4264 20806 4292 21490
rect 4448 21146 4476 22510
rect 4896 22500 4948 22506
rect 4896 22442 4948 22448
rect 4908 22234 4936 22442
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4632 21010 4660 21830
rect 4724 21690 4752 21966
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 5000 20942 5028 21830
rect 5276 21078 5304 21830
rect 5736 21690 5764 22374
rect 6104 21962 6132 22918
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 4264 19718 4292 20742
rect 5920 20482 5948 20878
rect 6196 20806 6224 21490
rect 6472 21486 6500 21966
rect 6656 21690 6684 23054
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 7116 22234 7144 22510
rect 9220 22432 9272 22438
rect 9220 22374 9272 22380
rect 8172 22332 8480 22341
rect 8172 22330 8178 22332
rect 8234 22330 8258 22332
rect 8314 22330 8338 22332
rect 8394 22330 8418 22332
rect 8474 22330 8480 22332
rect 8234 22278 8236 22330
rect 8416 22278 8418 22330
rect 8172 22276 8178 22278
rect 8234 22276 8258 22278
rect 8314 22276 8338 22278
rect 8394 22276 8418 22278
rect 8474 22276 8480 22278
rect 8172 22267 8480 22276
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 6644 21684 6696 21690
rect 6644 21626 6696 21632
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6104 20602 6132 20742
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 5828 20454 5948 20482
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4540 20058 4568 20334
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2424 17134 2452 19314
rect 2792 18970 2820 19314
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 4264 18698 4292 19654
rect 4816 19514 4844 19790
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 5092 19378 5120 20198
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 4816 18426 4844 18770
rect 5828 18766 5856 20454
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5920 18970 5948 20334
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6012 18834 6040 19110
rect 6104 18834 6132 19722
rect 6472 19718 6500 21422
rect 7116 21010 7144 22170
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7208 21690 7236 21830
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 7760 21146 7788 21966
rect 9048 21350 9076 21966
rect 9232 21622 9260 22374
rect 9784 22234 9812 22510
rect 9956 22500 10008 22506
rect 9956 22442 10008 22448
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9876 21622 9904 21830
rect 9220 21616 9272 21622
rect 9220 21558 9272 21564
rect 9864 21616 9916 21622
rect 9864 21558 9916 21564
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 7944 21146 7972 21286
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7024 20602 7052 20946
rect 9048 20942 9076 21286
rect 9036 20936 9088 20942
rect 9088 20884 9168 20890
rect 9036 20878 9168 20884
rect 9048 20862 9168 20878
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19378 6500 19654
rect 6564 19417 6592 20198
rect 6550 19408 6606 19417
rect 6460 19372 6512 19378
rect 6550 19343 6606 19352
rect 6460 19314 6512 19320
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5816 18760 5868 18766
rect 5868 18708 6040 18714
rect 5816 18702 6040 18708
rect 5828 18686 6040 18702
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 17338 3004 17478
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 1596 16658 1624 17070
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2516 16250 2544 16458
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2976 16250 3004 16390
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3068 16114 3096 16390
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 15162 2636 15438
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2884 15162 2912 15370
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 3056 15156 3108 15162
rect 3108 15116 3280 15144
rect 3056 15098 3108 15104
rect 3252 15026 3280 15116
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 2792 14890 2820 14962
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13394 2636 13670
rect 2792 13530 2820 14826
rect 3160 14618 3188 14962
rect 3344 14958 3372 16526
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16250 3464 16390
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3436 15638 3464 16186
rect 3528 15706 3556 17614
rect 3804 17338 3832 17614
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16726 3924 17070
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 4264 15502 4292 17478
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4540 16182 4568 16934
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4540 15638 4568 16118
rect 4632 16114 4660 16390
rect 4908 16250 4936 16458
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4356 15162 4384 15438
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 14618 3372 14894
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3344 14498 3372 14554
rect 3528 14550 3556 15098
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3516 14544 3568 14550
rect 3344 14470 3464 14498
rect 3516 14486 3568 14492
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 14074 3372 14214
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3436 13530 3464 14470
rect 3896 14414 3924 14894
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3988 14414 4016 14758
rect 4080 14618 4108 14758
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3620 13938 3648 14282
rect 3896 13938 3924 14350
rect 3988 14006 4016 14350
rect 4356 14074 4384 15098
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 13530 4108 13806
rect 4448 13530 4476 15438
rect 4632 15366 4660 16050
rect 5368 15706 5396 16050
rect 5552 15706 5580 16390
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 15162 4660 15302
rect 4724 15162 4752 15438
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14346 4568 14758
rect 4724 14618 4752 15098
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2608 12306 2636 13330
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2976 11898 3004 13262
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3436 12186 3464 12650
rect 3528 12374 3556 13262
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4080 12986 4108 13194
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3804 12238 3832 12718
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 3516 12232 3568 12238
rect 3436 12180 3516 12186
rect 3436 12174 3568 12180
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3436 12158 3556 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1412 800 1440 3431
rect 1596 3126 1624 10474
rect 2608 10470 2636 10950
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2424 10130 2452 10406
rect 2700 10266 2728 10474
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2044 9580 2096 9586
rect 2148 9568 2176 10066
rect 3068 9654 3096 10406
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 2096 9540 2176 9568
rect 2044 9522 2096 9528
rect 2148 7342 2176 9540
rect 3344 9450 3372 11698
rect 3528 10606 3556 12158
rect 3804 11898 3832 12174
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3896 11762 3924 12174
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4172 11558 4200 12038
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3528 10266 3556 10542
rect 3712 10266 3740 10542
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3804 9450 3832 11018
rect 4172 9654 4200 11222
rect 4264 11014 4292 12378
rect 4620 12096 4672 12102
rect 4724 12084 4752 13262
rect 5184 12442 5212 15370
rect 5552 15026 5580 15370
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5552 14634 5580 14962
rect 5644 14958 5672 16050
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15162 5764 15302
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5460 14606 5580 14634
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5460 12186 5488 14606
rect 5736 13002 5764 15098
rect 5184 12170 5488 12186
rect 5172 12164 5488 12170
rect 5224 12158 5488 12164
rect 5552 12974 5764 13002
rect 5172 12106 5224 12112
rect 4672 12056 4752 12084
rect 4620 12038 4672 12044
rect 4632 11354 4660 12038
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4264 10282 4292 10950
rect 4448 10470 4476 10950
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4264 10254 4476 10282
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4264 9722 4292 9998
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3804 8974 3832 9386
rect 4448 9382 4476 10254
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 8974 4476 9318
rect 4540 9042 4568 10134
rect 4632 9586 4660 11290
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10062 4752 11154
rect 5184 11014 5212 12106
rect 5552 11898 5580 12974
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12238 5764 12582
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5172 11008 5224 11014
rect 5224 10968 5304 10996
rect 5172 10950 5224 10956
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4816 9722 4844 10542
rect 4908 10266 4936 10610
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 5000 9654 5028 10406
rect 5184 9654 5212 10678
rect 5276 10470 5304 10968
rect 5368 10810 5396 11086
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 10130 5304 10406
rect 5460 10198 5488 10950
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5276 9586 5304 9930
rect 5460 9722 5488 10134
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2148 6798 2176 7278
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5914 1900 6054
rect 2148 5914 2176 6734
rect 2976 6730 3004 7686
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 3160 6458 3188 7346
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 7002 3648 7278
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3804 6322 3832 6598
rect 3896 6322 3924 7142
rect 4172 6746 4200 7686
rect 4264 7546 4292 7686
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4172 6718 4292 6746
rect 4264 6662 4292 6718
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4172 6458 4200 6598
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 2332 5914 2360 6190
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2148 4826 2176 5850
rect 3344 5846 3372 6054
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 4080 5710 4108 6190
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3068 5370 3096 5578
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 3534 1716 4626
rect 2332 4554 2360 4966
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3534 1900 3878
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1584 3120 1636 3126
rect 1584 3062 1636 3068
rect 1688 3058 1716 3470
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2240 800 2268 2994
rect 2700 2650 2728 4490
rect 2976 4282 3004 5102
rect 3620 4486 3648 5306
rect 3712 5166 3740 5510
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4826 3832 5102
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3896 4758 3924 5238
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3988 4622 4016 4927
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2792 3194 2820 4150
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3194 2912 3878
rect 3252 3738 3280 3946
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3620 3602 3648 4422
rect 4080 4078 4108 5646
rect 4264 5574 4292 6598
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4356 5574 4384 6326
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4264 4282 4292 5510
rect 4356 5250 4384 5510
rect 4448 5370 4476 8910
rect 4632 8838 4660 9522
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 5460 8634 5488 9318
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4356 5222 4476 5250
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4356 4282 4384 4966
rect 4448 4758 4476 5222
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3896 3738 3924 3946
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 4264 3398 4292 4218
rect 4540 4010 4568 8298
rect 5552 8294 5580 11834
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 4632 6934 4660 8230
rect 5000 7410 5028 8230
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 5092 6730 5120 7686
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5276 7342 5304 7482
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5184 6458 5212 7278
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5778 4660 6054
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4540 3602 4568 3946
rect 4632 3602 4660 5238
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4622 4752 4966
rect 4816 4690 4844 5578
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4146 4752 4558
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3738 4844 4082
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5000 3738 5028 4014
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2976 2774 3004 3334
rect 5092 3194 5120 5102
rect 5448 4072 5500 4078
rect 5354 4040 5410 4049
rect 5448 4014 5500 4020
rect 5354 3975 5410 3984
rect 5368 3534 5396 3975
rect 5460 3738 5488 4014
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 2976 2746 3188 2774
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 3160 2446 3188 2746
rect 4448 2650 4476 2994
rect 5276 2650 5304 3402
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2332 2106 2360 2382
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 3344 1170 3372 2450
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3068 1142 3372 1170
rect 3068 800 3096 1142
rect 3896 800 3924 2314
rect 4908 1306 4936 2382
rect 4724 1278 4936 1306
rect 4724 800 4752 1278
rect 5552 800 5580 2926
rect 5644 2854 5672 11698
rect 5736 11218 5764 12174
rect 5828 11898 5856 18566
rect 6012 15910 6040 18686
rect 6472 18290 6500 19314
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6472 17202 6500 18226
rect 6840 17814 6868 18838
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 17882 6960 18226
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16794 6960 17138
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6012 15162 6040 15846
rect 6564 15706 6592 15846
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6104 15162 6132 15438
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6472 14618 6500 15574
rect 6748 15502 6776 15982
rect 6840 15570 6868 16390
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 7024 15502 7052 20538
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7300 16046 7328 20198
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7944 18970 7972 19246
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8588 18834 8616 19110
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7484 18426 7512 18634
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7760 18290 7788 18770
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7392 15638 7420 17750
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 16046 7512 16526
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7484 15706 7512 15982
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 6736 15496 6788 15502
rect 7012 15496 7064 15502
rect 6788 15444 6868 15450
rect 6736 15438 6868 15444
rect 7012 15438 7064 15444
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 6552 15428 6604 15434
rect 6748 15422 6868 15438
rect 6552 15370 6604 15376
rect 6564 15026 6592 15370
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 14618 6592 14758
rect 6748 14618 6776 14962
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5920 13462 5948 13806
rect 6380 13530 6408 13874
rect 6840 13734 6868 15422
rect 7024 14958 7052 15438
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7024 14414 7052 14894
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 7208 14074 7236 15438
rect 7392 15434 7420 15574
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7286 15056 7342 15065
rect 7286 14991 7342 15000
rect 7300 14958 7328 14991
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 14074 7328 14214
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13530 6868 13670
rect 7392 13530 7420 15370
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6472 12374 6500 12854
rect 6656 12850 6684 13126
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 6472 11830 6500 12310
rect 6656 12238 6684 12786
rect 6840 12434 6868 13466
rect 6748 12406 6868 12434
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11830 6684 12174
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10538 5764 11154
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5736 10130 5764 10474
rect 5828 10266 5856 11018
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 10266 5948 10406
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5828 9654 5856 10202
rect 6012 10130 6040 10542
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6380 9178 6408 11494
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6472 10198 6500 11222
rect 6656 11150 6684 11766
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10810 6684 11086
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9586 6592 10066
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 5370 5764 7142
rect 5920 6118 5948 8230
rect 6104 7342 6132 9114
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6380 7954 6408 8502
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7342 6224 7686
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5736 3534 5764 5034
rect 5828 4622 5856 5170
rect 5920 4706 5948 6054
rect 6104 5846 6132 7278
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6104 5574 6132 5782
rect 6196 5710 6224 7278
rect 6380 6798 6408 7414
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 5846 6316 6598
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6380 5234 6408 6122
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 5920 4678 6132 4706
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5920 4554 5948 4678
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5906 4176 5962 4185
rect 5828 4134 5906 4162
rect 5828 3670 5856 4134
rect 5906 4111 5962 4120
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5724 3528 5776 3534
rect 5776 3488 5856 3516
rect 5724 3470 5776 3476
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 3058 5764 3334
rect 5828 3126 5856 3488
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5920 2378 5948 3402
rect 6012 3058 6040 4558
rect 6104 4554 6132 4678
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6472 4298 6500 8774
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6564 4622 6592 6190
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6380 4270 6500 4298
rect 6380 4146 6408 4270
rect 6656 4214 6684 9318
rect 6748 5370 6776 12406
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6840 11830 6868 12106
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 7010 11792 7066 11801
rect 7010 11727 7012 11736
rect 7064 11727 7066 11736
rect 7012 11698 7064 11704
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10266 6868 11154
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7024 9178 7052 11698
rect 7392 11558 7420 13466
rect 7562 12336 7618 12345
rect 7562 12271 7564 12280
rect 7616 12271 7618 12280
rect 7564 12242 7616 12248
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7102 11112 7158 11121
rect 7102 11047 7104 11056
rect 7156 11047 7158 11056
rect 7104 11018 7156 11024
rect 7116 9178 7144 11018
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6840 8566 6868 8842
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 7024 7886 7052 9114
rect 7116 8498 7144 9114
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7116 6458 7144 7958
rect 7392 7478 7420 8910
rect 7576 8634 7604 9454
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 8974 7696 9318
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7760 8430 7788 18226
rect 7852 17746 7880 18566
rect 8772 18086 8800 20742
rect 9140 19718 9168 20862
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 9324 19990 9352 20810
rect 9968 20482 9996 22442
rect 10060 21690 10088 22510
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22098 10180 22374
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10152 21962 10180 22034
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10704 21690 10732 22510
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 10888 21894 10916 22374
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 9968 20454 10088 20482
rect 10060 20398 10088 20454
rect 10152 20398 10180 21490
rect 10888 21078 10916 21830
rect 10980 21554 11008 21830
rect 11072 21690 11100 22918
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 11164 21010 11192 22170
rect 11348 21962 11376 22374
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11992 21690 12020 22510
rect 12084 22234 12112 23054
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12176 22098 12204 22714
rect 14108 22710 14136 23054
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12164 22092 12216 22098
rect 12636 22094 12664 22374
rect 12164 22034 12216 22040
rect 12452 22066 12664 22094
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10336 20466 10364 20742
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19990 9444 20198
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 10060 19786 10088 20334
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9140 18290 9168 19654
rect 9692 18970 9720 19722
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9784 18290 9812 19110
rect 10152 18850 10180 20334
rect 11256 19990 11284 20946
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20602 11652 20878
rect 11808 20602 11836 20946
rect 12176 20890 12204 22034
rect 12452 21894 12480 22066
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12452 21146 12480 21830
rect 12820 21690 12848 21830
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 13648 21554 13676 22578
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13832 22234 13860 22374
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12084 20862 12204 20890
rect 12084 20806 12112 20862
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11796 20596 11848 20602
rect 13556 20584 13584 21286
rect 13648 20754 13676 21490
rect 14292 21078 14320 21830
rect 14384 21690 14412 22986
rect 14568 22710 14596 23462
rect 15108 23180 15160 23186
rect 15108 23122 15160 23128
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 15120 22030 15148 23122
rect 15212 22778 15240 23598
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15304 22574 15332 23598
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 17408 23520 17460 23526
rect 17408 23462 17460 23468
rect 15394 22876 15702 22885
rect 15394 22874 15400 22876
rect 15456 22874 15480 22876
rect 15536 22874 15560 22876
rect 15616 22874 15640 22876
rect 15696 22874 15702 22876
rect 15456 22822 15458 22874
rect 15638 22822 15640 22874
rect 15394 22820 15400 22822
rect 15456 22820 15480 22822
rect 15536 22820 15560 22822
rect 15616 22820 15640 22822
rect 15696 22820 15702 22822
rect 15394 22811 15702 22820
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15384 22094 15436 22098
rect 15488 22094 15516 22578
rect 16120 22568 16172 22574
rect 16120 22510 16172 22516
rect 15384 22092 15516 22094
rect 15436 22066 15516 22092
rect 15384 22034 15436 22040
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14568 21554 14596 21830
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 13912 20800 13964 20806
rect 13648 20726 13860 20754
rect 13912 20742 13964 20748
rect 13556 20556 13676 20584
rect 11796 20538 11848 20544
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11256 19718 11284 19926
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10244 18970 10272 19246
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10152 18822 10272 18850
rect 10244 18630 10272 18822
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8172 17980 8480 17989
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 17270 8432 17478
rect 8392 17264 8444 17270
rect 8444 17224 8616 17252
rect 8392 17206 8444 17212
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 8588 16794 8616 17224
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16114 8248 16458
rect 8772 16114 8800 18022
rect 9140 17746 9168 18226
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9600 16794 9628 17546
rect 9876 17338 9904 18022
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7852 15026 7880 15302
rect 7930 15056 7986 15065
rect 7840 15020 7892 15026
rect 7930 14991 7986 15000
rect 7840 14962 7892 14968
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10810 7880 10950
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7760 8090 7788 8366
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 6458 7328 7346
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6458 7696 6734
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6458 7788 6598
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7116 6254 7144 6394
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 7024 5234 7052 5510
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6644 4208 6696 4214
rect 6642 4176 6644 4185
rect 6696 4176 6698 4185
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6460 4140 6512 4146
rect 6642 4111 6698 4120
rect 6460 4082 6512 4088
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6104 3516 6132 4014
rect 6104 3488 6224 3516
rect 6196 3482 6224 3488
rect 6196 3466 6316 3482
rect 6196 3460 6328 3466
rect 6196 3454 6276 3460
rect 6276 3402 6328 3408
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5998 2952 6054 2961
rect 5998 2887 6000 2896
rect 6052 2887 6054 2896
rect 6000 2858 6052 2864
rect 6472 2514 6500 4082
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3058 6684 3946
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6748 2378 6776 4966
rect 7208 4622 7236 5510
rect 7576 4826 7604 5646
rect 7760 5030 7788 5646
rect 7748 5024 7800 5030
rect 7746 4992 7748 5001
rect 7800 4992 7802 5001
rect 7746 4927 7802 4936
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7944 4706 7972 14991
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 8680 14414 8708 15370
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 14074 8708 14350
rect 9140 14278 9168 15370
rect 9232 15162 9260 15574
rect 9508 15502 9536 15914
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9600 15609 9628 15846
rect 9586 15600 9642 15609
rect 9586 15535 9642 15544
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9600 15162 9628 15535
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 9140 13870 9168 14214
rect 9692 13938 9720 17274
rect 10244 17134 10272 18566
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10336 17134 10364 17274
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16658 9812 16934
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9876 14958 9904 15302
rect 10336 15094 10364 15846
rect 10428 15570 10456 18770
rect 10612 18426 10640 19246
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17338 10548 17478
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 9864 14952 9916 14958
rect 10428 14906 10456 15506
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 9864 14894 9916 14900
rect 9876 14618 9904 14894
rect 10244 14878 10456 14906
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9876 14074 9904 14554
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 9968 14074 9996 14282
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9692 13802 9720 13874
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11898 8248 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8172 9211 8480 9220
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8498 8064 8774
rect 8588 8566 8616 9318
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8680 8498 8708 10134
rect 8772 9654 8800 13194
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12322 8984 12582
rect 9048 12434 9076 13126
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9232 12753 9260 12854
rect 9218 12744 9274 12753
rect 9218 12679 9274 12688
rect 9048 12406 9168 12434
rect 8956 12294 9076 12322
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8956 11626 8984 12174
rect 9048 12050 9076 12294
rect 9140 12170 9168 12406
rect 9128 12164 9180 12170
rect 9128 12106 9180 12112
rect 9048 12022 9168 12050
rect 9140 11898 9168 12022
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8956 10674 8984 11562
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9048 10266 9076 10678
rect 9232 10266 9260 12679
rect 9692 12434 9720 13738
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9784 12442 9812 12786
rect 9508 12406 9720 12434
rect 9772 12436 9824 12442
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9508 10198 9536 12406
rect 9772 12378 9824 12384
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9600 11082 9628 11630
rect 10152 11257 10180 12854
rect 10138 11248 10194 11257
rect 10138 11183 10194 11192
rect 10152 11150 10180 11183
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8956 9178 8984 9454
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8036 8090 8064 8434
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8220 7546 8248 7822
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8312 7478 8340 7822
rect 8588 7818 8616 8366
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8588 7342 8616 7754
rect 8680 7478 8708 8434
rect 8864 8430 8892 9046
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9232 8634 9260 8842
rect 9508 8838 9536 10134
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 9232 7546 9260 8570
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 9048 6730 9076 7346
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 7002 9168 7278
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9232 6338 9260 7482
rect 9232 6310 9352 6338
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 8680 5302 8708 6054
rect 9232 5914 9260 6190
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9324 5778 9352 6310
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 8668 5296 8720 5302
rect 9324 5250 9352 5714
rect 9508 5574 9536 6054
rect 9600 5914 9628 11018
rect 10152 10810 10180 11086
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10244 10452 10272 14878
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 14074 10640 14214
rect 10704 14074 10732 15302
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12889 10456 13126
rect 10414 12880 10470 12889
rect 10414 12815 10416 12824
rect 10468 12815 10470 12824
rect 10416 12786 10468 12792
rect 10520 12646 10548 13806
rect 10704 13530 10732 14010
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10612 12442 10640 13262
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10704 11830 10732 13466
rect 10796 11830 10824 19654
rect 11256 19514 11284 19654
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11072 18850 11100 19314
rect 10888 18822 11100 18850
rect 10888 18698 10916 18822
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 18290 11008 18566
rect 11072 18426 11100 18634
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10980 17814 11008 18226
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11072 17882 11100 18090
rect 11256 17882 11284 18158
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 11348 17746 11376 18634
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 18290 11744 18566
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15706 10916 15982
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10888 14074 10916 14282
rect 11348 14074 11376 17682
rect 11808 17338 11836 20538
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18290 11928 19110
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11900 17746 11928 18226
rect 12084 18222 12112 19246
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 12176 17542 12204 18702
rect 12268 18154 12296 19654
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12636 18970 12664 19246
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13096 18970 13124 19110
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11808 16998 11836 17274
rect 12176 17066 12204 17478
rect 12452 17338 12480 17546
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 17270 12572 18158
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11808 16794 11836 16934
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 11624 14958 11652 15846
rect 12084 15502 12112 15846
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 10876 14068 10928 14074
rect 11336 14068 11388 14074
rect 10876 14010 10928 14016
rect 11164 14028 11336 14056
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12918 11100 13126
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12306 11008 12718
rect 11164 12434 11192 14028
rect 11336 14010 11388 14016
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11072 12406 11192 12434
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 10810 10548 11698
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10612 10606 10640 11494
rect 10704 11098 10732 11766
rect 10796 11218 10824 11766
rect 10980 11762 11008 12242
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 11072 11098 11100 12406
rect 11152 12300 11204 12306
rect 11348 12288 11376 13670
rect 11532 13530 11560 14554
rect 11624 13734 11652 14894
rect 11716 14822 11744 15438
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 12084 14482 12112 15438
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 12176 13530 12204 17002
rect 12728 16998 12756 18158
rect 13004 17202 13032 18566
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12360 15502 12388 15846
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12268 14278 12296 14894
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12452 14074 12480 15982
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12268 13802 12296 14010
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11532 12850 11560 13194
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11204 12260 11376 12288
rect 11152 12242 11204 12248
rect 11164 11354 11192 12242
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11440 11898 11468 12174
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10704 11082 10916 11098
rect 10704 11076 10928 11082
rect 10704 11070 10876 11076
rect 11072 11070 11192 11098
rect 10876 11018 10928 11024
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10674 11100 10950
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10508 10464 10560 10470
rect 10244 10424 10508 10452
rect 10508 10406 10560 10412
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 7886 9720 9454
rect 9784 8974 9812 10202
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10336 9654 10364 9862
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10060 9466 10088 9522
rect 10060 9438 10180 9466
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 10152 8838 10180 9438
rect 10520 9110 10548 10406
rect 10612 9382 10640 10542
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8498 10180 8774
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 8090 10364 8230
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9692 7410 9720 7822
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 6322 9720 7346
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6458 10180 6598
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5574 10088 5714
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 8668 5238 8720 5244
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 9232 5222 9352 5250
rect 7852 4678 7972 4706
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6932 2514 6960 4150
rect 7852 4146 7880 4678
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7208 2446 7236 3334
rect 7300 3194 7328 3470
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6380 800 6408 2042
rect 7392 1714 7420 3538
rect 7944 3194 7972 4558
rect 8036 4282 8064 5170
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8036 3126 8064 4218
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8588 3058 8616 4422
rect 8864 4282 8892 4626
rect 9232 4282 9260 5222
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9324 4554 9352 5034
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9324 4282 9352 4490
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9232 4146 9260 4218
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9508 4078 9536 5510
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9692 5030 9720 5102
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9784 4622 9812 5102
rect 10060 4758 10088 5510
rect 10244 5098 10272 7754
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7342 10364 7686
rect 10428 7546 10456 8366
rect 10612 8362 10640 9318
rect 10888 9178 10916 9998
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11164 9042 11192 11070
rect 11348 10130 11376 11494
rect 11532 10606 11560 12786
rect 11624 12306 11652 13126
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 12424 11744 12582
rect 11796 12436 11848 12442
rect 11716 12396 11796 12424
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11716 11898 11744 12396
rect 12084 12434 12112 13194
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11796 12378 11848 12384
rect 11992 12406 12112 12434
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 9178 11560 9318
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10600 8356 10652 8362
rect 10704 8344 10732 8774
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10704 8316 11100 8344
rect 10600 8298 10652 8304
rect 10612 7750 10640 8298
rect 11072 7886 11100 8316
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10704 7206 10732 7482
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10520 5234 10548 5510
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9692 3534 9720 4422
rect 9784 3738 9812 4558
rect 10244 4282 10272 4626
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4282 10456 4422
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 7470 2952 7526 2961
rect 7470 2887 7526 2896
rect 7484 2774 7512 2887
rect 9968 2774 9996 4082
rect 10612 4010 10640 4626
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10704 3942 10732 7142
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 5914 10824 6734
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5710 10916 6598
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10888 5030 10916 5646
rect 10980 5370 11008 5646
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11072 5166 11100 7822
rect 11164 5370 11192 8570
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 11072 4842 11100 5102
rect 10980 4814 11100 4842
rect 10980 4758 11008 4814
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10796 3738 10824 4422
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3942 10916 4014
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10980 3738 11008 3946
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 10980 3126 11008 3402
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 11164 2854 11192 3334
rect 11256 3058 11284 4422
rect 11348 3738 11376 8842
rect 11532 8430 11560 9114
rect 11624 9110 11652 11018
rect 11716 9674 11744 11834
rect 11808 11626 11836 12242
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11716 9646 11928 9674
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11624 8430 11652 8842
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11624 8090 11652 8366
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11900 7478 11928 9646
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 6866 11560 7142
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 6458 11468 6734
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11900 6322 11928 7414
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5574 11836 6054
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11900 5098 11928 6258
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4826 11560 4966
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11900 3670 11928 3878
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11992 3194 12020 12406
rect 12176 12322 12204 12718
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12084 12294 12204 12322
rect 12084 11286 12112 12294
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12176 11218 12204 12174
rect 12268 11898 12296 12378
rect 12636 12306 12664 15098
rect 13188 15094 13216 15846
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12728 14074 12756 14826
rect 13188 14074 13216 15030
rect 13648 14822 13676 20556
rect 13832 19922 13860 20726
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13832 19378 13860 19858
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13740 17746 13768 18090
rect 13832 17882 13860 18702
rect 13924 18426 13952 20742
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14108 18698 14136 20198
rect 14292 19718 14320 21014
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14384 19854 14412 20742
rect 14936 20398 14964 21830
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15028 20602 15056 20878
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14936 19446 14964 20334
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14384 18970 14412 19314
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14108 18086 14136 18634
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13740 15706 13768 15982
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 13280 14074 13308 14282
rect 13464 14074 13492 14758
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12912 12850 12940 13330
rect 12990 13288 13046 13297
rect 12990 13223 12992 13232
rect 13044 13223 13046 13232
rect 12992 13194 13044 13200
rect 13372 12918 13400 13466
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12345 12940 12786
rect 13372 12434 13400 12854
rect 13648 12850 13676 14758
rect 13924 13938 13952 14894
rect 14108 14482 14136 14894
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13726 13424 13782 13433
rect 13726 13359 13728 13368
rect 13780 13359 13782 13368
rect 13728 13330 13780 13336
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13280 12406 13400 12434
rect 12898 12336 12954 12345
rect 12624 12300 12676 12306
rect 12898 12271 12954 12280
rect 12624 12242 12676 12248
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10690 12204 11154
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12084 10662 12204 10690
rect 12084 10266 12112 10662
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12176 10266 12204 10542
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12268 7546 12296 11018
rect 12636 10810 12664 11086
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 9586 12664 10542
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12360 6798 12388 8774
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12544 7954 12572 8298
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12360 6118 12388 6734
rect 12728 6440 12756 12038
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13004 9722 13032 9930
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 13188 9586 13216 11018
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 8090 12940 8366
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12992 7812 13044 7818
rect 12992 7754 13044 7760
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7546 12940 7686
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13004 6905 13032 7754
rect 12990 6896 13046 6905
rect 12990 6831 13046 6840
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12820 6458 12848 6666
rect 12452 6412 12756 6440
rect 12808 6452 12860 6458
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12452 5114 12480 6412
rect 12808 6394 12860 6400
rect 12532 6316 12584 6322
rect 12584 6276 12848 6304
rect 12532 6258 12584 6264
rect 12820 6118 12848 6276
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12268 5086 12480 5114
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 3194 12112 3878
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 7484 2746 7696 2774
rect 7208 1686 7420 1714
rect 7208 800 7236 1686
rect 1398 0 1454 800
rect 2226 0 2282 800
rect 3054 0 3110 800
rect 3882 0 3938 800
rect 4710 0 4766 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7194 0 7250 800
rect 7668 762 7696 2746
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 9876 2746 9996 2774
rect 9772 2644 9824 2650
rect 9876 2632 9904 2746
rect 9824 2604 9904 2632
rect 9772 2586 9824 2592
rect 11164 2446 11192 2790
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 10416 2372 10468 2378
rect 10468 2332 10548 2360
rect 10416 2314 10468 2320
rect 7944 870 8064 898
rect 7944 762 7972 870
rect 8036 800 8064 870
rect 8864 800 8892 2314
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10520 800 10548 2332
rect 11348 800 11376 2858
rect 11808 2650 11836 2994
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 12176 800 12204 4014
rect 12268 3398 12296 5086
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 3670 12388 4966
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12452 3670 12480 4626
rect 12544 4486 12572 6054
rect 13004 5914 13032 6831
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 6458 13216 6598
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13280 6254 13308 12406
rect 13832 12102 13860 12718
rect 13924 12306 13952 13874
rect 14200 12434 14228 18022
rect 15120 17626 15148 21966
rect 15394 21788 15702 21797
rect 15394 21786 15400 21788
rect 15456 21786 15480 21788
rect 15536 21786 15560 21788
rect 15616 21786 15640 21788
rect 15696 21786 15702 21788
rect 15456 21734 15458 21786
rect 15638 21734 15640 21786
rect 15394 21732 15400 21734
rect 15456 21732 15480 21734
rect 15536 21732 15560 21734
rect 15616 21732 15640 21734
rect 15696 21732 15702 21734
rect 15394 21723 15702 21732
rect 16132 21690 16160 22510
rect 16224 22094 16252 23462
rect 17420 23118 17448 23462
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16304 22976 16356 22982
rect 16356 22936 16436 22964
rect 16304 22918 16356 22924
rect 16408 22234 16436 22936
rect 16776 22710 16804 22986
rect 17972 22778 18000 23054
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16580 22500 16632 22506
rect 16580 22442 16632 22448
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16304 22094 16356 22098
rect 16224 22092 16356 22094
rect 16224 22066 16304 22092
rect 16408 22094 16436 22170
rect 16488 22094 16540 22098
rect 16408 22092 16540 22094
rect 16408 22066 16488 22092
rect 16304 22034 16356 22040
rect 16488 22034 16540 22040
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15396 21010 15424 21286
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15212 19514 15240 20334
rect 15304 19990 15332 20878
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15394 20700 15702 20709
rect 15394 20698 15400 20700
rect 15456 20698 15480 20700
rect 15536 20698 15560 20700
rect 15616 20698 15640 20700
rect 15696 20698 15702 20700
rect 15456 20646 15458 20698
rect 15638 20646 15640 20698
rect 15394 20644 15400 20646
rect 15456 20644 15480 20646
rect 15536 20644 15560 20646
rect 15616 20644 15640 20646
rect 15696 20644 15702 20646
rect 15394 20635 15702 20644
rect 15856 20466 15884 20742
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15292 19984 15344 19990
rect 15292 19926 15344 19932
rect 15856 19922 15884 20402
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15394 19612 15702 19621
rect 15394 19610 15400 19612
rect 15456 19610 15480 19612
rect 15536 19610 15560 19612
rect 15616 19610 15640 19612
rect 15696 19610 15702 19612
rect 15456 19558 15458 19610
rect 15638 19558 15640 19610
rect 15394 19556 15400 19558
rect 15456 19556 15480 19558
rect 15536 19556 15560 19558
rect 15616 19556 15640 19558
rect 15696 19556 15702 19558
rect 15394 19547 15702 19556
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 16040 19378 16068 20334
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 18834 15332 19110
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15856 18630 15884 19246
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15028 17598 15148 17626
rect 15028 17134 15056 17598
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15028 16998 15056 17070
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16046 14320 16526
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15434 14320 15982
rect 14844 15706 14872 16050
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14292 15162 14320 15370
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14292 14618 14320 15098
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14292 13394 14320 14554
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14200 12406 14320 12434
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13372 11354 13400 11494
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13556 10606 13584 11494
rect 13924 11354 13952 12106
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 11082 14044 12038
rect 14108 11762 14136 12038
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14200 10606 14228 11222
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13556 10266 13584 10542
rect 14200 10470 14228 10542
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 8090 14136 9998
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13280 5574 13308 6190
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5642 13400 6054
rect 13464 5914 13492 7822
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7274 13860 7346
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13280 5234 13308 5510
rect 13832 5302 13860 7210
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13924 5778 13952 7142
rect 14016 6458 14044 7482
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14016 5574 14044 6394
rect 14108 6390 14136 7686
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14200 6458 14228 6598
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4282 12572 4422
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12544 3534 12572 4218
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12544 3058 12572 3470
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12912 2854 12940 5102
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 3534 13124 4422
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13280 3058 13308 4558
rect 13464 4282 13492 4966
rect 14016 4622 14044 5510
rect 14292 5250 14320 12406
rect 14384 11286 14412 13806
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14476 11830 14504 12718
rect 14568 12442 14596 15302
rect 15028 14958 15056 16934
rect 15120 16590 15148 17478
rect 15212 17218 15240 18566
rect 15394 18524 15702 18533
rect 15394 18522 15400 18524
rect 15456 18522 15480 18524
rect 15536 18522 15560 18524
rect 15616 18522 15640 18524
rect 15696 18522 15702 18524
rect 15456 18470 15458 18522
rect 15638 18470 15640 18522
rect 15394 18468 15400 18470
rect 15456 18468 15480 18470
rect 15536 18468 15560 18470
rect 15616 18468 15640 18470
rect 15696 18468 15702 18470
rect 15394 18459 15702 18468
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15304 17338 15332 17614
rect 15394 17436 15702 17445
rect 15394 17434 15400 17436
rect 15456 17434 15480 17436
rect 15536 17434 15560 17436
rect 15616 17434 15640 17436
rect 15696 17434 15702 17436
rect 15456 17382 15458 17434
rect 15638 17382 15640 17434
rect 15394 17380 15400 17382
rect 15456 17380 15480 17382
rect 15536 17380 15560 17382
rect 15616 17380 15640 17382
rect 15696 17380 15702 17382
rect 15394 17371 15702 17380
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15844 17264 15896 17270
rect 15212 17190 15332 17218
rect 15844 17206 15896 17212
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14844 14618 14872 14894
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13326 14964 14214
rect 15028 13530 15056 14894
rect 15212 14890 15240 16934
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15212 14006 15240 14826
rect 15304 14346 15332 17190
rect 15394 16348 15702 16357
rect 15394 16346 15400 16348
rect 15456 16346 15480 16348
rect 15536 16346 15560 16348
rect 15616 16346 15640 16348
rect 15696 16346 15702 16348
rect 15456 16294 15458 16346
rect 15638 16294 15640 16346
rect 15394 16292 15400 16294
rect 15456 16292 15480 16294
rect 15536 16292 15560 16294
rect 15616 16292 15640 16294
rect 15696 16292 15702 16294
rect 15394 16283 15702 16292
rect 15856 16046 15884 17206
rect 15948 16794 15976 17614
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15580 15366 15608 15982
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15706 15792 15846
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15856 15366 15884 15982
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15948 15706 15976 15914
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15394 15260 15702 15269
rect 15394 15258 15400 15260
rect 15456 15258 15480 15260
rect 15536 15258 15560 15260
rect 15616 15258 15640 15260
rect 15696 15258 15702 15260
rect 15456 15206 15458 15258
rect 15638 15206 15640 15258
rect 15394 15204 15400 15206
rect 15456 15204 15480 15206
rect 15536 15204 15560 15206
rect 15616 15204 15640 15206
rect 15696 15204 15702 15206
rect 15394 15195 15702 15204
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15304 13870 15332 14282
rect 15394 14172 15702 14181
rect 15394 14170 15400 14172
rect 15456 14170 15480 14172
rect 15536 14170 15560 14172
rect 15616 14170 15640 14172
rect 15696 14170 15702 14172
rect 15456 14118 15458 14170
rect 15638 14118 15640 14170
rect 15394 14116 15400 14118
rect 15456 14116 15480 14118
rect 15536 14116 15560 14118
rect 15616 14116 15640 14118
rect 15696 14116 15702 14118
rect 15394 14107 15702 14116
rect 15752 13932 15804 13938
rect 15856 13920 15884 15302
rect 16040 14958 16068 19314
rect 16132 16114 16160 21626
rect 16224 21350 16252 21966
rect 16592 21350 16620 22442
rect 17144 22166 17172 22714
rect 17960 22636 18012 22642
rect 17880 22596 17960 22624
rect 17880 22166 17908 22596
rect 17960 22578 18012 22584
rect 17132 22160 17184 22166
rect 17132 22102 17184 22108
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16684 21078 16712 22034
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16868 21146 16896 21830
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16224 19174 16252 19790
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16224 17678 16252 19110
rect 16408 18970 16436 20946
rect 16488 20800 16540 20806
rect 16486 20768 16488 20777
rect 16540 20768 16542 20777
rect 16486 20703 16542 20712
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16500 19854 16528 20198
rect 16684 19990 16712 21014
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16500 19514 16528 19790
rect 16960 19718 16988 20742
rect 17144 20398 17172 22102
rect 17684 22092 17736 22098
rect 18064 22094 18092 22918
rect 18156 22778 18184 23598
rect 18248 23322 18276 23598
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 46848 23520 46900 23526
rect 46848 23462 46900 23468
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18892 22778 18920 23462
rect 22616 23420 22924 23429
rect 22616 23418 22622 23420
rect 22678 23418 22702 23420
rect 22758 23418 22782 23420
rect 22838 23418 22862 23420
rect 22918 23418 22924 23420
rect 22678 23366 22680 23418
rect 22860 23366 22862 23418
rect 22616 23364 22622 23366
rect 22678 23364 22702 23366
rect 22758 23364 22782 23366
rect 22838 23364 22862 23366
rect 22918 23364 22924 23366
rect 22616 23355 22924 23364
rect 37060 23420 37368 23429
rect 37060 23418 37066 23420
rect 37122 23418 37146 23420
rect 37202 23418 37226 23420
rect 37282 23418 37306 23420
rect 37362 23418 37368 23420
rect 37122 23366 37124 23418
rect 37304 23366 37306 23418
rect 37060 23364 37066 23366
rect 37122 23364 37146 23366
rect 37202 23364 37226 23366
rect 37282 23364 37306 23366
rect 37362 23364 37368 23366
rect 37060 23355 37368 23364
rect 46860 23322 46888 23462
rect 42524 23316 42576 23322
rect 42524 23258 42576 23264
rect 46848 23316 46900 23322
rect 46848 23258 46900 23264
rect 20444 23248 20496 23254
rect 20444 23190 20496 23196
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19800 22976 19852 22982
rect 19800 22918 19852 22924
rect 18144 22772 18196 22778
rect 18144 22714 18196 22720
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18708 22094 18736 22510
rect 17684 22034 17736 22040
rect 17972 22066 18092 22094
rect 18616 22066 18736 22094
rect 17696 21350 17724 22034
rect 17972 21962 18000 22066
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 18616 21894 18644 22066
rect 18892 22030 18920 22714
rect 19260 22030 19288 22918
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19536 22094 19564 22510
rect 19444 22066 19564 22094
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17420 20602 17448 20742
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17132 20392 17184 20398
rect 17132 20334 17184 20340
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 17144 19446 17172 20334
rect 17420 19990 17448 20538
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17972 19786 18000 20878
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 17880 19666 17908 19722
rect 17880 19638 18000 19666
rect 17972 19514 18000 19638
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16408 18222 16436 18906
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16776 17882 16804 18770
rect 17144 18630 17172 19382
rect 18064 19378 18092 19790
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17972 18970 18000 19314
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18156 18834 18184 19110
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16960 17338 16988 17614
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 16316 16658 16344 17002
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16028 14952 16080 14958
rect 16080 14912 16252 14940
rect 16028 14894 16080 14900
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 14074 15976 14214
rect 16040 14074 16068 14350
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 15804 13892 15884 13920
rect 15752 13874 15804 13880
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 9382 14412 11086
rect 14476 10130 14504 11766
rect 14568 11694 14596 12378
rect 15028 11898 15056 12786
rect 15120 12374 15148 12786
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11898 15240 12038
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 15304 11354 15332 13670
rect 15394 13084 15702 13093
rect 15394 13082 15400 13084
rect 15456 13082 15480 13084
rect 15536 13082 15560 13084
rect 15616 13082 15640 13084
rect 15696 13082 15702 13084
rect 15456 13030 15458 13082
rect 15638 13030 15640 13082
rect 15394 13028 15400 13030
rect 15456 13028 15480 13030
rect 15536 13028 15560 13030
rect 15616 13028 15640 13030
rect 15696 13028 15702 13030
rect 15394 13019 15702 13028
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 12238 15608 12718
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15764 12102 15792 13874
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 12434 16068 13670
rect 15948 12406 16068 12434
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15394 11996 15702 12005
rect 15394 11994 15400 11996
rect 15456 11994 15480 11996
rect 15536 11994 15560 11996
rect 15616 11994 15640 11996
rect 15696 11994 15702 11996
rect 15456 11942 15458 11994
rect 15638 11942 15640 11994
rect 15394 11940 15400 11942
rect 15456 11940 15480 11942
rect 15536 11940 15560 11942
rect 15616 11940 15640 11942
rect 15696 11940 15702 11942
rect 15394 11931 15702 11940
rect 15856 11626 15884 12242
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10810 15056 10950
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14476 9586 14504 10066
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14568 7546 14596 10610
rect 15028 10266 15056 10746
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 7546 14780 7822
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14844 6798 14872 8026
rect 15120 7750 15148 8230
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14936 5914 14964 6734
rect 15028 6186 15056 7278
rect 15212 6662 15240 11086
rect 15394 10908 15702 10917
rect 15394 10906 15400 10908
rect 15456 10906 15480 10908
rect 15536 10906 15560 10908
rect 15616 10906 15640 10908
rect 15696 10906 15702 10908
rect 15456 10854 15458 10906
rect 15638 10854 15640 10906
rect 15394 10852 15400 10854
rect 15456 10852 15480 10854
rect 15536 10852 15560 10854
rect 15616 10852 15640 10854
rect 15696 10852 15702 10854
rect 15394 10843 15702 10852
rect 15948 10690 15976 12406
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11354 16068 11494
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15856 10662 15976 10690
rect 15856 10470 15884 10662
rect 16040 10606 16068 11290
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15304 9654 15332 10406
rect 15396 10062 15424 10406
rect 15948 10266 15976 10542
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15394 9820 15702 9829
rect 15394 9818 15400 9820
rect 15456 9818 15480 9820
rect 15536 9818 15560 9820
rect 15616 9818 15640 9820
rect 15696 9818 15702 9820
rect 15456 9766 15458 9818
rect 15638 9766 15640 9818
rect 15394 9764 15400 9766
rect 15456 9764 15480 9766
rect 15536 9764 15560 9766
rect 15616 9764 15640 9766
rect 15696 9764 15702 9766
rect 15394 9755 15702 9764
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15394 8732 15702 8741
rect 15394 8730 15400 8732
rect 15456 8730 15480 8732
rect 15536 8730 15560 8732
rect 15616 8730 15640 8732
rect 15696 8730 15702 8732
rect 15456 8678 15458 8730
rect 15638 8678 15640 8730
rect 15394 8676 15400 8678
rect 15456 8676 15480 8678
rect 15536 8676 15560 8678
rect 15616 8676 15640 8678
rect 15696 8676 15702 8678
rect 15394 8667 15702 8676
rect 15394 7644 15702 7653
rect 15394 7642 15400 7644
rect 15456 7642 15480 7644
rect 15536 7642 15560 7644
rect 15616 7642 15640 7644
rect 15696 7642 15702 7644
rect 15456 7590 15458 7642
rect 15638 7590 15640 7642
rect 15394 7588 15400 7590
rect 15456 7588 15480 7590
rect 15536 7588 15560 7590
rect 15616 7588 15640 7590
rect 15696 7588 15702 7590
rect 15394 7579 15702 7588
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15384 6928 15436 6934
rect 15382 6896 15384 6905
rect 15436 6896 15438 6905
rect 15672 6866 15700 7414
rect 15382 6831 15438 6840
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 15212 5914 15240 6598
rect 15394 6556 15702 6565
rect 15394 6554 15400 6556
rect 15456 6554 15480 6556
rect 15536 6554 15560 6556
rect 15616 6554 15640 6556
rect 15696 6554 15702 6556
rect 15456 6502 15458 6554
rect 15638 6502 15640 6554
rect 15394 6500 15400 6502
rect 15456 6500 15480 6502
rect 15536 6500 15560 6502
rect 15616 6500 15640 6502
rect 15696 6500 15702 6502
rect 15394 6491 15702 6500
rect 15764 6390 15792 9862
rect 15856 9382 15884 10066
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 6934 15884 9318
rect 16040 8906 16068 10406
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14292 5222 14412 5250
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4826 14136 4966
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13924 3738 13952 4558
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 14292 3534 14320 5102
rect 14384 3534 14412 5222
rect 14844 5166 14872 5646
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14568 3602 14596 4966
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3738 14780 3878
rect 14936 3738 14964 4014
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15028 3602 15056 4762
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13004 800 13032 2450
rect 13832 800 13860 2450
rect 14016 2446 14044 3334
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15212 2774 15240 2994
rect 15304 2774 15332 5646
rect 15394 5468 15702 5477
rect 15394 5466 15400 5468
rect 15456 5466 15480 5468
rect 15536 5466 15560 5468
rect 15616 5466 15640 5468
rect 15696 5466 15702 5468
rect 15456 5414 15458 5466
rect 15638 5414 15640 5466
rect 15394 5412 15400 5414
rect 15456 5412 15480 5414
rect 15536 5412 15560 5414
rect 15616 5412 15640 5414
rect 15696 5412 15702 5414
rect 15394 5403 15702 5412
rect 15394 4380 15702 4389
rect 15394 4378 15400 4380
rect 15456 4378 15480 4380
rect 15536 4378 15560 4380
rect 15616 4378 15640 4380
rect 15696 4378 15702 4380
rect 15456 4326 15458 4378
rect 15638 4326 15640 4378
rect 15394 4324 15400 4326
rect 15456 4324 15480 4326
rect 15536 4324 15560 4326
rect 15616 4324 15640 4326
rect 15696 4324 15702 4326
rect 15394 4315 15702 4324
rect 15764 4282 15792 6054
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15394 3292 15702 3301
rect 15394 3290 15400 3292
rect 15456 3290 15480 3292
rect 15536 3290 15560 3292
rect 15616 3290 15640 3292
rect 15696 3290 15702 3292
rect 15456 3238 15458 3290
rect 15638 3238 15640 3290
rect 15394 3236 15400 3238
rect 15456 3236 15480 3238
rect 15536 3236 15560 3238
rect 15616 3236 15640 3238
rect 15696 3236 15702 3238
rect 15394 3227 15702 3236
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15212 2746 15332 2774
rect 15212 2446 15240 2746
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 7668 734 7972 762
rect 8022 0 8078 800
rect 8850 0 8906 800
rect 9678 0 9734 800
rect 10506 0 10562 800
rect 11334 0 11390 800
rect 12162 0 12218 800
rect 12990 0 13046 800
rect 13818 0 13874 800
rect 14292 762 14320 2314
rect 14476 2106 14504 2382
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 15304 1170 15332 2450
rect 15396 2446 15424 3130
rect 15764 3058 15792 3470
rect 15856 3126 15884 4966
rect 15948 4146 15976 7210
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 16040 5234 16068 5510
rect 16132 5370 16160 14486
rect 16224 14074 16252 14912
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16224 13870 16252 14010
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16316 13462 16344 16594
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17052 16250 17080 16526
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15162 16436 15846
rect 16592 15706 16620 16186
rect 17144 16130 17172 18566
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17236 17202 17264 17478
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16658 17264 17138
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17052 16102 17172 16130
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16408 13870 16436 15098
rect 16776 14822 16804 15506
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14482 16804 14758
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16316 12986 16344 13398
rect 16408 12986 16436 13806
rect 16592 13530 16620 13942
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16684 13410 16712 14350
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16960 14006 16988 14214
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16500 13394 16712 13410
rect 16488 13388 16712 13394
rect 16540 13382 16712 13388
rect 16488 13330 16540 13336
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12306 16252 12582
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16224 9178 16252 9998
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16224 8838 16252 9114
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7206 16252 7686
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6798 16252 7142
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 5710 16252 6734
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 4690 16068 5170
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16132 4282 16160 5306
rect 16224 5166 16252 5646
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16224 4826 16252 5102
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16224 4146 16252 4762
rect 16316 4758 16344 12922
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16408 8566 16436 11562
rect 16500 11558 16528 12242
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16500 6186 16528 11018
rect 17052 10810 17080 16102
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17328 13394 17356 14350
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12782 17172 13262
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17144 12374 17172 12718
rect 17512 12442 17540 14350
rect 17604 13462 17632 16594
rect 17788 16590 17816 17478
rect 18064 17134 18092 17478
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17788 15570 17816 16526
rect 17880 15706 17908 16662
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 18064 15502 18092 17070
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9382 16620 9998
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 9178 16712 9318
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16500 5642 16528 6122
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16408 3398 16436 3878
rect 16500 3738 16528 5102
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3194 16436 3334
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15394 2204 15702 2213
rect 15394 2202 15400 2204
rect 15456 2202 15480 2204
rect 15536 2202 15560 2204
rect 15616 2202 15640 2204
rect 15696 2202 15702 2204
rect 15456 2150 15458 2202
rect 15638 2150 15640 2202
rect 15394 2148 15400 2150
rect 15456 2148 15480 2150
rect 15536 2148 15560 2150
rect 15616 2148 15640 2150
rect 15696 2148 15702 2150
rect 15394 2139 15702 2148
rect 15304 1142 15516 1170
rect 14568 870 14688 898
rect 14568 762 14596 870
rect 14660 800 14688 870
rect 15488 800 15516 1142
rect 16316 800 16344 2790
rect 16592 2582 16620 4490
rect 16684 3602 16712 5510
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16684 2514 16712 3402
rect 16776 3194 16804 10610
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16868 9042 16896 10542
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 6458 16896 8978
rect 17328 8022 17356 12038
rect 17880 11150 17908 15030
rect 17972 14498 18000 15302
rect 18064 15162 18092 15438
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17972 14470 18092 14498
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17972 12986 18000 14350
rect 18064 13938 18092 14470
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 18064 11082 18092 13738
rect 18156 13190 18184 16730
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18248 15434 18276 16594
rect 18340 16182 18368 16934
rect 18432 16590 18460 21286
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 19786 18644 20198
rect 18696 20052 18748 20058
rect 18800 20040 18828 21490
rect 19076 21350 19104 21830
rect 19260 21350 19288 21966
rect 19444 21894 19472 22066
rect 19812 21962 19840 22918
rect 20364 22778 20392 23054
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20456 22574 20484 23190
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 34060 23112 34112 23118
rect 34060 23054 34112 23060
rect 36452 23112 36504 23118
rect 36452 23054 36504 23060
rect 40408 23112 40460 23118
rect 40408 23054 40460 23060
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22204 22778 22232 22918
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18748 20012 18828 20040
rect 18696 19994 18748 20000
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18328 15360 18380 15366
rect 18432 15348 18460 16526
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18616 16250 18644 16458
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18380 15320 18460 15348
rect 18328 15302 18380 15308
rect 18340 13802 18368 15302
rect 18800 15094 18828 20012
rect 18892 19854 18920 20878
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18892 16794 18920 17070
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18788 15088 18840 15094
rect 18788 15030 18840 15036
rect 18892 14618 18920 15098
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 14074 18644 14214
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18248 12306 18276 13262
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10062 17724 10950
rect 18248 10810 18276 11086
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9654 17724 9998
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17420 8498 17448 8774
rect 17972 8634 18000 9522
rect 18064 9178 18092 9930
rect 18248 9722 18276 10746
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18340 9586 18368 13466
rect 18616 13394 18644 14010
rect 18892 13530 18920 14554
rect 19076 14482 19104 21286
rect 19260 20942 19288 21286
rect 20640 21026 20668 22578
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20732 22234 20760 22510
rect 20812 22500 20864 22506
rect 20812 22442 20864 22448
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20824 22030 20852 22442
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20824 21622 20852 21966
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 21100 21026 21128 21626
rect 20640 21010 20760 21026
rect 21100 21010 21312 21026
rect 20640 21004 20772 21010
rect 20640 20998 20720 21004
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20602 20208 20810
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 19174 19380 19246
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19168 18426 19196 18702
rect 19352 18698 19380 19110
rect 19720 18698 19748 19654
rect 20272 19514 20300 19790
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20548 18970 20576 19790
rect 20640 19394 20668 20998
rect 20720 20946 20772 20952
rect 21100 21004 21324 21010
rect 21100 20998 21272 21004
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20466 20760 20742
rect 21100 20602 21128 20998
rect 21272 20946 21324 20952
rect 21284 20874 21312 20946
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 21744 20058 21772 22034
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 22112 20534 22140 21354
rect 22204 21146 22232 21966
rect 22296 21146 22324 23054
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22388 22098 22416 22578
rect 22616 22332 22924 22341
rect 22616 22330 22622 22332
rect 22678 22330 22702 22332
rect 22758 22330 22782 22332
rect 22838 22330 22862 22332
rect 22918 22330 22924 22332
rect 22678 22278 22680 22330
rect 22860 22278 22862 22330
rect 22616 22276 22622 22278
rect 22678 22276 22702 22278
rect 22758 22276 22782 22278
rect 22838 22276 22862 22278
rect 22918 22276 22924 22278
rect 22616 22267 22924 22276
rect 22376 22092 22428 22098
rect 22560 22092 22612 22098
rect 22376 22034 22428 22040
rect 22480 22052 22560 22080
rect 22480 21978 22508 22052
rect 22560 22034 22612 22040
rect 23216 22030 23244 22918
rect 23584 22778 23612 23054
rect 33416 22976 33468 22982
rect 33416 22918 33468 22924
rect 29838 22876 30146 22885
rect 29838 22874 29844 22876
rect 29900 22874 29924 22876
rect 29980 22874 30004 22876
rect 30060 22874 30084 22876
rect 30140 22874 30146 22876
rect 29900 22822 29902 22874
rect 30082 22822 30084 22874
rect 29838 22820 29844 22822
rect 29900 22820 29924 22822
rect 29980 22820 30004 22822
rect 30060 22820 30084 22822
rect 30140 22820 30146 22822
rect 29838 22811 30146 22820
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 32036 22704 32088 22710
rect 32036 22646 32088 22652
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 26332 22568 26384 22574
rect 26332 22510 26384 22516
rect 27896 22568 27948 22574
rect 27896 22510 27948 22516
rect 29184 22568 29236 22574
rect 29184 22510 29236 22516
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31668 22568 31720 22574
rect 31668 22510 31720 22516
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 22388 21950 22508 21978
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 22388 21690 22416 21950
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 21100 19514 21128 19722
rect 22284 19712 22336 19718
rect 22388 19700 22416 21626
rect 22480 20602 22508 21830
rect 22616 21244 22924 21253
rect 22616 21242 22622 21244
rect 22678 21242 22702 21244
rect 22758 21242 22782 21244
rect 22838 21242 22862 21244
rect 22918 21242 22924 21244
rect 22678 21190 22680 21242
rect 22860 21190 22862 21242
rect 22616 21188 22622 21190
rect 22678 21188 22702 21190
rect 22758 21188 22782 21190
rect 22838 21188 22862 21190
rect 22918 21188 22924 21190
rect 22616 21179 22924 21188
rect 23124 20806 23152 21830
rect 23216 20942 23244 21966
rect 23308 21554 23336 22374
rect 23400 22234 23428 22510
rect 24860 22500 24912 22506
rect 24860 22442 24912 22448
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 24872 22098 24900 22442
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 24044 21350 24072 22034
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24964 21690 24992 21966
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25608 21622 25636 22374
rect 26344 22234 26372 22510
rect 26792 22500 26844 22506
rect 26792 22442 26844 22448
rect 26804 22234 26832 22442
rect 27712 22432 27764 22438
rect 27712 22374 27764 22380
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 26332 22228 26384 22234
rect 26332 22170 26384 22176
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26700 22024 26752 22030
rect 26700 21966 26752 21972
rect 26976 22024 27028 22030
rect 26976 21966 27028 21972
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24044 21146 24072 21286
rect 25332 21146 25360 21490
rect 26712 21418 26740 21966
rect 26700 21412 26752 21418
rect 26700 21354 26752 21360
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22480 19922 22508 20334
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22616 20156 22924 20165
rect 22616 20154 22622 20156
rect 22678 20154 22702 20156
rect 22758 20154 22782 20156
rect 22838 20154 22862 20156
rect 22918 20154 22924 20156
rect 22678 20102 22680 20154
rect 22860 20102 22862 20154
rect 22616 20100 22622 20102
rect 22678 20100 22702 20102
rect 22758 20100 22782 20102
rect 22838 20100 22862 20102
rect 22918 20100 22924 20102
rect 22616 20091 22924 20100
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22336 19672 22416 19700
rect 22284 19654 22336 19660
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20640 19378 20760 19394
rect 20628 19372 20760 19378
rect 20680 19366 20760 19372
rect 20628 19314 20680 19320
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19352 17338 19380 18634
rect 20732 18358 20760 19366
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20824 18426 20852 19246
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18426 21128 19110
rect 21192 18426 21220 19178
rect 21548 19168 21600 19174
rect 21468 19128 21548 19156
rect 21468 18970 21496 19128
rect 21548 19110 21600 19116
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 21088 18420 21140 18426
rect 21088 18362 21140 18368
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19720 17882 19748 18226
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 20732 17746 20760 18022
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 21008 17542 21036 18158
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19260 16794 19288 17138
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19260 15502 19288 15982
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19812 15162 19840 15370
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19996 15026 20024 16390
rect 20364 16182 20392 16934
rect 20548 16658 20576 17274
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20732 16046 20760 17478
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20824 16250 20852 16526
rect 20916 16250 20944 17070
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 15026 20668 15302
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18892 12782 18920 13330
rect 18984 12918 19012 13670
rect 19812 13394 19840 13806
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19800 13252 19852 13258
rect 19800 13194 19852 13200
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 19720 12442 19748 12786
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19352 10248 19380 12242
rect 19812 12102 19840 13194
rect 19996 12850 20024 13806
rect 20088 13734 20116 14826
rect 20732 14346 20760 15982
rect 21100 15706 21128 17002
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21192 16046 21220 16458
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 16250 21312 16390
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21192 15162 21220 15982
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21284 15366 21312 15642
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20364 13462 20392 13806
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20732 13462 20760 13670
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20720 13456 20772 13462
rect 20720 13398 20772 13404
rect 20824 13394 20852 13670
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11558 19840 12038
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19616 10532 19668 10538
rect 19616 10474 19668 10480
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19260 10220 19380 10248
rect 19260 9654 19288 10220
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9178 18184 9318
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18800 8838 18828 9454
rect 19444 9382 19472 10406
rect 19628 9926 19656 10474
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19536 9654 19564 9862
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19628 9042 19656 9862
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19812 8906 19840 11494
rect 19904 11354 19932 12106
rect 20732 11626 20760 13126
rect 20916 12306 20944 13874
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21008 12986 21036 13806
rect 21192 13530 21220 14554
rect 21284 13802 21312 14758
rect 21376 14618 21404 15438
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21284 12306 21312 13738
rect 21468 12646 21496 18906
rect 21928 18698 21956 19314
rect 22296 19242 22324 19654
rect 22480 19334 22508 19858
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22848 19352 22876 19654
rect 22940 19514 22968 19722
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22388 19306 22508 19334
rect 22836 19346 22888 19352
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 21732 18284 21784 18290
rect 21732 18226 21784 18232
rect 21744 17542 21772 18226
rect 21928 18154 21956 18634
rect 22008 18624 22060 18630
rect 22008 18566 22060 18572
rect 22020 18222 22048 18566
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17746 21864 18022
rect 22112 17762 22140 18294
rect 22204 17882 22232 18634
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 21824 17740 21876 17746
rect 22112 17734 22324 17762
rect 21824 17682 21876 17688
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21744 17066 21772 17478
rect 21732 17060 21784 17066
rect 21732 17002 21784 17008
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 21836 15434 21864 16934
rect 22204 16658 22232 16934
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21732 15360 21784 15366
rect 21652 15320 21732 15348
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 13410 21588 14282
rect 21652 13512 21680 15320
rect 21732 15302 21784 15308
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 13938 21864 14214
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21652 13484 21864 13512
rect 21560 13382 21772 13410
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21652 12306 21680 13262
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20824 11830 20852 12038
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20088 11354 20116 11494
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20536 10736 20588 10742
rect 20536 10678 20588 10684
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 10130 20024 10542
rect 20548 10266 20576 10678
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 18800 8634 18828 8774
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 6662 17080 7142
rect 17328 7002 17356 7278
rect 17512 7041 17540 7754
rect 17604 7546 17632 7822
rect 17972 7818 18000 8298
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17498 7032 17554 7041
rect 17316 6996 17368 7002
rect 18064 7002 18092 7346
rect 18800 7342 18828 8570
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19260 8090 19288 8366
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19352 7546 19380 8366
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 17498 6967 17554 6976
rect 18052 6996 18104 7002
rect 17316 6938 17368 6944
rect 18052 6938 18104 6944
rect 18984 6866 19012 7142
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17052 6458 17080 6598
rect 18156 6458 18184 6734
rect 19260 6458 19288 7278
rect 19444 6866 19472 8774
rect 19536 8566 19564 8774
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19536 7410 19564 8502
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19524 7404 19576 7410
rect 19576 7364 19656 7392
rect 19524 7346 19576 7352
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19628 6730 19656 7364
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17052 4622 17080 5850
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17144 4146 17172 5510
rect 17604 4826 17632 5646
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17696 5302 17724 5510
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17972 4486 18000 5102
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16868 3534 16896 3975
rect 16960 3738 16988 4082
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17512 3670 17540 3878
rect 17880 3670 17908 4014
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 17880 3058 17908 3606
rect 17972 3126 18000 4422
rect 18064 3194 18092 6190
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 16960 2650 16988 2994
rect 18156 2774 18184 6190
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18248 5370 18276 5714
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 5370 18368 5646
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18696 5092 18748 5098
rect 18696 5034 18748 5040
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18432 4282 18460 4558
rect 18708 4554 18736 5034
rect 18696 4548 18748 4554
rect 18696 4490 18748 4496
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18708 2990 18736 4490
rect 18800 3534 18828 6054
rect 19260 5914 19288 6190
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19076 5234 19104 5510
rect 19352 5234 19380 6054
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19076 4078 19104 5170
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19260 4146 19288 4422
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19352 3942 19380 5170
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19444 3534 19472 6054
rect 19536 4146 19564 6598
rect 19628 5302 19656 6666
rect 19720 5370 19748 7890
rect 19904 7886 19932 8026
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7342 19840 7686
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19812 7002 19840 7278
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19904 6662 19932 7822
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19812 5642 19840 6054
rect 19800 5636 19852 5642
rect 19800 5578 19852 5584
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19812 5166 19840 5578
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 19536 3738 19564 3975
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19720 3534 19748 4762
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19904 3534 19932 4422
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19996 3058 20024 10066
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20088 9178 20116 9998
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20364 8566 20392 8842
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20088 7954 20116 8434
rect 20168 8288 20220 8294
rect 20168 8230 20220 8236
rect 20180 7954 20208 8230
rect 20364 8022 20392 8502
rect 20824 8090 20852 11018
rect 21100 10674 21128 12174
rect 21744 11778 21772 13382
rect 21836 12434 21864 13484
rect 21928 12986 21956 15846
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22112 13802 22140 14418
rect 22204 13938 22232 16390
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22204 13190 22232 13874
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 12434 22140 12582
rect 21836 12406 22048 12434
rect 22112 12406 22232 12434
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 22020 12220 22048 12406
rect 22100 12232 22152 12238
rect 22020 12192 22100 12220
rect 21928 11898 21956 12174
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21744 11750 21864 11778
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21100 10266 21128 10610
rect 21836 10538 21864 11750
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 21928 11150 21956 11222
rect 22020 11218 22048 12192
rect 22100 12174 22152 12180
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21928 10606 21956 11086
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21284 9042 21312 9318
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 21284 7954 21312 8978
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 20180 7546 20208 7890
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20732 7206 20760 7822
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 7410 21496 7686
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20272 6458 20300 6802
rect 20732 6798 20760 7142
rect 21008 7002 21036 7346
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20180 4282 20208 5170
rect 20640 4826 20668 5714
rect 20732 5166 20760 6258
rect 21928 6254 21956 10542
rect 22020 10062 22048 10950
rect 22112 10606 22140 11562
rect 22100 10600 22152 10606
rect 22100 10542 22152 10548
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22112 8922 22140 10542
rect 22020 8894 22140 8922
rect 22020 7970 22048 8894
rect 22020 7942 22140 7970
rect 22112 6866 22140 7942
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 5914 22048 6054
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21284 5370 21312 5646
rect 22020 5522 22048 5850
rect 22204 5658 22232 12406
rect 22296 11354 22324 17734
rect 22388 17338 22416 19306
rect 22836 19288 22888 19294
rect 22468 19236 22520 19242
rect 22468 19178 22520 19184
rect 22480 18850 22508 19178
rect 22616 19068 22924 19077
rect 22616 19066 22622 19068
rect 22678 19066 22702 19068
rect 22758 19066 22782 19068
rect 22838 19066 22862 19068
rect 22918 19066 22924 19068
rect 22678 19014 22680 19066
rect 22860 19014 22862 19066
rect 22616 19012 22622 19014
rect 22678 19012 22702 19014
rect 22758 19012 22782 19014
rect 22838 19012 22862 19014
rect 22918 19012 22924 19014
rect 22616 19003 22924 19012
rect 22480 18822 22600 18850
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 18086 22508 18702
rect 22572 18222 22600 18822
rect 23032 18698 23060 20198
rect 23124 19922 23152 20742
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23216 19310 23244 19858
rect 23308 19514 23336 20538
rect 23400 20534 23428 20946
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25976 20602 26004 20810
rect 26988 20806 27016 21966
rect 27436 21888 27488 21894
rect 27436 21830 27488 21836
rect 27448 21729 27476 21830
rect 27434 21720 27490 21729
rect 27434 21655 27490 21664
rect 27436 21480 27488 21486
rect 27724 21468 27752 22374
rect 27816 21962 27844 22374
rect 27804 21956 27856 21962
rect 27804 21898 27856 21904
rect 27488 21440 27752 21468
rect 27436 21422 27488 21428
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23400 19990 23428 20470
rect 26436 20466 26464 20742
rect 26528 20466 26556 20742
rect 26988 20534 27016 20742
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23492 20058 23520 20334
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23860 19310 23888 19654
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22480 17882 22508 18022
rect 22616 17980 22924 17989
rect 22616 17978 22622 17980
rect 22678 17978 22702 17980
rect 22758 17978 22782 17980
rect 22838 17978 22862 17980
rect 22918 17978 22924 17980
rect 22678 17926 22680 17978
rect 22860 17926 22862 17978
rect 22616 17924 22622 17926
rect 22678 17924 22702 17926
rect 22758 17924 22782 17926
rect 22838 17924 22862 17926
rect 22918 17924 22924 17926
rect 22616 17915 22924 17924
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22376 17332 22428 17338
rect 22428 17292 22508 17320
rect 22376 17274 22428 17280
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22388 16794 22416 17070
rect 22480 16794 22508 17292
rect 22616 16892 22924 16901
rect 22616 16890 22622 16892
rect 22678 16890 22702 16892
rect 22758 16890 22782 16892
rect 22838 16890 22862 16892
rect 22918 16890 22924 16892
rect 22678 16838 22680 16890
rect 22860 16838 22862 16890
rect 22616 16836 22622 16838
rect 22678 16836 22702 16838
rect 22758 16836 22782 16838
rect 22838 16836 22862 16838
rect 22918 16836 22924 16838
rect 22616 16827 22924 16836
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22572 16454 22600 16662
rect 22848 16658 22876 16730
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 16250 22784 16390
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22756 16114 22784 16186
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22480 15910 22508 16050
rect 22940 16046 22968 16526
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 23032 15978 23060 18158
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 16250 23152 16390
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23020 15972 23072 15978
rect 23020 15914 23072 15920
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15366 22508 15846
rect 22616 15804 22924 15813
rect 22616 15802 22622 15804
rect 22678 15802 22702 15804
rect 22758 15802 22782 15804
rect 22838 15802 22862 15804
rect 22918 15802 22924 15804
rect 22678 15750 22680 15802
rect 22860 15750 22862 15802
rect 22616 15748 22622 15750
rect 22678 15748 22702 15750
rect 22758 15748 22782 15750
rect 22838 15748 22862 15750
rect 22918 15748 22924 15750
rect 22616 15739 22924 15748
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 15026 22692 15302
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22616 14716 22924 14725
rect 22616 14714 22622 14716
rect 22678 14714 22702 14716
rect 22758 14714 22782 14716
rect 22838 14714 22862 14716
rect 22918 14714 22924 14716
rect 22678 14662 22680 14714
rect 22860 14662 22862 14714
rect 22616 14660 22622 14662
rect 22678 14660 22702 14662
rect 22758 14660 22782 14662
rect 22838 14660 22862 14662
rect 22918 14660 22924 14662
rect 22616 14651 22924 14660
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22388 13530 22416 14350
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22480 13326 22508 13738
rect 23032 13734 23060 15914
rect 23124 15162 23152 15982
rect 23216 15910 23244 19246
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23400 17202 23428 18022
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17338 24440 17478
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 23308 15434 23336 16390
rect 24412 16046 24440 16934
rect 24504 16590 24532 19110
rect 24872 18290 24900 19246
rect 24964 18970 24992 19790
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25608 19514 25636 19654
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 26252 18970 26280 19790
rect 26528 19514 26556 19790
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26988 18766 27016 20470
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 25596 18760 25648 18766
rect 25596 18702 25648 18708
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 25056 18358 25084 18566
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24872 17882 24900 18226
rect 25608 17882 25636 18702
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26252 18290 26280 18566
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24596 16522 24624 17478
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24872 16794 24900 16934
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24964 16522 24992 17614
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24308 16040 24360 16046
rect 24308 15982 24360 15988
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24320 15706 24348 15982
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23492 14822 23520 15438
rect 24596 15366 24624 16458
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 22616 13628 22924 13637
rect 22616 13626 22622 13628
rect 22678 13626 22702 13628
rect 22758 13626 22782 13628
rect 22838 13626 22862 13628
rect 22918 13626 22924 13628
rect 22678 13574 22680 13626
rect 22860 13574 22862 13626
rect 22616 13572 22622 13574
rect 22678 13572 22702 13574
rect 22758 13572 22782 13574
rect 22838 13572 22862 13574
rect 22918 13572 22924 13574
rect 22616 13563 22924 13572
rect 23308 13569 23336 13670
rect 23294 13560 23350 13569
rect 23492 13530 23520 13806
rect 23294 13495 23296 13504
rect 23348 13495 23350 13504
rect 23480 13524 23532 13530
rect 23296 13466 23348 13472
rect 23480 13466 23532 13472
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12986 22968 13126
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 12442 22508 12786
rect 23308 12646 23336 13194
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 22616 12540 22924 12549
rect 22616 12538 22622 12540
rect 22678 12538 22702 12540
rect 22758 12538 22782 12540
rect 22838 12538 22862 12540
rect 22918 12538 22924 12540
rect 22678 12486 22680 12538
rect 22860 12486 22862 12538
rect 22616 12484 22622 12486
rect 22678 12484 22702 12486
rect 22758 12484 22782 12486
rect 22838 12484 22862 12486
rect 22918 12484 22924 12486
rect 22616 12475 22924 12484
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 23308 11694 23336 12582
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 22616 11452 22924 11461
rect 22616 11450 22622 11452
rect 22678 11450 22702 11452
rect 22758 11450 22782 11452
rect 22838 11450 22862 11452
rect 22918 11450 22924 11452
rect 22678 11398 22680 11450
rect 22860 11398 22862 11450
rect 22616 11396 22622 11398
rect 22678 11396 22702 11398
rect 22758 11396 22782 11398
rect 22838 11396 22862 11398
rect 22918 11396 22924 11398
rect 22616 11387 22924 11396
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22572 10470 22600 11086
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22616 10364 22924 10373
rect 22616 10362 22622 10364
rect 22678 10362 22702 10364
rect 22758 10362 22782 10364
rect 22838 10362 22862 10364
rect 22918 10362 22924 10364
rect 22678 10310 22680 10362
rect 22860 10310 22862 10362
rect 22616 10308 22622 10310
rect 22678 10308 22702 10310
rect 22758 10308 22782 10310
rect 22838 10308 22862 10310
rect 22918 10308 22924 10310
rect 22616 10299 22924 10308
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22296 9654 22324 9998
rect 23032 9994 23060 11494
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 23020 9988 23072 9994
rect 23020 9930 23072 9936
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 22616 9276 22924 9285
rect 22616 9274 22622 9276
rect 22678 9274 22702 9276
rect 22758 9274 22782 9276
rect 22838 9274 22862 9276
rect 22918 9274 22924 9276
rect 22678 9222 22680 9274
rect 22860 9222 22862 9274
rect 22616 9220 22622 9222
rect 22678 9220 22702 9222
rect 22758 9220 22782 9222
rect 22838 9220 22862 9222
rect 22918 9220 22924 9222
rect 22616 9211 22924 9220
rect 23032 9178 23060 9522
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22388 7954 22416 8298
rect 22480 8022 22508 8774
rect 22616 8188 22924 8197
rect 22616 8186 22622 8188
rect 22678 8186 22702 8188
rect 22758 8186 22782 8188
rect 22838 8186 22862 8188
rect 22918 8186 22924 8188
rect 22678 8134 22680 8186
rect 22860 8134 22862 8186
rect 22616 8132 22622 8134
rect 22678 8132 22702 8134
rect 22758 8132 22782 8134
rect 22838 8132 22862 8134
rect 22918 8132 22924 8134
rect 22616 8123 22924 8132
rect 22468 8016 22520 8022
rect 22468 7958 22520 7964
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22480 7410 22508 7958
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 23032 7546 23060 7822
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22480 6866 22508 7346
rect 22616 7100 22924 7109
rect 22616 7098 22622 7100
rect 22678 7098 22702 7100
rect 22758 7098 22782 7100
rect 22838 7098 22862 7100
rect 22918 7098 22924 7100
rect 22678 7046 22680 7098
rect 22860 7046 22862 7098
rect 22616 7044 22622 7046
rect 22678 7044 22702 7046
rect 22758 7044 22782 7046
rect 22838 7044 22862 7046
rect 22918 7044 22924 7046
rect 22616 7035 22924 7044
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22388 5778 22416 6054
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22204 5630 22324 5658
rect 22192 5568 22244 5574
rect 22020 5494 22140 5522
rect 22192 5510 22244 5516
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 22112 5166 22140 5494
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 21088 5160 21140 5166
rect 22100 5160 22152 5166
rect 21140 5120 21312 5148
rect 21088 5102 21140 5108
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20456 4282 20484 4558
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4282 20668 4422
rect 20916 4282 20944 4966
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20824 3466 20852 3878
rect 21192 3738 21220 4558
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20824 3194 20852 3402
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 21100 2990 21128 3334
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 17972 2746 18184 2774
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17144 2514 17356 2530
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 17144 2508 17368 2514
rect 17144 2502 17316 2508
rect 17144 800 17172 2502
rect 17316 2450 17368 2456
rect 17972 800 18000 2746
rect 18800 800 18828 2926
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18892 2650 18920 2790
rect 21192 2774 21220 3674
rect 21008 2746 21220 2774
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 21008 2446 21036 2746
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19628 800 19656 2042
rect 20456 800 20484 2314
rect 21284 800 21312 5120
rect 22100 5102 22152 5108
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21468 3194 21496 4558
rect 21560 4282 21588 4626
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21468 2650 21496 2994
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21652 2446 21680 4966
rect 22112 4622 22140 5102
rect 22204 4622 22232 5510
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22112 3942 22140 4558
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22204 3534 22232 4422
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22296 3194 22324 5630
rect 22388 5098 22416 5714
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22480 4978 22508 6666
rect 22940 6458 22968 6666
rect 22928 6452 22980 6458
rect 22928 6394 22980 6400
rect 22616 6012 22924 6021
rect 22616 6010 22622 6012
rect 22678 6010 22702 6012
rect 22758 6010 22782 6012
rect 22838 6010 22862 6012
rect 22918 6010 22924 6012
rect 22678 5958 22680 6010
rect 22860 5958 22862 6010
rect 22616 5956 22622 5958
rect 22678 5956 22702 5958
rect 22758 5956 22782 5958
rect 22838 5956 22862 5958
rect 22918 5956 22924 5958
rect 22616 5947 22924 5956
rect 22388 4950 22508 4978
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 21640 2440 21692 2446
rect 21640 2382 21692 2388
rect 22112 800 22140 2450
rect 22204 2446 22232 2858
rect 22388 2650 22416 4950
rect 22616 4924 22924 4933
rect 22616 4922 22622 4924
rect 22678 4922 22702 4924
rect 22758 4922 22782 4924
rect 22838 4922 22862 4924
rect 22918 4922 22924 4924
rect 22678 4870 22680 4922
rect 22860 4870 22862 4922
rect 22616 4868 22622 4870
rect 22678 4868 22702 4870
rect 22758 4868 22782 4870
rect 22838 4868 22862 4870
rect 22918 4868 22924 4870
rect 22616 4859 22924 4868
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 22480 3534 22508 3878
rect 22616 3836 22924 3845
rect 22616 3834 22622 3836
rect 22678 3834 22702 3836
rect 22758 3834 22782 3836
rect 22838 3834 22862 3836
rect 22918 3834 22924 3836
rect 22678 3782 22680 3834
rect 22860 3782 22862 3834
rect 22616 3780 22622 3782
rect 22678 3780 22702 3782
rect 22758 3780 22782 3782
rect 22838 3780 22862 3782
rect 22918 3780 22924 3782
rect 22616 3771 22924 3780
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 23032 3466 23060 3878
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23124 3194 23152 11018
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23216 8838 23244 9998
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23308 7886 23336 10474
rect 23492 9586 23520 10610
rect 23584 10538 23612 11630
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23492 6322 23520 7958
rect 23584 7478 23612 8230
rect 23676 7954 23704 8910
rect 23768 8430 23796 15302
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24228 14278 24256 14758
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24228 14006 24256 14214
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24044 12850 24072 13670
rect 24228 13394 24256 13942
rect 24412 13938 24440 14214
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24688 13530 24716 14350
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24504 12442 24532 13262
rect 24964 12986 24992 13330
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24136 10606 24164 11154
rect 24872 11150 24900 12718
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24044 10266 24072 10542
rect 24136 10266 24164 10542
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24228 9518 24256 11086
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24596 10266 24624 10406
rect 24688 10266 24716 10610
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 9178 23888 9318
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 24412 8974 24440 9454
rect 24872 8974 24900 9998
rect 25056 9466 25084 16934
rect 25332 16658 25360 17818
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25884 17338 25912 17478
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 26068 17202 26096 17614
rect 26160 17202 26188 18022
rect 26436 17542 26464 18566
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25332 16250 25360 16594
rect 26068 16590 26096 17138
rect 26056 16584 26108 16590
rect 26056 16526 26108 16532
rect 25964 16516 26016 16522
rect 25964 16458 26016 16464
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25332 14074 25360 14350
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 25148 13462 25176 13738
rect 25136 13456 25188 13462
rect 25136 13398 25188 13404
rect 25136 13184 25188 13190
rect 25136 13126 25188 13132
rect 25148 12986 25176 13126
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25148 12782 25176 12922
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25148 12306 25176 12582
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25424 11354 25452 11630
rect 25516 11626 25544 15846
rect 25976 15706 26004 16458
rect 26436 16250 26464 17478
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 26068 14482 26096 16050
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26344 15706 26372 15982
rect 26332 15700 26384 15706
rect 26332 15642 26384 15648
rect 26330 15600 26386 15609
rect 26528 15586 26556 18566
rect 27080 18290 27108 19654
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27172 18970 27200 19246
rect 27448 18970 27476 19654
rect 27528 19372 27580 19378
rect 27528 19314 27580 19320
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 27172 18222 27200 18634
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 26896 16454 26924 18158
rect 27540 17678 27568 19314
rect 27632 18850 27660 21286
rect 27724 19334 27752 21440
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27816 20874 27844 21422
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27816 20602 27844 20810
rect 27908 20602 27936 22510
rect 28172 22432 28224 22438
rect 28172 22374 28224 22380
rect 28632 22432 28684 22438
rect 28632 22374 28684 22380
rect 28184 22094 28212 22374
rect 28644 22094 28672 22374
rect 29196 22234 29224 22510
rect 30564 22432 30616 22438
rect 30564 22374 30616 22380
rect 31024 22432 31076 22438
rect 31024 22374 31076 22380
rect 29184 22228 29236 22234
rect 29184 22170 29236 22176
rect 30576 22166 30604 22374
rect 30564 22160 30616 22166
rect 30564 22102 30616 22108
rect 28184 22066 28396 22094
rect 27988 21956 28040 21962
rect 27988 21898 28040 21904
rect 28000 21690 28028 21898
rect 28078 21720 28134 21729
rect 27988 21684 28040 21690
rect 28078 21655 28134 21664
rect 27988 21626 28040 21632
rect 28000 21010 28028 21626
rect 28092 21486 28120 21655
rect 28080 21480 28132 21486
rect 28080 21422 28132 21428
rect 28368 21418 28396 22066
rect 28460 22066 28672 22094
rect 28460 21554 28488 22066
rect 29368 22024 29420 22030
rect 29368 21966 29420 21972
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28356 21412 28408 21418
rect 28356 21354 28408 21360
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 28276 20534 28304 21286
rect 28264 20528 28316 20534
rect 28264 20470 28316 20476
rect 27724 19306 28028 19334
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 27632 18822 27752 18850
rect 27724 18766 27752 18822
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27804 18624 27856 18630
rect 27804 18566 27856 18572
rect 27618 18184 27674 18193
rect 27618 18119 27620 18128
rect 27672 18119 27674 18128
rect 27620 18090 27672 18096
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26804 15706 26832 15846
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26386 15558 26556 15586
rect 26896 15570 26924 16390
rect 27264 16182 27292 16934
rect 27632 16794 27660 17070
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27724 16794 27752 16934
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27816 16522 27844 18566
rect 27908 17882 27936 19110
rect 28000 18426 28028 19306
rect 27988 18420 28040 18426
rect 27988 18362 28040 18368
rect 28172 18420 28224 18426
rect 28172 18362 28224 18368
rect 28184 18290 28212 18362
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28368 18222 28396 21354
rect 28460 20602 28488 21490
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28736 20602 28764 20810
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 29288 20466 29316 21286
rect 29380 21146 29408 21966
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 30656 21888 30708 21894
rect 30656 21830 30708 21836
rect 29472 21622 29500 21830
rect 29564 21690 29592 21830
rect 29838 21788 30146 21797
rect 29838 21786 29844 21788
rect 29900 21786 29924 21788
rect 29980 21786 30004 21788
rect 30060 21786 30084 21788
rect 30140 21786 30146 21788
rect 29900 21734 29902 21786
rect 30082 21734 30084 21786
rect 29838 21732 29844 21734
rect 29900 21732 29924 21734
rect 29980 21732 30004 21734
rect 30060 21732 30084 21734
rect 30140 21732 30146 21734
rect 29838 21723 30146 21732
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29460 21616 29512 21622
rect 29460 21558 29512 21564
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 30116 20942 30144 21422
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28460 20058 28488 20334
rect 28448 20052 28500 20058
rect 28448 19994 28500 20000
rect 29276 19236 29328 19242
rect 29276 19178 29328 19184
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28828 18358 28856 18566
rect 28816 18352 28868 18358
rect 28816 18294 28868 18300
rect 27988 18216 28040 18222
rect 28356 18216 28408 18222
rect 27988 18158 28040 18164
rect 28354 18184 28356 18193
rect 28408 18184 28410 18193
rect 27896 17876 27948 17882
rect 27896 17818 27948 17824
rect 27896 17604 27948 17610
rect 27896 17546 27948 17552
rect 27908 17066 27936 17546
rect 28000 17338 28028 18158
rect 28354 18119 28410 18128
rect 29000 18148 29052 18154
rect 29000 18090 29052 18096
rect 28172 18080 28224 18086
rect 28172 18022 28224 18028
rect 28184 17882 28212 18022
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 28172 17876 28224 17882
rect 28172 17818 28224 17824
rect 27988 17332 28040 17338
rect 27988 17274 28040 17280
rect 28092 17270 28120 17818
rect 29012 17542 29040 18090
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17270 29040 17478
rect 28080 17264 28132 17270
rect 28080 17206 28132 17212
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 27896 17060 27948 17066
rect 27896 17002 27948 17008
rect 27908 16794 27936 17002
rect 28092 16794 28120 17206
rect 28172 17128 28224 17134
rect 28172 17070 28224 17076
rect 27896 16788 27948 16794
rect 27896 16730 27948 16736
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 27804 16516 27856 16522
rect 27804 16458 27856 16464
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26330 15535 26386 15544
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25884 13326 25912 13806
rect 26068 13546 26096 14214
rect 26160 14074 26188 14282
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26238 13560 26294 13569
rect 26068 13530 26188 13546
rect 26056 13524 26188 13530
rect 26108 13518 26188 13524
rect 26056 13466 26108 13472
rect 26160 13394 26188 13518
rect 26238 13495 26294 13504
rect 26252 13444 26280 13495
rect 26332 13456 26384 13462
rect 26252 13416 26332 13444
rect 26332 13398 26384 13404
rect 26148 13388 26200 13394
rect 26148 13330 26200 13336
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 12434 25912 13262
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26160 12730 26188 12786
rect 26436 12782 26464 13670
rect 26424 12776 26476 12782
rect 26160 12702 26280 12730
rect 26424 12718 26476 12724
rect 26252 12442 26280 12702
rect 25700 12406 25912 12434
rect 26240 12436 26292 12442
rect 25504 11620 25556 11626
rect 25504 11562 25556 11568
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 24964 9438 25084 9466
rect 25148 9450 25176 10066
rect 25516 10062 25544 10950
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25136 9444 25188 9450
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7546 23980 7822
rect 24044 7546 24072 8366
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 24136 6866 24164 8026
rect 24688 8022 24716 8230
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24412 7410 24440 7686
rect 24688 7478 24716 7958
rect 24872 7954 24900 8774
rect 24964 8514 24992 9438
rect 25136 9386 25188 9392
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 9178 25084 9318
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25148 8566 25176 9386
rect 25240 8634 25268 9658
rect 25516 9654 25544 9998
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25504 9512 25556 9518
rect 25608 9500 25636 11086
rect 25700 10674 25728 12406
rect 26240 12378 26292 12384
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26068 10674 26096 11494
rect 26160 11218 26188 11494
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 25700 10130 25728 10610
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 25556 9472 25636 9500
rect 25504 9454 25556 9460
rect 25516 8838 25544 9454
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25136 8560 25188 8566
rect 24964 8486 25084 8514
rect 25136 8502 25188 8508
rect 24860 7948 24912 7954
rect 24912 7908 24992 7936
rect 24860 7890 24912 7896
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 23940 6656 23992 6662
rect 23860 6604 23940 6610
rect 23860 6598 23992 6604
rect 23860 6582 23980 6598
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5302 23704 6054
rect 23860 5370 23888 6582
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 23952 5370 23980 6190
rect 24136 5914 24164 6802
rect 24412 6662 24440 7346
rect 24872 7002 24900 7754
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24964 6934 24992 7908
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24124 5908 24176 5914
rect 24412 5896 24440 6598
rect 24124 5850 24176 5856
rect 24320 5868 24440 5896
rect 24320 5642 24348 5868
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24216 5636 24268 5642
rect 24216 5578 24268 5584
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23768 4554 23796 4966
rect 23860 4826 23888 5306
rect 24228 4826 24256 5578
rect 24320 5370 24348 5578
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 24412 5370 24440 5510
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 23756 4548 23808 4554
rect 23756 4490 23808 4496
rect 24320 4282 24348 5306
rect 24412 4690 24440 5306
rect 24872 4758 24900 5510
rect 24964 5166 24992 5646
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 23492 3738 23520 4014
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 24872 3466 24900 3878
rect 24860 3460 24912 3466
rect 24860 3402 24912 3408
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 25056 3058 25084 8486
rect 25148 6730 25176 8502
rect 25240 7886 25268 8570
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25424 7954 25452 8230
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25516 6866 25544 8774
rect 25700 8106 25728 10066
rect 26160 9926 26188 11154
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26344 10606 26372 10950
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26436 10538 26464 11086
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26528 10130 26556 15558
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26620 10062 26648 13126
rect 26712 12918 26740 13806
rect 26804 13530 26832 13806
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 26988 12306 27016 12582
rect 26976 12300 27028 12306
rect 26976 12242 27028 12248
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26160 8974 26188 9862
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 25608 8078 25728 8106
rect 25608 7410 25636 8078
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25884 7546 25912 7686
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25884 7410 25912 7482
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 3738 25176 4626
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25240 3194 25268 4014
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 22616 2748 22924 2757
rect 22616 2746 22622 2748
rect 22678 2746 22702 2748
rect 22758 2746 22782 2748
rect 22838 2746 22862 2748
rect 22918 2746 22924 2748
rect 22678 2694 22680 2746
rect 22860 2694 22862 2746
rect 22616 2692 22622 2694
rect 22678 2692 22702 2694
rect 22758 2692 22782 2694
rect 22838 2692 22862 2694
rect 22918 2692 22924 2694
rect 22616 2683 22924 2692
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 23768 2446 23796 2790
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 14292 734 14596 762
rect 14646 0 14702 800
rect 15474 0 15530 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18786 0 18842 800
rect 19614 0 19670 800
rect 20442 0 20498 800
rect 21270 0 21326 800
rect 22098 0 22154 800
rect 22664 762 22692 2314
rect 22848 870 22968 898
rect 22848 762 22876 870
rect 22940 800 22968 870
rect 23768 870 23888 898
rect 23768 800 23796 870
rect 22664 734 22876 762
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 23860 762 23888 870
rect 24044 762 24072 2926
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 24596 800 24624 2858
rect 25332 2774 25360 6666
rect 25608 6458 25636 7346
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25700 7002 25728 7278
rect 26056 7268 26108 7274
rect 26056 7210 26108 7216
rect 25688 6996 25740 7002
rect 25688 6938 25740 6944
rect 26068 6798 26096 7210
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26160 6458 26188 8910
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 25608 4622 25636 6394
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 26160 5914 26188 6122
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25884 5370 25912 5646
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25596 4616 25648 4622
rect 25596 4558 25648 4564
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3534 25544 3878
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25608 3466 25636 4558
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 26068 3194 26096 3878
rect 26252 3194 26280 9862
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26528 9178 26556 9522
rect 26712 9518 26740 10406
rect 27080 9654 27108 16050
rect 28092 16046 28120 16730
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 28184 15910 28212 17070
rect 28724 16584 28776 16590
rect 28724 16526 28776 16532
rect 28540 16040 28592 16046
rect 28540 15982 28592 15988
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27264 14074 27292 14282
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27448 14074 27476 14214
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27264 13394 27292 14010
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27264 11286 27292 13330
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27344 13184 27396 13190
rect 27344 13126 27396 13132
rect 27356 12850 27384 13126
rect 27448 12850 27476 13262
rect 27540 13258 27568 13806
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27540 12442 27568 12718
rect 27804 12708 27856 12714
rect 27804 12650 27856 12656
rect 27528 12436 27580 12442
rect 27528 12378 27580 12384
rect 27816 12238 27844 12650
rect 28184 12434 28212 15846
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28276 15026 28304 15302
rect 28552 15026 28580 15982
rect 28736 15706 28764 16526
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28920 15706 28948 15846
rect 29288 15706 29316 19178
rect 29552 19168 29604 19174
rect 29552 19110 29604 19116
rect 29564 18766 29592 19110
rect 29656 18834 29684 20878
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 29838 20700 30146 20709
rect 29838 20698 29844 20700
rect 29900 20698 29924 20700
rect 29980 20698 30004 20700
rect 30060 20698 30084 20700
rect 30140 20698 30146 20700
rect 29900 20646 29902 20698
rect 30082 20646 30084 20698
rect 29838 20644 29844 20646
rect 29900 20644 29924 20646
rect 29980 20644 30004 20646
rect 30060 20644 30084 20646
rect 30140 20644 30146 20646
rect 29838 20635 30146 20644
rect 30576 20602 30604 20810
rect 30564 20596 30616 20602
rect 30564 20538 30616 20544
rect 30668 20466 30696 21830
rect 31036 21622 31064 22374
rect 31588 22234 31616 22510
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31484 21888 31536 21894
rect 31484 21830 31536 21836
rect 31496 21622 31524 21830
rect 31024 21616 31076 21622
rect 31024 21558 31076 21564
rect 31484 21616 31536 21622
rect 31484 21558 31536 21564
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29644 18828 29696 18834
rect 29644 18770 29696 18776
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29644 18692 29696 18698
rect 29644 18634 29696 18640
rect 29656 18426 29684 18634
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29748 18340 29776 19654
rect 29838 19612 30146 19621
rect 29838 19610 29844 19612
rect 29900 19610 29924 19612
rect 29980 19610 30004 19612
rect 30060 19610 30084 19612
rect 30140 19610 30146 19612
rect 29900 19558 29902 19610
rect 30082 19558 30084 19610
rect 29838 19556 29844 19558
rect 29900 19556 29924 19558
rect 29980 19556 30004 19558
rect 30060 19556 30084 19558
rect 30140 19556 30146 19558
rect 29838 19547 30146 19556
rect 30668 19514 30696 19790
rect 30840 19712 30892 19718
rect 30840 19654 30892 19660
rect 30852 19514 30880 19654
rect 30656 19508 30708 19514
rect 30656 19450 30708 19456
rect 30840 19508 30892 19514
rect 30840 19450 30892 19456
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 31300 19304 31352 19310
rect 31300 19246 31352 19252
rect 29838 18524 30146 18533
rect 29838 18522 29844 18524
rect 29900 18522 29924 18524
rect 29980 18522 30004 18524
rect 30060 18522 30084 18524
rect 30140 18522 30146 18524
rect 29900 18470 29902 18522
rect 30082 18470 30084 18522
rect 29838 18468 29844 18470
rect 29900 18468 29924 18470
rect 29980 18468 30004 18470
rect 30060 18468 30084 18470
rect 30140 18468 30146 18470
rect 29838 18459 30146 18468
rect 30208 18426 30236 19246
rect 31312 18970 31340 19246
rect 31300 18964 31352 18970
rect 31300 18906 31352 18912
rect 31404 18737 31432 19790
rect 31496 19378 31524 21558
rect 31484 19372 31536 19378
rect 31484 19314 31536 19320
rect 31588 19334 31616 21966
rect 31680 21690 31708 22510
rect 32048 22098 32076 22646
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33048 22432 33100 22438
rect 33048 22374 33100 22380
rect 32036 22092 32088 22098
rect 32036 22034 32088 22040
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32220 21956 32272 21962
rect 32220 21898 32272 21904
rect 31668 21684 31720 21690
rect 31668 21626 31720 21632
rect 32232 21457 32260 21898
rect 32218 21448 32274 21457
rect 32218 21383 32274 21392
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31864 21146 31892 21286
rect 32232 21146 32260 21383
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 32220 21140 32272 21146
rect 32220 21082 32272 21088
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31390 18728 31446 18737
rect 31390 18663 31446 18672
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 29828 18352 29880 18358
rect 29748 18312 29828 18340
rect 29828 18294 29880 18300
rect 30392 17542 30420 18566
rect 31404 18154 31432 18663
rect 31496 18222 31524 19314
rect 31588 19306 31708 19334
rect 31484 18216 31536 18222
rect 31484 18158 31536 18164
rect 31576 18216 31628 18222
rect 31576 18158 31628 18164
rect 31392 18148 31444 18154
rect 31392 18090 31444 18096
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 29838 17436 30146 17445
rect 29838 17434 29844 17436
rect 29900 17434 29924 17436
rect 29980 17434 30004 17436
rect 30060 17434 30084 17436
rect 30140 17434 30146 17436
rect 29900 17382 29902 17434
rect 30082 17382 30084 17434
rect 29838 17380 29844 17382
rect 29900 17380 29924 17382
rect 29980 17380 30004 17382
rect 30060 17380 30084 17382
rect 30140 17380 30146 17382
rect 29838 17371 30146 17380
rect 30392 16794 30420 17478
rect 31588 17338 31616 18158
rect 31576 17332 31628 17338
rect 31576 17274 31628 17280
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 29460 16516 29512 16522
rect 29460 16458 29512 16464
rect 29552 16516 29604 16522
rect 29552 16458 29604 16464
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29380 16250 29408 16390
rect 29368 16244 29420 16250
rect 29368 16186 29420 16192
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28552 14618 28580 14962
rect 28920 14618 28948 15642
rect 29472 15434 29500 16458
rect 29564 15638 29592 16458
rect 29838 16348 30146 16357
rect 29838 16346 29844 16348
rect 29900 16346 29924 16348
rect 29980 16346 30004 16348
rect 30060 16346 30084 16348
rect 30140 16346 30146 16348
rect 29900 16294 29902 16346
rect 30082 16294 30084 16346
rect 29838 16292 29844 16294
rect 29900 16292 29924 16294
rect 29980 16292 30004 16294
rect 30060 16292 30084 16294
rect 30140 16292 30146 16294
rect 29838 16283 30146 16292
rect 30208 16250 30236 16526
rect 30392 16250 30420 16730
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 31392 16448 31444 16454
rect 31392 16390 31444 16396
rect 31484 16448 31536 16454
rect 31484 16390 31536 16396
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30392 15706 30420 16186
rect 31312 16114 31340 16390
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 30472 15904 30524 15910
rect 30472 15846 30524 15852
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 29552 15632 29604 15638
rect 29552 15574 29604 15580
rect 30484 15502 30512 15846
rect 31404 15502 31432 16390
rect 31496 16250 31524 16390
rect 31484 16244 31536 16250
rect 31484 16186 31536 16192
rect 31588 15910 31616 17274
rect 31680 17202 31708 19306
rect 31772 19242 31800 19654
rect 31760 19236 31812 19242
rect 31760 19178 31812 19184
rect 31864 18902 31892 21082
rect 32600 21010 32628 21966
rect 33060 21894 33088 22374
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 33060 21554 33088 21830
rect 33336 21706 33364 22510
rect 33428 21962 33456 22918
rect 33784 22636 33836 22642
rect 33784 22578 33836 22584
rect 33416 21956 33468 21962
rect 33416 21898 33468 21904
rect 33336 21690 33640 21706
rect 33324 21684 33640 21690
rect 33376 21678 33640 21684
rect 33324 21626 33376 21632
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 32770 21448 32826 21457
rect 32968 21434 32996 21490
rect 33612 21486 33640 21678
rect 33796 21554 33824 22578
rect 33968 22568 34020 22574
rect 33968 22510 34020 22516
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 32826 21406 32996 21434
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33324 21412 33376 21418
rect 32770 21383 32826 21392
rect 33324 21354 33376 21360
rect 33336 21146 33364 21354
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33784 21344 33836 21350
rect 33784 21286 33836 21292
rect 33324 21140 33376 21146
rect 33324 21082 33376 21088
rect 32588 21004 32640 21010
rect 32588 20946 32640 20952
rect 32312 19712 32364 19718
rect 32312 19654 32364 19660
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31852 18896 31904 18902
rect 31852 18838 31904 18844
rect 31760 18692 31812 18698
rect 31760 18634 31812 18640
rect 31772 17338 31800 18634
rect 31760 17332 31812 17338
rect 31760 17274 31812 17280
rect 31668 17196 31720 17202
rect 31668 17138 31720 17144
rect 31576 15904 31628 15910
rect 31576 15846 31628 15852
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 31300 15496 31352 15502
rect 31300 15438 31352 15444
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31576 15496 31628 15502
rect 31576 15438 31628 15444
rect 29460 15428 29512 15434
rect 29460 15370 29512 15376
rect 29092 15360 29144 15366
rect 29092 15302 29144 15308
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29104 15162 29132 15302
rect 29092 15156 29144 15162
rect 29092 15098 29144 15104
rect 29184 15088 29236 15094
rect 29184 15030 29236 15036
rect 28540 14612 28592 14618
rect 28540 14554 28592 14560
rect 28908 14612 28960 14618
rect 28908 14554 28960 14560
rect 28816 13728 28868 13734
rect 28816 13670 28868 13676
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28552 12986 28580 13262
rect 28644 12986 28672 13262
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28632 12980 28684 12986
rect 28632 12922 28684 12928
rect 28828 12918 28856 13670
rect 28816 12912 28868 12918
rect 28816 12854 28868 12860
rect 28184 12406 28304 12434
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 28172 11552 28224 11558
rect 28172 11494 28224 11500
rect 27252 11280 27304 11286
rect 27252 11222 27304 11228
rect 27436 10124 27488 10130
rect 27436 10066 27488 10072
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 26712 8838 26740 9454
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26712 8498 26740 8774
rect 26700 8492 26752 8498
rect 26700 8434 26752 8440
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26436 7410 26464 7890
rect 26712 7750 26740 8434
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26344 6322 26372 6598
rect 26436 6458 26464 7346
rect 26712 7002 26740 7686
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 26896 6458 26924 8366
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 26976 6724 27028 6730
rect 26976 6666 27028 6672
rect 26988 6458 27016 6666
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 27080 6322 27108 7278
rect 26332 6316 26384 6322
rect 26332 6258 26384 6264
rect 27068 6316 27120 6322
rect 27068 6258 27120 6264
rect 26344 5778 26372 6258
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26896 5370 26924 5510
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 26700 4072 26752 4078
rect 26700 4014 26752 4020
rect 26620 3398 26648 4014
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26240 3188 26292 3194
rect 26240 3130 26292 3136
rect 25056 2746 25360 2774
rect 25056 2650 25084 2746
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 26620 2446 26648 3334
rect 26712 2990 26740 4014
rect 26804 3534 26832 4422
rect 27172 4026 27200 9522
rect 27252 7268 27304 7274
rect 27252 7210 27304 7216
rect 27264 5370 27292 7210
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27356 4826 27384 5170
rect 27448 5166 27476 10066
rect 28184 9926 28212 11494
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 28184 9674 28212 9862
rect 28092 9646 28212 9674
rect 28092 9518 28120 9646
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 28092 9178 28120 9454
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27540 7342 27568 7958
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27632 6322 27660 7142
rect 28276 6882 28304 12406
rect 28540 12096 28592 12102
rect 28540 12038 28592 12044
rect 29000 12096 29052 12102
rect 29000 12038 29052 12044
rect 28552 11898 28580 12038
rect 29012 11898 29040 12038
rect 28540 11892 28592 11898
rect 28540 11834 28592 11840
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 28448 9988 28500 9994
rect 28448 9930 28500 9936
rect 28460 8634 28488 9930
rect 28552 9654 28580 11018
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 28540 9648 28592 9654
rect 28540 9590 28592 9596
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28644 8634 28672 8774
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28920 8362 28948 8978
rect 29012 8906 29040 10542
rect 29104 10470 29132 11086
rect 29196 10588 29224 15030
rect 29288 13938 29316 15302
rect 29472 15094 29500 15370
rect 29838 15260 30146 15269
rect 29838 15258 29844 15260
rect 29900 15258 29924 15260
rect 29980 15258 30004 15260
rect 30060 15258 30084 15260
rect 30140 15258 30146 15260
rect 29900 15206 29902 15258
rect 30082 15206 30084 15258
rect 29838 15204 29844 15206
rect 29900 15204 29924 15206
rect 29980 15204 30004 15206
rect 30060 15204 30084 15206
rect 30140 15204 30146 15206
rect 29838 15195 30146 15204
rect 29460 15088 29512 15094
rect 29460 15030 29512 15036
rect 31312 14958 31340 15438
rect 31588 15026 31616 15438
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 31300 14952 31352 14958
rect 31300 14894 31352 14900
rect 31024 14544 31076 14550
rect 31024 14486 31076 14492
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29656 13938 29684 14214
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29288 12102 29316 13874
rect 29460 13864 29512 13870
rect 29460 13806 29512 13812
rect 29472 13530 29500 13806
rect 29460 13524 29512 13530
rect 29460 13466 29512 13472
rect 29552 13252 29604 13258
rect 29552 13194 29604 13200
rect 29276 12096 29328 12102
rect 29276 12038 29328 12044
rect 29276 10600 29328 10606
rect 29196 10560 29276 10588
rect 29276 10542 29328 10548
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29092 10464 29144 10470
rect 29092 10406 29144 10412
rect 29368 9920 29420 9926
rect 29368 9862 29420 9868
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29104 8634 29132 8774
rect 29092 8628 29144 8634
rect 29092 8570 29144 8576
rect 29380 8498 29408 9862
rect 29472 9722 29500 10542
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 28908 8356 28960 8362
rect 28908 8298 28960 8304
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 29368 7336 29420 7342
rect 29368 7278 29420 7284
rect 27896 6860 27948 6866
rect 27896 6802 27948 6808
rect 28184 6854 28304 6882
rect 27908 6458 27936 6802
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27908 5914 27936 6394
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 27908 5370 27936 5850
rect 27896 5364 27948 5370
rect 27896 5306 27948 5312
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27436 5160 27488 5166
rect 27436 5102 27488 5108
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 27540 4690 27568 5170
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27540 4570 27568 4626
rect 27448 4542 27568 4570
rect 27448 4078 27476 4542
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27540 4282 27568 4422
rect 27632 4282 27660 4966
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 27724 4282 27752 4558
rect 27528 4276 27580 4282
rect 27528 4218 27580 4224
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27712 4276 27764 4282
rect 27712 4218 27764 4224
rect 27080 3998 27200 4026
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 27080 3194 27108 3998
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27068 3188 27120 3194
rect 27068 3130 27120 3136
rect 26700 2984 26752 2990
rect 26700 2926 26752 2932
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 25596 2372 25648 2378
rect 25596 2314 25648 2320
rect 25608 1170 25636 2314
rect 26068 1442 26096 2382
rect 26068 1414 26280 1442
rect 25424 1142 25636 1170
rect 25424 800 25452 1142
rect 26252 800 26280 1414
rect 27080 800 27108 2926
rect 27172 2650 27200 3878
rect 28092 3738 28120 4558
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27908 3194 27936 3334
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 28000 1850 28028 3470
rect 28092 3058 28120 3674
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28184 2446 28212 6854
rect 28368 6730 28396 7278
rect 29276 7200 29328 7206
rect 29276 7142 29328 7148
rect 28264 6724 28316 6730
rect 28264 6666 28316 6672
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28276 6458 28304 6666
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 29288 6322 29316 7142
rect 29380 7002 29408 7278
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 29368 6996 29420 7002
rect 29368 6938 29420 6944
rect 29472 6730 29500 7142
rect 29460 6724 29512 6730
rect 29460 6666 29512 6672
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 28460 4826 28488 5306
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 28460 4282 28488 4762
rect 29368 4616 29420 4622
rect 29368 4558 29420 4564
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28460 3058 28488 4218
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28828 3194 28856 3470
rect 28816 3188 28868 3194
rect 28816 3130 28868 3136
rect 29012 3126 29040 4422
rect 29380 4282 29408 4558
rect 29368 4276 29420 4282
rect 29368 4218 29420 4224
rect 29472 4214 29500 4966
rect 29460 4208 29512 4214
rect 29460 4150 29512 4156
rect 29092 3528 29144 3534
rect 29564 3505 29592 13194
rect 29748 12986 29776 14350
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 29838 14172 30146 14181
rect 29838 14170 29844 14172
rect 29900 14170 29924 14172
rect 29980 14170 30004 14172
rect 30060 14170 30084 14172
rect 30140 14170 30146 14172
rect 29900 14118 29902 14170
rect 30082 14118 30084 14170
rect 29838 14116 29844 14118
rect 29900 14116 29924 14118
rect 29980 14116 30004 14118
rect 30060 14116 30084 14118
rect 30140 14116 30146 14118
rect 29838 14107 30146 14116
rect 30392 14074 30420 14282
rect 31036 14278 31064 14486
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 30932 14000 30984 14006
rect 30932 13942 30984 13948
rect 30748 13184 30800 13190
rect 30748 13126 30800 13132
rect 29838 13084 30146 13093
rect 29838 13082 29844 13084
rect 29900 13082 29924 13084
rect 29980 13082 30004 13084
rect 30060 13082 30084 13084
rect 30140 13082 30146 13084
rect 29900 13030 29902 13082
rect 30082 13030 30084 13082
rect 29838 13028 29844 13030
rect 29900 13028 29924 13030
rect 29980 13028 30004 13030
rect 30060 13028 30084 13030
rect 30140 13028 30146 13030
rect 29838 13019 30146 13028
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29748 12238 29776 12378
rect 30380 12368 30432 12374
rect 30380 12310 30432 12316
rect 30392 12238 30420 12310
rect 29736 12232 29788 12238
rect 30380 12232 30432 12238
rect 29736 12174 29788 12180
rect 30378 12200 30380 12209
rect 30432 12200 30434 12209
rect 30378 12135 30434 12144
rect 29838 11996 30146 12005
rect 29838 11994 29844 11996
rect 29900 11994 29924 11996
rect 29980 11994 30004 11996
rect 30060 11994 30084 11996
rect 30140 11994 30146 11996
rect 29900 11942 29902 11994
rect 30082 11942 30084 11994
rect 29838 11940 29844 11942
rect 29900 11940 29924 11942
rect 29980 11940 30004 11942
rect 30060 11940 30084 11942
rect 30140 11940 30146 11942
rect 29838 11931 30146 11940
rect 30392 11354 30420 12135
rect 30656 12096 30708 12102
rect 30656 12038 30708 12044
rect 30668 11898 30696 12038
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 29838 10908 30146 10917
rect 29838 10906 29844 10908
rect 29900 10906 29924 10908
rect 29980 10906 30004 10908
rect 30060 10906 30084 10908
rect 30140 10906 30146 10908
rect 29900 10854 29902 10906
rect 30082 10854 30084 10906
rect 29838 10852 29844 10854
rect 29900 10852 29924 10854
rect 29980 10852 30004 10854
rect 30060 10852 30084 10854
rect 30140 10852 30146 10854
rect 29838 10843 30146 10852
rect 30760 10742 30788 13126
rect 30840 12096 30892 12102
rect 30840 12038 30892 12044
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 29644 9920 29696 9926
rect 29644 9862 29696 9868
rect 29656 9586 29684 9862
rect 29838 9820 30146 9829
rect 29838 9818 29844 9820
rect 29900 9818 29924 9820
rect 29980 9818 30004 9820
rect 30060 9818 30084 9820
rect 30140 9818 30146 9820
rect 29900 9766 29902 9818
rect 30082 9766 30084 9818
rect 29838 9764 29844 9766
rect 29900 9764 29924 9766
rect 29980 9764 30004 9766
rect 30060 9764 30084 9766
rect 30140 9764 30146 9766
rect 29838 9755 30146 9764
rect 30576 9586 30604 10610
rect 30852 10470 30880 12038
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30748 9988 30800 9994
rect 30748 9930 30800 9936
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 30564 9580 30616 9586
rect 30564 9522 30616 9528
rect 30288 9512 30340 9518
rect 30472 9512 30524 9518
rect 30288 9454 30340 9460
rect 30392 9472 30472 9500
rect 30196 9444 30248 9450
rect 30196 9386 30248 9392
rect 30208 9110 30236 9386
rect 30196 9104 30248 9110
rect 30196 9046 30248 9052
rect 30300 8974 30328 9454
rect 30288 8968 30340 8974
rect 30288 8910 30340 8916
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 29838 8732 30146 8741
rect 29838 8730 29844 8732
rect 29900 8730 29924 8732
rect 29980 8730 30004 8732
rect 30060 8730 30084 8732
rect 30140 8730 30146 8732
rect 29900 8678 29902 8730
rect 30082 8678 30084 8730
rect 29838 8676 29844 8678
rect 29900 8676 29924 8678
rect 29980 8676 30004 8678
rect 30060 8676 30084 8678
rect 30140 8676 30146 8678
rect 29838 8667 30146 8676
rect 30208 8498 30236 8774
rect 30392 8634 30420 9472
rect 30472 9454 30524 9460
rect 30472 8832 30524 8838
rect 30472 8774 30524 8780
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 29838 7644 30146 7653
rect 29838 7642 29844 7644
rect 29900 7642 29924 7644
rect 29980 7642 30004 7644
rect 30060 7642 30084 7644
rect 30140 7642 30146 7644
rect 29900 7590 29902 7642
rect 30082 7590 30084 7642
rect 29838 7588 29844 7590
rect 29900 7588 29924 7590
rect 29980 7588 30004 7590
rect 30060 7588 30084 7590
rect 30140 7588 30146 7590
rect 29838 7579 30146 7588
rect 30484 7546 30512 8774
rect 30760 8634 30788 9930
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30852 8634 30880 9318
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 30852 7546 30880 8570
rect 30472 7540 30524 7546
rect 30392 7500 30472 7528
rect 30196 7336 30248 7342
rect 30196 7278 30248 7284
rect 29838 6556 30146 6565
rect 29838 6554 29844 6556
rect 29900 6554 29924 6556
rect 29980 6554 30004 6556
rect 30060 6554 30084 6556
rect 30140 6554 30146 6556
rect 29900 6502 29902 6554
rect 30082 6502 30084 6554
rect 29838 6500 29844 6502
rect 29900 6500 29924 6502
rect 29980 6500 30004 6502
rect 30060 6500 30084 6502
rect 30140 6500 30146 6502
rect 29838 6491 30146 6500
rect 30208 6458 30236 7278
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29656 4622 29684 6258
rect 30392 6254 30420 7500
rect 30472 7482 30524 7488
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30944 7342 30972 13942
rect 31128 13938 31156 14418
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31312 12238 31340 14894
rect 31576 14272 31628 14278
rect 31576 14214 31628 14220
rect 31588 12306 31616 14214
rect 31680 14006 31708 17138
rect 31772 16590 31800 17274
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 31864 15570 31892 18838
rect 31956 18834 31984 19110
rect 31944 18828 31996 18834
rect 31944 18770 31996 18776
rect 31956 18426 31984 18770
rect 31944 18420 31996 18426
rect 31944 18362 31996 18368
rect 32036 18352 32088 18358
rect 32036 18294 32088 18300
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 31956 17678 31984 18226
rect 32048 18154 32076 18294
rect 32140 18290 32168 19246
rect 32324 18766 32352 19654
rect 32600 19310 32628 20946
rect 32588 19304 32640 19310
rect 32588 19246 32640 19252
rect 32404 19168 32456 19174
rect 32404 19110 32456 19116
rect 32416 18970 32444 19110
rect 32404 18964 32456 18970
rect 32404 18906 32456 18912
rect 32772 18828 32824 18834
rect 32772 18770 32824 18776
rect 32312 18760 32364 18766
rect 32588 18760 32640 18766
rect 32508 18737 32588 18748
rect 32312 18702 32364 18708
rect 32494 18728 32588 18737
rect 32128 18284 32180 18290
rect 32128 18226 32180 18232
rect 32036 18148 32088 18154
rect 32036 18090 32088 18096
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 31944 17128 31996 17134
rect 31944 17070 31996 17076
rect 31956 16250 31984 17070
rect 31944 16244 31996 16250
rect 31944 16186 31996 16192
rect 31852 15564 31904 15570
rect 31852 15506 31904 15512
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31668 14000 31720 14006
rect 31668 13942 31720 13948
rect 31576 12300 31628 12306
rect 31576 12242 31628 12248
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31312 11558 31340 12174
rect 31772 11830 31800 15302
rect 31864 13870 31892 15506
rect 32048 15162 32076 18090
rect 32128 16584 32180 16590
rect 32128 16526 32180 16532
rect 32140 16250 32168 16526
rect 32128 16244 32180 16250
rect 32128 16186 32180 16192
rect 32036 15156 32088 15162
rect 32036 15098 32088 15104
rect 32324 14958 32352 18702
rect 32550 18720 32588 18728
rect 32588 18702 32640 18708
rect 32494 18663 32550 18672
rect 32784 18086 32812 18770
rect 33416 18760 33468 18766
rect 33416 18702 33468 18708
rect 32864 18624 32916 18630
rect 32864 18566 32916 18572
rect 32876 18426 32904 18566
rect 32864 18420 32916 18426
rect 32864 18362 32916 18368
rect 33428 18290 33456 18702
rect 33520 18290 33548 21286
rect 33796 20806 33824 21286
rect 33980 21146 34008 22510
rect 34072 21690 34100 23054
rect 35808 23044 35860 23050
rect 35808 22986 35860 22992
rect 34244 22976 34296 22982
rect 34244 22918 34296 22924
rect 34256 22438 34284 22918
rect 34336 22636 34388 22642
rect 34336 22578 34388 22584
rect 34244 22432 34296 22438
rect 34244 22374 34296 22380
rect 34256 22114 34284 22374
rect 34348 22234 34376 22578
rect 35256 22500 35308 22506
rect 35256 22442 35308 22448
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 34336 22228 34388 22234
rect 34336 22170 34388 22176
rect 34256 22086 34376 22114
rect 34152 21888 34204 21894
rect 34152 21830 34204 21836
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 34164 21434 34192 21830
rect 34072 21406 34192 21434
rect 34072 21350 34100 21406
rect 34060 21344 34112 21350
rect 34060 21286 34112 21292
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 33784 20800 33836 20806
rect 33784 20742 33836 20748
rect 33796 19786 33824 20742
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33692 19712 33744 19718
rect 33692 19654 33744 19660
rect 33704 18834 33732 19654
rect 33692 18828 33744 18834
rect 33692 18770 33744 18776
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32680 17740 32732 17746
rect 32680 17682 32732 17688
rect 32692 17338 32720 17682
rect 32784 17542 32812 18022
rect 33152 17882 33180 18226
rect 33140 17876 33192 17882
rect 33140 17818 33192 17824
rect 33428 17746 33456 18226
rect 33704 18086 33732 18770
rect 33600 18080 33652 18086
rect 33600 18022 33652 18028
rect 33692 18080 33744 18086
rect 33692 18022 33744 18028
rect 33508 17876 33560 17882
rect 33508 17818 33560 17824
rect 33416 17740 33468 17746
rect 33416 17682 33468 17688
rect 32772 17536 32824 17542
rect 32772 17478 32824 17484
rect 32680 17332 32732 17338
rect 32680 17274 32732 17280
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32508 15570 32536 16186
rect 32588 15972 32640 15978
rect 32588 15914 32640 15920
rect 32496 15564 32548 15570
rect 32496 15506 32548 15512
rect 32600 15502 32628 15914
rect 32588 15496 32640 15502
rect 32588 15438 32640 15444
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32600 14618 32628 15438
rect 32588 14612 32640 14618
rect 32588 14554 32640 14560
rect 32404 14408 32456 14414
rect 32404 14350 32456 14356
rect 32416 14074 32444 14350
rect 32404 14068 32456 14074
rect 32404 14010 32456 14016
rect 31852 13864 31904 13870
rect 31852 13806 31904 13812
rect 32588 13388 32640 13394
rect 32588 13330 32640 13336
rect 31852 12844 31904 12850
rect 31852 12786 31904 12792
rect 31760 11824 31812 11830
rect 31760 11766 31812 11772
rect 31864 11762 31892 12786
rect 32600 12434 32628 13330
rect 32600 12406 32720 12434
rect 32692 12374 32720 12406
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 31944 12300 31996 12306
rect 31944 12242 31996 12248
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 31956 11642 31984 12242
rect 31772 11620 31984 11642
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 31772 11614 31852 11620
rect 31300 11552 31352 11558
rect 31300 11494 31352 11500
rect 31208 10668 31260 10674
rect 31208 10610 31260 10616
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31128 9178 31156 10066
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 30932 7336 30984 7342
rect 30932 7278 30984 7284
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 30380 6248 30432 6254
rect 30380 6190 30432 6196
rect 30392 6118 30420 6190
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30392 5914 30420 6054
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 29736 5636 29788 5642
rect 29736 5578 29788 5584
rect 29644 4616 29696 4622
rect 29644 4558 29696 4564
rect 29748 3738 29776 5578
rect 29838 5468 30146 5477
rect 29838 5466 29844 5468
rect 29900 5466 29924 5468
rect 29980 5466 30004 5468
rect 30060 5466 30084 5468
rect 30140 5466 30146 5468
rect 29900 5414 29902 5466
rect 30082 5414 30084 5466
rect 29838 5412 29844 5414
rect 29900 5412 29924 5414
rect 29980 5412 30004 5414
rect 30060 5412 30084 5414
rect 30140 5412 30146 5414
rect 29838 5403 30146 5412
rect 30392 5250 30420 5850
rect 30300 5222 30420 5250
rect 30196 4752 30248 4758
rect 30194 4720 30196 4729
rect 30248 4720 30250 4729
rect 30194 4655 30250 4664
rect 30196 4480 30248 4486
rect 30196 4422 30248 4428
rect 29838 4380 30146 4389
rect 29838 4378 29844 4380
rect 29900 4378 29924 4380
rect 29980 4378 30004 4380
rect 30060 4378 30084 4380
rect 30140 4378 30146 4380
rect 29900 4326 29902 4378
rect 30082 4326 30084 4378
rect 29838 4324 29844 4326
rect 29900 4324 29924 4326
rect 29980 4324 30004 4326
rect 30060 4324 30084 4326
rect 30140 4324 30146 4326
rect 29838 4315 30146 4324
rect 30208 4146 30236 4422
rect 30300 4282 30328 5222
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30288 4276 30340 4282
rect 30288 4218 30340 4224
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 30392 4026 30420 5102
rect 30484 4826 30512 6326
rect 30944 5914 30972 7278
rect 31024 6656 31076 6662
rect 31024 6598 31076 6604
rect 31036 6390 31064 6598
rect 31024 6384 31076 6390
rect 31024 6326 31076 6332
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 30472 4820 30524 4826
rect 30472 4762 30524 4768
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30484 4282 30512 4558
rect 30472 4276 30524 4282
rect 30472 4218 30524 4224
rect 30208 4010 30420 4026
rect 30576 4010 30604 5170
rect 30196 4004 30420 4010
rect 30248 3998 30420 4004
rect 30564 4004 30616 4010
rect 30196 3946 30248 3952
rect 30564 3946 30616 3952
rect 30668 3942 30696 5510
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 29736 3732 29788 3738
rect 29736 3674 29788 3680
rect 29092 3470 29144 3476
rect 29550 3496 29606 3505
rect 29000 3120 29052 3126
rect 29000 3062 29052 3068
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 29104 2650 29132 3470
rect 29550 3431 29606 3440
rect 29838 3292 30146 3301
rect 29838 3290 29844 3292
rect 29900 3290 29924 3292
rect 29980 3290 30004 3292
rect 30060 3290 30084 3292
rect 30140 3290 30146 3292
rect 29900 3238 29902 3290
rect 30082 3238 30084 3290
rect 29838 3236 29844 3238
rect 29900 3236 29924 3238
rect 29980 3236 30004 3238
rect 30060 3236 30084 3238
rect 30140 3236 30146 3238
rect 29838 3227 30146 3236
rect 30944 2990 30972 5170
rect 31024 5024 31076 5030
rect 31024 4966 31076 4972
rect 31036 4282 31064 4966
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 31128 4078 31156 5850
rect 31116 4072 31168 4078
rect 31116 4014 31168 4020
rect 31220 3942 31248 10610
rect 31772 9178 31800 11614
rect 31904 11614 31984 11620
rect 31852 11562 31904 11568
rect 32036 11552 32088 11558
rect 32036 11494 32088 11500
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31760 9172 31812 9178
rect 31760 9114 31812 9120
rect 31772 8838 31800 9114
rect 31760 8832 31812 8838
rect 31760 8774 31812 8780
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31404 8090 31432 8366
rect 31864 8362 31892 10406
rect 31944 9512 31996 9518
rect 31944 9454 31996 9460
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31392 8084 31444 8090
rect 31392 8026 31444 8032
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31772 7546 31800 7822
rect 31760 7540 31812 7546
rect 31760 7482 31812 7488
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 31312 4826 31340 5102
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31588 4690 31616 4966
rect 31576 4684 31628 4690
rect 31576 4626 31628 4632
rect 31956 4622 31984 9454
rect 32048 9382 32076 11494
rect 32128 9512 32180 9518
rect 32128 9454 32180 9460
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 32048 8294 32076 9318
rect 32036 8288 32088 8294
rect 32036 8230 32088 8236
rect 32140 7954 32168 9454
rect 32404 9376 32456 9382
rect 32404 9318 32456 9324
rect 32416 8838 32444 9318
rect 32404 8832 32456 8838
rect 32404 8774 32456 8780
rect 32128 7948 32180 7954
rect 32128 7890 32180 7896
rect 32140 6798 32168 7890
rect 32128 6792 32180 6798
rect 32128 6734 32180 6740
rect 32140 6322 32168 6734
rect 32128 6316 32180 6322
rect 32128 6258 32180 6264
rect 32416 5030 32444 8774
rect 32404 5024 32456 5030
rect 32404 4966 32456 4972
rect 32416 4758 32444 4966
rect 32404 4752 32456 4758
rect 32402 4720 32404 4729
rect 32456 4720 32458 4729
rect 32402 4655 32458 4664
rect 31944 4616 31996 4622
rect 31944 4558 31996 4564
rect 31484 4480 31536 4486
rect 31484 4422 31536 4428
rect 31208 3936 31260 3942
rect 31208 3878 31260 3884
rect 31496 3194 31524 4422
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 31576 4072 31628 4078
rect 31576 4014 31628 4020
rect 31588 3194 31616 4014
rect 31484 3188 31536 3194
rect 31484 3130 31536 3136
rect 31576 3188 31628 3194
rect 31576 3130 31628 3136
rect 30932 2984 30984 2990
rect 30932 2926 30984 2932
rect 31680 2650 31708 4082
rect 31944 3392 31996 3398
rect 31944 3334 31996 3340
rect 31956 2990 31984 3334
rect 32508 3194 32536 11494
rect 32600 11354 32628 11630
rect 32784 11354 32812 17478
rect 33520 17338 33548 17818
rect 33508 17332 33560 17338
rect 33508 17274 33560 17280
rect 32956 16992 33008 16998
rect 32956 16934 33008 16940
rect 32968 16250 32996 16934
rect 33140 16652 33192 16658
rect 33140 16594 33192 16600
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 33152 16046 33180 16594
rect 33612 16538 33640 18022
rect 33704 17184 33732 18022
rect 33784 17196 33836 17202
rect 33704 17156 33784 17184
rect 33704 16658 33732 17156
rect 33784 17138 33836 17144
rect 33784 16992 33836 16998
rect 33784 16934 33836 16940
rect 33692 16652 33744 16658
rect 33692 16594 33744 16600
rect 33428 16510 33640 16538
rect 32956 16040 33008 16046
rect 32956 15982 33008 15988
rect 33140 16040 33192 16046
rect 33140 15982 33192 15988
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 32876 11626 32904 13806
rect 32968 12238 32996 15982
rect 33048 13456 33100 13462
rect 33048 13398 33100 13404
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32968 12102 32996 12174
rect 32956 12096 33008 12102
rect 32956 12038 33008 12044
rect 32864 11620 32916 11626
rect 32864 11562 32916 11568
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 32680 11008 32732 11014
rect 32680 10950 32732 10956
rect 32692 10062 32720 10950
rect 33060 10470 33088 13398
rect 33140 13252 33192 13258
rect 33140 13194 33192 13200
rect 33152 11694 33180 13194
rect 33232 12844 33284 12850
rect 33232 12786 33284 12792
rect 33244 11694 33272 12786
rect 33428 12434 33456 16510
rect 33600 16448 33652 16454
rect 33600 16390 33652 16396
rect 33612 15706 33640 16390
rect 33692 16108 33744 16114
rect 33692 16050 33744 16056
rect 33600 15700 33652 15706
rect 33600 15642 33652 15648
rect 33704 15502 33732 16050
rect 33796 16046 33824 16934
rect 33784 16040 33836 16046
rect 33784 15982 33836 15988
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33704 15162 33732 15438
rect 33968 15360 34020 15366
rect 33968 15302 34020 15308
rect 33692 15156 33744 15162
rect 33692 15098 33744 15104
rect 33980 15026 34008 15302
rect 33968 15020 34020 15026
rect 33968 14962 34020 14968
rect 34072 14906 34100 21286
rect 34244 17740 34296 17746
rect 34244 17682 34296 17688
rect 34152 16584 34204 16590
rect 34152 16526 34204 16532
rect 34164 16250 34192 16526
rect 34152 16244 34204 16250
rect 34152 16186 34204 16192
rect 33980 14878 34100 14906
rect 33508 13864 33560 13870
rect 33508 13806 33560 13812
rect 33520 12986 33548 13806
rect 33980 13802 34008 14878
rect 34060 14000 34112 14006
rect 34060 13942 34112 13948
rect 33968 13796 34020 13802
rect 33968 13738 34020 13744
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33600 12640 33652 12646
rect 33600 12582 33652 12588
rect 33428 12406 33548 12434
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33416 12096 33468 12102
rect 33416 12038 33468 12044
rect 33336 11898 33364 12038
rect 33428 11898 33456 12038
rect 33324 11892 33376 11898
rect 33324 11834 33376 11840
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33140 11688 33192 11694
rect 33140 11630 33192 11636
rect 33232 11688 33284 11694
rect 33232 11630 33284 11636
rect 33324 11076 33376 11082
rect 33324 11018 33376 11024
rect 33232 11008 33284 11014
rect 33232 10950 33284 10956
rect 33244 10538 33272 10950
rect 33232 10532 33284 10538
rect 33232 10474 33284 10480
rect 33048 10464 33100 10470
rect 33048 10406 33100 10412
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 33140 9580 33192 9586
rect 33140 9522 33192 9528
rect 33152 9178 33180 9522
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33140 7880 33192 7886
rect 33140 7822 33192 7828
rect 32588 7744 32640 7750
rect 32588 7686 32640 7692
rect 32600 6730 32628 7686
rect 33152 7546 33180 7822
rect 33140 7540 33192 7546
rect 33140 7482 33192 7488
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32956 6316 33008 6322
rect 32956 6258 33008 6264
rect 32968 5914 32996 6258
rect 32956 5908 33008 5914
rect 32956 5850 33008 5856
rect 33336 4826 33364 11018
rect 33520 7732 33548 12406
rect 33612 12306 33640 12582
rect 34072 12306 34100 13942
rect 34152 13864 34204 13870
rect 34152 13806 34204 13812
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 34060 12300 34112 12306
rect 34060 12242 34112 12248
rect 34072 11626 34100 12242
rect 34164 12170 34192 13806
rect 34256 13530 34284 17682
rect 34348 15502 34376 22086
rect 34440 21690 34468 22374
rect 35072 22228 35124 22234
rect 35072 22170 35124 22176
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34428 21684 34480 21690
rect 34428 21626 34480 21632
rect 34716 21146 34744 21830
rect 34704 21140 34756 21146
rect 34704 21082 34756 21088
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34716 18970 34744 19246
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34532 17882 34560 18158
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34532 16658 34560 16934
rect 34520 16652 34572 16658
rect 34520 16594 34572 16600
rect 34428 16108 34480 16114
rect 34428 16050 34480 16056
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 34348 14006 34376 15438
rect 34440 15162 34468 16050
rect 35084 15638 35112 22170
rect 35268 22030 35296 22442
rect 35820 22234 35848 22986
rect 35992 22976 36044 22982
rect 35992 22918 36044 22924
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 35256 22024 35308 22030
rect 35256 21966 35308 21972
rect 35452 21554 35480 22034
rect 36004 21554 36032 22918
rect 36464 22778 36492 23054
rect 39856 22976 39908 22982
rect 39856 22918 39908 22924
rect 39868 22778 39896 22918
rect 36452 22772 36504 22778
rect 36452 22714 36504 22720
rect 38660 22772 38712 22778
rect 38660 22714 38712 22720
rect 39856 22772 39908 22778
rect 39856 22714 39908 22720
rect 37464 22568 37516 22574
rect 37464 22510 37516 22516
rect 38568 22568 38620 22574
rect 38568 22510 38620 22516
rect 37060 22332 37368 22341
rect 37060 22330 37066 22332
rect 37122 22330 37146 22332
rect 37202 22330 37226 22332
rect 37282 22330 37306 22332
rect 37362 22330 37368 22332
rect 37122 22278 37124 22330
rect 37304 22278 37306 22330
rect 37060 22276 37066 22278
rect 37122 22276 37146 22278
rect 37202 22276 37226 22278
rect 37282 22276 37306 22278
rect 37362 22276 37368 22278
rect 37060 22267 37368 22276
rect 36360 21956 36412 21962
rect 36360 21898 36412 21904
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35992 21548 36044 21554
rect 35992 21490 36044 21496
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 35256 19508 35308 19514
rect 35256 19450 35308 19456
rect 35268 18834 35296 19450
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 35256 17196 35308 17202
rect 35256 17138 35308 17144
rect 35164 15904 35216 15910
rect 35164 15846 35216 15852
rect 35176 15706 35204 15846
rect 35164 15700 35216 15706
rect 35164 15642 35216 15648
rect 35072 15632 35124 15638
rect 35072 15574 35124 15580
rect 34612 15360 34664 15366
rect 34612 15302 34664 15308
rect 34704 15360 34756 15366
rect 34704 15302 34756 15308
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34624 14822 34652 15302
rect 34716 15026 34744 15302
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 34612 14816 34664 14822
rect 34612 14758 34664 14764
rect 35084 14618 35112 15574
rect 35268 15434 35296 17138
rect 35360 16794 35388 19654
rect 35452 19378 35480 21490
rect 36372 21146 36400 21898
rect 36820 21888 36872 21894
rect 36820 21830 36872 21836
rect 36912 21888 36964 21894
rect 36912 21830 36964 21836
rect 36832 21554 36860 21830
rect 36820 21548 36872 21554
rect 36820 21490 36872 21496
rect 36360 21140 36412 21146
rect 36360 21082 36412 21088
rect 36924 21010 36952 21830
rect 37476 21690 37504 22510
rect 37556 22432 37608 22438
rect 37556 22374 37608 22380
rect 37568 21894 37596 22374
rect 37832 22092 37884 22098
rect 37832 22034 37884 22040
rect 37556 21888 37608 21894
rect 37556 21830 37608 21836
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37568 21570 37596 21830
rect 37844 21690 37872 22034
rect 38384 22024 38436 22030
rect 38384 21966 38436 21972
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 37476 21542 37596 21570
rect 37060 21244 37368 21253
rect 37060 21242 37066 21244
rect 37122 21242 37146 21244
rect 37202 21242 37226 21244
rect 37282 21242 37306 21244
rect 37362 21242 37368 21244
rect 37122 21190 37124 21242
rect 37304 21190 37306 21242
rect 37060 21188 37066 21190
rect 37122 21188 37146 21190
rect 37202 21188 37226 21190
rect 37282 21188 37306 21190
rect 37362 21188 37368 21190
rect 37060 21179 37368 21188
rect 36912 21004 36964 21010
rect 36912 20946 36964 20952
rect 37060 20156 37368 20165
rect 37060 20154 37066 20156
rect 37122 20154 37146 20156
rect 37202 20154 37226 20156
rect 37282 20154 37306 20156
rect 37362 20154 37368 20156
rect 37122 20102 37124 20154
rect 37304 20102 37306 20154
rect 37060 20100 37066 20102
rect 37122 20100 37146 20102
rect 37202 20100 37226 20102
rect 37282 20100 37306 20102
rect 37362 20100 37368 20102
rect 37060 20091 37368 20100
rect 36912 19916 36964 19922
rect 36912 19858 36964 19864
rect 35992 19440 36044 19446
rect 35992 19382 36044 19388
rect 35440 19372 35492 19378
rect 35440 19314 35492 19320
rect 35440 18828 35492 18834
rect 35440 18770 35492 18776
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 35452 15978 35480 18770
rect 36004 18426 36032 19382
rect 36728 19168 36780 19174
rect 36728 19110 36780 19116
rect 36740 18834 36768 19110
rect 36924 18970 36952 19858
rect 37060 19068 37368 19077
rect 37060 19066 37066 19068
rect 37122 19066 37146 19068
rect 37202 19066 37226 19068
rect 37282 19066 37306 19068
rect 37362 19066 37368 19068
rect 37122 19014 37124 19066
rect 37304 19014 37306 19066
rect 37060 19012 37066 19014
rect 37122 19012 37146 19014
rect 37202 19012 37226 19014
rect 37282 19012 37306 19014
rect 37362 19012 37368 19014
rect 37060 19003 37368 19012
rect 36912 18964 36964 18970
rect 37476 18952 37504 21542
rect 38396 21078 38424 21966
rect 38580 21622 38608 22510
rect 38672 22098 38700 22714
rect 38936 22432 38988 22438
rect 38936 22374 38988 22380
rect 39212 22432 39264 22438
rect 39212 22374 39264 22380
rect 38948 22098 38976 22374
rect 39120 22160 39172 22166
rect 39120 22102 39172 22108
rect 38660 22092 38712 22098
rect 38660 22034 38712 22040
rect 38936 22092 38988 22098
rect 38936 22034 38988 22040
rect 39028 21888 39080 21894
rect 39028 21830 39080 21836
rect 38568 21616 38620 21622
rect 38568 21558 38620 21564
rect 38580 21146 38608 21558
rect 38568 21140 38620 21146
rect 38568 21082 38620 21088
rect 37648 21072 37700 21078
rect 37648 21014 37700 21020
rect 38384 21072 38436 21078
rect 38384 21014 38436 21020
rect 37660 20602 37688 21014
rect 37832 20800 37884 20806
rect 37832 20742 37884 20748
rect 37648 20596 37700 20602
rect 37648 20538 37700 20544
rect 37648 19848 37700 19854
rect 37648 19790 37700 19796
rect 37556 19712 37608 19718
rect 37556 19654 37608 19660
rect 36912 18906 36964 18912
rect 37292 18924 37504 18952
rect 36728 18828 36780 18834
rect 36728 18770 36780 18776
rect 36084 18624 36136 18630
rect 36084 18566 36136 18572
rect 36096 18426 36124 18566
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 36084 18420 36136 18426
rect 36084 18362 36136 18368
rect 36740 18290 36768 18770
rect 37292 18630 37320 18924
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 37292 18358 37320 18566
rect 37280 18352 37332 18358
rect 37280 18294 37332 18300
rect 36728 18284 36780 18290
rect 36728 18226 36780 18232
rect 35716 18148 35768 18154
rect 35716 18090 35768 18096
rect 35728 17882 35756 18090
rect 35716 17876 35768 17882
rect 35716 17818 35768 17824
rect 36084 17672 36136 17678
rect 36084 17614 36136 17620
rect 35808 17536 35860 17542
rect 35808 17478 35860 17484
rect 35820 17338 35848 17478
rect 35808 17332 35860 17338
rect 35808 17274 35860 17280
rect 35808 16992 35860 16998
rect 35808 16934 35860 16940
rect 35820 16590 35848 16934
rect 36096 16726 36124 17614
rect 36176 16992 36228 16998
rect 36176 16934 36228 16940
rect 36188 16794 36216 16934
rect 36176 16788 36228 16794
rect 36176 16730 36228 16736
rect 36084 16720 36136 16726
rect 36084 16662 36136 16668
rect 35808 16584 35860 16590
rect 35808 16526 35860 16532
rect 36096 16096 36124 16662
rect 36176 16108 36228 16114
rect 36096 16068 36176 16096
rect 36176 16050 36228 16056
rect 35716 16040 35768 16046
rect 35716 15982 35768 15988
rect 35992 16040 36044 16046
rect 35992 15982 36044 15988
rect 35440 15972 35492 15978
rect 35440 15914 35492 15920
rect 35256 15428 35308 15434
rect 35256 15370 35308 15376
rect 35072 14612 35124 14618
rect 35072 14554 35124 14560
rect 34428 14340 34480 14346
rect 34428 14282 34480 14288
rect 34336 14000 34388 14006
rect 34336 13942 34388 13948
rect 34440 13938 34468 14282
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34336 13796 34388 13802
rect 34336 13738 34388 13744
rect 34244 13524 34296 13530
rect 34244 13466 34296 13472
rect 34348 13394 34376 13738
rect 34336 13388 34388 13394
rect 34336 13330 34388 13336
rect 34348 12374 34376 13330
rect 34440 12850 34468 13874
rect 34796 13184 34848 13190
rect 34796 13126 34848 13132
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34612 12844 34664 12850
rect 34612 12786 34664 12792
rect 34624 12374 34652 12786
rect 34336 12368 34388 12374
rect 34336 12310 34388 12316
rect 34612 12368 34664 12374
rect 34612 12310 34664 12316
rect 34152 12164 34204 12170
rect 34152 12106 34204 12112
rect 34348 11762 34376 12310
rect 34808 12306 34836 13126
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 35084 12209 35112 14554
rect 35268 13394 35296 15370
rect 35452 14618 35480 15914
rect 35728 14958 35756 15982
rect 35808 15564 35860 15570
rect 35808 15506 35860 15512
rect 35716 14952 35768 14958
rect 35716 14894 35768 14900
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35452 13394 35480 14554
rect 35728 13734 35756 14894
rect 35820 14822 35848 15506
rect 36004 15502 36032 15982
rect 36360 15972 36412 15978
rect 36360 15914 36412 15920
rect 36084 15632 36136 15638
rect 36084 15574 36136 15580
rect 35992 15496 36044 15502
rect 35992 15438 36044 15444
rect 36096 15314 36124 15574
rect 36372 15570 36400 15914
rect 36544 15904 36596 15910
rect 36544 15846 36596 15852
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36004 15286 36124 15314
rect 35808 14816 35860 14822
rect 35808 14758 35860 14764
rect 35820 13818 35848 14758
rect 35820 13790 35940 13818
rect 35716 13728 35768 13734
rect 35716 13670 35768 13676
rect 35808 13728 35860 13734
rect 35808 13670 35860 13676
rect 35728 13394 35756 13670
rect 35256 13388 35308 13394
rect 35256 13330 35308 13336
rect 35440 13388 35492 13394
rect 35440 13330 35492 13336
rect 35716 13388 35768 13394
rect 35716 13330 35768 13336
rect 35164 13184 35216 13190
rect 35164 13126 35216 13132
rect 35176 12374 35204 13126
rect 35268 12986 35296 13330
rect 35256 12980 35308 12986
rect 35256 12922 35308 12928
rect 35164 12368 35216 12374
rect 35164 12310 35216 12316
rect 35070 12200 35126 12209
rect 35070 12135 35126 12144
rect 34336 11756 34388 11762
rect 34336 11698 34388 11704
rect 34060 11620 34112 11626
rect 34060 11562 34112 11568
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 34336 11144 34388 11150
rect 34336 11086 34388 11092
rect 33612 10538 33640 11086
rect 33784 11008 33836 11014
rect 33784 10950 33836 10956
rect 33796 10742 33824 10950
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 34244 10736 34296 10742
rect 34244 10678 34296 10684
rect 33968 10600 34020 10606
rect 33968 10542 34020 10548
rect 33600 10532 33652 10538
rect 33600 10474 33652 10480
rect 33980 10062 34008 10542
rect 34256 10130 34284 10678
rect 34348 10198 34376 11086
rect 34888 11008 34940 11014
rect 34888 10950 34940 10956
rect 34900 10674 34928 10950
rect 34888 10668 34940 10674
rect 34888 10610 34940 10616
rect 34900 10266 34928 10610
rect 34888 10260 34940 10266
rect 34888 10202 34940 10208
rect 34336 10192 34388 10198
rect 34336 10134 34388 10140
rect 34244 10124 34296 10130
rect 34244 10066 34296 10072
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 34428 10056 34480 10062
rect 34428 9998 34480 10004
rect 33600 9920 33652 9926
rect 33600 9862 33652 9868
rect 33612 9042 33640 9862
rect 33784 9376 33836 9382
rect 33784 9318 33836 9324
rect 33796 9178 33824 9318
rect 33784 9172 33836 9178
rect 33784 9114 33836 9120
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 34440 8922 34468 9998
rect 34520 9988 34572 9994
rect 34520 9930 34572 9936
rect 34532 9178 34560 9930
rect 34704 9920 34756 9926
rect 34704 9862 34756 9868
rect 34716 9722 34744 9862
rect 34704 9716 34756 9722
rect 35084 9674 35112 12135
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 35360 11150 35388 11494
rect 35348 11144 35400 11150
rect 35346 11112 35348 11121
rect 35400 11112 35402 11121
rect 35346 11047 35402 11056
rect 35452 11014 35480 13330
rect 35820 12782 35848 13670
rect 35808 12776 35860 12782
rect 35808 12718 35860 12724
rect 35716 12640 35768 12646
rect 35716 12582 35768 12588
rect 35728 12306 35756 12582
rect 35912 12306 35940 13790
rect 36004 13462 36032 15286
rect 36084 14408 36136 14414
rect 36084 14350 36136 14356
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 36096 14074 36124 14350
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 36084 13864 36136 13870
rect 36084 13806 36136 13812
rect 35992 13456 36044 13462
rect 35992 13398 36044 13404
rect 36096 12986 36124 13806
rect 36188 13308 36216 14350
rect 36556 14074 36584 15846
rect 36636 15564 36688 15570
rect 36636 15506 36688 15512
rect 36648 15366 36676 15506
rect 36636 15360 36688 15366
rect 36636 15302 36688 15308
rect 36544 14068 36596 14074
rect 36544 14010 36596 14016
rect 36636 13864 36688 13870
rect 36636 13806 36688 13812
rect 36648 13530 36676 13806
rect 36740 13734 36768 18226
rect 37060 17980 37368 17989
rect 37060 17978 37066 17980
rect 37122 17978 37146 17980
rect 37202 17978 37226 17980
rect 37282 17978 37306 17980
rect 37362 17978 37368 17980
rect 37122 17926 37124 17978
rect 37304 17926 37306 17978
rect 37060 17924 37066 17926
rect 37122 17924 37146 17926
rect 37202 17924 37226 17926
rect 37282 17924 37306 17926
rect 37362 17924 37368 17926
rect 37060 17915 37368 17924
rect 37476 17542 37504 18566
rect 37568 18290 37596 19654
rect 37660 19514 37688 19790
rect 37740 19712 37792 19718
rect 37740 19654 37792 19660
rect 37648 19508 37700 19514
rect 37648 19450 37700 19456
rect 37648 19168 37700 19174
rect 37648 19110 37700 19116
rect 37660 18970 37688 19110
rect 37648 18964 37700 18970
rect 37648 18906 37700 18912
rect 37556 18284 37608 18290
rect 37556 18226 37608 18232
rect 37464 17536 37516 17542
rect 37464 17478 37516 17484
rect 37476 17066 37504 17478
rect 37464 17060 37516 17066
rect 37464 17002 37516 17008
rect 37060 16892 37368 16901
rect 37060 16890 37066 16892
rect 37122 16890 37146 16892
rect 37202 16890 37226 16892
rect 37282 16890 37306 16892
rect 37362 16890 37368 16892
rect 37122 16838 37124 16890
rect 37304 16838 37306 16890
rect 37060 16836 37066 16838
rect 37122 16836 37146 16838
rect 37202 16836 37226 16838
rect 37282 16836 37306 16838
rect 37362 16836 37368 16838
rect 37060 16827 37368 16836
rect 37476 16794 37504 17002
rect 37556 16992 37608 16998
rect 37556 16934 37608 16940
rect 37464 16788 37516 16794
rect 37464 16730 37516 16736
rect 37568 16590 37596 16934
rect 37556 16584 37608 16590
rect 37556 16526 37608 16532
rect 37660 16538 37688 18906
rect 37752 18698 37780 19654
rect 37740 18692 37792 18698
rect 37740 18634 37792 18640
rect 37844 17610 37872 20742
rect 38108 20256 38160 20262
rect 38108 20198 38160 20204
rect 38120 19922 38148 20198
rect 38108 19916 38160 19922
rect 38108 19858 38160 19864
rect 37924 19168 37976 19174
rect 37924 19110 37976 19116
rect 37936 18834 37964 19110
rect 37924 18828 37976 18834
rect 37924 18770 37976 18776
rect 37936 18426 37964 18770
rect 37924 18420 37976 18426
rect 37924 18362 37976 18368
rect 38120 17746 38148 19858
rect 38396 19394 38424 21014
rect 38844 19984 38896 19990
rect 38844 19926 38896 19932
rect 38476 19712 38528 19718
rect 38476 19654 38528 19660
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 38212 19366 38424 19394
rect 38488 19378 38516 19654
rect 38476 19372 38528 19378
rect 38212 19334 38240 19366
rect 38212 19310 38424 19334
rect 38476 19314 38528 19320
rect 38212 19306 38436 19310
rect 38384 19304 38436 19306
rect 38384 19246 38436 19252
rect 38108 17740 38160 17746
rect 38108 17682 38160 17688
rect 37832 17604 37884 17610
rect 37832 17546 37884 17552
rect 37924 17128 37976 17134
rect 37924 17070 37976 17076
rect 37464 16516 37516 16522
rect 37660 16510 37780 16538
rect 37464 16458 37516 16464
rect 36820 16040 36872 16046
rect 36820 15982 36872 15988
rect 36832 15638 36860 15982
rect 37060 15804 37368 15813
rect 37060 15802 37066 15804
rect 37122 15802 37146 15804
rect 37202 15802 37226 15804
rect 37282 15802 37306 15804
rect 37362 15802 37368 15804
rect 37122 15750 37124 15802
rect 37304 15750 37306 15802
rect 37060 15748 37066 15750
rect 37122 15748 37146 15750
rect 37202 15748 37226 15750
rect 37282 15748 37306 15750
rect 37362 15748 37368 15750
rect 37060 15739 37368 15748
rect 36820 15632 36872 15638
rect 36820 15574 36872 15580
rect 37060 14716 37368 14725
rect 37060 14714 37066 14716
rect 37122 14714 37146 14716
rect 37202 14714 37226 14716
rect 37282 14714 37306 14716
rect 37362 14714 37368 14716
rect 37122 14662 37124 14714
rect 37304 14662 37306 14714
rect 37060 14660 37066 14662
rect 37122 14660 37146 14662
rect 37202 14660 37226 14662
rect 37282 14660 37306 14662
rect 37362 14660 37368 14662
rect 37060 14651 37368 14660
rect 37476 14618 37504 16458
rect 37648 16448 37700 16454
rect 37648 16390 37700 16396
rect 37660 16250 37688 16390
rect 37648 16244 37700 16250
rect 37648 16186 37700 16192
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37556 15904 37608 15910
rect 37556 15846 37608 15852
rect 37568 15706 37596 15846
rect 37556 15700 37608 15706
rect 37556 15642 37608 15648
rect 37660 15434 37688 16050
rect 37648 15428 37700 15434
rect 37648 15370 37700 15376
rect 37464 14612 37516 14618
rect 37464 14554 37516 14560
rect 36820 14272 36872 14278
rect 36820 14214 36872 14220
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 37004 14272 37056 14278
rect 37004 14214 37056 14220
rect 36728 13728 36780 13734
rect 36728 13670 36780 13676
rect 36636 13524 36688 13530
rect 36636 13466 36688 13472
rect 36728 13388 36780 13394
rect 36832 13376 36860 14214
rect 36780 13348 36860 13376
rect 36728 13330 36780 13336
rect 36636 13320 36688 13326
rect 36188 13280 36308 13308
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 35716 12300 35768 12306
rect 35716 12242 35768 12248
rect 35900 12300 35952 12306
rect 35900 12242 35952 12248
rect 35912 12102 35940 12242
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 35716 11552 35768 11558
rect 35716 11494 35768 11500
rect 35728 11286 35756 11494
rect 35716 11280 35768 11286
rect 35716 11222 35768 11228
rect 35440 11008 35492 11014
rect 35440 10950 35492 10956
rect 35452 10390 35664 10418
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 34704 9658 34756 9664
rect 34900 9646 35112 9674
rect 34612 9580 34664 9586
rect 34612 9522 34664 9528
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34440 8906 34560 8922
rect 34440 8900 34572 8906
rect 34440 8894 34520 8900
rect 34520 8842 34572 8848
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34152 8084 34204 8090
rect 34152 8026 34204 8032
rect 33428 7704 33548 7732
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 33048 4752 33100 4758
rect 33048 4694 33100 4700
rect 32864 3936 32916 3942
rect 32864 3878 32916 3884
rect 32876 3466 32904 3878
rect 32864 3460 32916 3466
rect 32864 3402 32916 3408
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 33060 2990 33088 4694
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 33152 3194 33180 4014
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 33244 3194 33272 3878
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33140 3188 33192 3194
rect 33140 3130 33192 3136
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 28724 2508 28776 2514
rect 28724 2450 28776 2456
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 27908 1822 28028 1850
rect 27908 800 27936 1822
rect 28736 800 28764 2450
rect 31956 2446 31984 2926
rect 33336 2446 33364 3674
rect 33428 3126 33456 7704
rect 33968 7472 34020 7478
rect 33968 7414 34020 7420
rect 33600 7336 33652 7342
rect 33600 7278 33652 7284
rect 33612 7002 33640 7278
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33692 6928 33744 6934
rect 33692 6870 33744 6876
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33520 5914 33548 6598
rect 33704 6458 33732 6870
rect 33980 6866 34008 7414
rect 34164 6866 34192 8026
rect 33968 6860 34020 6866
rect 33968 6802 34020 6808
rect 34152 6860 34204 6866
rect 34152 6802 34204 6808
rect 33876 6656 33928 6662
rect 33876 6598 33928 6604
rect 33692 6452 33744 6458
rect 33692 6394 33744 6400
rect 33784 6248 33836 6254
rect 33784 6190 33836 6196
rect 33692 6112 33744 6118
rect 33692 6054 33744 6060
rect 33704 5914 33732 6054
rect 33508 5908 33560 5914
rect 33508 5850 33560 5856
rect 33692 5908 33744 5914
rect 33692 5850 33744 5856
rect 33796 5098 33824 6190
rect 33888 5914 33916 6598
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 34164 5574 34192 6802
rect 34440 6254 34468 8230
rect 34520 7336 34572 7342
rect 34624 7324 34652 9522
rect 34808 8634 34836 9522
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 34900 8090 34928 9646
rect 35164 9580 35216 9586
rect 35164 9522 35216 9528
rect 35176 8906 35204 9522
rect 35164 8900 35216 8906
rect 35164 8842 35216 8848
rect 35176 8090 35204 8842
rect 35360 8294 35388 9998
rect 35452 9654 35480 10390
rect 35636 10266 35664 10390
rect 35624 10260 35676 10266
rect 35624 10202 35676 10208
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 35636 9926 35664 9998
rect 35624 9920 35676 9926
rect 35624 9862 35676 9868
rect 35728 9738 35756 11222
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35820 9926 35848 10950
rect 35912 10130 35940 12038
rect 36176 11756 36228 11762
rect 36176 11698 36228 11704
rect 36084 11212 36136 11218
rect 36084 11154 36136 11160
rect 35900 10124 35952 10130
rect 35900 10066 35952 10072
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 35728 9710 35848 9738
rect 35440 9648 35492 9654
rect 35440 9590 35492 9596
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35728 8634 35756 8774
rect 35716 8628 35768 8634
rect 35716 8570 35768 8576
rect 35348 8288 35400 8294
rect 35348 8230 35400 8236
rect 34888 8084 34940 8090
rect 34888 8026 34940 8032
rect 35164 8084 35216 8090
rect 35164 8026 35216 8032
rect 35176 7546 35204 8026
rect 35532 7744 35584 7750
rect 35532 7686 35584 7692
rect 35544 7546 35572 7686
rect 35164 7540 35216 7546
rect 35164 7482 35216 7488
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 35072 7404 35124 7410
rect 35072 7346 35124 7352
rect 34572 7296 34652 7324
rect 34520 7278 34572 7284
rect 34532 6798 34560 7278
rect 34704 7200 34756 7206
rect 34704 7142 34756 7148
rect 34520 6792 34572 6798
rect 34520 6734 34572 6740
rect 34716 6322 34744 7142
rect 35084 6458 35112 7346
rect 35176 6458 35204 7482
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35072 6452 35124 6458
rect 35072 6394 35124 6400
rect 35164 6452 35216 6458
rect 35164 6394 35216 6400
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34440 5778 34468 6190
rect 34624 5914 34652 6190
rect 34888 6180 34940 6186
rect 34888 6122 34940 6128
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34428 5772 34480 5778
rect 34428 5714 34480 5720
rect 34152 5568 34204 5574
rect 34152 5510 34204 5516
rect 34426 5536 34482 5545
rect 34426 5471 34482 5480
rect 33784 5092 33836 5098
rect 33784 5034 33836 5040
rect 34440 4826 34468 5471
rect 34900 5030 34928 6122
rect 34888 5024 34940 5030
rect 34888 4966 34940 4972
rect 34428 4820 34480 4826
rect 34428 4762 34480 4768
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 35532 4616 35584 4622
rect 35532 4558 35584 4564
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 3126 33640 3402
rect 33416 3120 33468 3126
rect 33416 3062 33468 3068
rect 33600 3120 33652 3126
rect 33600 3062 33652 3068
rect 33888 2774 33916 4558
rect 34980 4480 35032 4486
rect 34980 4422 35032 4428
rect 34152 4072 34204 4078
rect 34152 4014 34204 4020
rect 34888 4072 34940 4078
rect 34888 4014 34940 4020
rect 34164 3738 34192 4014
rect 34336 3936 34388 3942
rect 34336 3878 34388 3884
rect 34152 3732 34204 3738
rect 34152 3674 34204 3680
rect 34348 3194 34376 3878
rect 34900 3738 34928 4014
rect 34888 3732 34940 3738
rect 34888 3674 34940 3680
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34336 3188 34388 3194
rect 34336 3130 34388 3136
rect 34716 3058 34744 3470
rect 34704 3052 34756 3058
rect 34704 2994 34756 3000
rect 34900 2774 34928 3674
rect 34992 3126 35020 4422
rect 35544 4282 35572 4558
rect 35636 4282 35664 7142
rect 35820 6254 35848 9710
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35912 9042 35940 9318
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 36096 8906 36124 11154
rect 36188 10266 36216 11698
rect 36280 11694 36308 13280
rect 36636 13262 36688 13268
rect 36544 12912 36596 12918
rect 36544 12854 36596 12860
rect 36452 12776 36504 12782
rect 36452 12718 36504 12724
rect 36464 12102 36492 12718
rect 36556 12102 36584 12854
rect 36648 12374 36676 13262
rect 36740 12986 36768 13330
rect 36728 12980 36780 12986
rect 36728 12922 36780 12928
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 36832 12434 36860 12922
rect 36924 12782 36952 14214
rect 37016 13802 37044 14214
rect 37660 13802 37688 15370
rect 37004 13796 37056 13802
rect 37004 13738 37056 13744
rect 37648 13796 37700 13802
rect 37648 13738 37700 13744
rect 37060 13628 37368 13637
rect 37060 13626 37066 13628
rect 37122 13626 37146 13628
rect 37202 13626 37226 13628
rect 37282 13626 37306 13628
rect 37362 13626 37368 13628
rect 37122 13574 37124 13626
rect 37304 13574 37306 13626
rect 37060 13572 37066 13574
rect 37122 13572 37146 13574
rect 37202 13572 37226 13574
rect 37282 13572 37306 13574
rect 37362 13572 37368 13574
rect 37060 13563 37368 13572
rect 37752 13530 37780 16510
rect 37936 16250 37964 17070
rect 38016 16992 38068 16998
rect 38016 16934 38068 16940
rect 37924 16244 37976 16250
rect 37924 16186 37976 16192
rect 38028 16114 38056 16934
rect 38016 16108 38068 16114
rect 38016 16050 38068 16056
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37844 13870 37872 14350
rect 37924 14272 37976 14278
rect 37924 14214 37976 14220
rect 37936 13938 37964 14214
rect 37924 13932 37976 13938
rect 37924 13874 37976 13880
rect 37832 13864 37884 13870
rect 37832 13806 37884 13812
rect 37740 13524 37792 13530
rect 37740 13466 37792 13472
rect 37004 13456 37056 13462
rect 37004 13398 37056 13404
rect 37016 12986 37044 13398
rect 37936 13394 37964 13874
rect 38016 13864 38068 13870
rect 38016 13806 38068 13812
rect 37924 13388 37976 13394
rect 37924 13330 37976 13336
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 37004 12980 37056 12986
rect 37004 12922 37056 12928
rect 36912 12776 36964 12782
rect 36912 12718 36964 12724
rect 36740 12406 36860 12434
rect 36636 12368 36688 12374
rect 36636 12310 36688 12316
rect 36740 12306 36768 12406
rect 36728 12300 36780 12306
rect 36728 12242 36780 12248
rect 36820 12300 36872 12306
rect 36820 12242 36872 12248
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36544 12096 36596 12102
rect 36544 12038 36596 12044
rect 36268 11688 36320 11694
rect 36268 11630 36320 11636
rect 36176 10260 36228 10266
rect 36176 10202 36228 10208
rect 36176 9716 36228 9722
rect 36176 9658 36228 9664
rect 36084 8900 36136 8906
rect 36084 8842 36136 8848
rect 36096 8634 36124 8842
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 35992 8356 36044 8362
rect 35992 8298 36044 8304
rect 35900 7812 35952 7818
rect 35900 7754 35952 7760
rect 35808 6248 35860 6254
rect 35808 6190 35860 6196
rect 35820 5914 35848 6190
rect 35808 5908 35860 5914
rect 35808 5850 35860 5856
rect 35820 5370 35848 5850
rect 35808 5364 35860 5370
rect 35808 5306 35860 5312
rect 35716 5092 35768 5098
rect 35716 5034 35768 5040
rect 35728 4826 35756 5034
rect 35808 5024 35860 5030
rect 35808 4966 35860 4972
rect 35716 4820 35768 4826
rect 35716 4762 35768 4768
rect 35716 4480 35768 4486
rect 35716 4422 35768 4428
rect 35532 4276 35584 4282
rect 35532 4218 35584 4224
rect 35624 4276 35676 4282
rect 35624 4218 35676 4224
rect 35728 3466 35756 4422
rect 35820 4282 35848 4966
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35912 3942 35940 7754
rect 36004 6322 36032 8298
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 36096 6458 36124 7822
rect 36188 7478 36216 9658
rect 36280 7834 36308 11630
rect 36464 11150 36492 12038
rect 36452 11144 36504 11150
rect 36452 11086 36504 11092
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36464 10742 36492 10950
rect 36556 10742 36584 12038
rect 36832 11218 36860 12242
rect 36924 11898 36952 12718
rect 37060 12540 37368 12549
rect 37060 12538 37066 12540
rect 37122 12538 37146 12540
rect 37202 12538 37226 12540
rect 37282 12538 37306 12540
rect 37362 12538 37368 12540
rect 37122 12486 37124 12538
rect 37304 12486 37306 12538
rect 37060 12484 37066 12486
rect 37122 12484 37146 12486
rect 37202 12484 37226 12486
rect 37282 12484 37306 12486
rect 37362 12484 37368 12486
rect 37060 12475 37368 12484
rect 37660 12238 37688 13262
rect 38028 12434 38056 13806
rect 37936 12406 38056 12434
rect 37648 12232 37700 12238
rect 37648 12174 37700 12180
rect 36912 11892 36964 11898
rect 36912 11834 36964 11840
rect 36820 11212 36872 11218
rect 36820 11154 36872 11160
rect 36728 11144 36780 11150
rect 36728 11086 36780 11092
rect 36636 11008 36688 11014
rect 36636 10950 36688 10956
rect 36452 10736 36504 10742
rect 36452 10678 36504 10684
rect 36544 10736 36596 10742
rect 36544 10678 36596 10684
rect 36360 10668 36412 10674
rect 36360 10610 36412 10616
rect 36372 9761 36400 10610
rect 36452 10260 36504 10266
rect 36452 10202 36504 10208
rect 36358 9752 36414 9761
rect 36358 9687 36414 9696
rect 36280 7806 36400 7834
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 36176 7472 36228 7478
rect 36176 7414 36228 7420
rect 36280 6730 36308 7686
rect 36372 7274 36400 7806
rect 36360 7268 36412 7274
rect 36360 7210 36412 7216
rect 36464 6866 36492 10202
rect 36648 10130 36676 10950
rect 36636 10124 36688 10130
rect 36636 10066 36688 10072
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 36556 9178 36584 9998
rect 36648 9722 36676 10066
rect 36636 9716 36688 9722
rect 36636 9658 36688 9664
rect 36740 9382 36768 11086
rect 36820 11076 36872 11082
rect 36820 11018 36872 11024
rect 36832 10606 36860 11018
rect 36924 10742 36952 11834
rect 37060 11452 37368 11461
rect 37060 11450 37066 11452
rect 37122 11450 37146 11452
rect 37202 11450 37226 11452
rect 37282 11450 37306 11452
rect 37362 11450 37368 11452
rect 37122 11398 37124 11450
rect 37304 11398 37306 11450
rect 37060 11396 37066 11398
rect 37122 11396 37146 11398
rect 37202 11396 37226 11398
rect 37282 11396 37306 11398
rect 37362 11396 37368 11398
rect 37060 11387 37368 11396
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 36912 10736 36964 10742
rect 36912 10678 36964 10684
rect 36820 10600 36872 10606
rect 36820 10542 36872 10548
rect 36832 10062 36860 10542
rect 37292 10538 37320 11086
rect 37280 10532 37332 10538
rect 37280 10474 37332 10480
rect 37648 10464 37700 10470
rect 37648 10406 37700 10412
rect 37060 10364 37368 10373
rect 37060 10362 37066 10364
rect 37122 10362 37146 10364
rect 37202 10362 37226 10364
rect 37282 10362 37306 10364
rect 37362 10362 37368 10364
rect 37122 10310 37124 10362
rect 37304 10310 37306 10362
rect 37060 10308 37066 10310
rect 37122 10308 37146 10310
rect 37202 10308 37226 10310
rect 37282 10308 37306 10310
rect 37362 10308 37368 10310
rect 37060 10299 37368 10308
rect 36820 10056 36872 10062
rect 36820 9998 36872 10004
rect 37660 9994 37688 10406
rect 37004 9988 37056 9994
rect 37004 9930 37056 9936
rect 37556 9988 37608 9994
rect 37556 9930 37608 9936
rect 37648 9988 37700 9994
rect 37648 9930 37700 9936
rect 37016 9722 37044 9930
rect 37464 9920 37516 9926
rect 37464 9862 37516 9868
rect 37004 9716 37056 9722
rect 37004 9658 37056 9664
rect 37476 9586 37504 9862
rect 37464 9580 37516 9586
rect 37464 9522 37516 9528
rect 36728 9376 36780 9382
rect 36728 9318 36780 9324
rect 37060 9276 37368 9285
rect 37060 9274 37066 9276
rect 37122 9274 37146 9276
rect 37202 9274 37226 9276
rect 37282 9274 37306 9276
rect 37362 9274 37368 9276
rect 37122 9222 37124 9274
rect 37304 9222 37306 9274
rect 37060 9220 37066 9222
rect 37122 9220 37146 9222
rect 37202 9220 37226 9222
rect 37282 9220 37306 9222
rect 37362 9220 37368 9222
rect 37060 9211 37368 9220
rect 37568 9178 37596 9930
rect 37832 9716 37884 9722
rect 37832 9658 37884 9664
rect 37648 9376 37700 9382
rect 37648 9318 37700 9324
rect 37660 9178 37688 9318
rect 36544 9172 36596 9178
rect 36544 9114 36596 9120
rect 37556 9172 37608 9178
rect 37556 9114 37608 9120
rect 37648 9172 37700 9178
rect 37648 9114 37700 9120
rect 37844 8974 37872 9658
rect 37936 9654 37964 12406
rect 38120 12306 38148 17682
rect 38200 14612 38252 14618
rect 38200 14554 38252 14560
rect 38212 13870 38240 14554
rect 38396 14346 38424 19246
rect 38672 18766 38700 19654
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 38476 18692 38528 18698
rect 38476 18634 38528 18640
rect 38488 18426 38516 18634
rect 38476 18420 38528 18426
rect 38476 18362 38528 18368
rect 38856 18290 38884 19926
rect 39040 19854 39068 21830
rect 39028 19848 39080 19854
rect 39028 19790 39080 19796
rect 39132 19802 39160 22102
rect 39224 21554 39252 22374
rect 40040 22092 40092 22098
rect 40040 22034 40092 22040
rect 39580 21888 39632 21894
rect 39580 21830 39632 21836
rect 39592 21690 39620 21830
rect 39580 21684 39632 21690
rect 39580 21626 39632 21632
rect 40052 21554 40080 22034
rect 40132 21888 40184 21894
rect 40132 21830 40184 21836
rect 39212 21548 39264 21554
rect 39212 21490 39264 21496
rect 40040 21548 40092 21554
rect 40040 21490 40092 21496
rect 40144 21486 40172 21830
rect 40420 21690 40448 23054
rect 40592 22568 40644 22574
rect 40592 22510 40644 22516
rect 42064 22568 42116 22574
rect 42064 22510 42116 22516
rect 42432 22568 42484 22574
rect 42432 22510 42484 22516
rect 40604 22234 40632 22510
rect 40776 22432 40828 22438
rect 40776 22374 40828 22380
rect 41512 22432 41564 22438
rect 41512 22374 41564 22380
rect 40592 22228 40644 22234
rect 40592 22170 40644 22176
rect 40500 22092 40552 22098
rect 40500 22034 40552 22040
rect 40408 21684 40460 21690
rect 40408 21626 40460 21632
rect 40132 21480 40184 21486
rect 40512 21434 40540 22034
rect 40788 21554 40816 22374
rect 41144 22160 41196 22166
rect 41196 22108 41460 22114
rect 41144 22102 41460 22108
rect 41156 22086 41460 22102
rect 41432 22030 41460 22086
rect 41420 22024 41472 22030
rect 41420 21966 41472 21972
rect 41524 21554 41552 22374
rect 42076 22234 42104 22510
rect 42064 22228 42116 22234
rect 42064 22170 42116 22176
rect 40776 21548 40828 21554
rect 40776 21490 40828 21496
rect 41512 21548 41564 21554
rect 41512 21490 41564 21496
rect 40132 21422 40184 21428
rect 39764 20256 39816 20262
rect 39764 20198 39816 20204
rect 39776 19922 39804 20198
rect 39764 19916 39816 19922
rect 39764 19858 39816 19864
rect 39132 19774 39252 19802
rect 38936 19712 38988 19718
rect 38936 19654 38988 19660
rect 39028 19712 39080 19718
rect 39028 19654 39080 19660
rect 39120 19712 39172 19718
rect 39120 19654 39172 19660
rect 38948 18698 38976 19654
rect 38936 18692 38988 18698
rect 38936 18634 38988 18640
rect 38948 18426 38976 18634
rect 39040 18426 39068 19654
rect 39132 19514 39160 19654
rect 39120 19508 39172 19514
rect 39120 19450 39172 19456
rect 39224 19310 39252 19774
rect 39580 19780 39632 19786
rect 39580 19722 39632 19728
rect 39592 19446 39620 19722
rect 39580 19440 39632 19446
rect 39580 19382 39632 19388
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 39224 18970 39252 19246
rect 39212 18964 39264 18970
rect 39212 18906 39264 18912
rect 39592 18426 39620 19382
rect 38936 18420 38988 18426
rect 38936 18362 38988 18368
rect 39028 18420 39080 18426
rect 39028 18362 39080 18368
rect 39580 18420 39632 18426
rect 39580 18362 39632 18368
rect 38844 18284 38896 18290
rect 38844 18226 38896 18232
rect 39776 18154 39804 19858
rect 39856 19168 39908 19174
rect 39856 19110 39908 19116
rect 39868 18630 39896 19110
rect 39948 18760 40000 18766
rect 39948 18702 40000 18708
rect 39856 18624 39908 18630
rect 39856 18566 39908 18572
rect 39868 18290 39896 18566
rect 39856 18284 39908 18290
rect 39856 18226 39908 18232
rect 39764 18148 39816 18154
rect 39764 18090 39816 18096
rect 38660 17128 38712 17134
rect 38660 17070 38712 17076
rect 38672 16522 38700 17070
rect 38660 16516 38712 16522
rect 38660 16458 38712 16464
rect 38936 16516 38988 16522
rect 38936 16458 38988 16464
rect 38948 15706 38976 16458
rect 39028 16448 39080 16454
rect 39028 16390 39080 16396
rect 39040 15910 39068 16390
rect 39028 15904 39080 15910
rect 39028 15846 39080 15852
rect 39580 15904 39632 15910
rect 39580 15846 39632 15852
rect 38936 15700 38988 15706
rect 38936 15642 38988 15648
rect 38476 15360 38528 15366
rect 38476 15302 38528 15308
rect 38384 14340 38436 14346
rect 38384 14282 38436 14288
rect 38384 14068 38436 14074
rect 38384 14010 38436 14016
rect 38200 13864 38252 13870
rect 38200 13806 38252 13812
rect 38396 12434 38424 14010
rect 38488 12764 38516 15302
rect 39040 14958 39068 15846
rect 39592 15366 39620 15846
rect 39580 15360 39632 15366
rect 39580 15302 39632 15308
rect 39028 14952 39080 14958
rect 39028 14894 39080 14900
rect 38660 14408 38712 14414
rect 38660 14350 38712 14356
rect 38568 13184 38620 13190
rect 38568 13126 38620 13132
rect 38580 12866 38608 13126
rect 38672 12986 38700 14350
rect 38752 13728 38804 13734
rect 38752 13670 38804 13676
rect 38660 12980 38712 12986
rect 38660 12922 38712 12928
rect 38580 12838 38700 12866
rect 38764 12850 38792 13670
rect 39040 13326 39068 14894
rect 39776 14074 39804 18090
rect 39960 18086 39988 18702
rect 40144 18630 40172 21422
rect 40420 21406 40540 21434
rect 42444 21418 42472 22510
rect 42536 22098 42564 23258
rect 45560 23112 45612 23118
rect 45560 23054 45612 23060
rect 42708 23044 42760 23050
rect 42708 22986 42760 22992
rect 42720 22574 42748 22986
rect 45008 22976 45060 22982
rect 45008 22918 45060 22924
rect 44282 22876 44590 22885
rect 44282 22874 44288 22876
rect 44344 22874 44368 22876
rect 44424 22874 44448 22876
rect 44504 22874 44528 22876
rect 44584 22874 44590 22876
rect 44344 22822 44346 22874
rect 44526 22822 44528 22874
rect 44282 22820 44288 22822
rect 44344 22820 44368 22822
rect 44424 22820 44448 22822
rect 44504 22820 44528 22822
rect 44584 22820 44590 22822
rect 44282 22811 44590 22820
rect 45020 22642 45048 22918
rect 45008 22636 45060 22642
rect 45008 22578 45060 22584
rect 42708 22568 42760 22574
rect 42708 22510 42760 22516
rect 43444 22568 43496 22574
rect 43444 22510 43496 22516
rect 42616 22228 42668 22234
rect 42616 22170 42668 22176
rect 42524 22092 42576 22098
rect 42524 22034 42576 22040
rect 42524 21888 42576 21894
rect 42524 21830 42576 21836
rect 42432 21412 42484 21418
rect 40420 21350 40448 21406
rect 42432 21354 42484 21360
rect 40408 21344 40460 21350
rect 40408 21286 40460 21292
rect 40776 21344 40828 21350
rect 40776 21286 40828 21292
rect 40420 21146 40448 21286
rect 40408 21140 40460 21146
rect 40408 21082 40460 21088
rect 40788 20942 40816 21286
rect 40776 20936 40828 20942
rect 40776 20878 40828 20884
rect 42536 20890 42564 21830
rect 42628 21010 42656 22170
rect 42720 22098 42748 22510
rect 42708 22092 42760 22098
rect 42708 22034 42760 22040
rect 42720 21622 42748 22034
rect 43456 22030 43484 22510
rect 43628 22432 43680 22438
rect 43628 22374 43680 22380
rect 45284 22432 45336 22438
rect 45284 22374 45336 22380
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 43456 21690 43484 21966
rect 43640 21962 43668 22374
rect 45296 22094 45324 22374
rect 45204 22066 45324 22094
rect 43628 21956 43680 21962
rect 43628 21898 43680 21904
rect 43444 21684 43496 21690
rect 43444 21626 43496 21632
rect 42708 21616 42760 21622
rect 42708 21558 42760 21564
rect 42616 21004 42668 21010
rect 42616 20946 42668 20952
rect 42536 20862 42748 20890
rect 42720 19854 42748 20862
rect 41972 19848 42024 19854
rect 41972 19790 42024 19796
rect 42708 19848 42760 19854
rect 42708 19790 42760 19796
rect 40592 19712 40644 19718
rect 40592 19654 40644 19660
rect 41420 19712 41472 19718
rect 41420 19654 41472 19660
rect 40224 19508 40276 19514
rect 40224 19450 40276 19456
rect 40236 18766 40264 19450
rect 40224 18760 40276 18766
rect 40224 18702 40276 18708
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 39948 18080 40000 18086
rect 39948 18022 40000 18028
rect 40040 17128 40092 17134
rect 40040 17070 40092 17076
rect 40052 16658 40080 17070
rect 40040 16652 40092 16658
rect 40040 16594 40092 16600
rect 39856 15496 39908 15502
rect 39856 15438 39908 15444
rect 39868 14958 39896 15438
rect 39856 14952 39908 14958
rect 39856 14894 39908 14900
rect 39868 14618 39896 14894
rect 39856 14612 39908 14618
rect 39856 14554 39908 14560
rect 39764 14068 39816 14074
rect 39764 14010 39816 14016
rect 39120 13524 39172 13530
rect 39120 13466 39172 13472
rect 39028 13320 39080 13326
rect 38948 13280 39028 13308
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 38856 12986 38884 13194
rect 38844 12980 38896 12986
rect 38844 12922 38896 12928
rect 38948 12850 38976 13280
rect 39028 13262 39080 13268
rect 38488 12736 38608 12764
rect 38304 12406 38424 12434
rect 38108 12300 38160 12306
rect 38108 12242 38160 12248
rect 38120 11898 38148 12242
rect 38108 11892 38160 11898
rect 38108 11834 38160 11840
rect 38200 11008 38252 11014
rect 38200 10950 38252 10956
rect 38212 10742 38240 10950
rect 38200 10736 38252 10742
rect 38200 10678 38252 10684
rect 37924 9648 37976 9654
rect 37924 9590 37976 9596
rect 37936 9178 37964 9590
rect 38016 9580 38068 9586
rect 38016 9522 38068 9528
rect 38028 9178 38056 9522
rect 37924 9172 37976 9178
rect 37924 9114 37976 9120
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 36636 8424 36688 8430
rect 36636 8366 36688 8372
rect 36648 7546 36676 8366
rect 37464 8288 37516 8294
rect 37464 8230 37516 8236
rect 37060 8188 37368 8197
rect 37060 8186 37066 8188
rect 37122 8186 37146 8188
rect 37202 8186 37226 8188
rect 37282 8186 37306 8188
rect 37362 8186 37368 8188
rect 37122 8134 37124 8186
rect 37304 8134 37306 8186
rect 37060 8132 37066 8134
rect 37122 8132 37146 8134
rect 37202 8132 37226 8134
rect 37282 8132 37306 8134
rect 37362 8132 37368 8134
rect 37060 8123 37368 8132
rect 36820 7880 36872 7886
rect 36820 7822 36872 7828
rect 36728 7744 36780 7750
rect 36728 7686 36780 7692
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36452 6860 36504 6866
rect 36452 6802 36504 6808
rect 36268 6724 36320 6730
rect 36268 6666 36320 6672
rect 36740 6662 36768 7686
rect 36832 7002 36860 7822
rect 37060 7100 37368 7109
rect 37060 7098 37066 7100
rect 37122 7098 37146 7100
rect 37202 7098 37226 7100
rect 37282 7098 37306 7100
rect 37362 7098 37368 7100
rect 37122 7046 37124 7098
rect 37304 7046 37306 7098
rect 37060 7044 37066 7046
rect 37122 7044 37146 7046
rect 37202 7044 37226 7046
rect 37282 7044 37306 7046
rect 37362 7044 37368 7046
rect 37060 7035 37368 7044
rect 36820 6996 36872 7002
rect 36820 6938 36872 6944
rect 36820 6860 36872 6866
rect 36820 6802 36872 6808
rect 36832 6662 36860 6802
rect 36544 6656 36596 6662
rect 36544 6598 36596 6604
rect 36728 6656 36780 6662
rect 36728 6598 36780 6604
rect 36820 6656 36872 6662
rect 36820 6598 36872 6604
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36556 6390 36584 6598
rect 36544 6384 36596 6390
rect 36544 6326 36596 6332
rect 36740 6322 36768 6598
rect 36832 6458 36860 6598
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 36728 6316 36780 6322
rect 36728 6258 36780 6264
rect 36832 5642 36860 6394
rect 37476 6225 37504 8230
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 37568 6730 37596 7822
rect 37648 7404 37700 7410
rect 37648 7346 37700 7352
rect 37660 6798 37688 7346
rect 38120 7002 38148 7822
rect 38108 6996 38160 7002
rect 38108 6938 38160 6944
rect 38200 6996 38252 7002
rect 38200 6938 38252 6944
rect 37648 6792 37700 6798
rect 38212 6746 38240 6938
rect 37648 6734 37700 6740
rect 37556 6724 37608 6730
rect 37556 6666 37608 6672
rect 37462 6216 37518 6225
rect 37462 6151 37518 6160
rect 37476 6118 37504 6151
rect 37464 6112 37516 6118
rect 37464 6054 37516 6060
rect 37060 6012 37368 6021
rect 37060 6010 37066 6012
rect 37122 6010 37146 6012
rect 37202 6010 37226 6012
rect 37282 6010 37306 6012
rect 37362 6010 37368 6012
rect 37122 5958 37124 6010
rect 37304 5958 37306 6010
rect 37060 5956 37066 5958
rect 37122 5956 37146 5958
rect 37202 5956 37226 5958
rect 37282 5956 37306 5958
rect 37362 5956 37368 5958
rect 37060 5947 37368 5956
rect 36820 5636 36872 5642
rect 36820 5578 36872 5584
rect 37660 5574 37688 6734
rect 38028 6730 38240 6746
rect 38016 6724 38240 6730
rect 38068 6718 38240 6724
rect 38016 6666 38068 6672
rect 38108 6656 38160 6662
rect 38108 6598 38160 6604
rect 37832 6248 37884 6254
rect 37832 6190 37884 6196
rect 37844 5914 37872 6190
rect 38016 6180 38068 6186
rect 38016 6122 38068 6128
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 37740 5772 37792 5778
rect 37740 5714 37792 5720
rect 36912 5568 36964 5574
rect 36912 5510 36964 5516
rect 37648 5568 37700 5574
rect 37648 5510 37700 5516
rect 36924 5370 36952 5510
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 35992 5160 36044 5166
rect 35992 5102 36044 5108
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 35716 3460 35768 3466
rect 35716 3402 35768 3408
rect 36004 3194 36032 5102
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 36268 4616 36320 4622
rect 36268 4558 36320 4564
rect 36176 4548 36228 4554
rect 36176 4490 36228 4496
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 34980 3120 35032 3126
rect 34980 3062 35032 3068
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 33888 2746 34100 2774
rect 34072 2650 34100 2746
rect 34808 2746 34928 2774
rect 34060 2644 34112 2650
rect 34060 2586 34112 2592
rect 34060 2508 34112 2514
rect 34060 2450 34112 2456
rect 31208 2440 31260 2446
rect 30392 2378 30512 2394
rect 31208 2382 31260 2388
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 29368 2372 29420 2378
rect 29368 2314 29420 2320
rect 30392 2372 30524 2378
rect 30392 2366 30472 2372
rect 29380 1306 29408 2314
rect 29838 2204 30146 2213
rect 29838 2202 29844 2204
rect 29900 2202 29924 2204
rect 29980 2202 30004 2204
rect 30060 2202 30084 2204
rect 30140 2202 30146 2204
rect 29900 2150 29902 2202
rect 30082 2150 30084 2202
rect 29838 2148 29844 2150
rect 29900 2148 29924 2150
rect 29980 2148 30004 2150
rect 30060 2148 30084 2150
rect 30140 2148 30146 2150
rect 29838 2139 30146 2148
rect 29380 1278 29592 1306
rect 29564 800 29592 1278
rect 30392 800 30420 2366
rect 30472 2314 30524 2320
rect 31220 800 31248 2382
rect 32036 2372 32088 2378
rect 32036 2314 32088 2320
rect 32956 2372 33008 2378
rect 32956 2314 33008 2320
rect 32048 800 32076 2314
rect 32968 1306 32996 2314
rect 32876 1278 32996 1306
rect 32876 800 32904 1278
rect 33704 870 33824 898
rect 33704 800 33732 870
rect 23860 734 24072 762
rect 24582 0 24638 800
rect 25410 0 25466 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 33796 762 33824 870
rect 34072 762 34100 2450
rect 34808 2446 34836 2746
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 34532 870 34652 898
rect 34532 800 34560 870
rect 33796 734 34100 762
rect 34518 0 34574 800
rect 34624 762 34652 870
rect 34900 762 34928 2382
rect 35360 800 35388 3062
rect 36004 2922 36032 3130
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 36188 2650 36216 4490
rect 36280 4282 36308 4558
rect 36648 4486 36676 4966
rect 36924 4690 36952 5306
rect 37060 4924 37368 4933
rect 37060 4922 37066 4924
rect 37122 4922 37146 4924
rect 37202 4922 37226 4924
rect 37282 4922 37306 4924
rect 37362 4922 37368 4924
rect 37122 4870 37124 4922
rect 37304 4870 37306 4922
rect 37060 4868 37066 4870
rect 37122 4868 37146 4870
rect 37202 4868 37226 4870
rect 37282 4868 37306 4870
rect 37362 4868 37368 4870
rect 37060 4859 37368 4868
rect 36912 4684 36964 4690
rect 36912 4626 36964 4632
rect 36636 4480 36688 4486
rect 36636 4422 36688 4428
rect 36268 4276 36320 4282
rect 36268 4218 36320 4224
rect 36648 4078 36676 4422
rect 36912 4140 36964 4146
rect 36912 4082 36964 4088
rect 36360 4072 36412 4078
rect 36360 4014 36412 4020
rect 36636 4072 36688 4078
rect 36636 4014 36688 4020
rect 36372 3194 36400 4014
rect 36820 3392 36872 3398
rect 36820 3334 36872 3340
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 36832 3058 36860 3334
rect 36924 3194 36952 4082
rect 37660 3942 37688 5510
rect 37752 5302 37780 5714
rect 37740 5296 37792 5302
rect 37740 5238 37792 5244
rect 37740 5024 37792 5030
rect 37740 4966 37792 4972
rect 37752 4214 37780 4966
rect 38028 4554 38056 6122
rect 38120 5574 38148 6598
rect 38198 6216 38254 6225
rect 38198 6151 38200 6160
rect 38252 6151 38254 6160
rect 38200 6122 38252 6128
rect 38108 5568 38160 5574
rect 38108 5510 38160 5516
rect 38016 4548 38068 4554
rect 38016 4490 38068 4496
rect 37740 4208 37792 4214
rect 37740 4150 37792 4156
rect 38028 3942 38056 4490
rect 38120 4486 38148 5510
rect 38304 5250 38332 12406
rect 38476 9920 38528 9926
rect 38476 9862 38528 9868
rect 38488 9042 38516 9862
rect 38580 9518 38608 12736
rect 38672 12306 38700 12838
rect 38752 12844 38804 12850
rect 38752 12786 38804 12792
rect 38936 12844 38988 12850
rect 38936 12786 38988 12792
rect 38660 12300 38712 12306
rect 38660 12242 38712 12248
rect 38948 12102 38976 12786
rect 39132 12102 39160 13466
rect 39672 13252 39724 13258
rect 39672 13194 39724 13200
rect 39684 12986 39712 13194
rect 39672 12980 39724 12986
rect 39672 12922 39724 12928
rect 39304 12776 39356 12782
rect 39304 12718 39356 12724
rect 39316 12374 39344 12718
rect 39304 12368 39356 12374
rect 39304 12310 39356 12316
rect 39948 12232 40000 12238
rect 39948 12174 40000 12180
rect 38936 12096 38988 12102
rect 38936 12038 38988 12044
rect 39120 12096 39172 12102
rect 39120 12038 39172 12044
rect 38948 11626 38976 12038
rect 39960 11898 39988 12174
rect 39120 11892 39172 11898
rect 39120 11834 39172 11840
rect 39948 11892 40000 11898
rect 39948 11834 40000 11840
rect 38936 11620 38988 11626
rect 38936 11562 38988 11568
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38764 10266 38792 11086
rect 38948 10674 38976 11562
rect 39028 11008 39080 11014
rect 39028 10950 39080 10956
rect 38936 10668 38988 10674
rect 38936 10610 38988 10616
rect 38752 10260 38804 10266
rect 38752 10202 38804 10208
rect 39040 10130 39068 10950
rect 39132 10606 39160 11834
rect 40040 11552 40092 11558
rect 40040 11494 40092 11500
rect 40052 11257 40080 11494
rect 40144 11354 40172 18566
rect 40224 17128 40276 17134
rect 40224 17070 40276 17076
rect 40236 15910 40264 17070
rect 40316 17060 40368 17066
rect 40316 17002 40368 17008
rect 40224 15904 40276 15910
rect 40224 15846 40276 15852
rect 40132 11348 40184 11354
rect 40132 11290 40184 11296
rect 40038 11248 40094 11257
rect 40038 11183 40094 11192
rect 39580 11144 39632 11150
rect 39580 11086 39632 11092
rect 40132 11144 40184 11150
rect 40132 11086 40184 11092
rect 39304 10668 39356 10674
rect 39304 10610 39356 10616
rect 39120 10600 39172 10606
rect 39120 10542 39172 10548
rect 39028 10124 39080 10130
rect 39028 10066 39080 10072
rect 39132 9926 39160 10542
rect 39212 10124 39264 10130
rect 39212 10066 39264 10072
rect 38660 9920 38712 9926
rect 38660 9862 38712 9868
rect 39120 9920 39172 9926
rect 39120 9862 39172 9868
rect 38672 9654 38700 9862
rect 38660 9648 38712 9654
rect 38660 9590 38712 9596
rect 38568 9512 38620 9518
rect 38568 9454 38620 9460
rect 38580 9042 38608 9454
rect 38476 9036 38528 9042
rect 38476 8978 38528 8984
rect 38568 9036 38620 9042
rect 38568 8978 38620 8984
rect 38384 8900 38436 8906
rect 38384 8842 38436 8848
rect 38396 8294 38424 8842
rect 38384 8288 38436 8294
rect 38384 8230 38436 8236
rect 38568 6724 38620 6730
rect 38568 6666 38620 6672
rect 38384 6112 38436 6118
rect 38384 6054 38436 6060
rect 38396 5914 38424 6054
rect 38580 5930 38608 6666
rect 38672 6662 38700 9590
rect 39224 9178 39252 10066
rect 39316 9722 39344 10610
rect 39592 10470 39620 11086
rect 40144 10470 40172 11086
rect 39580 10464 39632 10470
rect 39580 10406 39632 10412
rect 40132 10464 40184 10470
rect 40132 10406 40184 10412
rect 39304 9716 39356 9722
rect 39304 9658 39356 9664
rect 39592 9586 39620 10406
rect 39304 9580 39356 9586
rect 39304 9522 39356 9528
rect 39580 9580 39632 9586
rect 39580 9522 39632 9528
rect 39316 9466 39344 9522
rect 39316 9438 39436 9466
rect 39304 9376 39356 9382
rect 39304 9318 39356 9324
rect 39212 9172 39264 9178
rect 39212 9114 39264 9120
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38844 7744 38896 7750
rect 38844 7686 38896 7692
rect 38764 6866 38792 7686
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38764 6458 38792 6802
rect 38752 6452 38804 6458
rect 38752 6394 38804 6400
rect 38752 6248 38804 6254
rect 38752 6190 38804 6196
rect 38580 5914 38654 5930
rect 38384 5908 38436 5914
rect 38580 5908 38666 5914
rect 38580 5902 38614 5908
rect 38384 5850 38436 5856
rect 38614 5850 38666 5856
rect 38212 5222 38332 5250
rect 38108 4480 38160 4486
rect 38108 4422 38160 4428
rect 38212 4282 38240 5222
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 38304 4826 38332 5102
rect 38568 5024 38620 5030
rect 38568 4966 38620 4972
rect 38292 4820 38344 4826
rect 38292 4762 38344 4768
rect 38200 4276 38252 4282
rect 38200 4218 38252 4224
rect 37648 3936 37700 3942
rect 38016 3936 38068 3942
rect 37700 3896 37780 3924
rect 37648 3878 37700 3884
rect 37060 3836 37368 3845
rect 37060 3834 37066 3836
rect 37122 3834 37146 3836
rect 37202 3834 37226 3836
rect 37282 3834 37306 3836
rect 37362 3834 37368 3836
rect 37122 3782 37124 3834
rect 37304 3782 37306 3834
rect 37060 3780 37066 3782
rect 37122 3780 37146 3782
rect 37202 3780 37226 3782
rect 37282 3780 37306 3782
rect 37362 3780 37368 3782
rect 37060 3771 37368 3780
rect 37752 3534 37780 3896
rect 38016 3878 38068 3884
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 37096 3460 37148 3466
rect 37096 3402 37148 3408
rect 36912 3188 36964 3194
rect 36912 3130 36964 3136
rect 37108 3126 37136 3402
rect 37752 3126 37780 3470
rect 37096 3120 37148 3126
rect 37096 3062 37148 3068
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 38580 3058 38608 4966
rect 38764 4826 38792 6190
rect 38856 6118 38884 7686
rect 39120 7336 39172 7342
rect 39120 7278 39172 7284
rect 38936 7200 38988 7206
rect 38936 7142 38988 7148
rect 38948 6798 38976 7142
rect 38936 6792 38988 6798
rect 38936 6734 38988 6740
rect 39028 6248 39080 6254
rect 39028 6190 39080 6196
rect 38844 6112 38896 6118
rect 38844 6054 38896 6060
rect 38856 5642 38884 6054
rect 39040 5778 39068 6190
rect 39132 5914 39160 7278
rect 39316 6458 39344 9318
rect 39408 8498 39436 9438
rect 39488 9376 39540 9382
rect 39488 9318 39540 9324
rect 39500 8974 39528 9318
rect 39488 8968 39540 8974
rect 39488 8910 39540 8916
rect 39396 8492 39448 8498
rect 39396 8434 39448 8440
rect 39396 7880 39448 7886
rect 39396 7822 39448 7828
rect 39408 7546 39436 7822
rect 39396 7540 39448 7546
rect 39396 7482 39448 7488
rect 39856 6792 39908 6798
rect 39856 6734 39908 6740
rect 39396 6656 39448 6662
rect 39396 6598 39448 6604
rect 39304 6452 39356 6458
rect 39304 6394 39356 6400
rect 39120 5908 39172 5914
rect 39120 5850 39172 5856
rect 39028 5772 39080 5778
rect 39028 5714 39080 5720
rect 39408 5710 39436 6598
rect 39868 6254 39896 6734
rect 39856 6248 39908 6254
rect 39856 6190 39908 6196
rect 39580 6112 39632 6118
rect 39580 6054 39632 6060
rect 39396 5704 39448 5710
rect 39396 5646 39448 5652
rect 38844 5636 38896 5642
rect 38844 5578 38896 5584
rect 39396 5568 39448 5574
rect 39396 5510 39448 5516
rect 38844 5024 38896 5030
rect 38844 4966 38896 4972
rect 39304 5024 39356 5030
rect 39304 4966 39356 4972
rect 38856 4826 38884 4966
rect 38752 4820 38804 4826
rect 38752 4762 38804 4768
rect 38844 4820 38896 4826
rect 38844 4762 38896 4768
rect 38660 4616 38712 4622
rect 38660 4558 38712 4564
rect 38672 4282 38700 4558
rect 39316 4282 39344 4966
rect 38660 4276 38712 4282
rect 38660 4218 38712 4224
rect 39304 4276 39356 4282
rect 39304 4218 39356 4224
rect 39028 4072 39080 4078
rect 39028 4014 39080 4020
rect 39040 3738 39068 4014
rect 39408 3738 39436 5510
rect 39488 5160 39540 5166
rect 39488 5102 39540 5108
rect 39500 4282 39528 5102
rect 39592 4282 39620 6054
rect 39868 5846 39896 6190
rect 39856 5840 39908 5846
rect 39856 5782 39908 5788
rect 39672 5160 39724 5166
rect 39672 5102 39724 5108
rect 39488 4276 39540 4282
rect 39488 4218 39540 4224
rect 39580 4276 39632 4282
rect 39580 4218 39632 4224
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39592 3738 39620 3878
rect 39028 3732 39080 3738
rect 39028 3674 39080 3680
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39120 3528 39172 3534
rect 39120 3470 39172 3476
rect 36820 3052 36872 3058
rect 36820 2994 36872 3000
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 36360 2984 36412 2990
rect 36360 2926 36412 2932
rect 36176 2644 36228 2650
rect 36176 2586 36228 2592
rect 36372 1578 36400 2926
rect 36820 2916 36872 2922
rect 36820 2858 36872 2864
rect 36832 2446 36860 2858
rect 37060 2748 37368 2757
rect 37060 2746 37066 2748
rect 37122 2746 37146 2748
rect 37202 2746 37226 2748
rect 37282 2746 37306 2748
rect 37362 2746 37368 2748
rect 37122 2694 37124 2746
rect 37304 2694 37306 2746
rect 37060 2692 37066 2694
rect 37122 2692 37146 2694
rect 37202 2692 37226 2694
rect 37282 2692 37306 2694
rect 37362 2692 37368 2694
rect 37060 2683 37368 2692
rect 39132 2650 39160 3470
rect 39684 3194 39712 5102
rect 40040 5024 40092 5030
rect 40040 4966 40092 4972
rect 40052 4690 40080 4966
rect 40132 4752 40184 4758
rect 40132 4694 40184 4700
rect 40040 4684 40092 4690
rect 40040 4626 40092 4632
rect 40144 4146 40172 4694
rect 39764 4140 39816 4146
rect 39764 4082 39816 4088
rect 40132 4140 40184 4146
rect 40132 4082 40184 4088
rect 39776 3602 39804 4082
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 39868 3194 39896 3470
rect 39672 3188 39724 3194
rect 39672 3130 39724 3136
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 37016 2514 37228 2530
rect 37016 2508 37240 2514
rect 37016 2502 37188 2508
rect 36820 2440 36872 2446
rect 36820 2382 36872 2388
rect 36188 1550 36400 1578
rect 36188 800 36216 1550
rect 37016 800 37044 2502
rect 37188 2450 37240 2456
rect 39028 2508 39080 2514
rect 39028 2450 39080 2456
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 37936 1306 37964 2382
rect 37844 1278 37964 1306
rect 37844 800 37872 1278
rect 38672 870 38792 898
rect 38672 800 38700 870
rect 34624 734 34928 762
rect 35346 0 35402 800
rect 36174 0 36230 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 38764 762 38792 870
rect 39040 762 39068 2450
rect 39500 800 39528 2926
rect 39684 2446 39712 3130
rect 40236 2446 40264 15846
rect 40328 14074 40356 17002
rect 40604 16590 40632 19654
rect 40960 19304 41012 19310
rect 40960 19246 41012 19252
rect 40972 18970 41000 19246
rect 41052 19168 41104 19174
rect 41052 19110 41104 19116
rect 40960 18964 41012 18970
rect 40960 18906 41012 18912
rect 41064 18834 41092 19110
rect 41052 18828 41104 18834
rect 41052 18770 41104 18776
rect 41432 18358 41460 19654
rect 41880 19168 41932 19174
rect 41880 19110 41932 19116
rect 41892 18834 41920 19110
rect 41984 18970 42012 19790
rect 42432 19304 42484 19310
rect 42432 19246 42484 19252
rect 41972 18964 42024 18970
rect 41972 18906 42024 18912
rect 41880 18828 41932 18834
rect 41880 18770 41932 18776
rect 41420 18352 41472 18358
rect 41420 18294 41472 18300
rect 40868 18284 40920 18290
rect 40868 18226 40920 18232
rect 40880 17882 40908 18226
rect 40868 17876 40920 17882
rect 40868 17818 40920 17824
rect 41144 17604 41196 17610
rect 41144 17546 41196 17552
rect 40684 16992 40736 16998
rect 40684 16934 40736 16940
rect 40696 16794 40724 16934
rect 40684 16788 40736 16794
rect 40684 16730 40736 16736
rect 40592 16584 40644 16590
rect 40592 16526 40644 16532
rect 40684 16448 40736 16454
rect 40684 16390 40736 16396
rect 40696 16250 40724 16390
rect 40684 16244 40736 16250
rect 40684 16186 40736 16192
rect 40776 15428 40828 15434
rect 40776 15370 40828 15376
rect 40788 15162 40816 15370
rect 40776 15156 40828 15162
rect 40776 15098 40828 15104
rect 40316 14068 40368 14074
rect 40316 14010 40368 14016
rect 41052 13864 41104 13870
rect 41052 13806 41104 13812
rect 41064 12986 41092 13806
rect 41156 13530 41184 17546
rect 41420 16652 41472 16658
rect 41420 16594 41472 16600
rect 41236 15904 41288 15910
rect 41236 15846 41288 15852
rect 41248 15094 41276 15846
rect 41236 15088 41288 15094
rect 41236 15030 41288 15036
rect 41432 14890 41460 16594
rect 41604 16040 41656 16046
rect 41604 15982 41656 15988
rect 41616 15502 41644 15982
rect 41604 15496 41656 15502
rect 41604 15438 41656 15444
rect 41512 14952 41564 14958
rect 41512 14894 41564 14900
rect 41696 14952 41748 14958
rect 41696 14894 41748 14900
rect 41420 14884 41472 14890
rect 41420 14826 41472 14832
rect 41524 14482 41552 14894
rect 41512 14476 41564 14482
rect 41512 14418 41564 14424
rect 41708 14346 41736 14894
rect 41696 14340 41748 14346
rect 41696 14282 41748 14288
rect 41788 14340 41840 14346
rect 41788 14282 41840 14288
rect 41604 13864 41656 13870
rect 41524 13824 41604 13852
rect 41144 13524 41196 13530
rect 41144 13466 41196 13472
rect 41052 12980 41104 12986
rect 41052 12922 41104 12928
rect 41156 12850 41184 13466
rect 41328 13252 41380 13258
rect 41328 13194 41380 13200
rect 40684 12844 40736 12850
rect 40684 12786 40736 12792
rect 41144 12844 41196 12850
rect 41144 12786 41196 12792
rect 40696 12434 40724 12786
rect 40696 12406 40908 12434
rect 40408 11076 40460 11082
rect 40408 11018 40460 11024
rect 40420 3738 40448 11018
rect 40500 10804 40552 10810
rect 40500 10746 40552 10752
rect 40512 9518 40540 10746
rect 40880 9625 40908 12406
rect 41340 12374 41368 13194
rect 41420 12776 41472 12782
rect 41420 12718 41472 12724
rect 41328 12368 41380 12374
rect 41328 12310 41380 12316
rect 40960 12164 41012 12170
rect 40960 12106 41012 12112
rect 40972 11830 41000 12106
rect 40960 11824 41012 11830
rect 40960 11766 41012 11772
rect 41432 11626 41460 12718
rect 41524 12306 41552 13824
rect 41604 13806 41656 13812
rect 41708 13530 41736 14282
rect 41696 13524 41748 13530
rect 41696 13466 41748 13472
rect 41800 13410 41828 14282
rect 41616 13382 41828 13410
rect 41616 12374 41644 13382
rect 41696 13184 41748 13190
rect 41696 13126 41748 13132
rect 41604 12368 41656 12374
rect 41604 12310 41656 12316
rect 41512 12300 41564 12306
rect 41512 12242 41564 12248
rect 41524 11762 41552 12242
rect 41708 11762 41736 13126
rect 41892 12753 41920 18770
rect 42444 18426 42472 19246
rect 42524 18964 42576 18970
rect 42524 18906 42576 18912
rect 42432 18420 42484 18426
rect 42432 18362 42484 18368
rect 42536 18222 42564 18906
rect 42616 18624 42668 18630
rect 42720 18578 42748 19790
rect 43456 19310 43484 21626
rect 43640 21554 43668 21898
rect 43812 21888 43864 21894
rect 43812 21830 43864 21836
rect 43824 21554 43852 21830
rect 44282 21788 44590 21797
rect 44282 21786 44288 21788
rect 44344 21786 44368 21788
rect 44424 21786 44448 21788
rect 44504 21786 44528 21788
rect 44584 21786 44590 21788
rect 44344 21734 44346 21786
rect 44526 21734 44528 21786
rect 44282 21732 44288 21734
rect 44344 21732 44368 21734
rect 44424 21732 44448 21734
rect 44504 21732 44528 21734
rect 44584 21732 44590 21734
rect 44282 21723 44590 21732
rect 45204 21690 45232 22066
rect 45284 21888 45336 21894
rect 45284 21830 45336 21836
rect 45376 21888 45428 21894
rect 45376 21830 45428 21836
rect 45468 21888 45520 21894
rect 45468 21830 45520 21836
rect 45192 21684 45244 21690
rect 45192 21626 45244 21632
rect 45296 21622 45324 21830
rect 45284 21616 45336 21622
rect 45284 21558 45336 21564
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 43812 21548 43864 21554
rect 43812 21490 43864 21496
rect 43824 21146 43852 21490
rect 45388 21486 45416 21830
rect 45480 21570 45508 21830
rect 45572 21690 45600 23054
rect 46204 22976 46256 22982
rect 46204 22918 46256 22924
rect 46216 22778 46244 22918
rect 47596 22778 47624 23598
rect 48136 23520 48188 23526
rect 48136 23462 48188 23468
rect 48228 23520 48280 23526
rect 48228 23462 48280 23468
rect 49332 23520 49384 23526
rect 49332 23462 49384 23468
rect 52736 23520 52788 23526
rect 52736 23462 52788 23468
rect 48148 23186 48176 23462
rect 48136 23180 48188 23186
rect 48136 23122 48188 23128
rect 48044 22976 48096 22982
rect 48044 22918 48096 22924
rect 46204 22772 46256 22778
rect 46204 22714 46256 22720
rect 47584 22772 47636 22778
rect 47584 22714 47636 22720
rect 48056 22658 48084 22918
rect 48148 22778 48176 23122
rect 48240 22982 48268 23462
rect 48596 23248 48648 23254
rect 48596 23190 48648 23196
rect 48228 22976 48280 22982
rect 48228 22918 48280 22924
rect 48136 22772 48188 22778
rect 48136 22714 48188 22720
rect 48056 22630 48176 22658
rect 46664 22432 46716 22438
rect 46664 22374 46716 22380
rect 47952 22432 48004 22438
rect 47952 22374 48004 22380
rect 46572 22160 46624 22166
rect 46572 22102 46624 22108
rect 45560 21684 45612 21690
rect 45560 21626 45612 21632
rect 45480 21554 45600 21570
rect 45480 21548 45612 21554
rect 45480 21542 45560 21548
rect 45560 21490 45612 21496
rect 44824 21480 44876 21486
rect 44824 21422 44876 21428
rect 44916 21480 44968 21486
rect 44916 21422 44968 21428
rect 45008 21480 45060 21486
rect 45008 21422 45060 21428
rect 45376 21480 45428 21486
rect 45376 21422 45428 21428
rect 44732 21344 44784 21350
rect 44732 21286 44784 21292
rect 43812 21140 43864 21146
rect 43812 21082 43864 21088
rect 44282 20700 44590 20709
rect 44282 20698 44288 20700
rect 44344 20698 44368 20700
rect 44424 20698 44448 20700
rect 44504 20698 44528 20700
rect 44584 20698 44590 20700
rect 44344 20646 44346 20698
rect 44526 20646 44528 20698
rect 44282 20644 44288 20646
rect 44344 20644 44368 20646
rect 44424 20644 44448 20646
rect 44504 20644 44528 20646
rect 44584 20644 44590 20646
rect 44282 20635 44590 20644
rect 44640 20528 44692 20534
rect 44640 20470 44692 20476
rect 44548 20256 44600 20262
rect 44548 20198 44600 20204
rect 44560 19922 44588 20198
rect 44652 19922 44680 20470
rect 44548 19916 44600 19922
rect 44548 19858 44600 19864
rect 44640 19916 44692 19922
rect 44640 19858 44692 19864
rect 44180 19712 44232 19718
rect 44180 19654 44232 19660
rect 44640 19712 44692 19718
rect 44640 19654 44692 19660
rect 44192 19310 44220 19654
rect 44282 19612 44590 19621
rect 44282 19610 44288 19612
rect 44344 19610 44368 19612
rect 44424 19610 44448 19612
rect 44504 19610 44528 19612
rect 44584 19610 44590 19612
rect 44344 19558 44346 19610
rect 44526 19558 44528 19610
rect 44282 19556 44288 19558
rect 44344 19556 44368 19558
rect 44424 19556 44448 19558
rect 44504 19556 44528 19558
rect 44584 19556 44590 19558
rect 44282 19547 44590 19556
rect 43444 19304 43496 19310
rect 43444 19246 43496 19252
rect 44180 19304 44232 19310
rect 44180 19246 44232 19252
rect 42892 19168 42944 19174
rect 42892 19110 42944 19116
rect 43260 19168 43312 19174
rect 43260 19110 43312 19116
rect 42904 18873 42932 19110
rect 42890 18864 42946 18873
rect 42890 18799 42946 18808
rect 42904 18766 42932 18799
rect 42892 18760 42944 18766
rect 42892 18702 42944 18708
rect 42668 18572 42748 18578
rect 42616 18566 42748 18572
rect 42628 18550 42748 18566
rect 42720 18358 42748 18550
rect 42708 18352 42760 18358
rect 42708 18294 42760 18300
rect 42524 18216 42576 18222
rect 42524 18158 42576 18164
rect 42156 16584 42208 16590
rect 42156 16526 42208 16532
rect 41972 16040 42024 16046
rect 41972 15982 42024 15988
rect 41984 15570 42012 15982
rect 42168 15910 42196 16526
rect 42340 16448 42392 16454
rect 42340 16390 42392 16396
rect 42352 15978 42380 16390
rect 42340 15972 42392 15978
rect 42340 15914 42392 15920
rect 42156 15904 42208 15910
rect 42156 15846 42208 15852
rect 42168 15570 42196 15846
rect 41972 15564 42024 15570
rect 41972 15506 42024 15512
rect 42156 15564 42208 15570
rect 42156 15506 42208 15512
rect 42064 15496 42116 15502
rect 42064 15438 42116 15444
rect 41972 15360 42024 15366
rect 41972 15302 42024 15308
rect 41984 15026 42012 15302
rect 41972 15020 42024 15026
rect 41972 14962 42024 14968
rect 42076 14090 42104 15438
rect 42168 14618 42196 15506
rect 42248 14884 42300 14890
rect 42248 14826 42300 14832
rect 42156 14612 42208 14618
rect 42156 14554 42208 14560
rect 42260 14482 42288 14826
rect 42352 14498 42380 15914
rect 42536 15706 42564 18158
rect 42524 15700 42576 15706
rect 42524 15642 42576 15648
rect 42432 14816 42484 14822
rect 42432 14758 42484 14764
rect 42444 14618 42472 14758
rect 42432 14612 42484 14618
rect 42432 14554 42484 14560
rect 42616 14612 42668 14618
rect 42616 14554 42668 14560
rect 42524 14544 42576 14550
rect 42248 14476 42300 14482
rect 42352 14470 42472 14498
rect 42524 14486 42576 14492
rect 42248 14418 42300 14424
rect 41984 14062 42104 14090
rect 42156 14068 42208 14074
rect 41984 13258 42012 14062
rect 42156 14010 42208 14016
rect 42064 13524 42116 13530
rect 42064 13466 42116 13472
rect 41972 13252 42024 13258
rect 41972 13194 42024 13200
rect 42076 12968 42104 13466
rect 42168 13394 42196 14010
rect 42260 13870 42288 14418
rect 42340 14272 42392 14278
rect 42340 14214 42392 14220
rect 42248 13864 42300 13870
rect 42352 13841 42380 14214
rect 42248 13806 42300 13812
rect 42338 13832 42394 13841
rect 42338 13767 42394 13776
rect 42444 13716 42472 14470
rect 42536 14074 42564 14486
rect 42524 14068 42576 14074
rect 42524 14010 42576 14016
rect 42524 13864 42576 13870
rect 42524 13806 42576 13812
rect 42260 13688 42472 13716
rect 42156 13388 42208 13394
rect 42156 13330 42208 13336
rect 41984 12940 42104 12968
rect 41878 12744 41934 12753
rect 41878 12679 41934 12688
rect 41984 12220 42012 12940
rect 42260 12900 42288 13688
rect 42536 13512 42564 13806
rect 42444 13484 42564 13512
rect 42340 13184 42392 13190
rect 42340 13126 42392 13132
rect 42168 12872 42288 12900
rect 42064 12232 42116 12238
rect 41984 12192 42064 12220
rect 42064 12174 42116 12180
rect 42076 11830 42104 12174
rect 42064 11824 42116 11830
rect 42064 11766 42116 11772
rect 41512 11756 41564 11762
rect 41512 11698 41564 11704
rect 41696 11756 41748 11762
rect 41696 11698 41748 11704
rect 42168 11676 42196 12872
rect 42352 12306 42380 13126
rect 42444 12646 42472 13484
rect 42628 13394 42656 14554
rect 42720 14090 42748 18294
rect 42800 18148 42852 18154
rect 42800 18090 42852 18096
rect 42812 17338 42840 18090
rect 43168 18080 43220 18086
rect 43168 18022 43220 18028
rect 43180 17746 43208 18022
rect 43168 17740 43220 17746
rect 43168 17682 43220 17688
rect 42800 17332 42852 17338
rect 42800 17274 42852 17280
rect 43168 16448 43220 16454
rect 43168 16390 43220 16396
rect 43180 16114 43208 16390
rect 43168 16108 43220 16114
rect 43168 16050 43220 16056
rect 42800 16040 42852 16046
rect 42800 15982 42852 15988
rect 42812 15366 42840 15982
rect 42800 15360 42852 15366
rect 42800 15302 42852 15308
rect 43180 15026 43208 16050
rect 43272 15162 43300 19110
rect 43352 18828 43404 18834
rect 43352 18770 43404 18776
rect 43364 18737 43392 18770
rect 43350 18728 43406 18737
rect 43350 18663 43406 18672
rect 43456 18170 43484 19246
rect 44088 19236 44140 19242
rect 44088 19178 44140 19184
rect 43536 19168 43588 19174
rect 43536 19110 43588 19116
rect 43548 18358 43576 19110
rect 43626 18864 43682 18873
rect 44100 18834 44128 19178
rect 44652 19174 44680 19654
rect 44640 19168 44692 19174
rect 44640 19110 44692 19116
rect 44652 18834 44680 19110
rect 43626 18799 43682 18808
rect 44088 18828 44140 18834
rect 43640 18748 43668 18799
rect 44088 18770 44140 18776
rect 44640 18828 44692 18834
rect 44640 18770 44692 18776
rect 43720 18760 43772 18766
rect 43640 18720 43720 18748
rect 43720 18702 43772 18708
rect 43812 18760 43864 18766
rect 43812 18702 43864 18708
rect 43536 18352 43588 18358
rect 43536 18294 43588 18300
rect 43628 18284 43680 18290
rect 43628 18226 43680 18232
rect 43640 18170 43668 18226
rect 43456 18142 43668 18170
rect 43824 17814 43852 18702
rect 44100 18086 44128 18770
rect 44180 18624 44232 18630
rect 44180 18566 44232 18572
rect 44088 18080 44140 18086
rect 44088 18022 44140 18028
rect 43812 17808 43864 17814
rect 43812 17750 43864 17756
rect 43824 17202 43852 17750
rect 44192 17746 44220 18566
rect 44282 18524 44590 18533
rect 44282 18522 44288 18524
rect 44344 18522 44368 18524
rect 44424 18522 44448 18524
rect 44504 18522 44528 18524
rect 44584 18522 44590 18524
rect 44344 18470 44346 18522
rect 44526 18470 44528 18522
rect 44282 18468 44288 18470
rect 44344 18468 44368 18470
rect 44424 18468 44448 18470
rect 44504 18468 44528 18470
rect 44584 18468 44590 18470
rect 44282 18459 44590 18468
rect 44180 17740 44232 17746
rect 44180 17682 44232 17688
rect 44744 17678 44772 21286
rect 44836 21146 44864 21422
rect 44824 21140 44876 21146
rect 44824 21082 44876 21088
rect 44928 21078 44956 21422
rect 44916 21072 44968 21078
rect 44916 21014 44968 21020
rect 44824 20256 44876 20262
rect 44824 20198 44876 20204
rect 44836 19922 44864 20198
rect 44916 19984 44968 19990
rect 44916 19926 44968 19932
rect 44824 19916 44876 19922
rect 44824 19858 44876 19864
rect 44836 18290 44864 19858
rect 44824 18284 44876 18290
rect 44824 18226 44876 18232
rect 44732 17672 44784 17678
rect 44732 17614 44784 17620
rect 43996 17536 44048 17542
rect 43996 17478 44048 17484
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 43536 16992 43588 16998
rect 43536 16934 43588 16940
rect 43548 16590 43576 16934
rect 43536 16584 43588 16590
rect 43536 16526 43588 16532
rect 44008 16250 44036 17478
rect 44282 17436 44590 17445
rect 44282 17434 44288 17436
rect 44344 17434 44368 17436
rect 44424 17434 44448 17436
rect 44504 17434 44528 17436
rect 44584 17434 44590 17436
rect 44344 17382 44346 17434
rect 44526 17382 44528 17434
rect 44282 17380 44288 17382
rect 44344 17380 44368 17382
rect 44424 17380 44448 17382
rect 44504 17380 44528 17382
rect 44584 17380 44590 17382
rect 44282 17371 44590 17380
rect 44088 17264 44140 17270
rect 44088 17206 44140 17212
rect 43996 16244 44048 16250
rect 43996 16186 44048 16192
rect 44100 16046 44128 17206
rect 44180 17128 44232 17134
rect 44180 17070 44232 17076
rect 44192 16046 44220 17070
rect 44282 16348 44590 16357
rect 44282 16346 44288 16348
rect 44344 16346 44368 16348
rect 44424 16346 44448 16348
rect 44504 16346 44528 16348
rect 44584 16346 44590 16348
rect 44344 16294 44346 16346
rect 44526 16294 44528 16346
rect 44282 16292 44288 16294
rect 44344 16292 44368 16294
rect 44424 16292 44448 16294
rect 44504 16292 44528 16294
rect 44584 16292 44590 16294
rect 44282 16283 44590 16292
rect 44088 16040 44140 16046
rect 44088 15982 44140 15988
rect 44180 16040 44232 16046
rect 44180 15982 44232 15988
rect 43720 15496 43772 15502
rect 43720 15438 43772 15444
rect 43352 15360 43404 15366
rect 43352 15302 43404 15308
rect 43260 15156 43312 15162
rect 43260 15098 43312 15104
rect 43364 15026 43392 15302
rect 43168 15020 43220 15026
rect 43168 14962 43220 14968
rect 43352 15020 43404 15026
rect 43352 14962 43404 14968
rect 43732 14482 43760 15438
rect 44732 15428 44784 15434
rect 44732 15370 44784 15376
rect 44180 15360 44232 15366
rect 44180 15302 44232 15308
rect 44640 15360 44692 15366
rect 44640 15302 44692 15308
rect 44192 15026 44220 15302
rect 44282 15260 44590 15269
rect 44282 15258 44288 15260
rect 44344 15258 44368 15260
rect 44424 15258 44448 15260
rect 44504 15258 44528 15260
rect 44584 15258 44590 15260
rect 44344 15206 44346 15258
rect 44526 15206 44528 15258
rect 44282 15204 44288 15206
rect 44344 15204 44368 15206
rect 44424 15204 44448 15206
rect 44504 15204 44528 15206
rect 44584 15204 44590 15206
rect 44282 15195 44590 15204
rect 44652 15026 44680 15302
rect 44744 15162 44772 15370
rect 44732 15156 44784 15162
rect 44732 15098 44784 15104
rect 44180 15020 44232 15026
rect 44180 14962 44232 14968
rect 44640 15020 44692 15026
rect 44640 14962 44692 14968
rect 43812 14816 43864 14822
rect 43812 14758 43864 14764
rect 43720 14476 43772 14482
rect 43720 14418 43772 14424
rect 43824 14278 43852 14758
rect 44836 14482 44864 18226
rect 44928 15570 44956 19926
rect 45020 19854 45048 21422
rect 45560 21412 45612 21418
rect 45560 21354 45612 21360
rect 45572 21146 45600 21354
rect 46584 21350 46612 22102
rect 46676 22030 46704 22374
rect 47964 22166 47992 22374
rect 47952 22160 48004 22166
rect 47952 22102 48004 22108
rect 46664 22024 46716 22030
rect 46664 21966 46716 21972
rect 47964 21978 47992 22102
rect 46572 21344 46624 21350
rect 46572 21286 46624 21292
rect 45192 21140 45244 21146
rect 45192 21082 45244 21088
rect 45560 21140 45612 21146
rect 45560 21082 45612 21088
rect 45008 19848 45060 19854
rect 45008 19790 45060 19796
rect 45204 19334 45232 21082
rect 45560 20392 45612 20398
rect 45560 20334 45612 20340
rect 45376 20256 45428 20262
rect 45376 20198 45428 20204
rect 45388 19718 45416 20198
rect 45376 19712 45428 19718
rect 45376 19654 45428 19660
rect 45204 19306 45324 19334
rect 45296 18737 45324 19306
rect 45388 18766 45416 19654
rect 45572 19514 45600 20334
rect 46676 19922 46704 21966
rect 47964 21950 48084 21978
rect 48148 21962 48176 22630
rect 48240 22574 48268 22918
rect 48228 22568 48280 22574
rect 48228 22510 48280 22516
rect 48608 22098 48636 23190
rect 49148 23112 49200 23118
rect 49148 23054 49200 23060
rect 49056 23044 49108 23050
rect 49056 22986 49108 22992
rect 48872 22636 48924 22642
rect 48872 22578 48924 22584
rect 48884 22234 48912 22578
rect 48872 22228 48924 22234
rect 48872 22170 48924 22176
rect 48596 22092 48648 22098
rect 48596 22034 48648 22040
rect 47952 21888 48004 21894
rect 47952 21830 48004 21836
rect 47964 21554 47992 21830
rect 47952 21548 48004 21554
rect 47952 21490 48004 21496
rect 48056 21434 48084 21950
rect 48136 21956 48188 21962
rect 48136 21898 48188 21904
rect 47964 21406 48084 21434
rect 47308 20256 47360 20262
rect 47308 20198 47360 20204
rect 46664 19916 46716 19922
rect 46664 19858 46716 19864
rect 47320 19854 47348 20198
rect 47308 19848 47360 19854
rect 47308 19790 47360 19796
rect 47860 19848 47912 19854
rect 47860 19790 47912 19796
rect 45836 19712 45888 19718
rect 45836 19654 45888 19660
rect 45848 19514 45876 19654
rect 45560 19508 45612 19514
rect 45560 19450 45612 19456
rect 45836 19508 45888 19514
rect 45836 19450 45888 19456
rect 47872 19446 47900 19790
rect 47860 19440 47912 19446
rect 47860 19382 47912 19388
rect 46296 19304 46348 19310
rect 46296 19246 46348 19252
rect 46756 19304 46808 19310
rect 46756 19246 46808 19252
rect 47768 19304 47820 19310
rect 47768 19246 47820 19252
rect 45836 19168 45888 19174
rect 45836 19110 45888 19116
rect 45848 18970 45876 19110
rect 45836 18964 45888 18970
rect 45836 18906 45888 18912
rect 45376 18760 45428 18766
rect 45282 18728 45338 18737
rect 45008 18692 45060 18698
rect 45376 18702 45428 18708
rect 45282 18663 45338 18672
rect 45008 18634 45060 18640
rect 45020 18426 45048 18634
rect 45296 18630 45324 18663
rect 45284 18624 45336 18630
rect 45284 18566 45336 18572
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 45296 18358 45324 18566
rect 46308 18426 46336 19246
rect 46768 18970 46796 19246
rect 46940 19168 46992 19174
rect 46940 19110 46992 19116
rect 46756 18964 46808 18970
rect 46756 18906 46808 18912
rect 46296 18420 46348 18426
rect 46296 18362 46348 18368
rect 45284 18352 45336 18358
rect 45284 18294 45336 18300
rect 45192 16788 45244 16794
rect 45192 16730 45244 16736
rect 45008 16448 45060 16454
rect 45008 16390 45060 16396
rect 45020 16046 45048 16390
rect 45204 16250 45232 16730
rect 45192 16244 45244 16250
rect 45192 16186 45244 16192
rect 45468 16108 45520 16114
rect 45468 16050 45520 16056
rect 45928 16108 45980 16114
rect 45928 16050 45980 16056
rect 45008 16040 45060 16046
rect 45008 15982 45060 15988
rect 44916 15564 44968 15570
rect 44916 15506 44968 15512
rect 44824 14476 44876 14482
rect 44824 14418 44876 14424
rect 44928 14414 44956 15506
rect 44916 14408 44968 14414
rect 44916 14350 44968 14356
rect 43812 14272 43864 14278
rect 43812 14214 43864 14220
rect 44180 14272 44232 14278
rect 44180 14214 44232 14220
rect 42720 14062 42840 14090
rect 43824 14074 43852 14214
rect 42708 14000 42760 14006
rect 42708 13942 42760 13948
rect 42616 13388 42668 13394
rect 42616 13330 42668 13336
rect 42616 13252 42668 13258
rect 42536 13212 42616 13240
rect 42432 12640 42484 12646
rect 42432 12582 42484 12588
rect 42340 12300 42392 12306
rect 42340 12242 42392 12248
rect 42444 12102 42472 12582
rect 42536 12102 42564 13212
rect 42616 13194 42668 13200
rect 42720 12986 42748 13942
rect 42708 12980 42760 12986
rect 42708 12922 42760 12928
rect 42812 12866 42840 14062
rect 43812 14068 43864 14074
rect 43812 14010 43864 14016
rect 44192 13938 44220 14214
rect 44282 14172 44590 14181
rect 44282 14170 44288 14172
rect 44344 14170 44368 14172
rect 44424 14170 44448 14172
rect 44504 14170 44528 14172
rect 44584 14170 44590 14172
rect 44344 14118 44346 14170
rect 44526 14118 44528 14170
rect 44282 14116 44288 14118
rect 44344 14116 44368 14118
rect 44424 14116 44448 14118
rect 44504 14116 44528 14118
rect 44584 14116 44590 14118
rect 44282 14107 44590 14116
rect 44088 13932 44140 13938
rect 44088 13874 44140 13880
rect 44180 13932 44232 13938
rect 44180 13874 44232 13880
rect 44100 13326 44128 13874
rect 44272 13728 44324 13734
rect 44272 13670 44324 13676
rect 43260 13320 43312 13326
rect 43260 13262 43312 13268
rect 44088 13320 44140 13326
rect 44088 13262 44140 13268
rect 43272 12986 43300 13262
rect 44284 13258 44312 13670
rect 44272 13252 44324 13258
rect 44272 13194 44324 13200
rect 44282 13084 44590 13093
rect 44282 13082 44288 13084
rect 44344 13082 44368 13084
rect 44424 13082 44448 13084
rect 44504 13082 44528 13084
rect 44584 13082 44590 13084
rect 44344 13030 44346 13082
rect 44526 13030 44528 13082
rect 44282 13028 44288 13030
rect 44344 13028 44368 13030
rect 44424 13028 44448 13030
rect 44504 13028 44528 13030
rect 44584 13028 44590 13030
rect 44282 13019 44590 13028
rect 43260 12980 43312 12986
rect 43260 12922 43312 12928
rect 42628 12838 42840 12866
rect 42892 12844 42944 12850
rect 42432 12096 42484 12102
rect 42432 12038 42484 12044
rect 42524 12096 42576 12102
rect 42524 12038 42576 12044
rect 42248 11892 42300 11898
rect 42248 11834 42300 11840
rect 41984 11648 42196 11676
rect 41420 11620 41472 11626
rect 41420 11562 41472 11568
rect 41236 11144 41288 11150
rect 41236 11086 41288 11092
rect 41144 11008 41196 11014
rect 41144 10950 41196 10956
rect 41156 10062 41184 10950
rect 41144 10056 41196 10062
rect 41144 9998 41196 10004
rect 40866 9616 40922 9625
rect 41248 9602 41276 11086
rect 41328 11008 41380 11014
rect 41328 10950 41380 10956
rect 41340 10674 41368 10950
rect 41328 10668 41380 10674
rect 41328 10610 41380 10616
rect 41604 10600 41656 10606
rect 41604 10542 41656 10548
rect 41788 10600 41840 10606
rect 41788 10542 41840 10548
rect 41328 10124 41380 10130
rect 41328 10066 41380 10072
rect 41512 10124 41564 10130
rect 41512 10066 41564 10072
rect 41340 9722 41368 10066
rect 41524 9994 41552 10066
rect 41616 10062 41644 10542
rect 41800 10266 41828 10542
rect 41880 10464 41932 10470
rect 41880 10406 41932 10412
rect 41788 10260 41840 10266
rect 41788 10202 41840 10208
rect 41892 10130 41920 10406
rect 41880 10124 41932 10130
rect 41880 10066 41932 10072
rect 41604 10056 41656 10062
rect 41604 9998 41656 10004
rect 41512 9988 41564 9994
rect 41512 9930 41564 9936
rect 41524 9722 41552 9930
rect 41616 9722 41644 9998
rect 41328 9716 41380 9722
rect 41328 9658 41380 9664
rect 41512 9716 41564 9722
rect 41512 9658 41564 9664
rect 41604 9716 41656 9722
rect 41604 9658 41656 9664
rect 41248 9574 41368 9602
rect 40866 9551 40922 9560
rect 40500 9512 40552 9518
rect 40500 9454 40552 9460
rect 40684 9512 40736 9518
rect 40684 9454 40736 9460
rect 40696 9110 40724 9454
rect 40684 9104 40736 9110
rect 40684 9046 40736 9052
rect 40592 9036 40644 9042
rect 40592 8978 40644 8984
rect 40604 8022 40632 8978
rect 40776 8288 40828 8294
rect 40776 8230 40828 8236
rect 40592 8016 40644 8022
rect 40592 7958 40644 7964
rect 40788 7478 40816 8230
rect 40776 7472 40828 7478
rect 40776 7414 40828 7420
rect 40880 5778 40908 9551
rect 41340 9382 41368 9574
rect 41328 9376 41380 9382
rect 41984 9330 42012 11648
rect 42260 11354 42288 11834
rect 42536 11694 42564 12038
rect 42524 11688 42576 11694
rect 42524 11630 42576 11636
rect 42248 11348 42300 11354
rect 42248 11290 42300 11296
rect 42064 11076 42116 11082
rect 42064 11018 42116 11024
rect 41328 9318 41380 9324
rect 41892 9302 42012 9330
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 41604 8424 41656 8430
rect 41604 8366 41656 8372
rect 41236 8288 41288 8294
rect 41236 8230 41288 8236
rect 41248 7886 41276 8230
rect 41432 8090 41460 8366
rect 41420 8084 41472 8090
rect 41420 8026 41472 8032
rect 41236 7880 41288 7886
rect 41236 7822 41288 7828
rect 41420 7880 41472 7886
rect 41472 7840 41552 7868
rect 41420 7822 41472 7828
rect 40960 6792 41012 6798
rect 40960 6734 41012 6740
rect 40868 5772 40920 5778
rect 40868 5714 40920 5720
rect 40868 5568 40920 5574
rect 40868 5510 40920 5516
rect 40880 4554 40908 5510
rect 40972 4622 41000 6734
rect 41420 5704 41472 5710
rect 41420 5646 41472 5652
rect 41432 5386 41460 5646
rect 41340 5370 41460 5386
rect 41524 5370 41552 7840
rect 41616 7546 41644 8366
rect 41696 7744 41748 7750
rect 41696 7686 41748 7692
rect 41604 7540 41656 7546
rect 41604 7482 41656 7488
rect 41708 6798 41736 7686
rect 41788 6928 41840 6934
rect 41788 6870 41840 6876
rect 41696 6792 41748 6798
rect 41696 6734 41748 6740
rect 41800 6458 41828 6870
rect 41788 6452 41840 6458
rect 41788 6394 41840 6400
rect 41788 5704 41840 5710
rect 41788 5646 41840 5652
rect 41696 5568 41748 5574
rect 41696 5510 41748 5516
rect 41328 5364 41460 5370
rect 41380 5358 41460 5364
rect 41512 5364 41564 5370
rect 41328 5306 41380 5312
rect 41512 5306 41564 5312
rect 41420 5024 41472 5030
rect 41420 4966 41472 4972
rect 40960 4616 41012 4622
rect 40960 4558 41012 4564
rect 40868 4548 40920 4554
rect 40868 4490 40920 4496
rect 40972 4214 41000 4558
rect 40960 4208 41012 4214
rect 40960 4150 41012 4156
rect 41432 4078 41460 4966
rect 41524 4146 41552 5306
rect 41708 4554 41736 5510
rect 41696 4548 41748 4554
rect 41696 4490 41748 4496
rect 41708 4282 41736 4490
rect 41696 4276 41748 4282
rect 41696 4218 41748 4224
rect 41512 4140 41564 4146
rect 41512 4082 41564 4088
rect 41420 4072 41472 4078
rect 41420 4014 41472 4020
rect 41800 3738 41828 5646
rect 41892 5302 41920 9302
rect 41972 9172 42024 9178
rect 41972 9114 42024 9120
rect 41984 8906 42012 9114
rect 41972 8900 42024 8906
rect 41972 8842 42024 8848
rect 41984 7954 42012 8842
rect 41972 7948 42024 7954
rect 41972 7890 42024 7896
rect 41984 7546 42012 7890
rect 41972 7540 42024 7546
rect 41972 7482 42024 7488
rect 41880 5296 41932 5302
rect 41880 5238 41932 5244
rect 41892 4570 41920 5238
rect 41892 4542 42012 4570
rect 41880 4480 41932 4486
rect 41880 4422 41932 4428
rect 40408 3732 40460 3738
rect 40408 3674 40460 3680
rect 41788 3732 41840 3738
rect 41788 3674 41840 3680
rect 41696 3664 41748 3670
rect 41696 3606 41748 3612
rect 41144 3460 41196 3466
rect 41144 3402 41196 3408
rect 40408 3392 40460 3398
rect 40408 3334 40460 3340
rect 40420 3058 40448 3334
rect 40408 3052 40460 3058
rect 40408 2994 40460 3000
rect 40960 3052 41012 3058
rect 40960 2994 41012 3000
rect 40972 2650 41000 2994
rect 40960 2644 41012 2650
rect 40960 2586 41012 2592
rect 40500 2576 40552 2582
rect 40328 2524 40500 2530
rect 40328 2518 40552 2524
rect 40328 2502 40540 2518
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 40224 2440 40276 2446
rect 40224 2382 40276 2388
rect 40328 800 40356 2502
rect 41156 800 41184 3402
rect 41708 3398 41736 3606
rect 41892 3534 41920 4422
rect 41984 3738 42012 4542
rect 42076 3942 42104 11018
rect 42260 10810 42288 11290
rect 42248 10804 42300 10810
rect 42248 10746 42300 10752
rect 42536 10062 42564 11630
rect 42628 11354 42656 12838
rect 42892 12786 42944 12792
rect 42708 12640 42760 12646
rect 42708 12582 42760 12588
rect 42720 12374 42748 12582
rect 42708 12368 42760 12374
rect 42708 12310 42760 12316
rect 42904 11898 42932 12786
rect 44456 12640 44508 12646
rect 44456 12582 44508 12588
rect 44468 12306 44496 12582
rect 44456 12300 44508 12306
rect 44456 12242 44508 12248
rect 43168 12232 43220 12238
rect 43168 12174 43220 12180
rect 43536 12232 43588 12238
rect 43536 12174 43588 12180
rect 42892 11892 42944 11898
rect 42892 11834 42944 11840
rect 42616 11348 42668 11354
rect 42616 11290 42668 11296
rect 43180 11014 43208 12174
rect 43548 11694 43576 12174
rect 44282 11996 44590 12005
rect 44282 11994 44288 11996
rect 44344 11994 44368 11996
rect 44424 11994 44448 11996
rect 44504 11994 44528 11996
rect 44584 11994 44590 11996
rect 44344 11942 44346 11994
rect 44526 11942 44528 11994
rect 44282 11940 44288 11942
rect 44344 11940 44368 11942
rect 44424 11940 44448 11942
rect 44504 11940 44528 11942
rect 44584 11940 44590 11942
rect 44282 11931 44590 11940
rect 43536 11688 43588 11694
rect 43536 11630 43588 11636
rect 43548 11354 43576 11630
rect 43536 11348 43588 11354
rect 43536 11290 43588 11296
rect 43812 11144 43864 11150
rect 43812 11086 43864 11092
rect 44180 11144 44232 11150
rect 44180 11086 44232 11092
rect 44824 11144 44876 11150
rect 44824 11086 44876 11092
rect 43168 11008 43220 11014
rect 43168 10950 43220 10956
rect 43180 10130 43208 10950
rect 43824 10810 43852 11086
rect 43904 11008 43956 11014
rect 43904 10950 43956 10956
rect 43812 10804 43864 10810
rect 43812 10746 43864 10752
rect 43916 10674 43944 10950
rect 43904 10668 43956 10674
rect 43904 10610 43956 10616
rect 44192 10266 44220 11086
rect 44640 11008 44692 11014
rect 44640 10950 44692 10956
rect 44282 10908 44590 10917
rect 44282 10906 44288 10908
rect 44344 10906 44368 10908
rect 44424 10906 44448 10908
rect 44504 10906 44528 10908
rect 44584 10906 44590 10908
rect 44344 10854 44346 10906
rect 44526 10854 44528 10906
rect 44282 10852 44288 10854
rect 44344 10852 44368 10854
rect 44424 10852 44448 10854
rect 44504 10852 44528 10854
rect 44584 10852 44590 10854
rect 44282 10843 44590 10852
rect 44652 10674 44680 10950
rect 44640 10668 44692 10674
rect 44640 10610 44692 10616
rect 44180 10260 44232 10266
rect 44180 10202 44232 10208
rect 43168 10124 43220 10130
rect 43168 10066 43220 10072
rect 42524 10056 42576 10062
rect 42444 10016 42524 10044
rect 42444 9178 42472 10016
rect 42524 9998 42576 10004
rect 44088 9988 44140 9994
rect 44088 9930 44140 9936
rect 42800 9920 42852 9926
rect 42800 9862 42852 9868
rect 42524 9716 42576 9722
rect 42524 9658 42576 9664
rect 42432 9172 42484 9178
rect 42432 9114 42484 9120
rect 42156 8900 42208 8906
rect 42156 8842 42208 8848
rect 42064 3936 42116 3942
rect 42064 3878 42116 3884
rect 41972 3732 42024 3738
rect 41972 3674 42024 3680
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 41696 3392 41748 3398
rect 41696 3334 41748 3340
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 41892 3074 41920 3334
rect 42168 3194 42196 8842
rect 42536 8498 42564 9658
rect 42812 9110 42840 9862
rect 44100 9722 44128 9930
rect 44282 9820 44590 9829
rect 44282 9818 44288 9820
rect 44344 9818 44368 9820
rect 44424 9818 44448 9820
rect 44504 9818 44528 9820
rect 44584 9818 44590 9820
rect 44344 9766 44346 9818
rect 44526 9766 44528 9818
rect 44282 9764 44288 9766
rect 44344 9764 44368 9766
rect 44424 9764 44448 9766
rect 44504 9764 44528 9766
rect 44584 9764 44590 9766
rect 44282 9755 44590 9764
rect 43996 9716 44048 9722
rect 43996 9658 44048 9664
rect 44088 9716 44140 9722
rect 44088 9658 44140 9664
rect 44008 9178 44036 9658
rect 44836 9450 44864 11086
rect 45020 10010 45048 15982
rect 45480 15706 45508 16050
rect 45468 15700 45520 15706
rect 45468 15642 45520 15648
rect 45940 15162 45968 16050
rect 46848 15564 46900 15570
rect 46848 15506 46900 15512
rect 46664 15496 46716 15502
rect 46664 15438 46716 15444
rect 46204 15360 46256 15366
rect 46204 15302 46256 15308
rect 45928 15156 45980 15162
rect 45928 15098 45980 15104
rect 46216 15026 46244 15302
rect 46204 15020 46256 15026
rect 46204 14962 46256 14968
rect 46676 14498 46704 15438
rect 46860 14822 46888 15506
rect 46848 14816 46900 14822
rect 46848 14758 46900 14764
rect 46676 14470 46796 14498
rect 46664 14408 46716 14414
rect 46664 14350 46716 14356
rect 45928 14272 45980 14278
rect 45928 14214 45980 14220
rect 46204 14272 46256 14278
rect 46204 14214 46256 14220
rect 45560 13864 45612 13870
rect 45560 13806 45612 13812
rect 45572 13530 45600 13806
rect 45560 13524 45612 13530
rect 45560 13466 45612 13472
rect 45940 13326 45968 14214
rect 46216 14074 46244 14214
rect 46676 14074 46704 14350
rect 46768 14074 46796 14470
rect 46204 14068 46256 14074
rect 46204 14010 46256 14016
rect 46664 14068 46716 14074
rect 46664 14010 46716 14016
rect 46756 14068 46808 14074
rect 46756 14010 46808 14016
rect 46216 13326 46244 14010
rect 46480 13728 46532 13734
rect 46480 13670 46532 13676
rect 45560 13320 45612 13326
rect 45560 13262 45612 13268
rect 45928 13320 45980 13326
rect 45928 13262 45980 13268
rect 46204 13320 46256 13326
rect 46204 13262 46256 13268
rect 45572 12986 45600 13262
rect 45560 12980 45612 12986
rect 45560 12922 45612 12928
rect 46020 12844 46072 12850
rect 46020 12786 46072 12792
rect 45100 12776 45152 12782
rect 45100 12718 45152 12724
rect 45744 12776 45796 12782
rect 45744 12718 45796 12724
rect 45112 12442 45140 12718
rect 45100 12436 45152 12442
rect 45756 12434 45784 12718
rect 45100 12378 45152 12384
rect 45664 12406 45784 12434
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 45192 10124 45244 10130
rect 45192 10066 45244 10072
rect 45020 9982 45140 10010
rect 45008 9920 45060 9926
rect 45008 9862 45060 9868
rect 45020 9586 45048 9862
rect 45008 9580 45060 9586
rect 45008 9522 45060 9528
rect 44824 9444 44876 9450
rect 44824 9386 44876 9392
rect 43996 9172 44048 9178
rect 43996 9114 44048 9120
rect 42800 9104 42852 9110
rect 42800 9046 42852 9052
rect 42524 8492 42576 8498
rect 42524 8434 42576 8440
rect 42616 8492 42668 8498
rect 42616 8434 42668 8440
rect 42628 7954 42656 8434
rect 42812 8090 42840 9046
rect 44916 9036 44968 9042
rect 44916 8978 44968 8984
rect 43444 8968 43496 8974
rect 43444 8910 43496 8916
rect 42892 8832 42944 8838
rect 42892 8774 42944 8780
rect 42904 8634 42932 8774
rect 42892 8628 42944 8634
rect 42892 8570 42944 8576
rect 43168 8288 43220 8294
rect 43168 8230 43220 8236
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 43076 8016 43128 8022
rect 43076 7958 43128 7964
rect 42616 7948 42668 7954
rect 42616 7890 42668 7896
rect 42892 7880 42944 7886
rect 42892 7822 42944 7828
rect 42904 6458 42932 7822
rect 43088 7410 43116 7958
rect 43180 7410 43208 8230
rect 43456 8090 43484 8910
rect 44282 8732 44590 8741
rect 44282 8730 44288 8732
rect 44344 8730 44368 8732
rect 44424 8730 44448 8732
rect 44504 8730 44528 8732
rect 44584 8730 44590 8732
rect 44344 8678 44346 8730
rect 44526 8678 44528 8730
rect 44282 8676 44288 8678
rect 44344 8676 44368 8678
rect 44424 8676 44448 8678
rect 44504 8676 44528 8678
rect 44584 8676 44590 8678
rect 44282 8667 44590 8676
rect 44180 8356 44232 8362
rect 44180 8298 44232 8304
rect 43996 8288 44048 8294
rect 43996 8230 44048 8236
rect 43444 8084 43496 8090
rect 43444 8026 43496 8032
rect 44008 7954 44036 8230
rect 43996 7948 44048 7954
rect 43996 7890 44048 7896
rect 43260 7880 43312 7886
rect 43260 7822 43312 7828
rect 43076 7404 43128 7410
rect 43076 7346 43128 7352
rect 43168 7404 43220 7410
rect 43272 7392 43300 7822
rect 43352 7744 43404 7750
rect 43352 7686 43404 7692
rect 43904 7744 43956 7750
rect 43904 7686 43956 7692
rect 43364 7546 43392 7686
rect 43352 7540 43404 7546
rect 43352 7482 43404 7488
rect 43352 7404 43404 7410
rect 43272 7364 43352 7392
rect 43168 7346 43220 7352
rect 43352 7346 43404 7352
rect 43916 6730 43944 7686
rect 44192 7342 44220 8298
rect 44640 7880 44692 7886
rect 44640 7822 44692 7828
rect 44282 7644 44590 7653
rect 44282 7642 44288 7644
rect 44344 7642 44368 7644
rect 44424 7642 44448 7644
rect 44504 7642 44528 7644
rect 44584 7642 44590 7644
rect 44344 7590 44346 7642
rect 44526 7590 44528 7642
rect 44282 7588 44288 7590
rect 44344 7588 44368 7590
rect 44424 7588 44448 7590
rect 44504 7588 44528 7590
rect 44584 7588 44590 7590
rect 44282 7579 44590 7588
rect 44652 7546 44680 7822
rect 44640 7540 44692 7546
rect 44640 7482 44692 7488
rect 44928 7342 44956 8978
rect 44180 7336 44232 7342
rect 44180 7278 44232 7284
rect 44916 7336 44968 7342
rect 44916 7278 44968 7284
rect 43996 7268 44048 7274
rect 43996 7210 44048 7216
rect 44008 6730 44036 7210
rect 43904 6724 43956 6730
rect 43904 6666 43956 6672
rect 43996 6724 44048 6730
rect 43996 6666 44048 6672
rect 43260 6656 43312 6662
rect 43260 6598 43312 6604
rect 42892 6452 42944 6458
rect 42892 6394 42944 6400
rect 43272 6338 43300 6598
rect 43272 6310 43392 6338
rect 42616 6180 42668 6186
rect 42616 6122 42668 6128
rect 42340 5704 42392 5710
rect 42340 5646 42392 5652
rect 42246 4040 42302 4049
rect 42246 3975 42302 3984
rect 42260 3534 42288 3975
rect 42352 3602 42380 5646
rect 42432 5160 42484 5166
rect 42432 5102 42484 5108
rect 42444 4826 42472 5102
rect 42628 5098 42656 6122
rect 42984 5704 43036 5710
rect 42984 5646 43036 5652
rect 43076 5704 43128 5710
rect 43076 5646 43128 5652
rect 42708 5636 42760 5642
rect 42708 5578 42760 5584
rect 42616 5092 42668 5098
rect 42616 5034 42668 5040
rect 42720 5030 42748 5578
rect 42892 5160 42944 5166
rect 42892 5102 42944 5108
rect 42708 5024 42760 5030
rect 42708 4966 42760 4972
rect 42800 5024 42852 5030
rect 42800 4966 42852 4972
rect 42432 4820 42484 4826
rect 42432 4762 42484 4768
rect 42812 4622 42840 4966
rect 42432 4616 42484 4622
rect 42432 4558 42484 4564
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 42444 4282 42472 4558
rect 42432 4276 42484 4282
rect 42432 4218 42484 4224
rect 42800 4140 42852 4146
rect 42800 4082 42852 4088
rect 42340 3596 42392 3602
rect 42340 3538 42392 3544
rect 42248 3528 42300 3534
rect 42248 3470 42300 3476
rect 42812 3194 42840 4082
rect 42904 3738 42932 5102
rect 42892 3732 42944 3738
rect 42892 3674 42944 3680
rect 42156 3188 42208 3194
rect 42156 3130 42208 3136
rect 42800 3188 42852 3194
rect 42800 3130 42852 3136
rect 41892 3046 42104 3074
rect 42996 3058 43024 5646
rect 43088 4758 43116 5646
rect 43260 5296 43312 5302
rect 43260 5238 43312 5244
rect 43168 5024 43220 5030
rect 43168 4966 43220 4972
rect 43076 4752 43128 4758
rect 43076 4694 43128 4700
rect 43180 4690 43208 4966
rect 43168 4684 43220 4690
rect 43168 4626 43220 4632
rect 43180 4282 43208 4626
rect 43168 4276 43220 4282
rect 43168 4218 43220 4224
rect 43272 4078 43300 5238
rect 43260 4072 43312 4078
rect 43260 4014 43312 4020
rect 43168 4004 43220 4010
rect 43168 3946 43220 3952
rect 43180 3738 43208 3946
rect 43364 3738 43392 6310
rect 44008 6100 44036 6666
rect 44282 6556 44590 6565
rect 44282 6554 44288 6556
rect 44344 6554 44368 6556
rect 44424 6554 44448 6556
rect 44504 6554 44528 6556
rect 44584 6554 44590 6556
rect 44344 6502 44346 6554
rect 44526 6502 44528 6554
rect 44282 6500 44288 6502
rect 44344 6500 44368 6502
rect 44424 6500 44448 6502
rect 44504 6500 44528 6502
rect 44584 6500 44590 6502
rect 44282 6491 44590 6500
rect 44928 6458 44956 7278
rect 45008 6792 45060 6798
rect 45008 6734 45060 6740
rect 44916 6452 44968 6458
rect 44916 6394 44968 6400
rect 45020 6322 45048 6734
rect 45008 6316 45060 6322
rect 45008 6258 45060 6264
rect 44088 6112 44140 6118
rect 44008 6072 44088 6100
rect 44088 6054 44140 6060
rect 44100 5778 44128 6054
rect 44088 5772 44140 5778
rect 44088 5714 44140 5720
rect 44180 5704 44232 5710
rect 44180 5646 44232 5652
rect 43628 5568 43680 5574
rect 43628 5510 43680 5516
rect 43536 4616 43588 4622
rect 43536 4558 43588 4564
rect 43548 4486 43576 4558
rect 43536 4480 43588 4486
rect 43536 4422 43588 4428
rect 43640 4146 43668 5510
rect 44192 5370 44220 5646
rect 44282 5468 44590 5477
rect 44282 5466 44288 5468
rect 44344 5466 44368 5468
rect 44424 5466 44448 5468
rect 44504 5466 44528 5468
rect 44584 5466 44590 5468
rect 44344 5414 44346 5466
rect 44526 5414 44528 5466
rect 44282 5412 44288 5414
rect 44344 5412 44368 5414
rect 44424 5412 44448 5414
rect 44504 5412 44528 5414
rect 44584 5412 44590 5414
rect 44282 5403 44590 5412
rect 44180 5364 44232 5370
rect 44180 5306 44232 5312
rect 43812 5228 43864 5234
rect 43812 5170 43864 5176
rect 43824 4706 43852 5170
rect 44732 5160 44784 5166
rect 44732 5102 44784 5108
rect 43732 4690 43852 4706
rect 43720 4684 43852 4690
rect 43772 4678 43852 4684
rect 43720 4626 43772 4632
rect 44282 4380 44590 4389
rect 44282 4378 44288 4380
rect 44344 4378 44368 4380
rect 44424 4378 44448 4380
rect 44504 4378 44528 4380
rect 44584 4378 44590 4380
rect 44344 4326 44346 4378
rect 44526 4326 44528 4378
rect 44282 4324 44288 4326
rect 44344 4324 44368 4326
rect 44424 4324 44448 4326
rect 44504 4324 44528 4326
rect 44584 4324 44590 4326
rect 44282 4315 44590 4324
rect 44744 4282 44772 5102
rect 45008 4480 45060 4486
rect 45008 4422 45060 4428
rect 45020 4282 45048 4422
rect 44732 4276 44784 4282
rect 44732 4218 44784 4224
rect 45008 4276 45060 4282
rect 45008 4218 45060 4224
rect 43628 4140 43680 4146
rect 43628 4082 43680 4088
rect 44916 4072 44968 4078
rect 44546 4040 44602 4049
rect 44916 4014 44968 4020
rect 44546 3975 44602 3984
rect 44272 3936 44324 3942
rect 44272 3878 44324 3884
rect 43168 3732 43220 3738
rect 43168 3674 43220 3680
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 44284 3602 44312 3878
rect 44560 3738 44588 3975
rect 44824 3936 44876 3942
rect 44824 3878 44876 3884
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 44836 3534 44864 3878
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 44928 3466 44956 4014
rect 43812 3460 43864 3466
rect 44916 3460 44968 3466
rect 43864 3420 44220 3448
rect 43812 3402 43864 3408
rect 41972 2916 42024 2922
rect 41972 2858 42024 2864
rect 41984 800 42012 2858
rect 42076 2514 42104 3046
rect 42984 3052 43036 3058
rect 42984 2994 43036 3000
rect 42800 2984 42852 2990
rect 42800 2926 42852 2932
rect 43628 2984 43680 2990
rect 43628 2926 43680 2932
rect 42812 2650 42840 2926
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 42800 2644 42852 2650
rect 42800 2586 42852 2592
rect 42064 2508 42116 2514
rect 42064 2450 42116 2456
rect 42996 1442 43024 2858
rect 42812 1414 43024 1442
rect 42812 800 42840 1414
rect 43640 800 43668 2926
rect 44192 2446 44220 3420
rect 44916 3402 44968 3408
rect 44282 3292 44590 3301
rect 44282 3290 44288 3292
rect 44344 3290 44368 3292
rect 44424 3290 44448 3292
rect 44504 3290 44528 3292
rect 44584 3290 44590 3292
rect 44344 3238 44346 3290
rect 44526 3238 44528 3290
rect 44282 3236 44288 3238
rect 44344 3236 44368 3238
rect 44424 3236 44448 3238
rect 44504 3236 44528 3238
rect 44584 3236 44590 3238
rect 44282 3227 44590 3236
rect 44640 3120 44692 3126
rect 44640 3062 44692 3068
rect 44180 2440 44232 2446
rect 44180 2382 44232 2388
rect 44282 2204 44590 2213
rect 44282 2202 44288 2204
rect 44344 2202 44368 2204
rect 44424 2202 44448 2204
rect 44504 2202 44528 2204
rect 44584 2202 44590 2204
rect 44344 2150 44346 2202
rect 44526 2150 44528 2202
rect 44282 2148 44288 2150
rect 44344 2148 44368 2150
rect 44424 2148 44448 2150
rect 44504 2148 44528 2150
rect 44584 2148 44590 2150
rect 44282 2139 44590 2148
rect 44652 1578 44680 3062
rect 45112 3058 45140 9982
rect 45204 9674 45232 10066
rect 45468 9920 45520 9926
rect 45468 9862 45520 9868
rect 45480 9722 45508 9862
rect 45468 9716 45520 9722
rect 45204 9646 45324 9674
rect 45468 9658 45520 9664
rect 45296 8974 45324 9646
rect 45284 8968 45336 8974
rect 45284 8910 45336 8916
rect 45296 8566 45324 8910
rect 45284 8560 45336 8566
rect 45284 8502 45336 8508
rect 45192 7200 45244 7206
rect 45192 7142 45244 7148
rect 45204 4486 45232 7142
rect 45480 6458 45508 9658
rect 45572 9450 45600 12038
rect 45664 11558 45692 12406
rect 46032 11898 46060 12786
rect 46492 12434 46520 13670
rect 46756 12640 46808 12646
rect 46860 12628 46888 14758
rect 46808 12600 46888 12628
rect 46756 12582 46808 12588
rect 46768 12434 46796 12582
rect 46952 12434 46980 19110
rect 47400 18624 47452 18630
rect 47400 18566 47452 18572
rect 47308 18080 47360 18086
rect 47308 18022 47360 18028
rect 47032 16448 47084 16454
rect 47032 16390 47084 16396
rect 47044 16250 47072 16390
rect 47032 16244 47084 16250
rect 47032 16186 47084 16192
rect 47320 16182 47348 18022
rect 47308 16176 47360 16182
rect 47308 16118 47360 16124
rect 47032 15904 47084 15910
rect 47032 15846 47084 15852
rect 47044 15026 47072 15846
rect 47320 15366 47348 16118
rect 47308 15360 47360 15366
rect 47308 15302 47360 15308
rect 47216 15156 47268 15162
rect 47216 15098 47268 15104
rect 47032 15020 47084 15026
rect 47032 14962 47084 14968
rect 47228 14618 47256 15098
rect 47216 14612 47268 14618
rect 47216 14554 47268 14560
rect 46400 12406 46520 12434
rect 46676 12406 46796 12434
rect 46860 12406 46980 12434
rect 47032 12436 47084 12442
rect 46020 11892 46072 11898
rect 46020 11834 46072 11840
rect 45652 11552 45704 11558
rect 45652 11494 45704 11500
rect 45664 11286 45692 11494
rect 45652 11280 45704 11286
rect 45652 11222 45704 11228
rect 45664 10742 45692 11222
rect 45836 11144 45888 11150
rect 45836 11086 45888 11092
rect 45848 10810 45876 11086
rect 46204 11008 46256 11014
rect 46204 10950 46256 10956
rect 45836 10804 45888 10810
rect 45836 10746 45888 10752
rect 45652 10736 45704 10742
rect 45652 10678 45704 10684
rect 46112 10668 46164 10674
rect 46112 10610 46164 10616
rect 46124 10198 46152 10610
rect 45652 10192 45704 10198
rect 45652 10134 45704 10140
rect 46112 10192 46164 10198
rect 46112 10134 46164 10140
rect 45664 9586 45692 10134
rect 46020 9988 46072 9994
rect 46020 9930 46072 9936
rect 46032 9722 46060 9930
rect 46020 9716 46072 9722
rect 46020 9658 46072 9664
rect 46216 9654 46244 10950
rect 46400 10266 46428 12406
rect 46676 12186 46704 12406
rect 46860 12322 46888 12406
rect 47032 12378 47084 12384
rect 46768 12306 46888 12322
rect 46756 12300 46888 12306
rect 46808 12294 46888 12300
rect 46756 12242 46808 12248
rect 46676 12158 46796 12186
rect 46480 11008 46532 11014
rect 46480 10950 46532 10956
rect 46492 10742 46520 10950
rect 46480 10736 46532 10742
rect 46480 10678 46532 10684
rect 46664 10736 46716 10742
rect 46664 10678 46716 10684
rect 46388 10260 46440 10266
rect 46388 10202 46440 10208
rect 46480 10260 46532 10266
rect 46480 10202 46532 10208
rect 46492 10146 46520 10202
rect 46400 10118 46520 10146
rect 46400 9722 46428 10118
rect 46570 9888 46626 9897
rect 46570 9823 46626 9832
rect 46388 9716 46440 9722
rect 46388 9658 46440 9664
rect 46480 9716 46532 9722
rect 46480 9658 46532 9664
rect 46204 9648 46256 9654
rect 46204 9590 46256 9596
rect 45652 9580 45704 9586
rect 45652 9522 45704 9528
rect 45560 9444 45612 9450
rect 45560 9386 45612 9392
rect 45572 8838 45600 9386
rect 46388 9376 46440 9382
rect 46388 9318 46440 9324
rect 45836 9172 45888 9178
rect 45836 9114 45888 9120
rect 45560 8832 45612 8838
rect 45560 8774 45612 8780
rect 45848 8090 45876 9114
rect 46400 9110 46428 9318
rect 46492 9178 46520 9658
rect 46584 9382 46612 9823
rect 46676 9722 46704 10678
rect 46664 9716 46716 9722
rect 46664 9658 46716 9664
rect 46572 9376 46624 9382
rect 46572 9318 46624 9324
rect 46480 9172 46532 9178
rect 46480 9114 46532 9120
rect 46388 9104 46440 9110
rect 46388 9046 46440 9052
rect 45836 8084 45888 8090
rect 45836 8026 45888 8032
rect 45744 7336 45796 7342
rect 45744 7278 45796 7284
rect 45652 7268 45704 7274
rect 45652 7210 45704 7216
rect 45560 7200 45612 7206
rect 45560 7142 45612 7148
rect 45572 6798 45600 7142
rect 45560 6792 45612 6798
rect 45560 6734 45612 6740
rect 45468 6452 45520 6458
rect 45468 6394 45520 6400
rect 45664 6322 45692 7210
rect 45756 6662 45784 7278
rect 45848 6769 45876 8026
rect 46480 7336 46532 7342
rect 46480 7278 46532 7284
rect 46664 7336 46716 7342
rect 46664 7278 46716 7284
rect 45834 6760 45890 6769
rect 45834 6695 45890 6704
rect 45744 6656 45796 6662
rect 45744 6598 45796 6604
rect 45652 6316 45704 6322
rect 45652 6258 45704 6264
rect 45848 5914 45876 6695
rect 46492 6458 46520 7278
rect 46676 7002 46704 7278
rect 46664 6996 46716 7002
rect 46664 6938 46716 6944
rect 46768 6882 46796 12158
rect 46860 11626 46888 12294
rect 47044 11898 47072 12378
rect 47032 11892 47084 11898
rect 47032 11834 47084 11840
rect 46848 11620 46900 11626
rect 46848 11562 46900 11568
rect 47032 11144 47084 11150
rect 47032 11086 47084 11092
rect 46848 10056 46900 10062
rect 46848 9998 46900 10004
rect 46860 9654 46888 9998
rect 47044 9897 47072 11086
rect 47030 9888 47086 9897
rect 47030 9823 47086 9832
rect 46848 9648 46900 9654
rect 46848 9590 46900 9596
rect 46940 8084 46992 8090
rect 46940 8026 46992 8032
rect 46676 6854 46796 6882
rect 46952 6866 46980 8026
rect 46940 6860 46992 6866
rect 46480 6452 46532 6458
rect 46480 6394 46532 6400
rect 46572 6316 46624 6322
rect 46572 6258 46624 6264
rect 46584 5914 46612 6258
rect 46676 6118 46704 6854
rect 46940 6802 46992 6808
rect 47124 6860 47176 6866
rect 47124 6802 47176 6808
rect 46756 6792 46808 6798
rect 46756 6734 46808 6740
rect 46664 6112 46716 6118
rect 46664 6054 46716 6060
rect 45836 5908 45888 5914
rect 45836 5850 45888 5856
rect 46572 5908 46624 5914
rect 46572 5850 46624 5856
rect 45376 5840 45428 5846
rect 45376 5782 45428 5788
rect 45284 5228 45336 5234
rect 45284 5170 45336 5176
rect 45192 4480 45244 4486
rect 45192 4422 45244 4428
rect 45100 3052 45152 3058
rect 45100 2994 45152 3000
rect 45296 2650 45324 5170
rect 45388 4690 45416 5782
rect 45848 4758 45876 5850
rect 46768 5370 46796 6734
rect 47136 6662 47164 6802
rect 47124 6656 47176 6662
rect 47124 6598 47176 6604
rect 47228 6254 47256 14554
rect 47320 12442 47348 15302
rect 47412 13462 47440 18566
rect 47780 18426 47808 19246
rect 47768 18420 47820 18426
rect 47768 18362 47820 18368
rect 47676 16584 47728 16590
rect 47676 16526 47728 16532
rect 47688 15706 47716 16526
rect 47676 15700 47728 15706
rect 47676 15642 47728 15648
rect 47584 15564 47636 15570
rect 47584 15506 47636 15512
rect 47596 15162 47624 15506
rect 47584 15156 47636 15162
rect 47584 15098 47636 15104
rect 47780 13870 47808 18362
rect 47964 18086 47992 21406
rect 48596 21344 48648 21350
rect 48596 21286 48648 21292
rect 48136 21004 48188 21010
rect 48136 20946 48188 20952
rect 48148 19174 48176 20946
rect 48608 20806 48636 21286
rect 48780 21004 48832 21010
rect 48780 20946 48832 20952
rect 48596 20800 48648 20806
rect 48596 20742 48648 20748
rect 48228 20392 48280 20398
rect 48228 20334 48280 20340
rect 48412 20392 48464 20398
rect 48412 20334 48464 20340
rect 48240 20058 48268 20334
rect 48424 20058 48452 20334
rect 48228 20052 48280 20058
rect 48228 19994 48280 20000
rect 48412 20052 48464 20058
rect 48412 19994 48464 20000
rect 48412 19780 48464 19786
rect 48412 19722 48464 19728
rect 48424 19446 48452 19722
rect 48412 19440 48464 19446
rect 48412 19382 48464 19388
rect 48136 19168 48188 19174
rect 48136 19110 48188 19116
rect 48320 19168 48372 19174
rect 48320 19110 48372 19116
rect 48228 18964 48280 18970
rect 48228 18906 48280 18912
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 47952 18080 48004 18086
rect 47952 18022 48004 18028
rect 48148 17202 48176 18770
rect 48136 17196 48188 17202
rect 48136 17138 48188 17144
rect 48148 16794 48176 17138
rect 48136 16788 48188 16794
rect 48136 16730 48188 16736
rect 48240 16454 48268 18906
rect 48332 18766 48360 19110
rect 48320 18760 48372 18766
rect 48320 18702 48372 18708
rect 48228 16448 48280 16454
rect 48228 16390 48280 16396
rect 48240 16130 48268 16390
rect 48148 16114 48268 16130
rect 48148 16108 48280 16114
rect 48148 16102 48228 16108
rect 48148 15706 48176 16102
rect 48228 16050 48280 16056
rect 48412 16040 48464 16046
rect 48240 15988 48412 15994
rect 48240 15982 48464 15988
rect 48240 15966 48452 15982
rect 48136 15700 48188 15706
rect 48136 15642 48188 15648
rect 48240 15434 48268 15966
rect 48608 15586 48636 20742
rect 48688 20256 48740 20262
rect 48688 20198 48740 20204
rect 48700 19922 48728 20198
rect 48792 19922 48820 20946
rect 48688 19916 48740 19922
rect 48688 19858 48740 19864
rect 48780 19916 48832 19922
rect 48780 19858 48832 19864
rect 48780 19712 48832 19718
rect 48780 19654 48832 19660
rect 48688 15972 48740 15978
rect 48688 15914 48740 15920
rect 48516 15570 48636 15586
rect 48504 15564 48636 15570
rect 48556 15558 48636 15564
rect 48504 15506 48556 15512
rect 48228 15428 48280 15434
rect 48228 15370 48280 15376
rect 48240 15162 48268 15370
rect 48228 15156 48280 15162
rect 48228 15098 48280 15104
rect 48516 15026 48544 15506
rect 48700 15450 48728 15914
rect 48608 15422 48728 15450
rect 48608 15366 48636 15422
rect 48596 15360 48648 15366
rect 48596 15302 48648 15308
rect 48504 15020 48556 15026
rect 48504 14962 48556 14968
rect 48596 14612 48648 14618
rect 48596 14554 48648 14560
rect 48608 14278 48636 14554
rect 48596 14272 48648 14278
rect 48596 14214 48648 14220
rect 48608 13938 48636 14214
rect 48320 13932 48372 13938
rect 48320 13874 48372 13880
rect 48596 13932 48648 13938
rect 48596 13874 48648 13880
rect 47584 13864 47636 13870
rect 47584 13806 47636 13812
rect 47768 13864 47820 13870
rect 47768 13806 47820 13812
rect 47596 13530 47624 13806
rect 47584 13524 47636 13530
rect 47584 13466 47636 13472
rect 47400 13456 47452 13462
rect 47400 13398 47452 13404
rect 48332 13394 48360 13874
rect 48228 13388 48280 13394
rect 48228 13330 48280 13336
rect 48320 13388 48372 13394
rect 48320 13330 48372 13336
rect 47584 13184 47636 13190
rect 47584 13126 47636 13132
rect 47596 12986 47624 13126
rect 47584 12980 47636 12986
rect 47584 12922 47636 12928
rect 47492 12776 47544 12782
rect 47492 12718 47544 12724
rect 47308 12436 47360 12442
rect 47504 12434 47532 12718
rect 47504 12406 47716 12434
rect 47308 12378 47360 12384
rect 47688 12306 47716 12406
rect 47676 12300 47728 12306
rect 47676 12242 47728 12248
rect 48240 10742 48268 13330
rect 48504 13320 48556 13326
rect 48332 13268 48504 13274
rect 48332 13262 48556 13268
rect 48332 13246 48544 13262
rect 48332 12918 48360 13246
rect 48412 13184 48464 13190
rect 48412 13126 48464 13132
rect 48320 12912 48372 12918
rect 48320 12854 48372 12860
rect 48424 12102 48452 13126
rect 48504 12300 48556 12306
rect 48504 12242 48556 12248
rect 48412 12096 48464 12102
rect 48412 12038 48464 12044
rect 48320 11008 48372 11014
rect 48320 10950 48372 10956
rect 48228 10736 48280 10742
rect 48228 10678 48280 10684
rect 48332 10606 48360 10950
rect 48320 10600 48372 10606
rect 48320 10542 48372 10548
rect 48228 10464 48280 10470
rect 48228 10406 48280 10412
rect 48240 10130 48268 10406
rect 47768 10124 47820 10130
rect 47768 10066 47820 10072
rect 48228 10124 48280 10130
rect 48228 10066 48280 10072
rect 47584 10056 47636 10062
rect 47584 9998 47636 10004
rect 47596 9382 47624 9998
rect 47780 9722 47808 10066
rect 48332 9994 48360 10542
rect 48424 10146 48452 12038
rect 48516 11014 48544 12242
rect 48504 11008 48556 11014
rect 48504 10950 48556 10956
rect 48516 10470 48544 10950
rect 48504 10464 48556 10470
rect 48504 10406 48556 10412
rect 48516 10266 48544 10406
rect 48504 10260 48556 10266
rect 48504 10202 48556 10208
rect 48424 10118 48544 10146
rect 48320 9988 48372 9994
rect 48320 9930 48372 9936
rect 47860 9920 47912 9926
rect 47860 9862 47912 9868
rect 47768 9716 47820 9722
rect 47768 9658 47820 9664
rect 47872 9586 47900 9862
rect 48332 9586 48360 9930
rect 48412 9920 48464 9926
rect 48412 9862 48464 9868
rect 47768 9580 47820 9586
rect 47768 9522 47820 9528
rect 47860 9580 47912 9586
rect 47860 9522 47912 9528
rect 48320 9580 48372 9586
rect 48320 9522 48372 9528
rect 47584 9376 47636 9382
rect 47584 9318 47636 9324
rect 47780 9042 47808 9522
rect 47952 9376 48004 9382
rect 47952 9318 48004 9324
rect 47768 9036 47820 9042
rect 47768 8978 47820 8984
rect 47584 8424 47636 8430
rect 47584 8366 47636 8372
rect 47596 8090 47624 8366
rect 47584 8084 47636 8090
rect 47584 8026 47636 8032
rect 47780 7546 47808 8978
rect 47964 8974 47992 9318
rect 47952 8968 48004 8974
rect 47952 8910 48004 8916
rect 48332 8634 48360 9522
rect 48320 8628 48372 8634
rect 48320 8570 48372 8576
rect 48228 8288 48280 8294
rect 48228 8230 48280 8236
rect 48240 7546 48268 8230
rect 48332 7954 48360 8570
rect 48320 7948 48372 7954
rect 48320 7890 48372 7896
rect 47768 7540 47820 7546
rect 47768 7482 47820 7488
rect 48228 7540 48280 7546
rect 48228 7482 48280 7488
rect 47952 7472 48004 7478
rect 47952 7414 48004 7420
rect 47400 7336 47452 7342
rect 47400 7278 47452 7284
rect 47216 6248 47268 6254
rect 47216 6190 47268 6196
rect 47032 5636 47084 5642
rect 47032 5578 47084 5584
rect 46756 5364 46808 5370
rect 46756 5306 46808 5312
rect 46020 5024 46072 5030
rect 46020 4966 46072 4972
rect 46572 5024 46624 5030
rect 46572 4966 46624 4972
rect 45836 4752 45888 4758
rect 45836 4694 45888 4700
rect 46032 4690 46060 4966
rect 45376 4684 45428 4690
rect 45376 4626 45428 4632
rect 46020 4684 46072 4690
rect 46020 4626 46072 4632
rect 45468 4616 45520 4622
rect 45468 4558 45520 4564
rect 46388 4616 46440 4622
rect 46388 4558 46440 4564
rect 45480 3466 45508 4558
rect 46400 4282 46428 4558
rect 46388 4276 46440 4282
rect 46388 4218 46440 4224
rect 46584 4010 46612 4966
rect 46768 4622 46796 5306
rect 46756 4616 46808 4622
rect 46756 4558 46808 4564
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 46572 4004 46624 4010
rect 46572 3946 46624 3952
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 46112 3392 46164 3398
rect 46112 3334 46164 3340
rect 45284 2644 45336 2650
rect 45284 2586 45336 2592
rect 45284 2372 45336 2378
rect 45284 2314 45336 2320
rect 44468 1550 44680 1578
rect 44468 800 44496 1550
rect 45296 800 45324 2314
rect 46124 800 46152 3334
rect 46296 3052 46348 3058
rect 46296 2994 46348 3000
rect 46308 2825 46336 2994
rect 46584 2990 46612 3946
rect 46676 3738 46704 4014
rect 46664 3732 46716 3738
rect 46664 3674 46716 3680
rect 46572 2984 46624 2990
rect 46572 2926 46624 2932
rect 46294 2816 46350 2825
rect 46294 2751 46350 2760
rect 46676 2446 46704 3674
rect 47044 2650 47072 5578
rect 47228 5574 47256 6190
rect 47216 5568 47268 5574
rect 47216 5510 47268 5516
rect 47412 4049 47440 7278
rect 47584 7200 47636 7206
rect 47584 7142 47636 7148
rect 47596 6866 47624 7142
rect 47492 6860 47544 6866
rect 47596 6860 47661 6866
rect 47596 6820 47609 6860
rect 47492 6802 47544 6808
rect 47609 6802 47661 6808
rect 47504 6474 47532 6802
rect 47768 6792 47820 6798
rect 47582 6760 47638 6769
rect 47688 6752 47768 6780
rect 47688 6746 47716 6752
rect 47638 6718 47716 6746
rect 47768 6734 47820 6740
rect 47582 6695 47638 6704
rect 47504 6458 47716 6474
rect 47504 6452 47728 6458
rect 47504 6446 47676 6452
rect 47676 6394 47728 6400
rect 47964 6390 47992 7414
rect 48424 6866 48452 9862
rect 48516 7478 48544 10118
rect 48504 7472 48556 7478
rect 48504 7414 48556 7420
rect 48412 6860 48464 6866
rect 48412 6802 48464 6808
rect 48320 6656 48372 6662
rect 48320 6598 48372 6604
rect 47952 6384 48004 6390
rect 47952 6326 48004 6332
rect 47584 6316 47636 6322
rect 47584 6258 47636 6264
rect 47596 5778 47624 6258
rect 47964 5914 47992 6326
rect 48136 6248 48188 6254
rect 48136 6190 48188 6196
rect 48148 5914 48176 6190
rect 47952 5908 48004 5914
rect 47952 5850 48004 5856
rect 48136 5908 48188 5914
rect 48136 5850 48188 5856
rect 47584 5772 47636 5778
rect 47584 5714 47636 5720
rect 47964 4486 47992 5850
rect 47952 4480 48004 4486
rect 47952 4422 48004 4428
rect 48136 4072 48188 4078
rect 47398 4040 47454 4049
rect 47308 4004 47360 4010
rect 48136 4014 48188 4020
rect 47398 3975 47454 3984
rect 47308 3946 47360 3952
rect 47216 3188 47268 3194
rect 47216 3130 47268 3136
rect 47228 3058 47256 3130
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 47320 2774 47348 3946
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47596 3466 47624 3878
rect 47584 3460 47636 3466
rect 47584 3402 47636 3408
rect 47676 3392 47728 3398
rect 47676 3334 47728 3340
rect 47688 3126 47716 3334
rect 47584 3120 47636 3126
rect 47584 3062 47636 3068
rect 47676 3120 47728 3126
rect 47676 3062 47728 3068
rect 47320 2746 47440 2774
rect 47412 2650 47440 2746
rect 47032 2644 47084 2650
rect 47032 2586 47084 2592
rect 47400 2644 47452 2650
rect 47400 2586 47452 2592
rect 46664 2440 46716 2446
rect 46664 2382 46716 2388
rect 46940 2372 46992 2378
rect 46940 2314 46992 2320
rect 46952 800 46980 2314
rect 47596 2310 47624 3062
rect 47780 2854 47808 3878
rect 48148 3194 48176 4014
rect 48136 3188 48188 3194
rect 48136 3130 48188 3136
rect 48332 3126 48360 6598
rect 48596 5908 48648 5914
rect 48596 5850 48648 5856
rect 48608 5574 48636 5850
rect 48596 5568 48648 5574
rect 48596 5510 48648 5516
rect 48688 5568 48740 5574
rect 48688 5510 48740 5516
rect 48700 4146 48728 5510
rect 48792 4282 48820 19654
rect 48884 18970 48912 22170
rect 49068 21690 49096 22986
rect 49160 22642 49188 23054
rect 49148 22636 49200 22642
rect 49148 22578 49200 22584
rect 49160 21690 49188 22578
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49056 21684 49108 21690
rect 49056 21626 49108 21632
rect 49148 21684 49200 21690
rect 49148 21626 49200 21632
rect 49252 21554 49280 21830
rect 49240 21548 49292 21554
rect 49240 21490 49292 21496
rect 49344 21418 49372 23462
rect 51504 23420 51812 23429
rect 51504 23418 51510 23420
rect 51566 23418 51590 23420
rect 51646 23418 51670 23420
rect 51726 23418 51750 23420
rect 51806 23418 51812 23420
rect 51566 23366 51568 23418
rect 51748 23366 51750 23418
rect 51504 23364 51510 23366
rect 51566 23364 51590 23366
rect 51646 23364 51670 23366
rect 51726 23364 51750 23366
rect 51806 23364 51812 23366
rect 51504 23355 51812 23364
rect 52552 23316 52604 23322
rect 52552 23258 52604 23264
rect 51540 23112 51592 23118
rect 51540 23054 51592 23060
rect 51908 23112 51960 23118
rect 51908 23054 51960 23060
rect 49976 22976 50028 22982
rect 49976 22918 50028 22924
rect 50068 22976 50120 22982
rect 50068 22918 50120 22924
rect 50252 22976 50304 22982
rect 50252 22918 50304 22924
rect 49988 22710 50016 22918
rect 49976 22704 50028 22710
rect 49976 22646 50028 22652
rect 50080 22642 50108 22918
rect 50264 22642 50292 22918
rect 51552 22778 51580 23054
rect 51540 22772 51592 22778
rect 51540 22714 51592 22720
rect 51080 22704 51132 22710
rect 51080 22646 51132 22652
rect 50068 22636 50120 22642
rect 50068 22578 50120 22584
rect 50252 22636 50304 22642
rect 50252 22578 50304 22584
rect 49424 22500 49476 22506
rect 49424 22442 49476 22448
rect 49436 22234 49464 22442
rect 49608 22432 49660 22438
rect 49608 22374 49660 22380
rect 49424 22228 49476 22234
rect 49424 22170 49476 22176
rect 49516 21956 49568 21962
rect 49516 21898 49568 21904
rect 49424 21888 49476 21894
rect 49424 21830 49476 21836
rect 48964 21412 49016 21418
rect 48964 21354 49016 21360
rect 49332 21412 49384 21418
rect 49332 21354 49384 21360
rect 48872 18964 48924 18970
rect 48872 18906 48924 18912
rect 48872 15972 48924 15978
rect 48872 15914 48924 15920
rect 48884 15706 48912 15914
rect 48872 15700 48924 15706
rect 48872 15642 48924 15648
rect 48872 14816 48924 14822
rect 48872 14758 48924 14764
rect 48884 13938 48912 14758
rect 48872 13932 48924 13938
rect 48872 13874 48924 13880
rect 48976 13462 49004 21354
rect 49056 21140 49108 21146
rect 49056 21082 49108 21088
rect 49068 20806 49096 21082
rect 49056 20800 49108 20806
rect 49056 20742 49108 20748
rect 49332 20324 49384 20330
rect 49332 20266 49384 20272
rect 49344 20058 49372 20266
rect 49332 20052 49384 20058
rect 49332 19994 49384 20000
rect 49436 19938 49464 21830
rect 49528 21146 49556 21898
rect 49516 21140 49568 21146
rect 49516 21082 49568 21088
rect 49252 19922 49464 19938
rect 49240 19916 49464 19922
rect 49292 19910 49464 19916
rect 49240 19858 49292 19864
rect 49332 19848 49384 19854
rect 49332 19790 49384 19796
rect 49148 19508 49200 19514
rect 49148 19450 49200 19456
rect 49160 19378 49188 19450
rect 49344 19378 49372 19790
rect 49436 19718 49464 19910
rect 49620 19854 49648 22374
rect 50080 22234 50108 22578
rect 50068 22228 50120 22234
rect 50068 22170 50120 22176
rect 50160 22092 50212 22098
rect 50160 22034 50212 22040
rect 50172 21350 50200 22034
rect 50264 21962 50292 22578
rect 51092 22234 51120 22646
rect 51172 22636 51224 22642
rect 51172 22578 51224 22584
rect 51080 22228 51132 22234
rect 51080 22170 51132 22176
rect 50252 21956 50304 21962
rect 50252 21898 50304 21904
rect 50896 21888 50948 21894
rect 50896 21830 50948 21836
rect 50908 21554 50936 21830
rect 51184 21690 51212 22578
rect 51504 22332 51812 22341
rect 51504 22330 51510 22332
rect 51566 22330 51590 22332
rect 51646 22330 51670 22332
rect 51726 22330 51750 22332
rect 51806 22330 51812 22332
rect 51566 22278 51568 22330
rect 51748 22278 51750 22330
rect 51504 22276 51510 22278
rect 51566 22276 51590 22278
rect 51646 22276 51670 22278
rect 51726 22276 51750 22278
rect 51806 22276 51812 22278
rect 51504 22267 51812 22276
rect 51920 22234 51948 23054
rect 51908 22228 51960 22234
rect 51908 22170 51960 22176
rect 51172 21684 51224 21690
rect 51172 21626 51224 21632
rect 50896 21548 50948 21554
rect 50896 21490 50948 21496
rect 50160 21344 50212 21350
rect 50160 21286 50212 21292
rect 49608 19848 49660 19854
rect 49608 19790 49660 19796
rect 49424 19712 49476 19718
rect 49424 19654 49476 19660
rect 49884 19712 49936 19718
rect 49884 19654 49936 19660
rect 49148 19372 49200 19378
rect 49148 19314 49200 19320
rect 49332 19372 49384 19378
rect 49332 19314 49384 19320
rect 49056 19304 49108 19310
rect 49056 19246 49108 19252
rect 49068 18698 49096 19246
rect 49608 19236 49660 19242
rect 49608 19178 49660 19184
rect 49056 18692 49108 18698
rect 49056 18634 49108 18640
rect 49620 18086 49648 19178
rect 49700 18964 49752 18970
rect 49700 18906 49752 18912
rect 49712 18086 49740 18906
rect 49896 18086 49924 19654
rect 50068 19304 50120 19310
rect 50068 19246 50120 19252
rect 50080 18970 50108 19246
rect 50068 18964 50120 18970
rect 50068 18906 50120 18912
rect 50080 18426 50108 18906
rect 50068 18420 50120 18426
rect 50068 18362 50120 18368
rect 49608 18080 49660 18086
rect 49608 18022 49660 18028
rect 49700 18080 49752 18086
rect 49700 18022 49752 18028
rect 49884 18080 49936 18086
rect 49884 18022 49936 18028
rect 49056 16652 49108 16658
rect 49056 16594 49108 16600
rect 49068 15706 49096 16594
rect 49240 16448 49292 16454
rect 49424 16448 49476 16454
rect 49240 16390 49292 16396
rect 49344 16396 49424 16402
rect 49344 16390 49476 16396
rect 49252 15706 49280 16390
rect 49344 16374 49464 16390
rect 49344 16046 49372 16374
rect 49332 16040 49384 16046
rect 49332 15982 49384 15988
rect 49424 16040 49476 16046
rect 49424 15982 49476 15988
rect 49056 15700 49108 15706
rect 49056 15642 49108 15648
rect 49240 15700 49292 15706
rect 49240 15642 49292 15648
rect 49436 15502 49464 15982
rect 49424 15496 49476 15502
rect 49424 15438 49476 15444
rect 49240 15428 49292 15434
rect 49240 15370 49292 15376
rect 49148 14544 49200 14550
rect 49148 14486 49200 14492
rect 49160 13938 49188 14486
rect 49252 14414 49280 15370
rect 49608 14952 49660 14958
rect 49608 14894 49660 14900
rect 49332 14816 49384 14822
rect 49332 14758 49384 14764
rect 49344 14414 49372 14758
rect 49620 14618 49648 14894
rect 49608 14612 49660 14618
rect 49608 14554 49660 14560
rect 49240 14408 49292 14414
rect 49240 14350 49292 14356
rect 49332 14408 49384 14414
rect 49332 14350 49384 14356
rect 49148 13932 49200 13938
rect 49148 13874 49200 13880
rect 48964 13456 49016 13462
rect 48964 13398 49016 13404
rect 48976 12306 49004 13398
rect 49252 13258 49280 14350
rect 49344 13394 49372 14350
rect 49712 14278 49740 18022
rect 49792 15904 49844 15910
rect 49792 15846 49844 15852
rect 49700 14272 49752 14278
rect 49700 14214 49752 14220
rect 49332 13388 49384 13394
rect 49332 13330 49384 13336
rect 49240 13252 49292 13258
rect 49240 13194 49292 13200
rect 49804 12850 49832 15846
rect 49792 12844 49844 12850
rect 49792 12786 49844 12792
rect 49700 12640 49752 12646
rect 49700 12582 49752 12588
rect 48964 12300 49016 12306
rect 48964 12242 49016 12248
rect 49240 11756 49292 11762
rect 49240 11698 49292 11704
rect 49056 10736 49108 10742
rect 49056 10678 49108 10684
rect 49068 10266 49096 10678
rect 49056 10260 49108 10266
rect 49056 10202 49108 10208
rect 49148 9988 49200 9994
rect 49148 9930 49200 9936
rect 49160 9178 49188 9930
rect 49148 9172 49200 9178
rect 49148 9114 49200 9120
rect 48964 7880 49016 7886
rect 48964 7822 49016 7828
rect 48976 7546 49004 7822
rect 48964 7540 49016 7546
rect 48964 7482 49016 7488
rect 48964 7404 49016 7410
rect 48964 7346 49016 7352
rect 48872 5228 48924 5234
rect 48872 5170 48924 5176
rect 48884 4758 48912 5170
rect 48872 4752 48924 4758
rect 48872 4694 48924 4700
rect 48780 4276 48832 4282
rect 48780 4218 48832 4224
rect 48688 4140 48740 4146
rect 48688 4082 48740 4088
rect 48976 3738 49004 7346
rect 49146 6896 49202 6905
rect 49068 6866 49146 6882
rect 49056 6860 49146 6866
rect 49108 6854 49146 6860
rect 49146 6831 49202 6840
rect 49056 6802 49108 6808
rect 49068 5914 49096 6802
rect 49056 5908 49108 5914
rect 49056 5850 49108 5856
rect 49056 4616 49108 4622
rect 49056 4558 49108 4564
rect 49068 4282 49096 4558
rect 49148 4480 49200 4486
rect 49148 4422 49200 4428
rect 49056 4276 49108 4282
rect 49056 4218 49108 4224
rect 48964 3732 49016 3738
rect 48964 3674 49016 3680
rect 49160 3534 49188 4422
rect 49252 3942 49280 11698
rect 49608 11076 49660 11082
rect 49608 11018 49660 11024
rect 49620 10810 49648 11018
rect 49608 10804 49660 10810
rect 49608 10746 49660 10752
rect 49332 9920 49384 9926
rect 49332 9862 49384 9868
rect 49344 9654 49372 9862
rect 49712 9704 49740 12582
rect 49896 12434 49924 18022
rect 50172 16658 50200 21286
rect 51504 21244 51812 21253
rect 51504 21242 51510 21244
rect 51566 21242 51590 21244
rect 51646 21242 51670 21244
rect 51726 21242 51750 21244
rect 51806 21242 51812 21244
rect 51566 21190 51568 21242
rect 51748 21190 51750 21242
rect 51504 21188 51510 21190
rect 51566 21188 51590 21190
rect 51646 21188 51670 21190
rect 51726 21188 51750 21190
rect 51806 21188 51812 21190
rect 51504 21179 51812 21188
rect 50252 20528 50304 20534
rect 50252 20470 50304 20476
rect 50264 20330 50292 20470
rect 50252 20324 50304 20330
rect 50252 20266 50304 20272
rect 50264 20058 50292 20266
rect 51504 20156 51812 20165
rect 51504 20154 51510 20156
rect 51566 20154 51590 20156
rect 51646 20154 51670 20156
rect 51726 20154 51750 20156
rect 51806 20154 51812 20156
rect 51566 20102 51568 20154
rect 51748 20102 51750 20154
rect 51504 20100 51510 20102
rect 51566 20100 51590 20102
rect 51646 20100 51670 20102
rect 51726 20100 51750 20102
rect 51806 20100 51812 20102
rect 51504 20091 51812 20100
rect 50252 20052 50304 20058
rect 50252 19994 50304 20000
rect 51920 19854 51948 22170
rect 52564 22166 52592 23258
rect 52748 23050 52776 23462
rect 52736 23044 52788 23050
rect 52736 22986 52788 22992
rect 53300 22778 53328 23598
rect 53472 23520 53524 23526
rect 53472 23462 53524 23468
rect 53484 22778 53512 23462
rect 54036 23322 54064 23598
rect 54484 23588 54536 23594
rect 54484 23530 54536 23536
rect 54024 23316 54076 23322
rect 54024 23258 54076 23264
rect 53288 22772 53340 22778
rect 53288 22714 53340 22720
rect 53472 22772 53524 22778
rect 53472 22714 53524 22720
rect 54036 22658 54064 23258
rect 54208 23044 54260 23050
rect 54208 22986 54260 22992
rect 53288 22636 53340 22642
rect 54036 22630 54156 22658
rect 53288 22578 53340 22584
rect 52552 22160 52604 22166
rect 52552 22102 52604 22108
rect 52564 21690 52592 22102
rect 53300 22094 53328 22578
rect 53932 22568 53984 22574
rect 53852 22516 53932 22522
rect 53852 22510 53984 22516
rect 54024 22568 54076 22574
rect 54024 22510 54076 22516
rect 53852 22494 53972 22510
rect 53300 22066 53512 22094
rect 53484 21962 53512 22066
rect 52736 21956 52788 21962
rect 52736 21898 52788 21904
rect 53472 21956 53524 21962
rect 53472 21898 53524 21904
rect 52748 21690 52776 21898
rect 52920 21888 52972 21894
rect 52920 21830 52972 21836
rect 53288 21888 53340 21894
rect 53288 21830 53340 21836
rect 52552 21684 52604 21690
rect 52552 21626 52604 21632
rect 52736 21684 52788 21690
rect 52736 21626 52788 21632
rect 52932 21622 52960 21830
rect 52920 21616 52972 21622
rect 52920 21558 52972 21564
rect 53300 21554 53328 21830
rect 53288 21548 53340 21554
rect 53288 21490 53340 21496
rect 53852 20806 53880 22494
rect 53932 22432 53984 22438
rect 53932 22374 53984 22380
rect 52460 20800 52512 20806
rect 52460 20742 52512 20748
rect 53840 20800 53892 20806
rect 53840 20742 53892 20748
rect 50344 19848 50396 19854
rect 50344 19790 50396 19796
rect 51908 19848 51960 19854
rect 51908 19790 51960 19796
rect 50356 19514 50384 19790
rect 51724 19712 51776 19718
rect 51724 19654 51776 19660
rect 51736 19514 51764 19654
rect 50344 19508 50396 19514
rect 50344 19450 50396 19456
rect 51724 19508 51776 19514
rect 51724 19450 51776 19456
rect 51920 19378 51948 19790
rect 51908 19372 51960 19378
rect 51908 19314 51960 19320
rect 51504 19068 51812 19077
rect 51504 19066 51510 19068
rect 51566 19066 51590 19068
rect 51646 19066 51670 19068
rect 51726 19066 51750 19068
rect 51806 19066 51812 19068
rect 51566 19014 51568 19066
rect 51748 19014 51750 19066
rect 51504 19012 51510 19014
rect 51566 19012 51590 19014
rect 51646 19012 51670 19014
rect 51726 19012 51750 19014
rect 51806 19012 51812 19014
rect 51504 19003 51812 19012
rect 51920 18766 51948 19314
rect 52472 19258 52500 20742
rect 53656 20256 53708 20262
rect 53656 20198 53708 20204
rect 53668 19854 53696 20198
rect 53944 19854 53972 22374
rect 54036 22030 54064 22510
rect 54128 22438 54156 22630
rect 54116 22432 54168 22438
rect 54116 22374 54168 22380
rect 54024 22024 54076 22030
rect 54024 21966 54076 21972
rect 54036 21690 54064 21966
rect 54116 21888 54168 21894
rect 54116 21830 54168 21836
rect 54024 21684 54076 21690
rect 54024 21626 54076 21632
rect 54128 21554 54156 21830
rect 54220 21690 54248 22986
rect 54496 22574 54524 23530
rect 55220 23112 55272 23118
rect 55220 23054 55272 23060
rect 56600 23112 56652 23118
rect 56600 23054 56652 23060
rect 55128 22976 55180 22982
rect 55128 22918 55180 22924
rect 55140 22574 55168 22918
rect 55232 22642 55260 23054
rect 56048 22976 56100 22982
rect 56048 22918 56100 22924
rect 56060 22710 56088 22918
rect 56612 22778 56640 23054
rect 58726 22876 59034 22885
rect 58726 22874 58732 22876
rect 58788 22874 58812 22876
rect 58868 22874 58892 22876
rect 58948 22874 58972 22876
rect 59028 22874 59034 22876
rect 58788 22822 58790 22874
rect 58970 22822 58972 22874
rect 58726 22820 58732 22822
rect 58788 22820 58812 22822
rect 58868 22820 58892 22822
rect 58948 22820 58972 22822
rect 59028 22820 59034 22822
rect 58726 22811 59034 22820
rect 56600 22772 56652 22778
rect 56600 22714 56652 22720
rect 56048 22704 56100 22710
rect 56048 22646 56100 22652
rect 55220 22636 55272 22642
rect 55220 22578 55272 22584
rect 54484 22568 54536 22574
rect 54484 22510 54536 22516
rect 54576 22568 54628 22574
rect 54576 22510 54628 22516
rect 55128 22568 55180 22574
rect 55128 22510 55180 22516
rect 54208 21684 54260 21690
rect 54208 21626 54260 21632
rect 54116 21548 54168 21554
rect 54116 21490 54168 21496
rect 54496 21078 54524 22510
rect 54588 22098 54616 22510
rect 54576 22092 54628 22098
rect 54576 22034 54628 22040
rect 54668 22092 54720 22098
rect 54668 22034 54720 22040
rect 55220 22092 55272 22098
rect 55220 22034 55272 22040
rect 54576 21888 54628 21894
rect 54576 21830 54628 21836
rect 54484 21072 54536 21078
rect 54484 21014 54536 21020
rect 54588 21026 54616 21830
rect 54680 21146 54708 22034
rect 55232 21418 55260 22034
rect 56060 22030 56088 22646
rect 57244 22568 57296 22574
rect 57244 22510 57296 22516
rect 56048 22024 56100 22030
rect 56048 21966 56100 21972
rect 57256 21894 57284 22510
rect 57244 21888 57296 21894
rect 57244 21830 57296 21836
rect 58726 21788 59034 21797
rect 58726 21786 58732 21788
rect 58788 21786 58812 21788
rect 58868 21786 58892 21788
rect 58948 21786 58972 21788
rect 59028 21786 59034 21788
rect 58788 21734 58790 21786
rect 58970 21734 58972 21786
rect 58726 21732 58732 21734
rect 58788 21732 58812 21734
rect 58868 21732 58892 21734
rect 58948 21732 58972 21734
rect 59028 21732 59034 21734
rect 58726 21723 59034 21732
rect 55220 21412 55272 21418
rect 55220 21354 55272 21360
rect 54668 21140 54720 21146
rect 54668 21082 54720 21088
rect 56508 21072 56560 21078
rect 54588 20998 54708 21026
rect 56508 21014 56560 21020
rect 54680 20602 54708 20998
rect 55220 21004 55272 21010
rect 55220 20946 55272 20952
rect 54668 20596 54720 20602
rect 54668 20538 54720 20544
rect 54576 20460 54628 20466
rect 54576 20402 54628 20408
rect 54208 20392 54260 20398
rect 54208 20334 54260 20340
rect 53656 19848 53708 19854
rect 53656 19790 53708 19796
rect 53932 19848 53984 19854
rect 53932 19790 53984 19796
rect 52380 19230 52500 19258
rect 52380 19174 52408 19230
rect 52368 19168 52420 19174
rect 52368 19110 52420 19116
rect 52460 19168 52512 19174
rect 52460 19110 52512 19116
rect 51908 18760 51960 18766
rect 51908 18702 51960 18708
rect 51172 18692 51224 18698
rect 51172 18634 51224 18640
rect 51632 18692 51684 18698
rect 51632 18634 51684 18640
rect 51184 17202 51212 18634
rect 51644 18426 51672 18634
rect 51632 18420 51684 18426
rect 51632 18362 51684 18368
rect 51504 17980 51812 17989
rect 51504 17978 51510 17980
rect 51566 17978 51590 17980
rect 51646 17978 51670 17980
rect 51726 17978 51750 17980
rect 51806 17978 51812 17980
rect 51566 17926 51568 17978
rect 51748 17926 51750 17978
rect 51504 17924 51510 17926
rect 51566 17924 51590 17926
rect 51646 17924 51670 17926
rect 51726 17924 51750 17926
rect 51806 17924 51812 17926
rect 51504 17915 51812 17924
rect 52184 17536 52236 17542
rect 52184 17478 52236 17484
rect 52368 17536 52420 17542
rect 52368 17478 52420 17484
rect 51172 17196 51224 17202
rect 51172 17138 51224 17144
rect 50896 17128 50948 17134
rect 50896 17070 50948 17076
rect 50252 16992 50304 16998
rect 50252 16934 50304 16940
rect 50160 16652 50212 16658
rect 50160 16594 50212 16600
rect 50172 15366 50200 16594
rect 50264 16454 50292 16934
rect 50908 16794 50936 17070
rect 50896 16788 50948 16794
rect 50896 16730 50948 16736
rect 51184 16658 51212 17138
rect 52196 17134 52224 17478
rect 52380 17338 52408 17478
rect 52368 17332 52420 17338
rect 52368 17274 52420 17280
rect 52184 17128 52236 17134
rect 52184 17070 52236 17076
rect 51504 16892 51812 16901
rect 51504 16890 51510 16892
rect 51566 16890 51590 16892
rect 51646 16890 51670 16892
rect 51726 16890 51750 16892
rect 51806 16890 51812 16892
rect 51566 16838 51568 16890
rect 51748 16838 51750 16890
rect 51504 16836 51510 16838
rect 51566 16836 51590 16838
rect 51646 16836 51670 16838
rect 51726 16836 51750 16838
rect 51806 16836 51812 16838
rect 51504 16827 51812 16836
rect 51172 16652 51224 16658
rect 51172 16594 51224 16600
rect 51724 16652 51776 16658
rect 51724 16594 51776 16600
rect 50988 16584 51040 16590
rect 50988 16526 51040 16532
rect 50252 16448 50304 16454
rect 50252 16390 50304 16396
rect 50620 16448 50672 16454
rect 50620 16390 50672 16396
rect 50632 15502 50660 16390
rect 51000 16250 51028 16526
rect 50988 16244 51040 16250
rect 50988 16186 51040 16192
rect 51736 16114 51764 16594
rect 51724 16108 51776 16114
rect 51724 16050 51776 16056
rect 51504 15804 51812 15813
rect 51504 15802 51510 15804
rect 51566 15802 51590 15804
rect 51646 15802 51670 15804
rect 51726 15802 51750 15804
rect 51806 15802 51812 15804
rect 51566 15750 51568 15802
rect 51748 15750 51750 15802
rect 51504 15748 51510 15750
rect 51566 15748 51590 15750
rect 51646 15748 51670 15750
rect 51726 15748 51750 15750
rect 51806 15748 51812 15750
rect 51504 15739 51812 15748
rect 50620 15496 50672 15502
rect 50620 15438 50672 15444
rect 50160 15360 50212 15366
rect 50160 15302 50212 15308
rect 50068 13864 50120 13870
rect 50068 13806 50120 13812
rect 50080 12986 50108 13806
rect 50068 12980 50120 12986
rect 50068 12922 50120 12928
rect 49804 12406 49924 12434
rect 49804 11898 49832 12406
rect 49884 12096 49936 12102
rect 49884 12038 49936 12044
rect 49792 11892 49844 11898
rect 49792 11834 49844 11840
rect 49896 10742 49924 12038
rect 50172 11898 50200 15302
rect 50252 14952 50304 14958
rect 50252 14894 50304 14900
rect 50264 14074 50292 14894
rect 51908 14884 51960 14890
rect 51908 14826 51960 14832
rect 51080 14816 51132 14822
rect 51080 14758 51132 14764
rect 50252 14068 50304 14074
rect 50252 14010 50304 14016
rect 50712 13728 50764 13734
rect 50712 13670 50764 13676
rect 50724 13394 50752 13670
rect 50712 13388 50764 13394
rect 50712 13330 50764 13336
rect 50988 13184 51040 13190
rect 50988 13126 51040 13132
rect 51000 12986 51028 13126
rect 50988 12980 51040 12986
rect 50988 12922 51040 12928
rect 50344 12776 50396 12782
rect 50344 12718 50396 12724
rect 50356 12442 50384 12718
rect 50344 12436 50396 12442
rect 50344 12378 50396 12384
rect 50160 11892 50212 11898
rect 50160 11834 50212 11840
rect 50356 11218 50384 12378
rect 51092 12238 51120 14758
rect 51504 14716 51812 14725
rect 51504 14714 51510 14716
rect 51566 14714 51590 14716
rect 51646 14714 51670 14716
rect 51726 14714 51750 14716
rect 51806 14714 51812 14716
rect 51566 14662 51568 14714
rect 51748 14662 51750 14714
rect 51504 14660 51510 14662
rect 51566 14660 51590 14662
rect 51646 14660 51670 14662
rect 51726 14660 51750 14662
rect 51806 14660 51812 14662
rect 51504 14651 51812 14660
rect 51920 14482 51948 14826
rect 51908 14476 51960 14482
rect 51908 14418 51960 14424
rect 51540 14340 51592 14346
rect 51540 14282 51592 14288
rect 51552 14074 51580 14282
rect 51908 14272 51960 14278
rect 51908 14214 51960 14220
rect 52092 14272 52144 14278
rect 52092 14214 52144 14220
rect 51540 14068 51592 14074
rect 51540 14010 51592 14016
rect 51504 13628 51812 13637
rect 51504 13626 51510 13628
rect 51566 13626 51590 13628
rect 51646 13626 51670 13628
rect 51726 13626 51750 13628
rect 51806 13626 51812 13628
rect 51566 13574 51568 13626
rect 51748 13574 51750 13626
rect 51504 13572 51510 13574
rect 51566 13572 51590 13574
rect 51646 13572 51670 13574
rect 51726 13572 51750 13574
rect 51806 13572 51812 13574
rect 51504 13563 51812 13572
rect 51920 13530 51948 14214
rect 52104 13938 52132 14214
rect 52092 13932 52144 13938
rect 52092 13874 52144 13880
rect 51908 13524 51960 13530
rect 51908 13466 51960 13472
rect 51356 13456 51408 13462
rect 52196 13433 52224 17070
rect 52368 16516 52420 16522
rect 52368 16458 52420 16464
rect 52380 15910 52408 16458
rect 52368 15904 52420 15910
rect 52368 15846 52420 15852
rect 52380 15570 52408 15846
rect 52368 15564 52420 15570
rect 52368 15506 52420 15512
rect 52380 15162 52408 15506
rect 52368 15156 52420 15162
rect 52368 15098 52420 15104
rect 52472 14006 52500 19110
rect 54220 18970 54248 20334
rect 54588 20058 54616 20402
rect 54576 20052 54628 20058
rect 54576 19994 54628 20000
rect 54392 19712 54444 19718
rect 54392 19654 54444 19660
rect 54208 18964 54260 18970
rect 54208 18906 54260 18912
rect 53656 18896 53708 18902
rect 53656 18838 53708 18844
rect 52736 18692 52788 18698
rect 52736 18634 52788 18640
rect 52748 18426 52776 18634
rect 53196 18624 53248 18630
rect 53196 18566 53248 18572
rect 53288 18624 53340 18630
rect 53288 18566 53340 18572
rect 52736 18420 52788 18426
rect 52736 18362 52788 18368
rect 53208 18222 53236 18566
rect 53300 18426 53328 18566
rect 53288 18420 53340 18426
rect 53288 18362 53340 18368
rect 52828 18216 52880 18222
rect 52828 18158 52880 18164
rect 53196 18216 53248 18222
rect 53196 18158 53248 18164
rect 52644 18080 52696 18086
rect 52644 18022 52696 18028
rect 52656 17270 52684 18022
rect 52644 17264 52696 17270
rect 52644 17206 52696 17212
rect 52552 16448 52604 16454
rect 52552 16390 52604 16396
rect 52564 16250 52592 16390
rect 52552 16244 52604 16250
rect 52604 16204 52684 16232
rect 52552 16186 52604 16192
rect 52656 15570 52684 16204
rect 52736 16108 52788 16114
rect 52736 16050 52788 16056
rect 52644 15564 52696 15570
rect 52644 15506 52696 15512
rect 52552 15496 52604 15502
rect 52552 15438 52604 15444
rect 52564 14550 52592 15438
rect 52552 14544 52604 14550
rect 52552 14486 52604 14492
rect 52460 14000 52512 14006
rect 52460 13942 52512 13948
rect 52368 13864 52420 13870
rect 52368 13806 52420 13812
rect 51356 13398 51408 13404
rect 52182 13424 52238 13433
rect 51172 12776 51224 12782
rect 51172 12718 51224 12724
rect 51184 12594 51212 12718
rect 51368 12646 51396 13398
rect 52182 13359 52238 13368
rect 51816 13184 51868 13190
rect 51816 13126 51868 13132
rect 51828 12986 51856 13126
rect 51816 12980 51868 12986
rect 51816 12922 51868 12928
rect 51356 12640 51408 12646
rect 51184 12566 51304 12594
rect 51356 12582 51408 12588
rect 51080 12232 51132 12238
rect 51080 12174 51132 12180
rect 51276 12102 51304 12566
rect 51368 12434 51396 12582
rect 51504 12540 51812 12549
rect 51504 12538 51510 12540
rect 51566 12538 51590 12540
rect 51646 12538 51670 12540
rect 51726 12538 51750 12540
rect 51806 12538 51812 12540
rect 51566 12486 51568 12538
rect 51748 12486 51750 12538
rect 51504 12484 51510 12486
rect 51566 12484 51590 12486
rect 51646 12484 51670 12486
rect 51726 12484 51750 12486
rect 51806 12484 51812 12486
rect 51504 12475 51812 12484
rect 51368 12406 51488 12434
rect 50896 12096 50948 12102
rect 50896 12038 50948 12044
rect 51264 12096 51316 12102
rect 51264 12038 51316 12044
rect 50908 11898 50936 12038
rect 50896 11892 50948 11898
rect 50896 11834 50948 11840
rect 51460 11694 51488 12406
rect 52380 12238 52408 13806
rect 52460 13320 52512 13326
rect 52460 13262 52512 13268
rect 52472 12986 52500 13262
rect 52460 12980 52512 12986
rect 52460 12922 52512 12928
rect 52748 12889 52776 16050
rect 52734 12880 52790 12889
rect 52734 12815 52790 12824
rect 52368 12232 52420 12238
rect 52368 12174 52420 12180
rect 51448 11688 51500 11694
rect 51448 11630 51500 11636
rect 52368 11688 52420 11694
rect 52368 11630 52420 11636
rect 51356 11552 51408 11558
rect 51356 11494 51408 11500
rect 50344 11212 50396 11218
rect 50344 11154 50396 11160
rect 50620 11212 50672 11218
rect 50620 11154 50672 11160
rect 50160 11008 50212 11014
rect 50160 10950 50212 10956
rect 50172 10742 50200 10950
rect 50632 10810 50660 11154
rect 50712 11144 50764 11150
rect 50712 11086 50764 11092
rect 50724 10810 50752 11086
rect 51080 11076 51132 11082
rect 51080 11018 51132 11024
rect 50620 10804 50672 10810
rect 50620 10746 50672 10752
rect 50712 10804 50764 10810
rect 50712 10746 50764 10752
rect 49884 10736 49936 10742
rect 49884 10678 49936 10684
rect 50160 10736 50212 10742
rect 50160 10678 50212 10684
rect 50436 10260 50488 10266
rect 50436 10202 50488 10208
rect 49976 10056 50028 10062
rect 49976 9998 50028 10004
rect 49712 9676 49832 9704
rect 49332 9648 49384 9654
rect 49332 9590 49384 9596
rect 49698 9616 49754 9625
rect 49698 9551 49700 9560
rect 49752 9551 49754 9560
rect 49700 9522 49752 9528
rect 49712 9178 49740 9522
rect 49700 9172 49752 9178
rect 49700 9114 49752 9120
rect 49712 8378 49740 9114
rect 49620 8350 49740 8378
rect 49332 7948 49384 7954
rect 49332 7890 49384 7896
rect 49344 6322 49372 7890
rect 49424 6656 49476 6662
rect 49424 6598 49476 6604
rect 49436 6458 49464 6598
rect 49424 6452 49476 6458
rect 49424 6394 49476 6400
rect 49332 6316 49384 6322
rect 49332 6258 49384 6264
rect 49620 5302 49648 8350
rect 49804 5658 49832 9676
rect 49988 8634 50016 9998
rect 50344 9988 50396 9994
rect 50344 9930 50396 9936
rect 50356 9382 50384 9930
rect 50448 9926 50476 10202
rect 50436 9920 50488 9926
rect 50436 9862 50488 9868
rect 50344 9376 50396 9382
rect 50344 9318 50396 9324
rect 50356 9178 50384 9318
rect 50344 9172 50396 9178
rect 50344 9114 50396 9120
rect 50356 8634 50384 9114
rect 49976 8628 50028 8634
rect 49976 8570 50028 8576
rect 50344 8628 50396 8634
rect 50344 8570 50396 8576
rect 50448 8090 50476 9862
rect 51092 8974 51120 11018
rect 51172 11008 51224 11014
rect 51172 10950 51224 10956
rect 51184 10810 51212 10950
rect 51172 10804 51224 10810
rect 51224 10764 51304 10792
rect 51172 10746 51224 10752
rect 51276 10130 51304 10764
rect 51368 10606 51396 11494
rect 51504 11452 51812 11461
rect 51504 11450 51510 11452
rect 51566 11450 51590 11452
rect 51646 11450 51670 11452
rect 51726 11450 51750 11452
rect 51806 11450 51812 11452
rect 51566 11398 51568 11450
rect 51748 11398 51750 11450
rect 51504 11396 51510 11398
rect 51566 11396 51590 11398
rect 51646 11396 51670 11398
rect 51726 11396 51750 11398
rect 51806 11396 51812 11398
rect 51504 11387 51812 11396
rect 52092 11212 52144 11218
rect 52092 11154 52144 11160
rect 51816 10736 51868 10742
rect 51816 10678 51868 10684
rect 51356 10600 51408 10606
rect 51356 10542 51408 10548
rect 51828 10470 51856 10678
rect 51908 10668 51960 10674
rect 51908 10610 51960 10616
rect 51816 10464 51868 10470
rect 51816 10406 51868 10412
rect 51504 10364 51812 10373
rect 51504 10362 51510 10364
rect 51566 10362 51590 10364
rect 51646 10362 51670 10364
rect 51726 10362 51750 10364
rect 51806 10362 51812 10364
rect 51566 10310 51568 10362
rect 51748 10310 51750 10362
rect 51504 10308 51510 10310
rect 51566 10308 51590 10310
rect 51646 10308 51670 10310
rect 51726 10308 51750 10310
rect 51806 10308 51812 10310
rect 51504 10299 51812 10308
rect 51264 10124 51316 10130
rect 51264 10066 51316 10072
rect 51448 10056 51500 10062
rect 51448 9998 51500 10004
rect 51632 10056 51684 10062
rect 51632 9998 51684 10004
rect 51920 10010 51948 10610
rect 52000 10464 52052 10470
rect 52000 10406 52052 10412
rect 52012 10198 52040 10406
rect 52000 10192 52052 10198
rect 52000 10134 52052 10140
rect 51460 9926 51488 9998
rect 51448 9920 51500 9926
rect 51448 9862 51500 9868
rect 51644 9382 51672 9998
rect 51920 9982 52040 10010
rect 52012 9586 52040 9982
rect 52000 9580 52052 9586
rect 52000 9522 52052 9528
rect 51356 9376 51408 9382
rect 51356 9318 51408 9324
rect 51632 9376 51684 9382
rect 51632 9318 51684 9324
rect 51080 8968 51132 8974
rect 51080 8910 51132 8916
rect 51368 8566 51396 9318
rect 51504 9276 51812 9285
rect 51504 9274 51510 9276
rect 51566 9274 51590 9276
rect 51646 9274 51670 9276
rect 51726 9274 51750 9276
rect 51806 9274 51812 9276
rect 51566 9222 51568 9274
rect 51748 9222 51750 9274
rect 51504 9220 51510 9222
rect 51566 9220 51590 9222
rect 51646 9220 51670 9222
rect 51726 9220 51750 9222
rect 51806 9220 51812 9222
rect 51504 9211 51812 9220
rect 51356 8560 51408 8566
rect 51356 8502 51408 8508
rect 52012 8498 52040 9522
rect 52000 8492 52052 8498
rect 52000 8434 52052 8440
rect 51172 8288 51224 8294
rect 51172 8230 51224 8236
rect 50436 8084 50488 8090
rect 50436 8026 50488 8032
rect 50804 7948 50856 7954
rect 50804 7890 50856 7896
rect 50620 7880 50672 7886
rect 50620 7822 50672 7828
rect 50632 7206 50660 7822
rect 50816 7546 50844 7890
rect 50804 7540 50856 7546
rect 50804 7482 50856 7488
rect 50712 7404 50764 7410
rect 50712 7346 50764 7352
rect 50724 7206 50752 7346
rect 49884 7200 49936 7206
rect 49884 7142 49936 7148
rect 50620 7200 50672 7206
rect 50620 7142 50672 7148
rect 50712 7200 50764 7206
rect 50712 7142 50764 7148
rect 49896 6662 49924 7142
rect 50632 6866 50660 7142
rect 51184 6934 51212 8230
rect 51504 8188 51812 8197
rect 51504 8186 51510 8188
rect 51566 8186 51590 8188
rect 51646 8186 51670 8188
rect 51726 8186 51750 8188
rect 51806 8186 51812 8188
rect 51566 8134 51568 8186
rect 51748 8134 51750 8186
rect 51504 8132 51510 8134
rect 51566 8132 51590 8134
rect 51646 8132 51670 8134
rect 51726 8132 51750 8134
rect 51806 8132 51812 8134
rect 51504 8123 51812 8132
rect 51264 7812 51316 7818
rect 51264 7754 51316 7760
rect 51276 7410 51304 7754
rect 51632 7744 51684 7750
rect 51632 7686 51684 7692
rect 51644 7546 51672 7686
rect 51632 7540 51684 7546
rect 51632 7482 51684 7488
rect 52012 7410 52040 8434
rect 52104 8362 52132 11154
rect 52184 11144 52236 11150
rect 52184 11086 52236 11092
rect 52196 10810 52224 11086
rect 52184 10804 52236 10810
rect 52184 10746 52236 10752
rect 52380 10606 52408 11630
rect 52644 10668 52696 10674
rect 52644 10610 52696 10616
rect 52368 10600 52420 10606
rect 52368 10542 52420 10548
rect 52552 10600 52604 10606
rect 52552 10542 52604 10548
rect 52460 10260 52512 10266
rect 52460 10202 52512 10208
rect 52184 8492 52236 8498
rect 52184 8434 52236 8440
rect 52092 8356 52144 8362
rect 52092 8298 52144 8304
rect 51264 7404 51316 7410
rect 51264 7346 51316 7352
rect 52000 7404 52052 7410
rect 52000 7346 52052 7352
rect 51504 7100 51812 7109
rect 51504 7098 51510 7100
rect 51566 7098 51590 7100
rect 51646 7098 51670 7100
rect 51726 7098 51750 7100
rect 51806 7098 51812 7100
rect 51566 7046 51568 7098
rect 51748 7046 51750 7098
rect 51504 7044 51510 7046
rect 51566 7044 51590 7046
rect 51646 7044 51670 7046
rect 51726 7044 51750 7046
rect 51806 7044 51812 7046
rect 51504 7035 51812 7044
rect 51172 6928 51224 6934
rect 51172 6870 51224 6876
rect 50620 6860 50672 6866
rect 50620 6802 50672 6808
rect 49976 6792 50028 6798
rect 49976 6734 50028 6740
rect 50804 6792 50856 6798
rect 50804 6734 50856 6740
rect 49884 6656 49936 6662
rect 49884 6598 49936 6604
rect 49988 6458 50016 6734
rect 50816 6458 50844 6734
rect 51184 6662 51212 6870
rect 51356 6860 51408 6866
rect 51276 6820 51356 6848
rect 51172 6656 51224 6662
rect 51172 6598 51224 6604
rect 49976 6452 50028 6458
rect 49976 6394 50028 6400
rect 50804 6452 50856 6458
rect 50804 6394 50856 6400
rect 51172 6452 51224 6458
rect 51172 6394 51224 6400
rect 51184 6322 51212 6394
rect 51172 6316 51224 6322
rect 51172 6258 51224 6264
rect 50252 6112 50304 6118
rect 50252 6054 50304 6060
rect 50712 6112 50764 6118
rect 50712 6054 50764 6060
rect 49712 5630 49832 5658
rect 49884 5704 49936 5710
rect 49884 5646 49936 5652
rect 49608 5296 49660 5302
rect 49608 5238 49660 5244
rect 49620 4826 49648 5238
rect 49608 4820 49660 4826
rect 49608 4762 49660 4768
rect 49712 4282 49740 5630
rect 49792 5568 49844 5574
rect 49792 5510 49844 5516
rect 49700 4276 49752 4282
rect 49700 4218 49752 4224
rect 49804 4146 49832 5510
rect 49792 4140 49844 4146
rect 49792 4082 49844 4088
rect 49240 3936 49292 3942
rect 49240 3878 49292 3884
rect 49896 3738 49924 5646
rect 50264 4078 50292 6054
rect 50724 5914 50752 6054
rect 50712 5908 50764 5914
rect 50712 5850 50764 5856
rect 50528 5704 50580 5710
rect 50528 5646 50580 5652
rect 50436 4480 50488 4486
rect 50436 4422 50488 4428
rect 50252 4072 50304 4078
rect 50304 4020 50384 4026
rect 50252 4014 50384 4020
rect 50264 3998 50384 4014
rect 49884 3732 49936 3738
rect 49884 3674 49936 3680
rect 49896 3618 49924 3674
rect 50356 3641 50384 3998
rect 50342 3632 50398 3641
rect 49896 3590 50200 3618
rect 48504 3528 48556 3534
rect 48504 3470 48556 3476
rect 49148 3528 49200 3534
rect 49148 3470 49200 3476
rect 48320 3120 48372 3126
rect 48320 3062 48372 3068
rect 48516 3058 48544 3470
rect 48780 3392 48832 3398
rect 48780 3334 48832 3340
rect 48504 3052 48556 3058
rect 48504 2994 48556 3000
rect 48320 2916 48372 2922
rect 48320 2858 48372 2864
rect 47768 2848 47820 2854
rect 47768 2790 47820 2796
rect 47860 2848 47912 2854
rect 47860 2790 47912 2796
rect 47584 2304 47636 2310
rect 47584 2246 47636 2252
rect 47872 1306 47900 2790
rect 48332 2650 48360 2858
rect 48320 2644 48372 2650
rect 48320 2586 48372 2592
rect 48688 2508 48740 2514
rect 48688 2450 48740 2456
rect 47780 1278 47900 1306
rect 47780 800 47808 1278
rect 48700 1170 48728 2450
rect 48792 2446 48820 3334
rect 49422 2952 49478 2961
rect 49422 2887 49478 2896
rect 48780 2440 48832 2446
rect 48780 2382 48832 2388
rect 48608 1142 48728 1170
rect 48608 800 48636 1142
rect 49436 800 49464 2887
rect 49976 2848 50028 2854
rect 49976 2790 50028 2796
rect 49988 2650 50016 2790
rect 49976 2644 50028 2650
rect 49976 2586 50028 2592
rect 50172 2446 50200 3590
rect 50252 3596 50304 3602
rect 50342 3567 50398 3576
rect 50252 3538 50304 3544
rect 50160 2440 50212 2446
rect 50160 2382 50212 2388
rect 50264 800 50292 3538
rect 50448 3126 50476 4422
rect 50540 3534 50568 5646
rect 51184 5370 51212 6258
rect 51276 6118 51304 6820
rect 51356 6802 51408 6808
rect 51724 6792 51776 6798
rect 51776 6752 51948 6780
rect 51724 6734 51776 6740
rect 51264 6112 51316 6118
rect 51264 6054 51316 6060
rect 51276 5914 51304 6054
rect 51504 6012 51812 6021
rect 51504 6010 51510 6012
rect 51566 6010 51590 6012
rect 51646 6010 51670 6012
rect 51726 6010 51750 6012
rect 51806 6010 51812 6012
rect 51566 5958 51568 6010
rect 51748 5958 51750 6010
rect 51504 5956 51510 5958
rect 51566 5956 51590 5958
rect 51646 5956 51670 5958
rect 51726 5956 51750 5958
rect 51806 5956 51812 5958
rect 51504 5947 51812 5956
rect 51264 5908 51316 5914
rect 51264 5850 51316 5856
rect 51172 5364 51224 5370
rect 51172 5306 51224 5312
rect 51080 5160 51132 5166
rect 51080 5102 51132 5108
rect 50712 5024 50764 5030
rect 50712 4966 50764 4972
rect 50724 4622 50752 4966
rect 50712 4616 50764 4622
rect 50712 4558 50764 4564
rect 50988 4276 51040 4282
rect 51092 4264 51120 5102
rect 51040 4236 51120 4264
rect 50988 4218 51040 4224
rect 51184 4146 51212 5306
rect 51264 5296 51316 5302
rect 51264 5238 51316 5244
rect 51276 4826 51304 5238
rect 51920 5234 51948 6752
rect 52012 6458 52040 7346
rect 52104 6905 52132 8298
rect 52196 8022 52224 8434
rect 52184 8016 52236 8022
rect 52184 7958 52236 7964
rect 52090 6896 52146 6905
rect 52196 6866 52224 7958
rect 52276 7880 52328 7886
rect 52276 7822 52328 7828
rect 52288 7546 52316 7822
rect 52276 7540 52328 7546
rect 52276 7482 52328 7488
rect 52090 6831 52146 6840
rect 52184 6860 52236 6866
rect 52000 6452 52052 6458
rect 52000 6394 52052 6400
rect 52104 6254 52132 6831
rect 52184 6802 52236 6808
rect 52472 6746 52500 10202
rect 52564 9178 52592 10542
rect 52656 10266 52684 10610
rect 52644 10260 52696 10266
rect 52644 10202 52696 10208
rect 52736 10056 52788 10062
rect 52736 9998 52788 10004
rect 52748 9178 52776 9998
rect 52552 9172 52604 9178
rect 52552 9114 52604 9120
rect 52736 9172 52788 9178
rect 52736 9114 52788 9120
rect 52748 8634 52776 9114
rect 52736 8628 52788 8634
rect 52736 8570 52788 8576
rect 52748 8090 52776 8570
rect 52736 8084 52788 8090
rect 52736 8026 52788 8032
rect 52840 7562 52868 18158
rect 53668 18086 53696 18838
rect 54404 18766 54432 19654
rect 54576 19372 54628 19378
rect 54576 19314 54628 19320
rect 54484 18896 54536 18902
rect 54484 18838 54536 18844
rect 54392 18760 54444 18766
rect 54392 18702 54444 18708
rect 53748 18624 53800 18630
rect 53748 18566 53800 18572
rect 53760 18426 53788 18566
rect 53748 18420 53800 18426
rect 53748 18362 53800 18368
rect 54496 18086 54524 18838
rect 53656 18080 53708 18086
rect 53656 18022 53708 18028
rect 54484 18080 54536 18086
rect 54484 18022 54536 18028
rect 53668 17882 53696 18022
rect 53656 17876 53708 17882
rect 53656 17818 53708 17824
rect 53472 17808 53524 17814
rect 53472 17750 53524 17756
rect 53012 17672 53064 17678
rect 53012 17614 53064 17620
rect 53104 17672 53156 17678
rect 53104 17614 53156 17620
rect 52920 17128 52972 17134
rect 52920 17070 52972 17076
rect 52932 16674 52960 17070
rect 53024 16794 53052 17614
rect 53116 17338 53144 17614
rect 53484 17338 53512 17750
rect 53840 17672 53892 17678
rect 53840 17614 53892 17620
rect 53656 17536 53708 17542
rect 53656 17478 53708 17484
rect 53104 17332 53156 17338
rect 53104 17274 53156 17280
rect 53472 17332 53524 17338
rect 53472 17274 53524 17280
rect 53012 16788 53064 16794
rect 53012 16730 53064 16736
rect 52932 16646 53052 16674
rect 53024 16182 53052 16646
rect 53012 16176 53064 16182
rect 53012 16118 53064 16124
rect 53024 14346 53052 16118
rect 53484 15570 53512 17274
rect 53564 16992 53616 16998
rect 53564 16934 53616 16940
rect 53576 16590 53604 16934
rect 53668 16658 53696 17478
rect 53852 16658 53880 17614
rect 53656 16652 53708 16658
rect 53656 16594 53708 16600
rect 53748 16652 53800 16658
rect 53748 16594 53800 16600
rect 53840 16652 53892 16658
rect 53840 16594 53892 16600
rect 54208 16652 54260 16658
rect 54208 16594 54260 16600
rect 53564 16584 53616 16590
rect 53564 16526 53616 16532
rect 53564 16448 53616 16454
rect 53564 16390 53616 16396
rect 53576 16250 53604 16390
rect 53564 16244 53616 16250
rect 53564 16186 53616 16192
rect 53668 15570 53696 16594
rect 53472 15564 53524 15570
rect 53472 15506 53524 15512
rect 53656 15564 53708 15570
rect 53656 15506 53708 15512
rect 53012 14340 53064 14346
rect 53012 14282 53064 14288
rect 53288 13864 53340 13870
rect 53288 13806 53340 13812
rect 53472 13864 53524 13870
rect 53472 13806 53524 13812
rect 53104 13796 53156 13802
rect 53104 13738 53156 13744
rect 53116 13394 53144 13738
rect 53300 13462 53328 13806
rect 53288 13456 53340 13462
rect 53288 13398 53340 13404
rect 53104 13388 53156 13394
rect 53104 13330 53156 13336
rect 53196 13252 53248 13258
rect 53196 13194 53248 13200
rect 53208 12850 53236 13194
rect 53196 12844 53248 12850
rect 53196 12786 53248 12792
rect 53484 12714 53512 13806
rect 53760 13297 53788 16594
rect 53932 15428 53984 15434
rect 53932 15370 53984 15376
rect 53746 13288 53802 13297
rect 53746 13223 53802 13232
rect 53748 13184 53800 13190
rect 53748 13126 53800 13132
rect 53760 12918 53788 13126
rect 53944 13002 53972 15370
rect 54116 15020 54168 15026
rect 54116 14962 54168 14968
rect 54128 14618 54156 14962
rect 54116 14612 54168 14618
rect 54116 14554 54168 14560
rect 54128 13870 54156 14554
rect 54116 13864 54168 13870
rect 54116 13806 54168 13812
rect 54024 13728 54076 13734
rect 54024 13670 54076 13676
rect 53852 12974 53972 13002
rect 54036 12986 54064 13670
rect 54024 12980 54076 12986
rect 53748 12912 53800 12918
rect 53748 12854 53800 12860
rect 53472 12708 53524 12714
rect 53472 12650 53524 12656
rect 53104 11756 53156 11762
rect 53104 11698 53156 11704
rect 52920 9376 52972 9382
rect 52920 9318 52972 9324
rect 52932 8906 52960 9318
rect 52920 8900 52972 8906
rect 52920 8842 52972 8848
rect 52920 8356 52972 8362
rect 52920 8298 52972 8304
rect 52656 7534 52868 7562
rect 52472 6718 52592 6746
rect 52460 6656 52512 6662
rect 52460 6598 52512 6604
rect 52472 6458 52500 6598
rect 52460 6452 52512 6458
rect 52460 6394 52512 6400
rect 52564 6322 52592 6718
rect 52552 6316 52604 6322
rect 52552 6258 52604 6264
rect 52000 6248 52052 6254
rect 52000 6190 52052 6196
rect 52092 6248 52144 6254
rect 52092 6190 52144 6196
rect 52012 5914 52040 6190
rect 52368 6112 52420 6118
rect 52368 6054 52420 6060
rect 52000 5908 52052 5914
rect 52000 5850 52052 5856
rect 52380 5642 52408 6054
rect 52368 5636 52420 5642
rect 52368 5578 52420 5584
rect 52000 5568 52052 5574
rect 52000 5510 52052 5516
rect 51908 5228 51960 5234
rect 51908 5170 51960 5176
rect 51356 5160 51408 5166
rect 51356 5102 51408 5108
rect 51264 4820 51316 4826
rect 51264 4762 51316 4768
rect 51172 4140 51224 4146
rect 51172 4082 51224 4088
rect 50986 4040 51042 4049
rect 50986 3975 51042 3984
rect 50528 3528 50580 3534
rect 50528 3470 50580 3476
rect 50540 3194 50568 3470
rect 51000 3194 51028 3975
rect 51172 3528 51224 3534
rect 51276 3516 51304 4762
rect 51368 4010 51396 5102
rect 51504 4924 51812 4933
rect 51504 4922 51510 4924
rect 51566 4922 51590 4924
rect 51646 4922 51670 4924
rect 51726 4922 51750 4924
rect 51806 4922 51812 4924
rect 51566 4870 51568 4922
rect 51748 4870 51750 4922
rect 51504 4868 51510 4870
rect 51566 4868 51590 4870
rect 51646 4868 51670 4870
rect 51726 4868 51750 4870
rect 51806 4868 51812 4870
rect 51504 4859 51812 4868
rect 51540 4616 51592 4622
rect 51540 4558 51592 4564
rect 51552 4078 51580 4558
rect 52012 4146 52040 5510
rect 52380 5250 52408 5578
rect 52288 5222 52408 5250
rect 52288 4758 52316 5222
rect 52368 5160 52420 5166
rect 52368 5102 52420 5108
rect 52380 4826 52408 5102
rect 52368 4820 52420 4826
rect 52368 4762 52420 4768
rect 52276 4752 52328 4758
rect 52276 4694 52328 4700
rect 52276 4616 52328 4622
rect 52276 4558 52328 4564
rect 52288 4282 52316 4558
rect 52368 4480 52420 4486
rect 52368 4422 52420 4428
rect 52276 4276 52328 4282
rect 52276 4218 52328 4224
rect 52000 4140 52052 4146
rect 52000 4082 52052 4088
rect 51540 4072 51592 4078
rect 51540 4014 51592 4020
rect 51356 4004 51408 4010
rect 51356 3946 51408 3952
rect 51504 3836 51812 3845
rect 51504 3834 51510 3836
rect 51566 3834 51590 3836
rect 51646 3834 51670 3836
rect 51726 3834 51750 3836
rect 51806 3834 51812 3836
rect 51566 3782 51568 3834
rect 51748 3782 51750 3834
rect 51504 3780 51510 3782
rect 51566 3780 51590 3782
rect 51646 3780 51670 3782
rect 51726 3780 51750 3782
rect 51806 3780 51812 3782
rect 51504 3771 51812 3780
rect 51224 3488 51304 3516
rect 51172 3470 51224 3476
rect 51184 3194 51212 3470
rect 50528 3188 50580 3194
rect 50528 3130 50580 3136
rect 50988 3188 51040 3194
rect 50988 3130 51040 3136
rect 51172 3188 51224 3194
rect 51172 3130 51224 3136
rect 50436 3120 50488 3126
rect 50436 3062 50488 3068
rect 52380 3058 52408 4422
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 51080 2916 51132 2922
rect 51080 2858 51132 2864
rect 51092 2446 51120 2858
rect 51356 2848 51408 2854
rect 51170 2816 51226 2825
rect 51356 2790 51408 2796
rect 51170 2751 51226 2760
rect 51184 2650 51212 2751
rect 51172 2644 51224 2650
rect 51172 2586 51224 2592
rect 51080 2440 51132 2446
rect 51080 2382 51132 2388
rect 51092 870 51212 898
rect 51092 800 51120 870
rect 38764 734 39068 762
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43626 0 43682 800
rect 44454 0 44510 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46938 0 46994 800
rect 47766 0 47822 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51078 0 51134 800
rect 51184 762 51212 870
rect 51368 762 51396 2790
rect 51504 2748 51812 2757
rect 51504 2746 51510 2748
rect 51566 2746 51590 2748
rect 51646 2746 51670 2748
rect 51726 2746 51750 2748
rect 51806 2746 51812 2748
rect 51566 2694 51568 2746
rect 51748 2694 51750 2746
rect 51504 2692 51510 2694
rect 51566 2692 51590 2694
rect 51646 2692 51670 2694
rect 51726 2692 51750 2694
rect 51806 2692 51812 2694
rect 51504 2683 51812 2692
rect 52656 2446 52684 7534
rect 52736 7200 52788 7206
rect 52736 7142 52788 7148
rect 52748 6390 52776 7142
rect 52736 6384 52788 6390
rect 52736 6326 52788 6332
rect 52736 6112 52788 6118
rect 52736 6054 52788 6060
rect 52748 4282 52776 6054
rect 52932 5914 52960 8298
rect 52920 5908 52972 5914
rect 52972 5868 53052 5896
rect 52920 5850 52972 5856
rect 52828 5704 52880 5710
rect 52828 5646 52880 5652
rect 52736 4276 52788 4282
rect 52736 4218 52788 4224
rect 52736 4072 52788 4078
rect 52736 4014 52788 4020
rect 52748 3738 52776 4014
rect 52736 3732 52788 3738
rect 52736 3674 52788 3680
rect 52748 3641 52776 3674
rect 52734 3632 52790 3641
rect 52734 3567 52790 3576
rect 52840 2854 52868 5646
rect 52920 5024 52972 5030
rect 52920 4966 52972 4972
rect 52932 4758 52960 4966
rect 52920 4752 52972 4758
rect 52920 4694 52972 4700
rect 52932 3738 52960 4694
rect 52920 3732 52972 3738
rect 52920 3674 52972 3680
rect 53024 2990 53052 5868
rect 53116 4049 53144 11698
rect 53472 10464 53524 10470
rect 53472 10406 53524 10412
rect 53484 9994 53512 10406
rect 53852 9994 53880 12974
rect 54024 12922 54076 12928
rect 53932 12912 53984 12918
rect 53932 12854 53984 12860
rect 53944 12442 53972 12854
rect 53932 12436 53984 12442
rect 53932 12378 53984 12384
rect 54220 10810 54248 16594
rect 54392 16108 54444 16114
rect 54392 16050 54444 16056
rect 54404 15162 54432 16050
rect 54496 15570 54524 18022
rect 54588 17746 54616 19314
rect 54680 18630 54708 20538
rect 55232 20482 55260 20946
rect 55864 20936 55916 20942
rect 55864 20878 55916 20884
rect 56048 20936 56100 20942
rect 56048 20878 56100 20884
rect 55404 20868 55456 20874
rect 55404 20810 55456 20816
rect 55312 20800 55364 20806
rect 55312 20742 55364 20748
rect 55140 20466 55260 20482
rect 55128 20460 55260 20466
rect 55180 20454 55260 20460
rect 55128 20402 55180 20408
rect 55220 19780 55272 19786
rect 55220 19722 55272 19728
rect 55232 18834 55260 19722
rect 55324 19378 55352 20742
rect 55416 20466 55444 20810
rect 55876 20602 55904 20878
rect 55864 20596 55916 20602
rect 55864 20538 55916 20544
rect 55404 20460 55456 20466
rect 55404 20402 55456 20408
rect 55416 19922 55444 20402
rect 55404 19916 55456 19922
rect 55404 19858 55456 19864
rect 56060 19514 56088 20878
rect 56324 20392 56376 20398
rect 56324 20334 56376 20340
rect 56140 19848 56192 19854
rect 56140 19790 56192 19796
rect 56048 19508 56100 19514
rect 56048 19450 56100 19456
rect 55312 19372 55364 19378
rect 55312 19314 55364 19320
rect 56152 18970 56180 19790
rect 56336 19378 56364 20334
rect 56520 19990 56548 21014
rect 57336 20936 57388 20942
rect 57336 20878 57388 20884
rect 56692 20800 56744 20806
rect 56692 20742 56744 20748
rect 56784 20800 56836 20806
rect 56784 20742 56836 20748
rect 56704 20262 56732 20742
rect 56796 20534 56824 20742
rect 56784 20528 56836 20534
rect 56784 20470 56836 20476
rect 56876 20460 56928 20466
rect 56876 20402 56928 20408
rect 56692 20256 56744 20262
rect 56692 20198 56744 20204
rect 56704 20058 56732 20198
rect 56888 20058 56916 20402
rect 57244 20256 57296 20262
rect 57244 20198 57296 20204
rect 56692 20052 56744 20058
rect 56692 19994 56744 20000
rect 56876 20052 56928 20058
rect 56876 19994 56928 20000
rect 56508 19984 56560 19990
rect 56508 19926 56560 19932
rect 56324 19372 56376 19378
rect 56324 19314 56376 19320
rect 56140 18964 56192 18970
rect 56140 18906 56192 18912
rect 55220 18828 55272 18834
rect 55220 18770 55272 18776
rect 54668 18624 54720 18630
rect 54668 18566 54720 18572
rect 54576 17740 54628 17746
rect 54576 17682 54628 17688
rect 54588 17202 54616 17682
rect 54576 17196 54628 17202
rect 54576 17138 54628 17144
rect 54588 16250 54616 17138
rect 54576 16244 54628 16250
rect 54576 16186 54628 16192
rect 54680 16130 54708 18566
rect 55864 17672 55916 17678
rect 55864 17614 55916 17620
rect 56048 17672 56100 17678
rect 56048 17614 56100 17620
rect 55312 17536 55364 17542
rect 55312 17478 55364 17484
rect 55324 17338 55352 17478
rect 55312 17332 55364 17338
rect 55312 17274 55364 17280
rect 55876 16794 55904 17614
rect 56060 17338 56088 17614
rect 56048 17332 56100 17338
rect 56048 17274 56100 17280
rect 56520 16998 56548 19926
rect 57256 19922 57284 20198
rect 57244 19916 57296 19922
rect 57244 19858 57296 19864
rect 57256 18766 57284 19858
rect 57348 18970 57376 20878
rect 58726 20700 59034 20709
rect 58726 20698 58732 20700
rect 58788 20698 58812 20700
rect 58868 20698 58892 20700
rect 58948 20698 58972 20700
rect 59028 20698 59034 20700
rect 58788 20646 58790 20698
rect 58970 20646 58972 20698
rect 58726 20644 58732 20646
rect 58788 20644 58812 20646
rect 58868 20644 58892 20646
rect 58948 20644 58972 20646
rect 59028 20644 59034 20646
rect 58726 20635 59034 20644
rect 57428 19916 57480 19922
rect 57428 19858 57480 19864
rect 57336 18964 57388 18970
rect 57336 18906 57388 18912
rect 57244 18760 57296 18766
rect 57244 18702 57296 18708
rect 57060 17876 57112 17882
rect 57060 17818 57112 17824
rect 56600 17536 56652 17542
rect 56600 17478 56652 17484
rect 56324 16992 56376 16998
rect 56324 16934 56376 16940
rect 56508 16992 56560 16998
rect 56508 16934 56560 16940
rect 55864 16788 55916 16794
rect 55864 16730 55916 16736
rect 56336 16590 56364 16934
rect 56324 16584 56376 16590
rect 56324 16526 56376 16532
rect 56416 16584 56468 16590
rect 56416 16526 56468 16532
rect 55220 16448 55272 16454
rect 55220 16390 55272 16396
rect 54588 16102 54708 16130
rect 54484 15564 54536 15570
rect 54484 15506 54536 15512
rect 54392 15156 54444 15162
rect 54392 15098 54444 15104
rect 54300 14272 54352 14278
rect 54300 14214 54352 14220
rect 54312 13258 54340 14214
rect 54300 13252 54352 13258
rect 54300 13194 54352 13200
rect 54392 12096 54444 12102
rect 54392 12038 54444 12044
rect 54404 11082 54432 12038
rect 54588 11898 54616 16102
rect 55232 15366 55260 16390
rect 55312 16244 55364 16250
rect 55312 16186 55364 16192
rect 55324 15638 55352 16186
rect 56336 15910 56364 16526
rect 55496 15904 55548 15910
rect 55496 15846 55548 15852
rect 56324 15904 56376 15910
rect 56324 15846 56376 15852
rect 55508 15706 55536 15846
rect 56428 15706 56456 16526
rect 56520 16250 56548 16934
rect 56612 16794 56640 17478
rect 56876 17196 56928 17202
rect 56876 17138 56928 17144
rect 56784 16992 56836 16998
rect 56784 16934 56836 16940
rect 56796 16794 56824 16934
rect 56888 16794 56916 17138
rect 56600 16788 56652 16794
rect 56600 16730 56652 16736
rect 56784 16788 56836 16794
rect 56784 16730 56836 16736
rect 56876 16788 56928 16794
rect 56876 16730 56928 16736
rect 56612 16590 56640 16730
rect 56784 16652 56836 16658
rect 56784 16594 56836 16600
rect 56600 16584 56652 16590
rect 56600 16526 56652 16532
rect 56508 16244 56560 16250
rect 56508 16186 56560 16192
rect 56796 15706 56824 16594
rect 56888 16454 56916 16730
rect 56876 16448 56928 16454
rect 56876 16390 56928 16396
rect 55496 15700 55548 15706
rect 55496 15642 55548 15648
rect 56416 15700 56468 15706
rect 56416 15642 56468 15648
rect 56784 15700 56836 15706
rect 56784 15642 56836 15648
rect 55312 15632 55364 15638
rect 55312 15574 55364 15580
rect 54668 15360 54720 15366
rect 54668 15302 54720 15308
rect 55220 15360 55272 15366
rect 55220 15302 55272 15308
rect 54680 15026 54708 15302
rect 54668 15020 54720 15026
rect 54668 14962 54720 14968
rect 54852 14408 54904 14414
rect 54852 14350 54904 14356
rect 54864 14074 54892 14350
rect 54852 14068 54904 14074
rect 54852 14010 54904 14016
rect 55128 14000 55180 14006
rect 55324 13954 55352 15574
rect 56784 15564 56836 15570
rect 56784 15506 56836 15512
rect 56796 15366 56824 15506
rect 55772 15360 55824 15366
rect 55772 15302 55824 15308
rect 56784 15360 56836 15366
rect 56784 15302 56836 15308
rect 55128 13942 55180 13948
rect 55140 13190 55168 13942
rect 55232 13926 55352 13954
rect 55128 13184 55180 13190
rect 55128 13126 55180 13132
rect 54760 12980 54812 12986
rect 54760 12922 54812 12928
rect 54772 12850 54800 12922
rect 54760 12844 54812 12850
rect 54760 12786 54812 12792
rect 55140 12782 55168 13126
rect 54668 12776 54720 12782
rect 54668 12718 54720 12724
rect 54944 12776 54996 12782
rect 54944 12718 54996 12724
rect 55128 12776 55180 12782
rect 55128 12718 55180 12724
rect 54680 12102 54708 12718
rect 54956 12442 54984 12718
rect 55232 12714 55260 13926
rect 55312 13864 55364 13870
rect 55312 13806 55364 13812
rect 55324 13530 55352 13806
rect 55312 13524 55364 13530
rect 55312 13466 55364 13472
rect 55312 13320 55364 13326
rect 55312 13262 55364 13268
rect 55220 12708 55272 12714
rect 55220 12650 55272 12656
rect 54944 12436 54996 12442
rect 54944 12378 54996 12384
rect 55232 12170 55260 12650
rect 55324 12434 55352 13262
rect 55496 12436 55548 12442
rect 55324 12406 55496 12434
rect 55496 12378 55548 12384
rect 55220 12164 55272 12170
rect 55220 12106 55272 12112
rect 54668 12096 54720 12102
rect 54668 12038 54720 12044
rect 54576 11892 54628 11898
rect 54576 11834 54628 11840
rect 54392 11076 54444 11082
rect 54392 11018 54444 11024
rect 54208 10804 54260 10810
rect 54208 10746 54260 10752
rect 54116 10600 54168 10606
rect 54116 10542 54168 10548
rect 54128 10266 54156 10542
rect 54208 10464 54260 10470
rect 54208 10406 54260 10412
rect 54220 10266 54248 10406
rect 54116 10260 54168 10266
rect 54116 10202 54168 10208
rect 54208 10260 54260 10266
rect 54208 10202 54260 10208
rect 53472 9988 53524 9994
rect 53472 9930 53524 9936
rect 53840 9988 53892 9994
rect 53840 9930 53892 9936
rect 53484 9722 53512 9930
rect 53472 9716 53524 9722
rect 53472 9658 53524 9664
rect 53748 9512 53800 9518
rect 53748 9454 53800 9460
rect 53760 9178 53788 9454
rect 53748 9172 53800 9178
rect 53748 9114 53800 9120
rect 53852 9110 53880 9930
rect 53840 9104 53892 9110
rect 53840 9046 53892 9052
rect 54024 9104 54076 9110
rect 54024 9046 54076 9052
rect 54036 8430 54064 9046
rect 54024 8424 54076 8430
rect 54024 8366 54076 8372
rect 53932 8288 53984 8294
rect 53932 8230 53984 8236
rect 53840 7880 53892 7886
rect 53840 7822 53892 7828
rect 53852 7546 53880 7822
rect 53840 7540 53892 7546
rect 53840 7482 53892 7488
rect 53288 7336 53340 7342
rect 53288 7278 53340 7284
rect 53300 7002 53328 7278
rect 53288 6996 53340 7002
rect 53288 6938 53340 6944
rect 53852 6798 53880 7482
rect 53944 7478 53972 8230
rect 53932 7472 53984 7478
rect 53932 7414 53984 7420
rect 54036 6866 54064 8366
rect 54404 8294 54432 11018
rect 54760 10600 54812 10606
rect 54760 10542 54812 10548
rect 55496 10600 55548 10606
rect 55496 10542 55548 10548
rect 54668 10532 54720 10538
rect 54668 10474 54720 10480
rect 54680 9722 54708 10474
rect 54668 9716 54720 9722
rect 54668 9658 54720 9664
rect 54680 9110 54708 9658
rect 54772 9382 54800 10542
rect 54944 10464 54996 10470
rect 54944 10406 54996 10412
rect 54956 9654 54984 10406
rect 55508 10266 55536 10542
rect 55496 10260 55548 10266
rect 55496 10202 55548 10208
rect 55128 10056 55180 10062
rect 55128 9998 55180 10004
rect 54944 9648 54996 9654
rect 54944 9590 54996 9596
rect 54760 9376 54812 9382
rect 54760 9318 54812 9324
rect 55140 9178 55168 9998
rect 55404 9988 55456 9994
rect 55404 9930 55456 9936
rect 55416 9586 55444 9930
rect 55404 9580 55456 9586
rect 55404 9522 55456 9528
rect 55588 9444 55640 9450
rect 55588 9386 55640 9392
rect 55312 9376 55364 9382
rect 55312 9318 55364 9324
rect 55324 9178 55352 9318
rect 55128 9172 55180 9178
rect 55128 9114 55180 9120
rect 55312 9172 55364 9178
rect 55312 9114 55364 9120
rect 54668 9104 54720 9110
rect 54668 9046 54720 9052
rect 54576 8424 54628 8430
rect 54576 8366 54628 8372
rect 54392 8288 54444 8294
rect 54392 8230 54444 8236
rect 54208 7200 54260 7206
rect 54260 7148 54340 7154
rect 54208 7142 54340 7148
rect 54220 7126 54340 7142
rect 54024 6860 54076 6866
rect 54024 6802 54076 6808
rect 53840 6792 53892 6798
rect 53840 6734 53892 6740
rect 54208 6724 54260 6730
rect 54208 6666 54260 6672
rect 54220 6458 54248 6666
rect 54208 6452 54260 6458
rect 54208 6394 54260 6400
rect 53748 5704 53800 5710
rect 53748 5646 53800 5652
rect 53564 5568 53616 5574
rect 53564 5510 53616 5516
rect 53288 5228 53340 5234
rect 53288 5170 53340 5176
rect 53196 5160 53248 5166
rect 53196 5102 53248 5108
rect 53102 4040 53158 4049
rect 53102 3975 53158 3984
rect 53104 3936 53156 3942
rect 53104 3878 53156 3884
rect 53116 3058 53144 3878
rect 53208 3738 53236 5102
rect 53300 4826 53328 5170
rect 53288 4820 53340 4826
rect 53288 4762 53340 4768
rect 53472 4480 53524 4486
rect 53472 4422 53524 4428
rect 53484 4214 53512 4422
rect 53472 4208 53524 4214
rect 53472 4150 53524 4156
rect 53288 4072 53340 4078
rect 53288 4014 53340 4020
rect 53196 3732 53248 3738
rect 53196 3674 53248 3680
rect 53300 3346 53328 4014
rect 53380 3936 53432 3942
rect 53380 3878 53432 3884
rect 53392 3534 53420 3878
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 53208 3318 53328 3346
rect 53484 3346 53512 4150
rect 53576 3534 53604 5510
rect 53656 4616 53708 4622
rect 53656 4558 53708 4564
rect 53564 3528 53616 3534
rect 53564 3470 53616 3476
rect 53562 3360 53618 3369
rect 53484 3318 53562 3346
rect 53208 3058 53236 3318
rect 53562 3295 53618 3304
rect 53104 3052 53156 3058
rect 53104 2994 53156 3000
rect 53196 3052 53248 3058
rect 53196 2994 53248 3000
rect 53012 2984 53064 2990
rect 53012 2926 53064 2932
rect 53564 2984 53616 2990
rect 53564 2926 53616 2932
rect 52828 2848 52880 2854
rect 52734 2816 52790 2825
rect 52828 2790 52880 2796
rect 52734 2751 52790 2760
rect 52644 2440 52696 2446
rect 52644 2382 52696 2388
rect 52092 2372 52144 2378
rect 51920 2332 52092 2360
rect 51920 800 51948 2332
rect 52092 2314 52144 2320
rect 52748 800 52776 2751
rect 53576 800 53604 2926
rect 53668 2378 53696 4558
rect 53760 2922 53788 5646
rect 54208 5568 54260 5574
rect 54208 5510 54260 5516
rect 54024 5228 54076 5234
rect 54024 5170 54076 5176
rect 53932 4480 53984 4486
rect 53932 4422 53984 4428
rect 53944 3738 53972 4422
rect 54036 4078 54064 5170
rect 54220 4146 54248 5510
rect 54208 4140 54260 4146
rect 54208 4082 54260 4088
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 53932 3732 53984 3738
rect 53932 3674 53984 3680
rect 54312 3602 54340 7126
rect 54588 6662 54616 8366
rect 54760 8288 54812 8294
rect 54760 8230 54812 8236
rect 54772 7206 54800 8230
rect 55496 7744 55548 7750
rect 55496 7686 55548 7692
rect 55312 7540 55364 7546
rect 55312 7482 55364 7488
rect 54760 7200 54812 7206
rect 54760 7142 54812 7148
rect 54392 6656 54444 6662
rect 54392 6598 54444 6604
rect 54576 6656 54628 6662
rect 54576 6598 54628 6604
rect 54404 6458 54432 6598
rect 54392 6452 54444 6458
rect 54392 6394 54444 6400
rect 54484 5636 54536 5642
rect 54484 5578 54536 5584
rect 54496 5166 54524 5578
rect 54668 5568 54720 5574
rect 54668 5510 54720 5516
rect 54680 5370 54708 5510
rect 54668 5364 54720 5370
rect 54668 5306 54720 5312
rect 54484 5160 54536 5166
rect 54484 5102 54536 5108
rect 54680 4146 54708 5306
rect 54668 4140 54720 4146
rect 54668 4082 54720 4088
rect 54772 4010 54800 7142
rect 55220 6656 55272 6662
rect 55220 6598 55272 6604
rect 54852 5704 54904 5710
rect 54852 5646 54904 5652
rect 54760 4004 54812 4010
rect 54760 3946 54812 3952
rect 54864 3670 54892 5646
rect 55232 5234 55260 6598
rect 55324 6322 55352 7482
rect 55508 6322 55536 7686
rect 55600 6866 55628 9386
rect 55784 8634 55812 15302
rect 56598 15056 56654 15065
rect 56598 14991 56654 15000
rect 56612 14618 56640 14991
rect 56600 14612 56652 14618
rect 56600 14554 56652 14560
rect 56612 14074 56640 14554
rect 56600 14068 56652 14074
rect 56600 14010 56652 14016
rect 55864 13932 55916 13938
rect 55864 13874 55916 13880
rect 55876 12782 55904 13874
rect 56600 13864 56652 13870
rect 56600 13806 56652 13812
rect 56048 13728 56100 13734
rect 56048 13670 56100 13676
rect 56060 13258 56088 13670
rect 56048 13252 56100 13258
rect 56048 13194 56100 13200
rect 56612 12986 56640 13806
rect 56692 13184 56744 13190
rect 56692 13126 56744 13132
rect 56704 12986 56732 13126
rect 56600 12980 56652 12986
rect 56600 12922 56652 12928
rect 56692 12980 56744 12986
rect 56692 12922 56744 12928
rect 55864 12776 55916 12782
rect 55864 12718 55916 12724
rect 56508 12776 56560 12782
rect 56508 12718 56560 12724
rect 56140 12640 56192 12646
rect 56140 12582 56192 12588
rect 56048 12232 56100 12238
rect 56048 12174 56100 12180
rect 56060 11898 56088 12174
rect 56048 11892 56100 11898
rect 56048 11834 56100 11840
rect 56152 11150 56180 12582
rect 56232 12096 56284 12102
rect 56232 12038 56284 12044
rect 56140 11144 56192 11150
rect 56140 11086 56192 11092
rect 56244 11014 56272 12038
rect 56520 11762 56548 12718
rect 56692 12232 56744 12238
rect 56692 12174 56744 12180
rect 56704 11898 56732 12174
rect 56692 11892 56744 11898
rect 56692 11834 56744 11840
rect 56508 11756 56560 11762
rect 56508 11698 56560 11704
rect 56232 11008 56284 11014
rect 56232 10950 56284 10956
rect 56244 10588 56272 10950
rect 56324 10600 56376 10606
rect 56244 10560 56324 10588
rect 56048 9988 56100 9994
rect 56048 9930 56100 9936
rect 56060 9722 56088 9930
rect 56048 9716 56100 9722
rect 56048 9658 56100 9664
rect 55772 8628 55824 8634
rect 55772 8570 55824 8576
rect 55772 8424 55824 8430
rect 55772 8366 55824 8372
rect 55680 8356 55732 8362
rect 55680 8298 55732 8304
rect 55588 6860 55640 6866
rect 55588 6802 55640 6808
rect 55600 6458 55628 6802
rect 55588 6452 55640 6458
rect 55588 6394 55640 6400
rect 55312 6316 55364 6322
rect 55312 6258 55364 6264
rect 55496 6316 55548 6322
rect 55496 6258 55548 6264
rect 55404 6112 55456 6118
rect 55404 6054 55456 6060
rect 55220 5228 55272 5234
rect 55220 5170 55272 5176
rect 55128 5092 55180 5098
rect 55128 5034 55180 5040
rect 55036 4684 55088 4690
rect 55036 4626 55088 4632
rect 54944 4548 54996 4554
rect 54944 4490 54996 4496
rect 54956 3670 54984 4490
rect 55048 4434 55076 4626
rect 55140 4622 55168 5034
rect 55232 4690 55260 5170
rect 55312 5024 55364 5030
rect 55312 4966 55364 4972
rect 55220 4684 55272 4690
rect 55220 4626 55272 4632
rect 55128 4616 55180 4622
rect 55128 4558 55180 4564
rect 55048 4406 55168 4434
rect 55140 4282 55168 4406
rect 55036 4276 55088 4282
rect 55036 4218 55088 4224
rect 55128 4276 55180 4282
rect 55128 4218 55180 4224
rect 55048 4162 55076 4218
rect 55324 4162 55352 4966
rect 55416 4758 55444 6054
rect 55404 4752 55456 4758
rect 55404 4694 55456 4700
rect 55496 4684 55548 4690
rect 55496 4626 55548 4632
rect 55048 4146 55352 4162
rect 55048 4140 55364 4146
rect 55048 4134 55312 4140
rect 55312 4082 55364 4088
rect 54852 3664 54904 3670
rect 54852 3606 54904 3612
rect 54944 3664 54996 3670
rect 54944 3606 54996 3612
rect 54300 3596 54352 3602
rect 54300 3538 54352 3544
rect 54208 3460 54260 3466
rect 54208 3402 54260 3408
rect 53748 2916 53800 2922
rect 53748 2858 53800 2864
rect 54220 2650 54248 3402
rect 55508 3398 55536 4626
rect 55588 3936 55640 3942
rect 55588 3878 55640 3884
rect 55600 3670 55628 3878
rect 55588 3664 55640 3670
rect 55588 3606 55640 3612
rect 55496 3392 55548 3398
rect 55496 3334 55548 3340
rect 55692 3194 55720 8298
rect 55680 3188 55732 3194
rect 55680 3130 55732 3136
rect 54758 2952 54814 2961
rect 54392 2916 54444 2922
rect 54758 2887 54814 2896
rect 54392 2858 54444 2864
rect 54208 2644 54260 2650
rect 54208 2586 54260 2592
rect 53656 2372 53708 2378
rect 53656 2314 53708 2320
rect 54404 800 54432 2858
rect 54772 2446 54800 2887
rect 55784 2774 55812 8366
rect 56244 8294 56272 10560
rect 56324 10542 56376 10548
rect 56416 10600 56468 10606
rect 56416 10542 56468 10548
rect 56600 10600 56652 10606
rect 56600 10542 56652 10548
rect 56428 9926 56456 10542
rect 56416 9920 56468 9926
rect 56416 9862 56468 9868
rect 56428 9110 56456 9862
rect 56612 9654 56640 10542
rect 56704 10130 56732 11834
rect 56796 11218 56824 15302
rect 56876 14272 56928 14278
rect 56876 14214 56928 14220
rect 56888 13326 56916 14214
rect 56876 13320 56928 13326
rect 56876 13262 56928 13268
rect 56968 11756 57020 11762
rect 56968 11698 57020 11704
rect 56784 11212 56836 11218
rect 56784 11154 56836 11160
rect 56784 11076 56836 11082
rect 56784 11018 56836 11024
rect 56796 10606 56824 11018
rect 56876 11008 56928 11014
rect 56876 10950 56928 10956
rect 56888 10810 56916 10950
rect 56876 10804 56928 10810
rect 56876 10746 56928 10752
rect 56784 10600 56836 10606
rect 56784 10542 56836 10548
rect 56692 10124 56744 10130
rect 56692 10066 56744 10072
rect 56692 9920 56744 9926
rect 56692 9862 56744 9868
rect 56600 9648 56652 9654
rect 56600 9590 56652 9596
rect 56612 9178 56640 9590
rect 56600 9172 56652 9178
rect 56600 9114 56652 9120
rect 56416 9104 56468 9110
rect 56416 9046 56468 9052
rect 56704 9042 56732 9862
rect 56980 9586 57008 11698
rect 57072 11354 57100 17818
rect 57440 17338 57468 19858
rect 57520 19712 57572 19718
rect 57520 19654 57572 19660
rect 57612 19712 57664 19718
rect 57612 19654 57664 19660
rect 57980 19712 58032 19718
rect 57980 19654 58032 19660
rect 57532 18970 57560 19654
rect 57520 18964 57572 18970
rect 57520 18906 57572 18912
rect 57624 18630 57652 19654
rect 57992 19378 58020 19654
rect 58726 19612 59034 19621
rect 58726 19610 58732 19612
rect 58788 19610 58812 19612
rect 58868 19610 58892 19612
rect 58948 19610 58972 19612
rect 59028 19610 59034 19612
rect 58788 19558 58790 19610
rect 58970 19558 58972 19610
rect 58726 19556 58732 19558
rect 58788 19556 58812 19558
rect 58868 19556 58892 19558
rect 58948 19556 58972 19558
rect 59028 19556 59034 19558
rect 58726 19547 59034 19556
rect 58256 19508 58308 19514
rect 58256 19450 58308 19456
rect 57980 19372 58032 19378
rect 57980 19314 58032 19320
rect 58268 18834 58296 19450
rect 58256 18828 58308 18834
rect 58256 18770 58308 18776
rect 57612 18624 57664 18630
rect 57612 18566 57664 18572
rect 58726 18524 59034 18533
rect 58726 18522 58732 18524
rect 58788 18522 58812 18524
rect 58868 18522 58892 18524
rect 58948 18522 58972 18524
rect 59028 18522 59034 18524
rect 58788 18470 58790 18522
rect 58970 18470 58972 18522
rect 58726 18468 58732 18470
rect 58788 18468 58812 18470
rect 58868 18468 58892 18470
rect 58948 18468 58972 18470
rect 59028 18468 59034 18470
rect 58726 18459 59034 18468
rect 58072 18216 58124 18222
rect 58072 18158 58124 18164
rect 57888 18080 57940 18086
rect 57888 18022 57940 18028
rect 57520 17604 57572 17610
rect 57520 17546 57572 17552
rect 57428 17332 57480 17338
rect 57428 17274 57480 17280
rect 57336 17060 57388 17066
rect 57336 17002 57388 17008
rect 57348 16182 57376 17002
rect 57336 16176 57388 16182
rect 57336 16118 57388 16124
rect 57440 15994 57468 17274
rect 57532 16250 57560 17546
rect 57900 17270 57928 18022
rect 57888 17264 57940 17270
rect 57888 17206 57940 17212
rect 57900 16658 57928 17206
rect 57888 16652 57940 16658
rect 57888 16594 57940 16600
rect 57612 16448 57664 16454
rect 57612 16390 57664 16396
rect 57888 16448 57940 16454
rect 57888 16390 57940 16396
rect 57624 16250 57652 16390
rect 57520 16244 57572 16250
rect 57520 16186 57572 16192
rect 57612 16244 57664 16250
rect 57612 16186 57664 16192
rect 57348 15966 57468 15994
rect 57244 14272 57296 14278
rect 57244 14214 57296 14220
rect 57256 14074 57284 14214
rect 57244 14068 57296 14074
rect 57244 14010 57296 14016
rect 57152 12776 57204 12782
rect 57152 12718 57204 12724
rect 57164 11762 57192 12718
rect 57152 11756 57204 11762
rect 57152 11698 57204 11704
rect 57348 11642 57376 15966
rect 57900 15706 57928 16390
rect 58084 16046 58112 18158
rect 58256 17536 58308 17542
rect 58256 17478 58308 17484
rect 58164 16652 58216 16658
rect 58164 16594 58216 16600
rect 58072 16040 58124 16046
rect 58072 15982 58124 15988
rect 57888 15700 57940 15706
rect 57888 15642 57940 15648
rect 57520 15360 57572 15366
rect 57520 15302 57572 15308
rect 57428 14816 57480 14822
rect 57428 14758 57480 14764
rect 57440 11801 57468 14758
rect 57532 14074 57560 15302
rect 58176 14822 58204 16594
rect 58268 15570 58296 17478
rect 58726 17436 59034 17445
rect 58726 17434 58732 17436
rect 58788 17434 58812 17436
rect 58868 17434 58892 17436
rect 58948 17434 58972 17436
rect 59028 17434 59034 17436
rect 58788 17382 58790 17434
rect 58970 17382 58972 17434
rect 58726 17380 58732 17382
rect 58788 17380 58812 17382
rect 58868 17380 58892 17382
rect 58948 17380 58972 17382
rect 59028 17380 59034 17382
rect 58726 17371 59034 17380
rect 58726 16348 59034 16357
rect 58726 16346 58732 16348
rect 58788 16346 58812 16348
rect 58868 16346 58892 16348
rect 58948 16346 58972 16348
rect 59028 16346 59034 16348
rect 58788 16294 58790 16346
rect 58970 16294 58972 16346
rect 58726 16292 58732 16294
rect 58788 16292 58812 16294
rect 58868 16292 58892 16294
rect 58948 16292 58972 16294
rect 59028 16292 59034 16294
rect 58726 16283 59034 16292
rect 58256 15564 58308 15570
rect 58256 15506 58308 15512
rect 58726 15260 59034 15269
rect 58726 15258 58732 15260
rect 58788 15258 58812 15260
rect 58868 15258 58892 15260
rect 58948 15258 58972 15260
rect 59028 15258 59034 15260
rect 58788 15206 58790 15258
rect 58970 15206 58972 15258
rect 58726 15204 58732 15206
rect 58788 15204 58812 15206
rect 58868 15204 58892 15206
rect 58948 15204 58972 15206
rect 59028 15204 59034 15206
rect 58726 15195 59034 15204
rect 58164 14816 58216 14822
rect 58164 14758 58216 14764
rect 58440 14408 58492 14414
rect 58440 14350 58492 14356
rect 57520 14068 57572 14074
rect 57520 14010 57572 14016
rect 57888 13728 57940 13734
rect 57888 13670 57940 13676
rect 57900 13326 57928 13670
rect 58452 13530 58480 14350
rect 58726 14172 59034 14181
rect 58726 14170 58732 14172
rect 58788 14170 58812 14172
rect 58868 14170 58892 14172
rect 58948 14170 58972 14172
rect 59028 14170 59034 14172
rect 58788 14118 58790 14170
rect 58970 14118 58972 14170
rect 58726 14116 58732 14118
rect 58788 14116 58812 14118
rect 58868 14116 58892 14118
rect 58948 14116 58972 14118
rect 59028 14116 59034 14118
rect 58726 14107 59034 14116
rect 58440 13524 58492 13530
rect 58440 13466 58492 13472
rect 57888 13320 57940 13326
rect 57888 13262 57940 13268
rect 58452 12434 58480 13466
rect 58726 13084 59034 13093
rect 58726 13082 58732 13084
rect 58788 13082 58812 13084
rect 58868 13082 58892 13084
rect 58948 13082 58972 13084
rect 59028 13082 59034 13084
rect 58788 13030 58790 13082
rect 58970 13030 58972 13082
rect 58726 13028 58732 13030
rect 58788 13028 58812 13030
rect 58868 13028 58892 13030
rect 58948 13028 58972 13030
rect 59028 13028 59034 13030
rect 58726 13019 59034 13028
rect 57992 12406 58480 12434
rect 57520 12096 57572 12102
rect 57520 12038 57572 12044
rect 57426 11792 57482 11801
rect 57426 11727 57482 11736
rect 57532 11694 57560 12038
rect 57428 11688 57480 11694
rect 57348 11636 57428 11642
rect 57348 11630 57480 11636
rect 57520 11688 57572 11694
rect 57520 11630 57572 11636
rect 57348 11614 57468 11630
rect 57060 11348 57112 11354
rect 57060 11290 57112 11296
rect 57336 11008 57388 11014
rect 57336 10950 57388 10956
rect 57348 10690 57376 10950
rect 57164 10662 57376 10690
rect 56968 9580 57020 9586
rect 56968 9522 57020 9528
rect 56876 9376 56928 9382
rect 56876 9318 56928 9324
rect 56888 9178 56916 9318
rect 56876 9172 56928 9178
rect 56876 9114 56928 9120
rect 56692 9036 56744 9042
rect 56692 8978 56744 8984
rect 56600 8900 56652 8906
rect 56600 8842 56652 8848
rect 56612 8430 56640 8842
rect 57060 8560 57112 8566
rect 57060 8502 57112 8508
rect 56692 8492 56744 8498
rect 56692 8434 56744 8440
rect 56600 8424 56652 8430
rect 56600 8366 56652 8372
rect 56232 8288 56284 8294
rect 56232 8230 56284 8236
rect 55956 7880 56008 7886
rect 55956 7822 56008 7828
rect 55968 7002 55996 7822
rect 56244 7410 56272 8230
rect 56612 8090 56640 8366
rect 56600 8084 56652 8090
rect 56600 8026 56652 8032
rect 56416 7880 56468 7886
rect 56416 7822 56468 7828
rect 56324 7540 56376 7546
rect 56324 7482 56376 7488
rect 56336 7410 56364 7482
rect 56232 7404 56284 7410
rect 56232 7346 56284 7352
rect 56324 7404 56376 7410
rect 56324 7346 56376 7352
rect 55956 6996 56008 7002
rect 55956 6938 56008 6944
rect 56140 6792 56192 6798
rect 56140 6734 56192 6740
rect 55864 5704 55916 5710
rect 55864 5646 55916 5652
rect 55956 5704 56008 5710
rect 55956 5646 56008 5652
rect 55876 5370 55904 5646
rect 55968 5370 55996 5646
rect 56048 5568 56100 5574
rect 56048 5510 56100 5516
rect 55864 5364 55916 5370
rect 55864 5306 55916 5312
rect 55956 5364 56008 5370
rect 55956 5306 56008 5312
rect 56060 5302 56088 5510
rect 56152 5370 56180 6734
rect 56140 5364 56192 5370
rect 56140 5306 56192 5312
rect 56048 5296 56100 5302
rect 56048 5238 56100 5244
rect 56244 5114 56272 7346
rect 56324 7200 56376 7206
rect 56324 7142 56376 7148
rect 56060 5086 56272 5114
rect 56060 4078 56088 5086
rect 56336 4690 56364 7142
rect 56428 6798 56456 7822
rect 56508 7404 56560 7410
rect 56508 7346 56560 7352
rect 56416 6792 56468 6798
rect 56416 6734 56468 6740
rect 56520 6730 56548 7346
rect 56508 6724 56560 6730
rect 56508 6666 56560 6672
rect 56416 6452 56468 6458
rect 56520 6440 56548 6666
rect 56468 6412 56548 6440
rect 56416 6394 56468 6400
rect 56704 5370 56732 8434
rect 56784 8288 56836 8294
rect 56784 8230 56836 8236
rect 56796 7886 56824 8230
rect 56784 7880 56836 7886
rect 56784 7822 56836 7828
rect 56876 7200 56928 7206
rect 56876 7142 56928 7148
rect 56888 6254 56916 7142
rect 57072 6662 57100 8502
rect 57164 6882 57192 10662
rect 57336 10600 57388 10606
rect 57336 10542 57388 10548
rect 57348 9722 57376 10542
rect 57440 10418 57468 11614
rect 57532 10674 57560 11630
rect 57520 10668 57572 10674
rect 57520 10610 57572 10616
rect 57888 10464 57940 10470
rect 57440 10390 57560 10418
rect 57888 10406 57940 10412
rect 57336 9716 57388 9722
rect 57336 9658 57388 9664
rect 57336 9512 57388 9518
rect 57336 9454 57388 9460
rect 57428 9512 57480 9518
rect 57428 9454 57480 9460
rect 57244 8492 57296 8498
rect 57244 8434 57296 8440
rect 57256 7410 57284 8434
rect 57348 7478 57376 9454
rect 57440 8430 57468 9454
rect 57428 8424 57480 8430
rect 57428 8366 57480 8372
rect 57440 7886 57468 8366
rect 57428 7880 57480 7886
rect 57428 7822 57480 7828
rect 57336 7472 57388 7478
rect 57336 7414 57388 7420
rect 57244 7404 57296 7410
rect 57244 7346 57296 7352
rect 57336 7336 57388 7342
rect 57336 7278 57388 7284
rect 57164 6854 57284 6882
rect 57060 6656 57112 6662
rect 57060 6598 57112 6604
rect 57072 6458 57100 6598
rect 57060 6452 57112 6458
rect 57060 6394 57112 6400
rect 56876 6248 56928 6254
rect 56876 6190 56928 6196
rect 56784 5568 56836 5574
rect 56784 5510 56836 5516
rect 56692 5364 56744 5370
rect 56692 5306 56744 5312
rect 56508 5228 56560 5234
rect 56508 5170 56560 5176
rect 56324 4684 56376 4690
rect 56324 4626 56376 4632
rect 56140 4548 56192 4554
rect 56140 4490 56192 4496
rect 56152 4282 56180 4490
rect 56140 4276 56192 4282
rect 56140 4218 56192 4224
rect 56048 4072 56100 4078
rect 56048 4014 56100 4020
rect 56140 4004 56192 4010
rect 56140 3946 56192 3952
rect 56152 3194 56180 3946
rect 56520 3738 56548 5170
rect 56692 5160 56744 5166
rect 56692 5102 56744 5108
rect 56508 3732 56560 3738
rect 56508 3674 56560 3680
rect 56520 3194 56548 3674
rect 56704 3466 56732 5102
rect 56600 3460 56652 3466
rect 56600 3402 56652 3408
rect 56692 3460 56744 3466
rect 56692 3402 56744 3408
rect 56140 3188 56192 3194
rect 56140 3130 56192 3136
rect 56508 3188 56560 3194
rect 56612 3176 56640 3402
rect 56692 3188 56744 3194
rect 56612 3148 56692 3176
rect 56508 3130 56560 3136
rect 56692 3130 56744 3136
rect 56796 3126 56824 5510
rect 57152 4548 57204 4554
rect 57152 4490 57204 4496
rect 56784 3120 56836 3126
rect 56784 3062 56836 3068
rect 55784 2746 56088 2774
rect 54760 2440 54812 2446
rect 54760 2382 54812 2388
rect 55220 2372 55272 2378
rect 55220 2314 55272 2320
rect 55232 800 55260 2314
rect 56060 800 56088 2746
rect 56888 870 57008 898
rect 56888 800 56916 870
rect 51184 734 51396 762
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53562 0 53618 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56874 0 56930 800
rect 56980 762 57008 870
rect 57164 762 57192 4490
rect 57256 2446 57284 6854
rect 57348 6254 57376 7278
rect 57532 7206 57560 10390
rect 57612 9988 57664 9994
rect 57612 9930 57664 9936
rect 57624 9178 57652 9930
rect 57612 9172 57664 9178
rect 57612 9114 57664 9120
rect 57704 8832 57756 8838
rect 57704 8774 57756 8780
rect 57520 7200 57572 7206
rect 57520 7142 57572 7148
rect 57428 6792 57480 6798
rect 57428 6734 57480 6740
rect 57440 6458 57468 6734
rect 57428 6452 57480 6458
rect 57428 6394 57480 6400
rect 57336 6248 57388 6254
rect 57336 6190 57388 6196
rect 57716 5794 57744 8774
rect 57796 6656 57848 6662
rect 57796 6598 57848 6604
rect 57808 6458 57836 6598
rect 57796 6452 57848 6458
rect 57796 6394 57848 6400
rect 57624 5766 57744 5794
rect 57336 5704 57388 5710
rect 57336 5646 57388 5652
rect 57348 2650 57376 5646
rect 57428 3460 57480 3466
rect 57428 3402 57480 3408
rect 57440 3369 57468 3402
rect 57426 3360 57482 3369
rect 57426 3295 57482 3304
rect 57336 2644 57388 2650
rect 57336 2586 57388 2592
rect 57440 2514 57468 3295
rect 57624 2514 57652 5766
rect 57796 5704 57848 5710
rect 57796 5646 57848 5652
rect 57704 5024 57756 5030
rect 57704 4966 57756 4972
rect 57716 3534 57744 4966
rect 57808 3670 57836 5646
rect 57900 5370 57928 10406
rect 57888 5364 57940 5370
rect 57888 5306 57940 5312
rect 57888 5160 57940 5166
rect 57888 5102 57940 5108
rect 57900 3738 57928 5102
rect 57992 4146 58020 12406
rect 58726 11996 59034 12005
rect 58726 11994 58732 11996
rect 58788 11994 58812 11996
rect 58868 11994 58892 11996
rect 58948 11994 58972 11996
rect 59028 11994 59034 11996
rect 58788 11942 58790 11994
rect 58970 11942 58972 11994
rect 58726 11940 58732 11942
rect 58788 11940 58812 11942
rect 58868 11940 58892 11942
rect 58948 11940 58972 11942
rect 59028 11940 59034 11942
rect 58726 11931 59034 11940
rect 58726 10908 59034 10917
rect 58726 10906 58732 10908
rect 58788 10906 58812 10908
rect 58868 10906 58892 10908
rect 58948 10906 58972 10908
rect 59028 10906 59034 10908
rect 58788 10854 58790 10906
rect 58970 10854 58972 10906
rect 58726 10852 58732 10854
rect 58788 10852 58812 10854
rect 58868 10852 58892 10854
rect 58948 10852 58972 10854
rect 59028 10852 59034 10854
rect 58726 10843 59034 10852
rect 58440 10600 58492 10606
rect 58492 10560 58572 10588
rect 58440 10542 58492 10548
rect 58164 9920 58216 9926
rect 58164 9862 58216 9868
rect 58176 9586 58204 9862
rect 58164 9580 58216 9586
rect 58164 9522 58216 9528
rect 58256 8968 58308 8974
rect 58256 8910 58308 8916
rect 58164 5568 58216 5574
rect 58164 5510 58216 5516
rect 58072 4480 58124 4486
rect 58072 4422 58124 4428
rect 57980 4140 58032 4146
rect 57980 4082 58032 4088
rect 57888 3732 57940 3738
rect 57888 3674 57940 3680
rect 57796 3664 57848 3670
rect 57796 3606 57848 3612
rect 57704 3528 57756 3534
rect 57704 3470 57756 3476
rect 57704 3392 57756 3398
rect 57704 3334 57756 3340
rect 57428 2508 57480 2514
rect 57428 2450 57480 2456
rect 57612 2508 57664 2514
rect 57612 2450 57664 2456
rect 57244 2440 57296 2446
rect 57244 2382 57296 2388
rect 57716 800 57744 3334
rect 57808 2650 57836 3606
rect 58084 3534 58112 4422
rect 58176 3602 58204 5510
rect 58268 4622 58296 8910
rect 58440 8424 58492 8430
rect 58440 8366 58492 8372
rect 58452 8090 58480 8366
rect 58440 8084 58492 8090
rect 58440 8026 58492 8032
rect 58440 7404 58492 7410
rect 58440 7346 58492 7352
rect 58256 4616 58308 4622
rect 58256 4558 58308 4564
rect 58164 3596 58216 3602
rect 58164 3538 58216 3544
rect 58072 3528 58124 3534
rect 58072 3470 58124 3476
rect 58268 2990 58296 4558
rect 58348 4072 58400 4078
rect 58348 4014 58400 4020
rect 58256 2984 58308 2990
rect 58256 2926 58308 2932
rect 57796 2644 57848 2650
rect 57796 2586 57848 2592
rect 58360 2122 58388 4014
rect 58452 4010 58480 7346
rect 58440 4004 58492 4010
rect 58440 3946 58492 3952
rect 58544 3398 58572 10560
rect 58726 9820 59034 9829
rect 58726 9818 58732 9820
rect 58788 9818 58812 9820
rect 58868 9818 58892 9820
rect 58948 9818 58972 9820
rect 59028 9818 59034 9820
rect 58788 9766 58790 9818
rect 58970 9766 58972 9818
rect 58726 9764 58732 9766
rect 58788 9764 58812 9766
rect 58868 9764 58892 9766
rect 58948 9764 58972 9766
rect 59028 9764 59034 9766
rect 58726 9755 59034 9764
rect 58726 8732 59034 8741
rect 58726 8730 58732 8732
rect 58788 8730 58812 8732
rect 58868 8730 58892 8732
rect 58948 8730 58972 8732
rect 59028 8730 59034 8732
rect 58788 8678 58790 8730
rect 58970 8678 58972 8730
rect 58726 8676 58732 8678
rect 58788 8676 58812 8678
rect 58868 8676 58892 8678
rect 58948 8676 58972 8678
rect 59028 8676 59034 8678
rect 58726 8667 59034 8676
rect 58726 7644 59034 7653
rect 58726 7642 58732 7644
rect 58788 7642 58812 7644
rect 58868 7642 58892 7644
rect 58948 7642 58972 7644
rect 59028 7642 59034 7644
rect 58788 7590 58790 7642
rect 58970 7590 58972 7642
rect 58726 7588 58732 7590
rect 58788 7588 58812 7590
rect 58868 7588 58892 7590
rect 58948 7588 58972 7590
rect 59028 7588 59034 7590
rect 58726 7579 59034 7588
rect 58726 6556 59034 6565
rect 58726 6554 58732 6556
rect 58788 6554 58812 6556
rect 58868 6554 58892 6556
rect 58948 6554 58972 6556
rect 59028 6554 59034 6556
rect 58788 6502 58790 6554
rect 58970 6502 58972 6554
rect 58726 6500 58732 6502
rect 58788 6500 58812 6502
rect 58868 6500 58892 6502
rect 58948 6500 58972 6502
rect 59028 6500 59034 6502
rect 58726 6491 59034 6500
rect 58726 5468 59034 5477
rect 58726 5466 58732 5468
rect 58788 5466 58812 5468
rect 58868 5466 58892 5468
rect 58948 5466 58972 5468
rect 59028 5466 59034 5468
rect 58788 5414 58790 5466
rect 58970 5414 58972 5466
rect 58726 5412 58732 5414
rect 58788 5412 58812 5414
rect 58868 5412 58892 5414
rect 58948 5412 58972 5414
rect 59028 5412 59034 5414
rect 58726 5403 59034 5412
rect 58726 4380 59034 4389
rect 58726 4378 58732 4380
rect 58788 4378 58812 4380
rect 58868 4378 58892 4380
rect 58948 4378 58972 4380
rect 59028 4378 59034 4380
rect 58788 4326 58790 4378
rect 58970 4326 58972 4378
rect 58726 4324 58732 4326
rect 58788 4324 58812 4326
rect 58868 4324 58892 4326
rect 58948 4324 58972 4326
rect 59028 4324 59034 4326
rect 58726 4315 59034 4324
rect 58532 3392 58584 3398
rect 58532 3334 58584 3340
rect 58726 3292 59034 3301
rect 58726 3290 58732 3292
rect 58788 3290 58812 3292
rect 58868 3290 58892 3292
rect 58948 3290 58972 3292
rect 59028 3290 59034 3292
rect 58788 3238 58790 3290
rect 58970 3238 58972 3290
rect 58726 3236 58732 3238
rect 58788 3236 58812 3238
rect 58868 3236 58892 3238
rect 58948 3236 58972 3238
rect 59028 3236 59034 3238
rect 58726 3227 59034 3236
rect 58438 2816 58494 2825
rect 58438 2751 58494 2760
rect 58452 2514 58480 2751
rect 58440 2508 58492 2514
rect 58440 2450 58492 2456
rect 58726 2204 59034 2213
rect 58726 2202 58732 2204
rect 58788 2202 58812 2204
rect 58868 2202 58892 2204
rect 58948 2202 58972 2204
rect 59028 2202 59034 2204
rect 58788 2150 58790 2202
rect 58970 2150 58972 2202
rect 58726 2148 58732 2150
rect 58788 2148 58812 2150
rect 58868 2148 58892 2150
rect 58948 2148 58972 2150
rect 59028 2148 59034 2150
rect 58726 2139 59034 2148
rect 58360 2094 58572 2122
rect 58544 800 58572 2094
rect 56980 734 57192 762
rect 57702 0 57758 800
rect 58530 0 58586 800
<< via2 >>
rect 8178 27770 8234 27772
rect 8258 27770 8314 27772
rect 8338 27770 8394 27772
rect 8418 27770 8474 27772
rect 8178 27718 8224 27770
rect 8224 27718 8234 27770
rect 8258 27718 8288 27770
rect 8288 27718 8300 27770
rect 8300 27718 8314 27770
rect 8338 27718 8352 27770
rect 8352 27718 8364 27770
rect 8364 27718 8394 27770
rect 8418 27718 8428 27770
rect 8428 27718 8474 27770
rect 8178 27716 8234 27718
rect 8258 27716 8314 27718
rect 8338 27716 8394 27718
rect 8418 27716 8474 27718
rect 22622 27770 22678 27772
rect 22702 27770 22758 27772
rect 22782 27770 22838 27772
rect 22862 27770 22918 27772
rect 22622 27718 22668 27770
rect 22668 27718 22678 27770
rect 22702 27718 22732 27770
rect 22732 27718 22744 27770
rect 22744 27718 22758 27770
rect 22782 27718 22796 27770
rect 22796 27718 22808 27770
rect 22808 27718 22838 27770
rect 22862 27718 22872 27770
rect 22872 27718 22918 27770
rect 22622 27716 22678 27718
rect 22702 27716 22758 27718
rect 22782 27716 22838 27718
rect 22862 27716 22918 27718
rect 37066 27770 37122 27772
rect 37146 27770 37202 27772
rect 37226 27770 37282 27772
rect 37306 27770 37362 27772
rect 37066 27718 37112 27770
rect 37112 27718 37122 27770
rect 37146 27718 37176 27770
rect 37176 27718 37188 27770
rect 37188 27718 37202 27770
rect 37226 27718 37240 27770
rect 37240 27718 37252 27770
rect 37252 27718 37282 27770
rect 37306 27718 37316 27770
rect 37316 27718 37362 27770
rect 37066 27716 37122 27718
rect 37146 27716 37202 27718
rect 37226 27716 37282 27718
rect 37306 27716 37362 27718
rect 51510 27770 51566 27772
rect 51590 27770 51646 27772
rect 51670 27770 51726 27772
rect 51750 27770 51806 27772
rect 51510 27718 51556 27770
rect 51556 27718 51566 27770
rect 51590 27718 51620 27770
rect 51620 27718 51632 27770
rect 51632 27718 51646 27770
rect 51670 27718 51684 27770
rect 51684 27718 51696 27770
rect 51696 27718 51726 27770
rect 51750 27718 51760 27770
rect 51760 27718 51806 27770
rect 51510 27716 51566 27718
rect 51590 27716 51646 27718
rect 51670 27716 51726 27718
rect 51750 27716 51806 27718
rect 15400 27226 15456 27228
rect 15480 27226 15536 27228
rect 15560 27226 15616 27228
rect 15640 27226 15696 27228
rect 15400 27174 15446 27226
rect 15446 27174 15456 27226
rect 15480 27174 15510 27226
rect 15510 27174 15522 27226
rect 15522 27174 15536 27226
rect 15560 27174 15574 27226
rect 15574 27174 15586 27226
rect 15586 27174 15616 27226
rect 15640 27174 15650 27226
rect 15650 27174 15696 27226
rect 15400 27172 15456 27174
rect 15480 27172 15536 27174
rect 15560 27172 15616 27174
rect 15640 27172 15696 27174
rect 29844 27226 29900 27228
rect 29924 27226 29980 27228
rect 30004 27226 30060 27228
rect 30084 27226 30140 27228
rect 29844 27174 29890 27226
rect 29890 27174 29900 27226
rect 29924 27174 29954 27226
rect 29954 27174 29966 27226
rect 29966 27174 29980 27226
rect 30004 27174 30018 27226
rect 30018 27174 30030 27226
rect 30030 27174 30060 27226
rect 30084 27174 30094 27226
rect 30094 27174 30140 27226
rect 29844 27172 29900 27174
rect 29924 27172 29980 27174
rect 30004 27172 30060 27174
rect 30084 27172 30140 27174
rect 44288 27226 44344 27228
rect 44368 27226 44424 27228
rect 44448 27226 44504 27228
rect 44528 27226 44584 27228
rect 44288 27174 44334 27226
rect 44334 27174 44344 27226
rect 44368 27174 44398 27226
rect 44398 27174 44410 27226
rect 44410 27174 44424 27226
rect 44448 27174 44462 27226
rect 44462 27174 44474 27226
rect 44474 27174 44504 27226
rect 44528 27174 44538 27226
rect 44538 27174 44584 27226
rect 44288 27172 44344 27174
rect 44368 27172 44424 27174
rect 44448 27172 44504 27174
rect 44528 27172 44584 27174
rect 58732 27226 58788 27228
rect 58812 27226 58868 27228
rect 58892 27226 58948 27228
rect 58972 27226 59028 27228
rect 58732 27174 58778 27226
rect 58778 27174 58788 27226
rect 58812 27174 58842 27226
rect 58842 27174 58854 27226
rect 58854 27174 58868 27226
rect 58892 27174 58906 27226
rect 58906 27174 58918 27226
rect 58918 27174 58948 27226
rect 58972 27174 58982 27226
rect 58982 27174 59028 27226
rect 58732 27172 58788 27174
rect 58812 27172 58868 27174
rect 58892 27172 58948 27174
rect 58972 27172 59028 27174
rect 8178 26682 8234 26684
rect 8258 26682 8314 26684
rect 8338 26682 8394 26684
rect 8418 26682 8474 26684
rect 8178 26630 8224 26682
rect 8224 26630 8234 26682
rect 8258 26630 8288 26682
rect 8288 26630 8300 26682
rect 8300 26630 8314 26682
rect 8338 26630 8352 26682
rect 8352 26630 8364 26682
rect 8364 26630 8394 26682
rect 8418 26630 8428 26682
rect 8428 26630 8474 26682
rect 8178 26628 8234 26630
rect 8258 26628 8314 26630
rect 8338 26628 8394 26630
rect 8418 26628 8474 26630
rect 22622 26682 22678 26684
rect 22702 26682 22758 26684
rect 22782 26682 22838 26684
rect 22862 26682 22918 26684
rect 22622 26630 22668 26682
rect 22668 26630 22678 26682
rect 22702 26630 22732 26682
rect 22732 26630 22744 26682
rect 22744 26630 22758 26682
rect 22782 26630 22796 26682
rect 22796 26630 22808 26682
rect 22808 26630 22838 26682
rect 22862 26630 22872 26682
rect 22872 26630 22918 26682
rect 22622 26628 22678 26630
rect 22702 26628 22758 26630
rect 22782 26628 22838 26630
rect 22862 26628 22918 26630
rect 37066 26682 37122 26684
rect 37146 26682 37202 26684
rect 37226 26682 37282 26684
rect 37306 26682 37362 26684
rect 37066 26630 37112 26682
rect 37112 26630 37122 26682
rect 37146 26630 37176 26682
rect 37176 26630 37188 26682
rect 37188 26630 37202 26682
rect 37226 26630 37240 26682
rect 37240 26630 37252 26682
rect 37252 26630 37282 26682
rect 37306 26630 37316 26682
rect 37316 26630 37362 26682
rect 37066 26628 37122 26630
rect 37146 26628 37202 26630
rect 37226 26628 37282 26630
rect 37306 26628 37362 26630
rect 51510 26682 51566 26684
rect 51590 26682 51646 26684
rect 51670 26682 51726 26684
rect 51750 26682 51806 26684
rect 51510 26630 51556 26682
rect 51556 26630 51566 26682
rect 51590 26630 51620 26682
rect 51620 26630 51632 26682
rect 51632 26630 51646 26682
rect 51670 26630 51684 26682
rect 51684 26630 51696 26682
rect 51696 26630 51726 26682
rect 51750 26630 51760 26682
rect 51760 26630 51806 26682
rect 51510 26628 51566 26630
rect 51590 26628 51646 26630
rect 51670 26628 51726 26630
rect 51750 26628 51806 26630
rect 15400 26138 15456 26140
rect 15480 26138 15536 26140
rect 15560 26138 15616 26140
rect 15640 26138 15696 26140
rect 15400 26086 15446 26138
rect 15446 26086 15456 26138
rect 15480 26086 15510 26138
rect 15510 26086 15522 26138
rect 15522 26086 15536 26138
rect 15560 26086 15574 26138
rect 15574 26086 15586 26138
rect 15586 26086 15616 26138
rect 15640 26086 15650 26138
rect 15650 26086 15696 26138
rect 15400 26084 15456 26086
rect 15480 26084 15536 26086
rect 15560 26084 15616 26086
rect 15640 26084 15696 26086
rect 29844 26138 29900 26140
rect 29924 26138 29980 26140
rect 30004 26138 30060 26140
rect 30084 26138 30140 26140
rect 29844 26086 29890 26138
rect 29890 26086 29900 26138
rect 29924 26086 29954 26138
rect 29954 26086 29966 26138
rect 29966 26086 29980 26138
rect 30004 26086 30018 26138
rect 30018 26086 30030 26138
rect 30030 26086 30060 26138
rect 30084 26086 30094 26138
rect 30094 26086 30140 26138
rect 29844 26084 29900 26086
rect 29924 26084 29980 26086
rect 30004 26084 30060 26086
rect 30084 26084 30140 26086
rect 44288 26138 44344 26140
rect 44368 26138 44424 26140
rect 44448 26138 44504 26140
rect 44528 26138 44584 26140
rect 44288 26086 44334 26138
rect 44334 26086 44344 26138
rect 44368 26086 44398 26138
rect 44398 26086 44410 26138
rect 44410 26086 44424 26138
rect 44448 26086 44462 26138
rect 44462 26086 44474 26138
rect 44474 26086 44504 26138
rect 44528 26086 44538 26138
rect 44538 26086 44584 26138
rect 44288 26084 44344 26086
rect 44368 26084 44424 26086
rect 44448 26084 44504 26086
rect 44528 26084 44584 26086
rect 58732 26138 58788 26140
rect 58812 26138 58868 26140
rect 58892 26138 58948 26140
rect 58972 26138 59028 26140
rect 58732 26086 58778 26138
rect 58778 26086 58788 26138
rect 58812 26086 58842 26138
rect 58842 26086 58854 26138
rect 58854 26086 58868 26138
rect 58892 26086 58906 26138
rect 58906 26086 58918 26138
rect 58918 26086 58948 26138
rect 58972 26086 58982 26138
rect 58982 26086 59028 26138
rect 58732 26084 58788 26086
rect 58812 26084 58868 26086
rect 58892 26084 58948 26086
rect 58972 26084 59028 26086
rect 8178 25594 8234 25596
rect 8258 25594 8314 25596
rect 8338 25594 8394 25596
rect 8418 25594 8474 25596
rect 8178 25542 8224 25594
rect 8224 25542 8234 25594
rect 8258 25542 8288 25594
rect 8288 25542 8300 25594
rect 8300 25542 8314 25594
rect 8338 25542 8352 25594
rect 8352 25542 8364 25594
rect 8364 25542 8394 25594
rect 8418 25542 8428 25594
rect 8428 25542 8474 25594
rect 8178 25540 8234 25542
rect 8258 25540 8314 25542
rect 8338 25540 8394 25542
rect 8418 25540 8474 25542
rect 22622 25594 22678 25596
rect 22702 25594 22758 25596
rect 22782 25594 22838 25596
rect 22862 25594 22918 25596
rect 22622 25542 22668 25594
rect 22668 25542 22678 25594
rect 22702 25542 22732 25594
rect 22732 25542 22744 25594
rect 22744 25542 22758 25594
rect 22782 25542 22796 25594
rect 22796 25542 22808 25594
rect 22808 25542 22838 25594
rect 22862 25542 22872 25594
rect 22872 25542 22918 25594
rect 22622 25540 22678 25542
rect 22702 25540 22758 25542
rect 22782 25540 22838 25542
rect 22862 25540 22918 25542
rect 37066 25594 37122 25596
rect 37146 25594 37202 25596
rect 37226 25594 37282 25596
rect 37306 25594 37362 25596
rect 37066 25542 37112 25594
rect 37112 25542 37122 25594
rect 37146 25542 37176 25594
rect 37176 25542 37188 25594
rect 37188 25542 37202 25594
rect 37226 25542 37240 25594
rect 37240 25542 37252 25594
rect 37252 25542 37282 25594
rect 37306 25542 37316 25594
rect 37316 25542 37362 25594
rect 37066 25540 37122 25542
rect 37146 25540 37202 25542
rect 37226 25540 37282 25542
rect 37306 25540 37362 25542
rect 51510 25594 51566 25596
rect 51590 25594 51646 25596
rect 51670 25594 51726 25596
rect 51750 25594 51806 25596
rect 51510 25542 51556 25594
rect 51556 25542 51566 25594
rect 51590 25542 51620 25594
rect 51620 25542 51632 25594
rect 51632 25542 51646 25594
rect 51670 25542 51684 25594
rect 51684 25542 51696 25594
rect 51696 25542 51726 25594
rect 51750 25542 51760 25594
rect 51760 25542 51806 25594
rect 51510 25540 51566 25542
rect 51590 25540 51646 25542
rect 51670 25540 51726 25542
rect 51750 25540 51806 25542
rect 15400 25050 15456 25052
rect 15480 25050 15536 25052
rect 15560 25050 15616 25052
rect 15640 25050 15696 25052
rect 15400 24998 15446 25050
rect 15446 24998 15456 25050
rect 15480 24998 15510 25050
rect 15510 24998 15522 25050
rect 15522 24998 15536 25050
rect 15560 24998 15574 25050
rect 15574 24998 15586 25050
rect 15586 24998 15616 25050
rect 15640 24998 15650 25050
rect 15650 24998 15696 25050
rect 15400 24996 15456 24998
rect 15480 24996 15536 24998
rect 15560 24996 15616 24998
rect 15640 24996 15696 24998
rect 29844 25050 29900 25052
rect 29924 25050 29980 25052
rect 30004 25050 30060 25052
rect 30084 25050 30140 25052
rect 29844 24998 29890 25050
rect 29890 24998 29900 25050
rect 29924 24998 29954 25050
rect 29954 24998 29966 25050
rect 29966 24998 29980 25050
rect 30004 24998 30018 25050
rect 30018 24998 30030 25050
rect 30030 24998 30060 25050
rect 30084 24998 30094 25050
rect 30094 24998 30140 25050
rect 29844 24996 29900 24998
rect 29924 24996 29980 24998
rect 30004 24996 30060 24998
rect 30084 24996 30140 24998
rect 44288 25050 44344 25052
rect 44368 25050 44424 25052
rect 44448 25050 44504 25052
rect 44528 25050 44584 25052
rect 44288 24998 44334 25050
rect 44334 24998 44344 25050
rect 44368 24998 44398 25050
rect 44398 24998 44410 25050
rect 44410 24998 44424 25050
rect 44448 24998 44462 25050
rect 44462 24998 44474 25050
rect 44474 24998 44504 25050
rect 44528 24998 44538 25050
rect 44538 24998 44584 25050
rect 44288 24996 44344 24998
rect 44368 24996 44424 24998
rect 44448 24996 44504 24998
rect 44528 24996 44584 24998
rect 58732 25050 58788 25052
rect 58812 25050 58868 25052
rect 58892 25050 58948 25052
rect 58972 25050 59028 25052
rect 58732 24998 58778 25050
rect 58778 24998 58788 25050
rect 58812 24998 58842 25050
rect 58842 24998 58854 25050
rect 58854 24998 58868 25050
rect 58892 24998 58906 25050
rect 58906 24998 58918 25050
rect 58918 24998 58948 25050
rect 58972 24998 58982 25050
rect 58982 24998 59028 25050
rect 58732 24996 58788 24998
rect 58812 24996 58868 24998
rect 58892 24996 58948 24998
rect 58972 24996 59028 24998
rect 8178 24506 8234 24508
rect 8258 24506 8314 24508
rect 8338 24506 8394 24508
rect 8418 24506 8474 24508
rect 8178 24454 8224 24506
rect 8224 24454 8234 24506
rect 8258 24454 8288 24506
rect 8288 24454 8300 24506
rect 8300 24454 8314 24506
rect 8338 24454 8352 24506
rect 8352 24454 8364 24506
rect 8364 24454 8394 24506
rect 8418 24454 8428 24506
rect 8428 24454 8474 24506
rect 8178 24452 8234 24454
rect 8258 24452 8314 24454
rect 8338 24452 8394 24454
rect 8418 24452 8474 24454
rect 22622 24506 22678 24508
rect 22702 24506 22758 24508
rect 22782 24506 22838 24508
rect 22862 24506 22918 24508
rect 22622 24454 22668 24506
rect 22668 24454 22678 24506
rect 22702 24454 22732 24506
rect 22732 24454 22744 24506
rect 22744 24454 22758 24506
rect 22782 24454 22796 24506
rect 22796 24454 22808 24506
rect 22808 24454 22838 24506
rect 22862 24454 22872 24506
rect 22872 24454 22918 24506
rect 22622 24452 22678 24454
rect 22702 24452 22758 24454
rect 22782 24452 22838 24454
rect 22862 24452 22918 24454
rect 37066 24506 37122 24508
rect 37146 24506 37202 24508
rect 37226 24506 37282 24508
rect 37306 24506 37362 24508
rect 37066 24454 37112 24506
rect 37112 24454 37122 24506
rect 37146 24454 37176 24506
rect 37176 24454 37188 24506
rect 37188 24454 37202 24506
rect 37226 24454 37240 24506
rect 37240 24454 37252 24506
rect 37252 24454 37282 24506
rect 37306 24454 37316 24506
rect 37316 24454 37362 24506
rect 37066 24452 37122 24454
rect 37146 24452 37202 24454
rect 37226 24452 37282 24454
rect 37306 24452 37362 24454
rect 51510 24506 51566 24508
rect 51590 24506 51646 24508
rect 51670 24506 51726 24508
rect 51750 24506 51806 24508
rect 51510 24454 51556 24506
rect 51556 24454 51566 24506
rect 51590 24454 51620 24506
rect 51620 24454 51632 24506
rect 51632 24454 51646 24506
rect 51670 24454 51684 24506
rect 51684 24454 51696 24506
rect 51696 24454 51726 24506
rect 51750 24454 51760 24506
rect 51760 24454 51806 24506
rect 51510 24452 51566 24454
rect 51590 24452 51646 24454
rect 51670 24452 51726 24454
rect 51750 24452 51806 24454
rect 15400 23962 15456 23964
rect 15480 23962 15536 23964
rect 15560 23962 15616 23964
rect 15640 23962 15696 23964
rect 15400 23910 15446 23962
rect 15446 23910 15456 23962
rect 15480 23910 15510 23962
rect 15510 23910 15522 23962
rect 15522 23910 15536 23962
rect 15560 23910 15574 23962
rect 15574 23910 15586 23962
rect 15586 23910 15616 23962
rect 15640 23910 15650 23962
rect 15650 23910 15696 23962
rect 15400 23908 15456 23910
rect 15480 23908 15536 23910
rect 15560 23908 15616 23910
rect 15640 23908 15696 23910
rect 29844 23962 29900 23964
rect 29924 23962 29980 23964
rect 30004 23962 30060 23964
rect 30084 23962 30140 23964
rect 29844 23910 29890 23962
rect 29890 23910 29900 23962
rect 29924 23910 29954 23962
rect 29954 23910 29966 23962
rect 29966 23910 29980 23962
rect 30004 23910 30018 23962
rect 30018 23910 30030 23962
rect 30030 23910 30060 23962
rect 30084 23910 30094 23962
rect 30094 23910 30140 23962
rect 29844 23908 29900 23910
rect 29924 23908 29980 23910
rect 30004 23908 30060 23910
rect 30084 23908 30140 23910
rect 44288 23962 44344 23964
rect 44368 23962 44424 23964
rect 44448 23962 44504 23964
rect 44528 23962 44584 23964
rect 44288 23910 44334 23962
rect 44334 23910 44344 23962
rect 44368 23910 44398 23962
rect 44398 23910 44410 23962
rect 44410 23910 44424 23962
rect 44448 23910 44462 23962
rect 44462 23910 44474 23962
rect 44474 23910 44504 23962
rect 44528 23910 44538 23962
rect 44538 23910 44584 23962
rect 44288 23908 44344 23910
rect 44368 23908 44424 23910
rect 44448 23908 44504 23910
rect 44528 23908 44584 23910
rect 58732 23962 58788 23964
rect 58812 23962 58868 23964
rect 58892 23962 58948 23964
rect 58972 23962 59028 23964
rect 58732 23910 58778 23962
rect 58778 23910 58788 23962
rect 58812 23910 58842 23962
rect 58842 23910 58854 23962
rect 58854 23910 58868 23962
rect 58892 23910 58906 23962
rect 58906 23910 58918 23962
rect 58918 23910 58948 23962
rect 58972 23910 58982 23962
rect 58982 23910 59028 23962
rect 58732 23908 58788 23910
rect 58812 23908 58868 23910
rect 58892 23908 58948 23910
rect 58972 23908 59028 23910
rect 8178 23418 8234 23420
rect 8258 23418 8314 23420
rect 8338 23418 8394 23420
rect 8418 23418 8474 23420
rect 8178 23366 8224 23418
rect 8224 23366 8234 23418
rect 8258 23366 8288 23418
rect 8288 23366 8300 23418
rect 8300 23366 8314 23418
rect 8338 23366 8352 23418
rect 8352 23366 8364 23418
rect 8364 23366 8394 23418
rect 8418 23366 8428 23418
rect 8428 23366 8474 23418
rect 8178 23364 8234 23366
rect 8258 23364 8314 23366
rect 8338 23364 8394 23366
rect 8418 23364 8474 23366
rect 8178 22330 8234 22332
rect 8258 22330 8314 22332
rect 8338 22330 8394 22332
rect 8418 22330 8474 22332
rect 8178 22278 8224 22330
rect 8224 22278 8234 22330
rect 8258 22278 8288 22330
rect 8288 22278 8300 22330
rect 8300 22278 8314 22330
rect 8338 22278 8352 22330
rect 8352 22278 8364 22330
rect 8364 22278 8394 22330
rect 8418 22278 8428 22330
rect 8428 22278 8474 22330
rect 8178 22276 8234 22278
rect 8258 22276 8314 22278
rect 8338 22276 8394 22278
rect 8418 22276 8474 22278
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 6550 19352 6606 19408
rect 1398 3440 1454 3496
rect 3974 4936 4030 4992
rect 5354 3984 5410 4040
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 7286 15000 7342 15056
rect 5906 4120 5962 4176
rect 7010 11756 7066 11792
rect 7010 11736 7012 11756
rect 7012 11736 7064 11756
rect 7064 11736 7066 11756
rect 7562 12300 7618 12336
rect 7562 12280 7564 12300
rect 7564 12280 7616 12300
rect 7616 12280 7618 12300
rect 7102 11076 7158 11112
rect 7102 11056 7104 11076
rect 7104 11056 7156 11076
rect 7156 11056 7158 11076
rect 15400 22874 15456 22876
rect 15480 22874 15536 22876
rect 15560 22874 15616 22876
rect 15640 22874 15696 22876
rect 15400 22822 15446 22874
rect 15446 22822 15456 22874
rect 15480 22822 15510 22874
rect 15510 22822 15522 22874
rect 15522 22822 15536 22874
rect 15560 22822 15574 22874
rect 15574 22822 15586 22874
rect 15586 22822 15616 22874
rect 15640 22822 15650 22874
rect 15650 22822 15696 22874
rect 15400 22820 15456 22822
rect 15480 22820 15536 22822
rect 15560 22820 15616 22822
rect 15640 22820 15696 22822
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 7930 15000 7986 15056
rect 6642 4156 6644 4176
rect 6644 4156 6696 4176
rect 6696 4156 6698 4176
rect 6642 4120 6698 4156
rect 5998 2916 6054 2952
rect 5998 2896 6000 2916
rect 6000 2896 6052 2916
rect 6052 2896 6054 2916
rect 7746 4972 7748 4992
rect 7748 4972 7800 4992
rect 7800 4972 7802 4992
rect 7746 4936 7802 4972
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 9586 15544 9642 15600
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 9218 12688 9274 12744
rect 10138 11192 10194 11248
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 10414 12844 10470 12880
rect 10414 12824 10416 12844
rect 10416 12824 10468 12844
rect 10468 12824 10470 12844
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 7470 2896 7526 2952
rect 12990 13252 13046 13288
rect 12990 13232 12992 13252
rect 12992 13232 13044 13252
rect 13044 13232 13046 13252
rect 13726 13388 13782 13424
rect 13726 13368 13728 13388
rect 13728 13368 13780 13388
rect 13780 13368 13782 13388
rect 12898 12280 12954 12336
rect 12990 6840 13046 6896
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 15400 21786 15456 21788
rect 15480 21786 15536 21788
rect 15560 21786 15616 21788
rect 15640 21786 15696 21788
rect 15400 21734 15446 21786
rect 15446 21734 15456 21786
rect 15480 21734 15510 21786
rect 15510 21734 15522 21786
rect 15522 21734 15536 21786
rect 15560 21734 15574 21786
rect 15574 21734 15586 21786
rect 15586 21734 15616 21786
rect 15640 21734 15650 21786
rect 15650 21734 15696 21786
rect 15400 21732 15456 21734
rect 15480 21732 15536 21734
rect 15560 21732 15616 21734
rect 15640 21732 15696 21734
rect 15400 20698 15456 20700
rect 15480 20698 15536 20700
rect 15560 20698 15616 20700
rect 15640 20698 15696 20700
rect 15400 20646 15446 20698
rect 15446 20646 15456 20698
rect 15480 20646 15510 20698
rect 15510 20646 15522 20698
rect 15522 20646 15536 20698
rect 15560 20646 15574 20698
rect 15574 20646 15586 20698
rect 15586 20646 15616 20698
rect 15640 20646 15650 20698
rect 15650 20646 15696 20698
rect 15400 20644 15456 20646
rect 15480 20644 15536 20646
rect 15560 20644 15616 20646
rect 15640 20644 15696 20646
rect 15400 19610 15456 19612
rect 15480 19610 15536 19612
rect 15560 19610 15616 19612
rect 15640 19610 15696 19612
rect 15400 19558 15446 19610
rect 15446 19558 15456 19610
rect 15480 19558 15510 19610
rect 15510 19558 15522 19610
rect 15522 19558 15536 19610
rect 15560 19558 15574 19610
rect 15574 19558 15586 19610
rect 15586 19558 15616 19610
rect 15640 19558 15650 19610
rect 15650 19558 15696 19610
rect 15400 19556 15456 19558
rect 15480 19556 15536 19558
rect 15560 19556 15616 19558
rect 15640 19556 15696 19558
rect 15400 18522 15456 18524
rect 15480 18522 15536 18524
rect 15560 18522 15616 18524
rect 15640 18522 15696 18524
rect 15400 18470 15446 18522
rect 15446 18470 15456 18522
rect 15480 18470 15510 18522
rect 15510 18470 15522 18522
rect 15522 18470 15536 18522
rect 15560 18470 15574 18522
rect 15574 18470 15586 18522
rect 15586 18470 15616 18522
rect 15640 18470 15650 18522
rect 15650 18470 15696 18522
rect 15400 18468 15456 18470
rect 15480 18468 15536 18470
rect 15560 18468 15616 18470
rect 15640 18468 15696 18470
rect 15400 17434 15456 17436
rect 15480 17434 15536 17436
rect 15560 17434 15616 17436
rect 15640 17434 15696 17436
rect 15400 17382 15446 17434
rect 15446 17382 15456 17434
rect 15480 17382 15510 17434
rect 15510 17382 15522 17434
rect 15522 17382 15536 17434
rect 15560 17382 15574 17434
rect 15574 17382 15586 17434
rect 15586 17382 15616 17434
rect 15640 17382 15650 17434
rect 15650 17382 15696 17434
rect 15400 17380 15456 17382
rect 15480 17380 15536 17382
rect 15560 17380 15616 17382
rect 15640 17380 15696 17382
rect 15400 16346 15456 16348
rect 15480 16346 15536 16348
rect 15560 16346 15616 16348
rect 15640 16346 15696 16348
rect 15400 16294 15446 16346
rect 15446 16294 15456 16346
rect 15480 16294 15510 16346
rect 15510 16294 15522 16346
rect 15522 16294 15536 16346
rect 15560 16294 15574 16346
rect 15574 16294 15586 16346
rect 15586 16294 15616 16346
rect 15640 16294 15650 16346
rect 15650 16294 15696 16346
rect 15400 16292 15456 16294
rect 15480 16292 15536 16294
rect 15560 16292 15616 16294
rect 15640 16292 15696 16294
rect 15400 15258 15456 15260
rect 15480 15258 15536 15260
rect 15560 15258 15616 15260
rect 15640 15258 15696 15260
rect 15400 15206 15446 15258
rect 15446 15206 15456 15258
rect 15480 15206 15510 15258
rect 15510 15206 15522 15258
rect 15522 15206 15536 15258
rect 15560 15206 15574 15258
rect 15574 15206 15586 15258
rect 15586 15206 15616 15258
rect 15640 15206 15650 15258
rect 15650 15206 15696 15258
rect 15400 15204 15456 15206
rect 15480 15204 15536 15206
rect 15560 15204 15616 15206
rect 15640 15204 15696 15206
rect 15400 14170 15456 14172
rect 15480 14170 15536 14172
rect 15560 14170 15616 14172
rect 15640 14170 15696 14172
rect 15400 14118 15446 14170
rect 15446 14118 15456 14170
rect 15480 14118 15510 14170
rect 15510 14118 15522 14170
rect 15522 14118 15536 14170
rect 15560 14118 15574 14170
rect 15574 14118 15586 14170
rect 15586 14118 15616 14170
rect 15640 14118 15650 14170
rect 15650 14118 15696 14170
rect 15400 14116 15456 14118
rect 15480 14116 15536 14118
rect 15560 14116 15616 14118
rect 15640 14116 15696 14118
rect 16486 20748 16488 20768
rect 16488 20748 16540 20768
rect 16540 20748 16542 20768
rect 16486 20712 16542 20748
rect 22622 23418 22678 23420
rect 22702 23418 22758 23420
rect 22782 23418 22838 23420
rect 22862 23418 22918 23420
rect 22622 23366 22668 23418
rect 22668 23366 22678 23418
rect 22702 23366 22732 23418
rect 22732 23366 22744 23418
rect 22744 23366 22758 23418
rect 22782 23366 22796 23418
rect 22796 23366 22808 23418
rect 22808 23366 22838 23418
rect 22862 23366 22872 23418
rect 22872 23366 22918 23418
rect 22622 23364 22678 23366
rect 22702 23364 22758 23366
rect 22782 23364 22838 23366
rect 22862 23364 22918 23366
rect 37066 23418 37122 23420
rect 37146 23418 37202 23420
rect 37226 23418 37282 23420
rect 37306 23418 37362 23420
rect 37066 23366 37112 23418
rect 37112 23366 37122 23418
rect 37146 23366 37176 23418
rect 37176 23366 37188 23418
rect 37188 23366 37202 23418
rect 37226 23366 37240 23418
rect 37240 23366 37252 23418
rect 37252 23366 37282 23418
rect 37306 23366 37316 23418
rect 37316 23366 37362 23418
rect 37066 23364 37122 23366
rect 37146 23364 37202 23366
rect 37226 23364 37282 23366
rect 37306 23364 37362 23366
rect 15400 13082 15456 13084
rect 15480 13082 15536 13084
rect 15560 13082 15616 13084
rect 15640 13082 15696 13084
rect 15400 13030 15446 13082
rect 15446 13030 15456 13082
rect 15480 13030 15510 13082
rect 15510 13030 15522 13082
rect 15522 13030 15536 13082
rect 15560 13030 15574 13082
rect 15574 13030 15586 13082
rect 15586 13030 15616 13082
rect 15640 13030 15650 13082
rect 15650 13030 15696 13082
rect 15400 13028 15456 13030
rect 15480 13028 15536 13030
rect 15560 13028 15616 13030
rect 15640 13028 15696 13030
rect 15400 11994 15456 11996
rect 15480 11994 15536 11996
rect 15560 11994 15616 11996
rect 15640 11994 15696 11996
rect 15400 11942 15446 11994
rect 15446 11942 15456 11994
rect 15480 11942 15510 11994
rect 15510 11942 15522 11994
rect 15522 11942 15536 11994
rect 15560 11942 15574 11994
rect 15574 11942 15586 11994
rect 15586 11942 15616 11994
rect 15640 11942 15650 11994
rect 15650 11942 15696 11994
rect 15400 11940 15456 11942
rect 15480 11940 15536 11942
rect 15560 11940 15616 11942
rect 15640 11940 15696 11942
rect 15400 10906 15456 10908
rect 15480 10906 15536 10908
rect 15560 10906 15616 10908
rect 15640 10906 15696 10908
rect 15400 10854 15446 10906
rect 15446 10854 15456 10906
rect 15480 10854 15510 10906
rect 15510 10854 15522 10906
rect 15522 10854 15536 10906
rect 15560 10854 15574 10906
rect 15574 10854 15586 10906
rect 15586 10854 15616 10906
rect 15640 10854 15650 10906
rect 15650 10854 15696 10906
rect 15400 10852 15456 10854
rect 15480 10852 15536 10854
rect 15560 10852 15616 10854
rect 15640 10852 15696 10854
rect 15400 9818 15456 9820
rect 15480 9818 15536 9820
rect 15560 9818 15616 9820
rect 15640 9818 15696 9820
rect 15400 9766 15446 9818
rect 15446 9766 15456 9818
rect 15480 9766 15510 9818
rect 15510 9766 15522 9818
rect 15522 9766 15536 9818
rect 15560 9766 15574 9818
rect 15574 9766 15586 9818
rect 15586 9766 15616 9818
rect 15640 9766 15650 9818
rect 15650 9766 15696 9818
rect 15400 9764 15456 9766
rect 15480 9764 15536 9766
rect 15560 9764 15616 9766
rect 15640 9764 15696 9766
rect 15400 8730 15456 8732
rect 15480 8730 15536 8732
rect 15560 8730 15616 8732
rect 15640 8730 15696 8732
rect 15400 8678 15446 8730
rect 15446 8678 15456 8730
rect 15480 8678 15510 8730
rect 15510 8678 15522 8730
rect 15522 8678 15536 8730
rect 15560 8678 15574 8730
rect 15574 8678 15586 8730
rect 15586 8678 15616 8730
rect 15640 8678 15650 8730
rect 15650 8678 15696 8730
rect 15400 8676 15456 8678
rect 15480 8676 15536 8678
rect 15560 8676 15616 8678
rect 15640 8676 15696 8678
rect 15400 7642 15456 7644
rect 15480 7642 15536 7644
rect 15560 7642 15616 7644
rect 15640 7642 15696 7644
rect 15400 7590 15446 7642
rect 15446 7590 15456 7642
rect 15480 7590 15510 7642
rect 15510 7590 15522 7642
rect 15522 7590 15536 7642
rect 15560 7590 15574 7642
rect 15574 7590 15586 7642
rect 15586 7590 15616 7642
rect 15640 7590 15650 7642
rect 15650 7590 15696 7642
rect 15400 7588 15456 7590
rect 15480 7588 15536 7590
rect 15560 7588 15616 7590
rect 15640 7588 15696 7590
rect 15382 6876 15384 6896
rect 15384 6876 15436 6896
rect 15436 6876 15438 6896
rect 15382 6840 15438 6876
rect 15400 6554 15456 6556
rect 15480 6554 15536 6556
rect 15560 6554 15616 6556
rect 15640 6554 15696 6556
rect 15400 6502 15446 6554
rect 15446 6502 15456 6554
rect 15480 6502 15510 6554
rect 15510 6502 15522 6554
rect 15522 6502 15536 6554
rect 15560 6502 15574 6554
rect 15574 6502 15586 6554
rect 15586 6502 15616 6554
rect 15640 6502 15650 6554
rect 15650 6502 15696 6554
rect 15400 6500 15456 6502
rect 15480 6500 15536 6502
rect 15560 6500 15616 6502
rect 15640 6500 15696 6502
rect 15400 5466 15456 5468
rect 15480 5466 15536 5468
rect 15560 5466 15616 5468
rect 15640 5466 15696 5468
rect 15400 5414 15446 5466
rect 15446 5414 15456 5466
rect 15480 5414 15510 5466
rect 15510 5414 15522 5466
rect 15522 5414 15536 5466
rect 15560 5414 15574 5466
rect 15574 5414 15586 5466
rect 15586 5414 15616 5466
rect 15640 5414 15650 5466
rect 15650 5414 15696 5466
rect 15400 5412 15456 5414
rect 15480 5412 15536 5414
rect 15560 5412 15616 5414
rect 15640 5412 15696 5414
rect 15400 4378 15456 4380
rect 15480 4378 15536 4380
rect 15560 4378 15616 4380
rect 15640 4378 15696 4380
rect 15400 4326 15446 4378
rect 15446 4326 15456 4378
rect 15480 4326 15510 4378
rect 15510 4326 15522 4378
rect 15522 4326 15536 4378
rect 15560 4326 15574 4378
rect 15574 4326 15586 4378
rect 15586 4326 15616 4378
rect 15640 4326 15650 4378
rect 15650 4326 15696 4378
rect 15400 4324 15456 4326
rect 15480 4324 15536 4326
rect 15560 4324 15616 4326
rect 15640 4324 15696 4326
rect 15400 3290 15456 3292
rect 15480 3290 15536 3292
rect 15560 3290 15616 3292
rect 15640 3290 15696 3292
rect 15400 3238 15446 3290
rect 15446 3238 15456 3290
rect 15480 3238 15510 3290
rect 15510 3238 15522 3290
rect 15522 3238 15536 3290
rect 15560 3238 15574 3290
rect 15574 3238 15586 3290
rect 15586 3238 15616 3290
rect 15640 3238 15650 3290
rect 15650 3238 15696 3290
rect 15400 3236 15456 3238
rect 15480 3236 15536 3238
rect 15560 3236 15616 3238
rect 15640 3236 15696 3238
rect 15400 2202 15456 2204
rect 15480 2202 15536 2204
rect 15560 2202 15616 2204
rect 15640 2202 15696 2204
rect 15400 2150 15446 2202
rect 15446 2150 15456 2202
rect 15480 2150 15510 2202
rect 15510 2150 15522 2202
rect 15522 2150 15536 2202
rect 15560 2150 15574 2202
rect 15574 2150 15586 2202
rect 15586 2150 15616 2202
rect 15640 2150 15650 2202
rect 15650 2150 15696 2202
rect 15400 2148 15456 2150
rect 15480 2148 15536 2150
rect 15560 2148 15616 2150
rect 15640 2148 15696 2150
rect 22622 22330 22678 22332
rect 22702 22330 22758 22332
rect 22782 22330 22838 22332
rect 22862 22330 22918 22332
rect 22622 22278 22668 22330
rect 22668 22278 22678 22330
rect 22702 22278 22732 22330
rect 22732 22278 22744 22330
rect 22744 22278 22758 22330
rect 22782 22278 22796 22330
rect 22796 22278 22808 22330
rect 22808 22278 22838 22330
rect 22862 22278 22872 22330
rect 22872 22278 22918 22330
rect 22622 22276 22678 22278
rect 22702 22276 22758 22278
rect 22782 22276 22838 22278
rect 22862 22276 22918 22278
rect 29844 22874 29900 22876
rect 29924 22874 29980 22876
rect 30004 22874 30060 22876
rect 30084 22874 30140 22876
rect 29844 22822 29890 22874
rect 29890 22822 29900 22874
rect 29924 22822 29954 22874
rect 29954 22822 29966 22874
rect 29966 22822 29980 22874
rect 30004 22822 30018 22874
rect 30018 22822 30030 22874
rect 30030 22822 30060 22874
rect 30084 22822 30094 22874
rect 30094 22822 30140 22874
rect 29844 22820 29900 22822
rect 29924 22820 29980 22822
rect 30004 22820 30060 22822
rect 30084 22820 30140 22822
rect 22622 21242 22678 21244
rect 22702 21242 22758 21244
rect 22782 21242 22838 21244
rect 22862 21242 22918 21244
rect 22622 21190 22668 21242
rect 22668 21190 22678 21242
rect 22702 21190 22732 21242
rect 22732 21190 22744 21242
rect 22744 21190 22758 21242
rect 22782 21190 22796 21242
rect 22796 21190 22808 21242
rect 22808 21190 22838 21242
rect 22862 21190 22872 21242
rect 22872 21190 22918 21242
rect 22622 21188 22678 21190
rect 22702 21188 22758 21190
rect 22782 21188 22838 21190
rect 22862 21188 22918 21190
rect 22622 20154 22678 20156
rect 22702 20154 22758 20156
rect 22782 20154 22838 20156
rect 22862 20154 22918 20156
rect 22622 20102 22668 20154
rect 22668 20102 22678 20154
rect 22702 20102 22732 20154
rect 22732 20102 22744 20154
rect 22744 20102 22758 20154
rect 22782 20102 22796 20154
rect 22796 20102 22808 20154
rect 22808 20102 22838 20154
rect 22862 20102 22872 20154
rect 22872 20102 22918 20154
rect 22622 20100 22678 20102
rect 22702 20100 22758 20102
rect 22782 20100 22838 20102
rect 22862 20100 22918 20102
rect 17498 6976 17554 7032
rect 16854 3984 16910 4040
rect 19522 3984 19578 4040
rect 22622 19066 22678 19068
rect 22702 19066 22758 19068
rect 22782 19066 22838 19068
rect 22862 19066 22918 19068
rect 22622 19014 22668 19066
rect 22668 19014 22678 19066
rect 22702 19014 22732 19066
rect 22732 19014 22744 19066
rect 22744 19014 22758 19066
rect 22782 19014 22796 19066
rect 22796 19014 22808 19066
rect 22808 19014 22838 19066
rect 22862 19014 22872 19066
rect 22872 19014 22918 19066
rect 22622 19012 22678 19014
rect 22702 19012 22758 19014
rect 22782 19012 22838 19014
rect 22862 19012 22918 19014
rect 27434 21664 27490 21720
rect 22622 17978 22678 17980
rect 22702 17978 22758 17980
rect 22782 17978 22838 17980
rect 22862 17978 22918 17980
rect 22622 17926 22668 17978
rect 22668 17926 22678 17978
rect 22702 17926 22732 17978
rect 22732 17926 22744 17978
rect 22744 17926 22758 17978
rect 22782 17926 22796 17978
rect 22796 17926 22808 17978
rect 22808 17926 22838 17978
rect 22862 17926 22872 17978
rect 22872 17926 22918 17978
rect 22622 17924 22678 17926
rect 22702 17924 22758 17926
rect 22782 17924 22838 17926
rect 22862 17924 22918 17926
rect 22622 16890 22678 16892
rect 22702 16890 22758 16892
rect 22782 16890 22838 16892
rect 22862 16890 22918 16892
rect 22622 16838 22668 16890
rect 22668 16838 22678 16890
rect 22702 16838 22732 16890
rect 22732 16838 22744 16890
rect 22744 16838 22758 16890
rect 22782 16838 22796 16890
rect 22796 16838 22808 16890
rect 22808 16838 22838 16890
rect 22862 16838 22872 16890
rect 22872 16838 22918 16890
rect 22622 16836 22678 16838
rect 22702 16836 22758 16838
rect 22782 16836 22838 16838
rect 22862 16836 22918 16838
rect 22622 15802 22678 15804
rect 22702 15802 22758 15804
rect 22782 15802 22838 15804
rect 22862 15802 22918 15804
rect 22622 15750 22668 15802
rect 22668 15750 22678 15802
rect 22702 15750 22732 15802
rect 22732 15750 22744 15802
rect 22744 15750 22758 15802
rect 22782 15750 22796 15802
rect 22796 15750 22808 15802
rect 22808 15750 22838 15802
rect 22862 15750 22872 15802
rect 22872 15750 22918 15802
rect 22622 15748 22678 15750
rect 22702 15748 22758 15750
rect 22782 15748 22838 15750
rect 22862 15748 22918 15750
rect 22622 14714 22678 14716
rect 22702 14714 22758 14716
rect 22782 14714 22838 14716
rect 22862 14714 22918 14716
rect 22622 14662 22668 14714
rect 22668 14662 22678 14714
rect 22702 14662 22732 14714
rect 22732 14662 22744 14714
rect 22744 14662 22758 14714
rect 22782 14662 22796 14714
rect 22796 14662 22808 14714
rect 22808 14662 22838 14714
rect 22862 14662 22872 14714
rect 22872 14662 22918 14714
rect 22622 14660 22678 14662
rect 22702 14660 22758 14662
rect 22782 14660 22838 14662
rect 22862 14660 22918 14662
rect 22622 13626 22678 13628
rect 22702 13626 22758 13628
rect 22782 13626 22838 13628
rect 22862 13626 22918 13628
rect 22622 13574 22668 13626
rect 22668 13574 22678 13626
rect 22702 13574 22732 13626
rect 22732 13574 22744 13626
rect 22744 13574 22758 13626
rect 22782 13574 22796 13626
rect 22796 13574 22808 13626
rect 22808 13574 22838 13626
rect 22862 13574 22872 13626
rect 22872 13574 22918 13626
rect 22622 13572 22678 13574
rect 22702 13572 22758 13574
rect 22782 13572 22838 13574
rect 22862 13572 22918 13574
rect 23294 13524 23350 13560
rect 23294 13504 23296 13524
rect 23296 13504 23348 13524
rect 23348 13504 23350 13524
rect 22622 12538 22678 12540
rect 22702 12538 22758 12540
rect 22782 12538 22838 12540
rect 22862 12538 22918 12540
rect 22622 12486 22668 12538
rect 22668 12486 22678 12538
rect 22702 12486 22732 12538
rect 22732 12486 22744 12538
rect 22744 12486 22758 12538
rect 22782 12486 22796 12538
rect 22796 12486 22808 12538
rect 22808 12486 22838 12538
rect 22862 12486 22872 12538
rect 22872 12486 22918 12538
rect 22622 12484 22678 12486
rect 22702 12484 22758 12486
rect 22782 12484 22838 12486
rect 22862 12484 22918 12486
rect 22622 11450 22678 11452
rect 22702 11450 22758 11452
rect 22782 11450 22838 11452
rect 22862 11450 22918 11452
rect 22622 11398 22668 11450
rect 22668 11398 22678 11450
rect 22702 11398 22732 11450
rect 22732 11398 22744 11450
rect 22744 11398 22758 11450
rect 22782 11398 22796 11450
rect 22796 11398 22808 11450
rect 22808 11398 22838 11450
rect 22862 11398 22872 11450
rect 22872 11398 22918 11450
rect 22622 11396 22678 11398
rect 22702 11396 22758 11398
rect 22782 11396 22838 11398
rect 22862 11396 22918 11398
rect 22622 10362 22678 10364
rect 22702 10362 22758 10364
rect 22782 10362 22838 10364
rect 22862 10362 22918 10364
rect 22622 10310 22668 10362
rect 22668 10310 22678 10362
rect 22702 10310 22732 10362
rect 22732 10310 22744 10362
rect 22744 10310 22758 10362
rect 22782 10310 22796 10362
rect 22796 10310 22808 10362
rect 22808 10310 22838 10362
rect 22862 10310 22872 10362
rect 22872 10310 22918 10362
rect 22622 10308 22678 10310
rect 22702 10308 22758 10310
rect 22782 10308 22838 10310
rect 22862 10308 22918 10310
rect 22622 9274 22678 9276
rect 22702 9274 22758 9276
rect 22782 9274 22838 9276
rect 22862 9274 22918 9276
rect 22622 9222 22668 9274
rect 22668 9222 22678 9274
rect 22702 9222 22732 9274
rect 22732 9222 22744 9274
rect 22744 9222 22758 9274
rect 22782 9222 22796 9274
rect 22796 9222 22808 9274
rect 22808 9222 22838 9274
rect 22862 9222 22872 9274
rect 22872 9222 22918 9274
rect 22622 9220 22678 9222
rect 22702 9220 22758 9222
rect 22782 9220 22838 9222
rect 22862 9220 22918 9222
rect 22622 8186 22678 8188
rect 22702 8186 22758 8188
rect 22782 8186 22838 8188
rect 22862 8186 22918 8188
rect 22622 8134 22668 8186
rect 22668 8134 22678 8186
rect 22702 8134 22732 8186
rect 22732 8134 22744 8186
rect 22744 8134 22758 8186
rect 22782 8134 22796 8186
rect 22796 8134 22808 8186
rect 22808 8134 22838 8186
rect 22862 8134 22872 8186
rect 22872 8134 22918 8186
rect 22622 8132 22678 8134
rect 22702 8132 22758 8134
rect 22782 8132 22838 8134
rect 22862 8132 22918 8134
rect 22622 7098 22678 7100
rect 22702 7098 22758 7100
rect 22782 7098 22838 7100
rect 22862 7098 22918 7100
rect 22622 7046 22668 7098
rect 22668 7046 22678 7098
rect 22702 7046 22732 7098
rect 22732 7046 22744 7098
rect 22744 7046 22758 7098
rect 22782 7046 22796 7098
rect 22796 7046 22808 7098
rect 22808 7046 22838 7098
rect 22862 7046 22872 7098
rect 22872 7046 22918 7098
rect 22622 7044 22678 7046
rect 22702 7044 22758 7046
rect 22782 7044 22838 7046
rect 22862 7044 22918 7046
rect 22622 6010 22678 6012
rect 22702 6010 22758 6012
rect 22782 6010 22838 6012
rect 22862 6010 22918 6012
rect 22622 5958 22668 6010
rect 22668 5958 22678 6010
rect 22702 5958 22732 6010
rect 22732 5958 22744 6010
rect 22744 5958 22758 6010
rect 22782 5958 22796 6010
rect 22796 5958 22808 6010
rect 22808 5958 22838 6010
rect 22862 5958 22872 6010
rect 22872 5958 22918 6010
rect 22622 5956 22678 5958
rect 22702 5956 22758 5958
rect 22782 5956 22838 5958
rect 22862 5956 22918 5958
rect 22622 4922 22678 4924
rect 22702 4922 22758 4924
rect 22782 4922 22838 4924
rect 22862 4922 22918 4924
rect 22622 4870 22668 4922
rect 22668 4870 22678 4922
rect 22702 4870 22732 4922
rect 22732 4870 22744 4922
rect 22744 4870 22758 4922
rect 22782 4870 22796 4922
rect 22796 4870 22808 4922
rect 22808 4870 22838 4922
rect 22862 4870 22872 4922
rect 22872 4870 22918 4922
rect 22622 4868 22678 4870
rect 22702 4868 22758 4870
rect 22782 4868 22838 4870
rect 22862 4868 22918 4870
rect 22622 3834 22678 3836
rect 22702 3834 22758 3836
rect 22782 3834 22838 3836
rect 22862 3834 22918 3836
rect 22622 3782 22668 3834
rect 22668 3782 22678 3834
rect 22702 3782 22732 3834
rect 22732 3782 22744 3834
rect 22744 3782 22758 3834
rect 22782 3782 22796 3834
rect 22796 3782 22808 3834
rect 22808 3782 22838 3834
rect 22862 3782 22872 3834
rect 22872 3782 22918 3834
rect 22622 3780 22678 3782
rect 22702 3780 22758 3782
rect 22782 3780 22838 3782
rect 22862 3780 22918 3782
rect 26330 15544 26386 15600
rect 28078 21664 28134 21720
rect 27618 18148 27674 18184
rect 27618 18128 27620 18148
rect 27620 18128 27672 18148
rect 27672 18128 27674 18148
rect 29844 21786 29900 21788
rect 29924 21786 29980 21788
rect 30004 21786 30060 21788
rect 30084 21786 30140 21788
rect 29844 21734 29890 21786
rect 29890 21734 29900 21786
rect 29924 21734 29954 21786
rect 29954 21734 29966 21786
rect 29966 21734 29980 21786
rect 30004 21734 30018 21786
rect 30018 21734 30030 21786
rect 30030 21734 30060 21786
rect 30084 21734 30094 21786
rect 30094 21734 30140 21786
rect 29844 21732 29900 21734
rect 29924 21732 29980 21734
rect 30004 21732 30060 21734
rect 30084 21732 30140 21734
rect 28354 18164 28356 18184
rect 28356 18164 28408 18184
rect 28408 18164 28410 18184
rect 28354 18128 28410 18164
rect 26238 13504 26294 13560
rect 22622 2746 22678 2748
rect 22702 2746 22758 2748
rect 22782 2746 22838 2748
rect 22862 2746 22918 2748
rect 22622 2694 22668 2746
rect 22668 2694 22678 2746
rect 22702 2694 22732 2746
rect 22732 2694 22744 2746
rect 22744 2694 22758 2746
rect 22782 2694 22796 2746
rect 22796 2694 22808 2746
rect 22808 2694 22838 2746
rect 22862 2694 22872 2746
rect 22872 2694 22918 2746
rect 22622 2692 22678 2694
rect 22702 2692 22758 2694
rect 22782 2692 22838 2694
rect 22862 2692 22918 2694
rect 29844 20698 29900 20700
rect 29924 20698 29980 20700
rect 30004 20698 30060 20700
rect 30084 20698 30140 20700
rect 29844 20646 29890 20698
rect 29890 20646 29900 20698
rect 29924 20646 29954 20698
rect 29954 20646 29966 20698
rect 29966 20646 29980 20698
rect 30004 20646 30018 20698
rect 30018 20646 30030 20698
rect 30030 20646 30060 20698
rect 30084 20646 30094 20698
rect 30094 20646 30140 20698
rect 29844 20644 29900 20646
rect 29924 20644 29980 20646
rect 30004 20644 30060 20646
rect 30084 20644 30140 20646
rect 29844 19610 29900 19612
rect 29924 19610 29980 19612
rect 30004 19610 30060 19612
rect 30084 19610 30140 19612
rect 29844 19558 29890 19610
rect 29890 19558 29900 19610
rect 29924 19558 29954 19610
rect 29954 19558 29966 19610
rect 29966 19558 29980 19610
rect 30004 19558 30018 19610
rect 30018 19558 30030 19610
rect 30030 19558 30060 19610
rect 30084 19558 30094 19610
rect 30094 19558 30140 19610
rect 29844 19556 29900 19558
rect 29924 19556 29980 19558
rect 30004 19556 30060 19558
rect 30084 19556 30140 19558
rect 29844 18522 29900 18524
rect 29924 18522 29980 18524
rect 30004 18522 30060 18524
rect 30084 18522 30140 18524
rect 29844 18470 29890 18522
rect 29890 18470 29900 18522
rect 29924 18470 29954 18522
rect 29954 18470 29966 18522
rect 29966 18470 29980 18522
rect 30004 18470 30018 18522
rect 30018 18470 30030 18522
rect 30030 18470 30060 18522
rect 30084 18470 30094 18522
rect 30094 18470 30140 18522
rect 29844 18468 29900 18470
rect 29924 18468 29980 18470
rect 30004 18468 30060 18470
rect 30084 18468 30140 18470
rect 32218 21392 32274 21448
rect 31390 18672 31446 18728
rect 29844 17434 29900 17436
rect 29924 17434 29980 17436
rect 30004 17434 30060 17436
rect 30084 17434 30140 17436
rect 29844 17382 29890 17434
rect 29890 17382 29900 17434
rect 29924 17382 29954 17434
rect 29954 17382 29966 17434
rect 29966 17382 29980 17434
rect 30004 17382 30018 17434
rect 30018 17382 30030 17434
rect 30030 17382 30060 17434
rect 30084 17382 30094 17434
rect 30094 17382 30140 17434
rect 29844 17380 29900 17382
rect 29924 17380 29980 17382
rect 30004 17380 30060 17382
rect 30084 17380 30140 17382
rect 29844 16346 29900 16348
rect 29924 16346 29980 16348
rect 30004 16346 30060 16348
rect 30084 16346 30140 16348
rect 29844 16294 29890 16346
rect 29890 16294 29900 16346
rect 29924 16294 29954 16346
rect 29954 16294 29966 16346
rect 29966 16294 29980 16346
rect 30004 16294 30018 16346
rect 30018 16294 30030 16346
rect 30030 16294 30060 16346
rect 30084 16294 30094 16346
rect 30094 16294 30140 16346
rect 29844 16292 29900 16294
rect 29924 16292 29980 16294
rect 30004 16292 30060 16294
rect 30084 16292 30140 16294
rect 32770 21392 32826 21448
rect 29844 15258 29900 15260
rect 29924 15258 29980 15260
rect 30004 15258 30060 15260
rect 30084 15258 30140 15260
rect 29844 15206 29890 15258
rect 29890 15206 29900 15258
rect 29924 15206 29954 15258
rect 29954 15206 29966 15258
rect 29966 15206 29980 15258
rect 30004 15206 30018 15258
rect 30018 15206 30030 15258
rect 30030 15206 30060 15258
rect 30084 15206 30094 15258
rect 30094 15206 30140 15258
rect 29844 15204 29900 15206
rect 29924 15204 29980 15206
rect 30004 15204 30060 15206
rect 30084 15204 30140 15206
rect 29844 14170 29900 14172
rect 29924 14170 29980 14172
rect 30004 14170 30060 14172
rect 30084 14170 30140 14172
rect 29844 14118 29890 14170
rect 29890 14118 29900 14170
rect 29924 14118 29954 14170
rect 29954 14118 29966 14170
rect 29966 14118 29980 14170
rect 30004 14118 30018 14170
rect 30018 14118 30030 14170
rect 30030 14118 30060 14170
rect 30084 14118 30094 14170
rect 30094 14118 30140 14170
rect 29844 14116 29900 14118
rect 29924 14116 29980 14118
rect 30004 14116 30060 14118
rect 30084 14116 30140 14118
rect 29844 13082 29900 13084
rect 29924 13082 29980 13084
rect 30004 13082 30060 13084
rect 30084 13082 30140 13084
rect 29844 13030 29890 13082
rect 29890 13030 29900 13082
rect 29924 13030 29954 13082
rect 29954 13030 29966 13082
rect 29966 13030 29980 13082
rect 30004 13030 30018 13082
rect 30018 13030 30030 13082
rect 30030 13030 30060 13082
rect 30084 13030 30094 13082
rect 30094 13030 30140 13082
rect 29844 13028 29900 13030
rect 29924 13028 29980 13030
rect 30004 13028 30060 13030
rect 30084 13028 30140 13030
rect 30378 12180 30380 12200
rect 30380 12180 30432 12200
rect 30432 12180 30434 12200
rect 30378 12144 30434 12180
rect 29844 11994 29900 11996
rect 29924 11994 29980 11996
rect 30004 11994 30060 11996
rect 30084 11994 30140 11996
rect 29844 11942 29890 11994
rect 29890 11942 29900 11994
rect 29924 11942 29954 11994
rect 29954 11942 29966 11994
rect 29966 11942 29980 11994
rect 30004 11942 30018 11994
rect 30018 11942 30030 11994
rect 30030 11942 30060 11994
rect 30084 11942 30094 11994
rect 30094 11942 30140 11994
rect 29844 11940 29900 11942
rect 29924 11940 29980 11942
rect 30004 11940 30060 11942
rect 30084 11940 30140 11942
rect 29844 10906 29900 10908
rect 29924 10906 29980 10908
rect 30004 10906 30060 10908
rect 30084 10906 30140 10908
rect 29844 10854 29890 10906
rect 29890 10854 29900 10906
rect 29924 10854 29954 10906
rect 29954 10854 29966 10906
rect 29966 10854 29980 10906
rect 30004 10854 30018 10906
rect 30018 10854 30030 10906
rect 30030 10854 30060 10906
rect 30084 10854 30094 10906
rect 30094 10854 30140 10906
rect 29844 10852 29900 10854
rect 29924 10852 29980 10854
rect 30004 10852 30060 10854
rect 30084 10852 30140 10854
rect 29844 9818 29900 9820
rect 29924 9818 29980 9820
rect 30004 9818 30060 9820
rect 30084 9818 30140 9820
rect 29844 9766 29890 9818
rect 29890 9766 29900 9818
rect 29924 9766 29954 9818
rect 29954 9766 29966 9818
rect 29966 9766 29980 9818
rect 30004 9766 30018 9818
rect 30018 9766 30030 9818
rect 30030 9766 30060 9818
rect 30084 9766 30094 9818
rect 30094 9766 30140 9818
rect 29844 9764 29900 9766
rect 29924 9764 29980 9766
rect 30004 9764 30060 9766
rect 30084 9764 30140 9766
rect 29844 8730 29900 8732
rect 29924 8730 29980 8732
rect 30004 8730 30060 8732
rect 30084 8730 30140 8732
rect 29844 8678 29890 8730
rect 29890 8678 29900 8730
rect 29924 8678 29954 8730
rect 29954 8678 29966 8730
rect 29966 8678 29980 8730
rect 30004 8678 30018 8730
rect 30018 8678 30030 8730
rect 30030 8678 30060 8730
rect 30084 8678 30094 8730
rect 30094 8678 30140 8730
rect 29844 8676 29900 8678
rect 29924 8676 29980 8678
rect 30004 8676 30060 8678
rect 30084 8676 30140 8678
rect 29844 7642 29900 7644
rect 29924 7642 29980 7644
rect 30004 7642 30060 7644
rect 30084 7642 30140 7644
rect 29844 7590 29890 7642
rect 29890 7590 29900 7642
rect 29924 7590 29954 7642
rect 29954 7590 29966 7642
rect 29966 7590 29980 7642
rect 30004 7590 30018 7642
rect 30018 7590 30030 7642
rect 30030 7590 30060 7642
rect 30084 7590 30094 7642
rect 30094 7590 30140 7642
rect 29844 7588 29900 7590
rect 29924 7588 29980 7590
rect 30004 7588 30060 7590
rect 30084 7588 30140 7590
rect 29844 6554 29900 6556
rect 29924 6554 29980 6556
rect 30004 6554 30060 6556
rect 30084 6554 30140 6556
rect 29844 6502 29890 6554
rect 29890 6502 29900 6554
rect 29924 6502 29954 6554
rect 29954 6502 29966 6554
rect 29966 6502 29980 6554
rect 30004 6502 30018 6554
rect 30018 6502 30030 6554
rect 30030 6502 30060 6554
rect 30084 6502 30094 6554
rect 30094 6502 30140 6554
rect 29844 6500 29900 6502
rect 29924 6500 29980 6502
rect 30004 6500 30060 6502
rect 30084 6500 30140 6502
rect 32494 18672 32550 18728
rect 29844 5466 29900 5468
rect 29924 5466 29980 5468
rect 30004 5466 30060 5468
rect 30084 5466 30140 5468
rect 29844 5414 29890 5466
rect 29890 5414 29900 5466
rect 29924 5414 29954 5466
rect 29954 5414 29966 5466
rect 29966 5414 29980 5466
rect 30004 5414 30018 5466
rect 30018 5414 30030 5466
rect 30030 5414 30060 5466
rect 30084 5414 30094 5466
rect 30094 5414 30140 5466
rect 29844 5412 29900 5414
rect 29924 5412 29980 5414
rect 30004 5412 30060 5414
rect 30084 5412 30140 5414
rect 30194 4700 30196 4720
rect 30196 4700 30248 4720
rect 30248 4700 30250 4720
rect 30194 4664 30250 4700
rect 29844 4378 29900 4380
rect 29924 4378 29980 4380
rect 30004 4378 30060 4380
rect 30084 4378 30140 4380
rect 29844 4326 29890 4378
rect 29890 4326 29900 4378
rect 29924 4326 29954 4378
rect 29954 4326 29966 4378
rect 29966 4326 29980 4378
rect 30004 4326 30018 4378
rect 30018 4326 30030 4378
rect 30030 4326 30060 4378
rect 30084 4326 30094 4378
rect 30094 4326 30140 4378
rect 29844 4324 29900 4326
rect 29924 4324 29980 4326
rect 30004 4324 30060 4326
rect 30084 4324 30140 4326
rect 29550 3440 29606 3496
rect 29844 3290 29900 3292
rect 29924 3290 29980 3292
rect 30004 3290 30060 3292
rect 30084 3290 30140 3292
rect 29844 3238 29890 3290
rect 29890 3238 29900 3290
rect 29924 3238 29954 3290
rect 29954 3238 29966 3290
rect 29966 3238 29980 3290
rect 30004 3238 30018 3290
rect 30018 3238 30030 3290
rect 30030 3238 30060 3290
rect 30084 3238 30094 3290
rect 30094 3238 30140 3290
rect 29844 3236 29900 3238
rect 29924 3236 29980 3238
rect 30004 3236 30060 3238
rect 30084 3236 30140 3238
rect 32402 4700 32404 4720
rect 32404 4700 32456 4720
rect 32456 4700 32458 4720
rect 32402 4664 32458 4700
rect 37066 22330 37122 22332
rect 37146 22330 37202 22332
rect 37226 22330 37282 22332
rect 37306 22330 37362 22332
rect 37066 22278 37112 22330
rect 37112 22278 37122 22330
rect 37146 22278 37176 22330
rect 37176 22278 37188 22330
rect 37188 22278 37202 22330
rect 37226 22278 37240 22330
rect 37240 22278 37252 22330
rect 37252 22278 37282 22330
rect 37306 22278 37316 22330
rect 37316 22278 37362 22330
rect 37066 22276 37122 22278
rect 37146 22276 37202 22278
rect 37226 22276 37282 22278
rect 37306 22276 37362 22278
rect 37066 21242 37122 21244
rect 37146 21242 37202 21244
rect 37226 21242 37282 21244
rect 37306 21242 37362 21244
rect 37066 21190 37112 21242
rect 37112 21190 37122 21242
rect 37146 21190 37176 21242
rect 37176 21190 37188 21242
rect 37188 21190 37202 21242
rect 37226 21190 37240 21242
rect 37240 21190 37252 21242
rect 37252 21190 37282 21242
rect 37306 21190 37316 21242
rect 37316 21190 37362 21242
rect 37066 21188 37122 21190
rect 37146 21188 37202 21190
rect 37226 21188 37282 21190
rect 37306 21188 37362 21190
rect 37066 20154 37122 20156
rect 37146 20154 37202 20156
rect 37226 20154 37282 20156
rect 37306 20154 37362 20156
rect 37066 20102 37112 20154
rect 37112 20102 37122 20154
rect 37146 20102 37176 20154
rect 37176 20102 37188 20154
rect 37188 20102 37202 20154
rect 37226 20102 37240 20154
rect 37240 20102 37252 20154
rect 37252 20102 37282 20154
rect 37306 20102 37316 20154
rect 37316 20102 37362 20154
rect 37066 20100 37122 20102
rect 37146 20100 37202 20102
rect 37226 20100 37282 20102
rect 37306 20100 37362 20102
rect 37066 19066 37122 19068
rect 37146 19066 37202 19068
rect 37226 19066 37282 19068
rect 37306 19066 37362 19068
rect 37066 19014 37112 19066
rect 37112 19014 37122 19066
rect 37146 19014 37176 19066
rect 37176 19014 37188 19066
rect 37188 19014 37202 19066
rect 37226 19014 37240 19066
rect 37240 19014 37252 19066
rect 37252 19014 37282 19066
rect 37306 19014 37316 19066
rect 37316 19014 37362 19066
rect 37066 19012 37122 19014
rect 37146 19012 37202 19014
rect 37226 19012 37282 19014
rect 37306 19012 37362 19014
rect 35070 12144 35126 12200
rect 35346 11092 35348 11112
rect 35348 11092 35400 11112
rect 35400 11092 35402 11112
rect 35346 11056 35402 11092
rect 37066 17978 37122 17980
rect 37146 17978 37202 17980
rect 37226 17978 37282 17980
rect 37306 17978 37362 17980
rect 37066 17926 37112 17978
rect 37112 17926 37122 17978
rect 37146 17926 37176 17978
rect 37176 17926 37188 17978
rect 37188 17926 37202 17978
rect 37226 17926 37240 17978
rect 37240 17926 37252 17978
rect 37252 17926 37282 17978
rect 37306 17926 37316 17978
rect 37316 17926 37362 17978
rect 37066 17924 37122 17926
rect 37146 17924 37202 17926
rect 37226 17924 37282 17926
rect 37306 17924 37362 17926
rect 37066 16890 37122 16892
rect 37146 16890 37202 16892
rect 37226 16890 37282 16892
rect 37306 16890 37362 16892
rect 37066 16838 37112 16890
rect 37112 16838 37122 16890
rect 37146 16838 37176 16890
rect 37176 16838 37188 16890
rect 37188 16838 37202 16890
rect 37226 16838 37240 16890
rect 37240 16838 37252 16890
rect 37252 16838 37282 16890
rect 37306 16838 37316 16890
rect 37316 16838 37362 16890
rect 37066 16836 37122 16838
rect 37146 16836 37202 16838
rect 37226 16836 37282 16838
rect 37306 16836 37362 16838
rect 37066 15802 37122 15804
rect 37146 15802 37202 15804
rect 37226 15802 37282 15804
rect 37306 15802 37362 15804
rect 37066 15750 37112 15802
rect 37112 15750 37122 15802
rect 37146 15750 37176 15802
rect 37176 15750 37188 15802
rect 37188 15750 37202 15802
rect 37226 15750 37240 15802
rect 37240 15750 37252 15802
rect 37252 15750 37282 15802
rect 37306 15750 37316 15802
rect 37316 15750 37362 15802
rect 37066 15748 37122 15750
rect 37146 15748 37202 15750
rect 37226 15748 37282 15750
rect 37306 15748 37362 15750
rect 37066 14714 37122 14716
rect 37146 14714 37202 14716
rect 37226 14714 37282 14716
rect 37306 14714 37362 14716
rect 37066 14662 37112 14714
rect 37112 14662 37122 14714
rect 37146 14662 37176 14714
rect 37176 14662 37188 14714
rect 37188 14662 37202 14714
rect 37226 14662 37240 14714
rect 37240 14662 37252 14714
rect 37252 14662 37282 14714
rect 37306 14662 37316 14714
rect 37316 14662 37362 14714
rect 37066 14660 37122 14662
rect 37146 14660 37202 14662
rect 37226 14660 37282 14662
rect 37306 14660 37362 14662
rect 34426 5480 34482 5536
rect 37066 13626 37122 13628
rect 37146 13626 37202 13628
rect 37226 13626 37282 13628
rect 37306 13626 37362 13628
rect 37066 13574 37112 13626
rect 37112 13574 37122 13626
rect 37146 13574 37176 13626
rect 37176 13574 37188 13626
rect 37188 13574 37202 13626
rect 37226 13574 37240 13626
rect 37240 13574 37252 13626
rect 37252 13574 37282 13626
rect 37306 13574 37316 13626
rect 37316 13574 37362 13626
rect 37066 13572 37122 13574
rect 37146 13572 37202 13574
rect 37226 13572 37282 13574
rect 37306 13572 37362 13574
rect 37066 12538 37122 12540
rect 37146 12538 37202 12540
rect 37226 12538 37282 12540
rect 37306 12538 37362 12540
rect 37066 12486 37112 12538
rect 37112 12486 37122 12538
rect 37146 12486 37176 12538
rect 37176 12486 37188 12538
rect 37188 12486 37202 12538
rect 37226 12486 37240 12538
rect 37240 12486 37252 12538
rect 37252 12486 37282 12538
rect 37306 12486 37316 12538
rect 37316 12486 37362 12538
rect 37066 12484 37122 12486
rect 37146 12484 37202 12486
rect 37226 12484 37282 12486
rect 37306 12484 37362 12486
rect 36358 9696 36414 9752
rect 37066 11450 37122 11452
rect 37146 11450 37202 11452
rect 37226 11450 37282 11452
rect 37306 11450 37362 11452
rect 37066 11398 37112 11450
rect 37112 11398 37122 11450
rect 37146 11398 37176 11450
rect 37176 11398 37188 11450
rect 37188 11398 37202 11450
rect 37226 11398 37240 11450
rect 37240 11398 37252 11450
rect 37252 11398 37282 11450
rect 37306 11398 37316 11450
rect 37316 11398 37362 11450
rect 37066 11396 37122 11398
rect 37146 11396 37202 11398
rect 37226 11396 37282 11398
rect 37306 11396 37362 11398
rect 37066 10362 37122 10364
rect 37146 10362 37202 10364
rect 37226 10362 37282 10364
rect 37306 10362 37362 10364
rect 37066 10310 37112 10362
rect 37112 10310 37122 10362
rect 37146 10310 37176 10362
rect 37176 10310 37188 10362
rect 37188 10310 37202 10362
rect 37226 10310 37240 10362
rect 37240 10310 37252 10362
rect 37252 10310 37282 10362
rect 37306 10310 37316 10362
rect 37316 10310 37362 10362
rect 37066 10308 37122 10310
rect 37146 10308 37202 10310
rect 37226 10308 37282 10310
rect 37306 10308 37362 10310
rect 37066 9274 37122 9276
rect 37146 9274 37202 9276
rect 37226 9274 37282 9276
rect 37306 9274 37362 9276
rect 37066 9222 37112 9274
rect 37112 9222 37122 9274
rect 37146 9222 37176 9274
rect 37176 9222 37188 9274
rect 37188 9222 37202 9274
rect 37226 9222 37240 9274
rect 37240 9222 37252 9274
rect 37252 9222 37282 9274
rect 37306 9222 37316 9274
rect 37316 9222 37362 9274
rect 37066 9220 37122 9222
rect 37146 9220 37202 9222
rect 37226 9220 37282 9222
rect 37306 9220 37362 9222
rect 44288 22874 44344 22876
rect 44368 22874 44424 22876
rect 44448 22874 44504 22876
rect 44528 22874 44584 22876
rect 44288 22822 44334 22874
rect 44334 22822 44344 22874
rect 44368 22822 44398 22874
rect 44398 22822 44410 22874
rect 44410 22822 44424 22874
rect 44448 22822 44462 22874
rect 44462 22822 44474 22874
rect 44474 22822 44504 22874
rect 44528 22822 44538 22874
rect 44538 22822 44584 22874
rect 44288 22820 44344 22822
rect 44368 22820 44424 22822
rect 44448 22820 44504 22822
rect 44528 22820 44584 22822
rect 37066 8186 37122 8188
rect 37146 8186 37202 8188
rect 37226 8186 37282 8188
rect 37306 8186 37362 8188
rect 37066 8134 37112 8186
rect 37112 8134 37122 8186
rect 37146 8134 37176 8186
rect 37176 8134 37188 8186
rect 37188 8134 37202 8186
rect 37226 8134 37240 8186
rect 37240 8134 37252 8186
rect 37252 8134 37282 8186
rect 37306 8134 37316 8186
rect 37316 8134 37362 8186
rect 37066 8132 37122 8134
rect 37146 8132 37202 8134
rect 37226 8132 37282 8134
rect 37306 8132 37362 8134
rect 37066 7098 37122 7100
rect 37146 7098 37202 7100
rect 37226 7098 37282 7100
rect 37306 7098 37362 7100
rect 37066 7046 37112 7098
rect 37112 7046 37122 7098
rect 37146 7046 37176 7098
rect 37176 7046 37188 7098
rect 37188 7046 37202 7098
rect 37226 7046 37240 7098
rect 37240 7046 37252 7098
rect 37252 7046 37282 7098
rect 37306 7046 37316 7098
rect 37316 7046 37362 7098
rect 37066 7044 37122 7046
rect 37146 7044 37202 7046
rect 37226 7044 37282 7046
rect 37306 7044 37362 7046
rect 37462 6160 37518 6216
rect 37066 6010 37122 6012
rect 37146 6010 37202 6012
rect 37226 6010 37282 6012
rect 37306 6010 37362 6012
rect 37066 5958 37112 6010
rect 37112 5958 37122 6010
rect 37146 5958 37176 6010
rect 37176 5958 37188 6010
rect 37188 5958 37202 6010
rect 37226 5958 37240 6010
rect 37240 5958 37252 6010
rect 37252 5958 37282 6010
rect 37306 5958 37316 6010
rect 37316 5958 37362 6010
rect 37066 5956 37122 5958
rect 37146 5956 37202 5958
rect 37226 5956 37282 5958
rect 37306 5956 37362 5958
rect 29844 2202 29900 2204
rect 29924 2202 29980 2204
rect 30004 2202 30060 2204
rect 30084 2202 30140 2204
rect 29844 2150 29890 2202
rect 29890 2150 29900 2202
rect 29924 2150 29954 2202
rect 29954 2150 29966 2202
rect 29966 2150 29980 2202
rect 30004 2150 30018 2202
rect 30018 2150 30030 2202
rect 30030 2150 30060 2202
rect 30084 2150 30094 2202
rect 30094 2150 30140 2202
rect 29844 2148 29900 2150
rect 29924 2148 29980 2150
rect 30004 2148 30060 2150
rect 30084 2148 30140 2150
rect 37066 4922 37122 4924
rect 37146 4922 37202 4924
rect 37226 4922 37282 4924
rect 37306 4922 37362 4924
rect 37066 4870 37112 4922
rect 37112 4870 37122 4922
rect 37146 4870 37176 4922
rect 37176 4870 37188 4922
rect 37188 4870 37202 4922
rect 37226 4870 37240 4922
rect 37240 4870 37252 4922
rect 37252 4870 37282 4922
rect 37306 4870 37316 4922
rect 37316 4870 37362 4922
rect 37066 4868 37122 4870
rect 37146 4868 37202 4870
rect 37226 4868 37282 4870
rect 37306 4868 37362 4870
rect 38198 6180 38254 6216
rect 38198 6160 38200 6180
rect 38200 6160 38252 6180
rect 38252 6160 38254 6180
rect 40038 11192 40094 11248
rect 37066 3834 37122 3836
rect 37146 3834 37202 3836
rect 37226 3834 37282 3836
rect 37306 3834 37362 3836
rect 37066 3782 37112 3834
rect 37112 3782 37122 3834
rect 37146 3782 37176 3834
rect 37176 3782 37188 3834
rect 37188 3782 37202 3834
rect 37226 3782 37240 3834
rect 37240 3782 37252 3834
rect 37252 3782 37282 3834
rect 37306 3782 37316 3834
rect 37316 3782 37362 3834
rect 37066 3780 37122 3782
rect 37146 3780 37202 3782
rect 37226 3780 37282 3782
rect 37306 3780 37362 3782
rect 37066 2746 37122 2748
rect 37146 2746 37202 2748
rect 37226 2746 37282 2748
rect 37306 2746 37362 2748
rect 37066 2694 37112 2746
rect 37112 2694 37122 2746
rect 37146 2694 37176 2746
rect 37176 2694 37188 2746
rect 37188 2694 37202 2746
rect 37226 2694 37240 2746
rect 37240 2694 37252 2746
rect 37252 2694 37282 2746
rect 37306 2694 37316 2746
rect 37316 2694 37362 2746
rect 37066 2692 37122 2694
rect 37146 2692 37202 2694
rect 37226 2692 37282 2694
rect 37306 2692 37362 2694
rect 44288 21786 44344 21788
rect 44368 21786 44424 21788
rect 44448 21786 44504 21788
rect 44528 21786 44584 21788
rect 44288 21734 44334 21786
rect 44334 21734 44344 21786
rect 44368 21734 44398 21786
rect 44398 21734 44410 21786
rect 44410 21734 44424 21786
rect 44448 21734 44462 21786
rect 44462 21734 44474 21786
rect 44474 21734 44504 21786
rect 44528 21734 44538 21786
rect 44538 21734 44584 21786
rect 44288 21732 44344 21734
rect 44368 21732 44424 21734
rect 44448 21732 44504 21734
rect 44528 21732 44584 21734
rect 44288 20698 44344 20700
rect 44368 20698 44424 20700
rect 44448 20698 44504 20700
rect 44528 20698 44584 20700
rect 44288 20646 44334 20698
rect 44334 20646 44344 20698
rect 44368 20646 44398 20698
rect 44398 20646 44410 20698
rect 44410 20646 44424 20698
rect 44448 20646 44462 20698
rect 44462 20646 44474 20698
rect 44474 20646 44504 20698
rect 44528 20646 44538 20698
rect 44538 20646 44584 20698
rect 44288 20644 44344 20646
rect 44368 20644 44424 20646
rect 44448 20644 44504 20646
rect 44528 20644 44584 20646
rect 44288 19610 44344 19612
rect 44368 19610 44424 19612
rect 44448 19610 44504 19612
rect 44528 19610 44584 19612
rect 44288 19558 44334 19610
rect 44334 19558 44344 19610
rect 44368 19558 44398 19610
rect 44398 19558 44410 19610
rect 44410 19558 44424 19610
rect 44448 19558 44462 19610
rect 44462 19558 44474 19610
rect 44474 19558 44504 19610
rect 44528 19558 44538 19610
rect 44538 19558 44584 19610
rect 44288 19556 44344 19558
rect 44368 19556 44424 19558
rect 44448 19556 44504 19558
rect 44528 19556 44584 19558
rect 42890 18808 42946 18864
rect 42338 13776 42394 13832
rect 41878 12688 41934 12744
rect 43350 18672 43406 18728
rect 43626 18808 43682 18864
rect 44288 18522 44344 18524
rect 44368 18522 44424 18524
rect 44448 18522 44504 18524
rect 44528 18522 44584 18524
rect 44288 18470 44334 18522
rect 44334 18470 44344 18522
rect 44368 18470 44398 18522
rect 44398 18470 44410 18522
rect 44410 18470 44424 18522
rect 44448 18470 44462 18522
rect 44462 18470 44474 18522
rect 44474 18470 44504 18522
rect 44528 18470 44538 18522
rect 44538 18470 44584 18522
rect 44288 18468 44344 18470
rect 44368 18468 44424 18470
rect 44448 18468 44504 18470
rect 44528 18468 44584 18470
rect 44288 17434 44344 17436
rect 44368 17434 44424 17436
rect 44448 17434 44504 17436
rect 44528 17434 44584 17436
rect 44288 17382 44334 17434
rect 44334 17382 44344 17434
rect 44368 17382 44398 17434
rect 44398 17382 44410 17434
rect 44410 17382 44424 17434
rect 44448 17382 44462 17434
rect 44462 17382 44474 17434
rect 44474 17382 44504 17434
rect 44528 17382 44538 17434
rect 44538 17382 44584 17434
rect 44288 17380 44344 17382
rect 44368 17380 44424 17382
rect 44448 17380 44504 17382
rect 44528 17380 44584 17382
rect 44288 16346 44344 16348
rect 44368 16346 44424 16348
rect 44448 16346 44504 16348
rect 44528 16346 44584 16348
rect 44288 16294 44334 16346
rect 44334 16294 44344 16346
rect 44368 16294 44398 16346
rect 44398 16294 44410 16346
rect 44410 16294 44424 16346
rect 44448 16294 44462 16346
rect 44462 16294 44474 16346
rect 44474 16294 44504 16346
rect 44528 16294 44538 16346
rect 44538 16294 44584 16346
rect 44288 16292 44344 16294
rect 44368 16292 44424 16294
rect 44448 16292 44504 16294
rect 44528 16292 44584 16294
rect 44288 15258 44344 15260
rect 44368 15258 44424 15260
rect 44448 15258 44504 15260
rect 44528 15258 44584 15260
rect 44288 15206 44334 15258
rect 44334 15206 44344 15258
rect 44368 15206 44398 15258
rect 44398 15206 44410 15258
rect 44410 15206 44424 15258
rect 44448 15206 44462 15258
rect 44462 15206 44474 15258
rect 44474 15206 44504 15258
rect 44528 15206 44538 15258
rect 44538 15206 44584 15258
rect 44288 15204 44344 15206
rect 44368 15204 44424 15206
rect 44448 15204 44504 15206
rect 44528 15204 44584 15206
rect 45282 18672 45338 18728
rect 44288 14170 44344 14172
rect 44368 14170 44424 14172
rect 44448 14170 44504 14172
rect 44528 14170 44584 14172
rect 44288 14118 44334 14170
rect 44334 14118 44344 14170
rect 44368 14118 44398 14170
rect 44398 14118 44410 14170
rect 44410 14118 44424 14170
rect 44448 14118 44462 14170
rect 44462 14118 44474 14170
rect 44474 14118 44504 14170
rect 44528 14118 44538 14170
rect 44538 14118 44584 14170
rect 44288 14116 44344 14118
rect 44368 14116 44424 14118
rect 44448 14116 44504 14118
rect 44528 14116 44584 14118
rect 44288 13082 44344 13084
rect 44368 13082 44424 13084
rect 44448 13082 44504 13084
rect 44528 13082 44584 13084
rect 44288 13030 44334 13082
rect 44334 13030 44344 13082
rect 44368 13030 44398 13082
rect 44398 13030 44410 13082
rect 44410 13030 44424 13082
rect 44448 13030 44462 13082
rect 44462 13030 44474 13082
rect 44474 13030 44504 13082
rect 44528 13030 44538 13082
rect 44538 13030 44584 13082
rect 44288 13028 44344 13030
rect 44368 13028 44424 13030
rect 44448 13028 44504 13030
rect 44528 13028 44584 13030
rect 40866 9560 40922 9616
rect 44288 11994 44344 11996
rect 44368 11994 44424 11996
rect 44448 11994 44504 11996
rect 44528 11994 44584 11996
rect 44288 11942 44334 11994
rect 44334 11942 44344 11994
rect 44368 11942 44398 11994
rect 44398 11942 44410 11994
rect 44410 11942 44424 11994
rect 44448 11942 44462 11994
rect 44462 11942 44474 11994
rect 44474 11942 44504 11994
rect 44528 11942 44538 11994
rect 44538 11942 44584 11994
rect 44288 11940 44344 11942
rect 44368 11940 44424 11942
rect 44448 11940 44504 11942
rect 44528 11940 44584 11942
rect 44288 10906 44344 10908
rect 44368 10906 44424 10908
rect 44448 10906 44504 10908
rect 44528 10906 44584 10908
rect 44288 10854 44334 10906
rect 44334 10854 44344 10906
rect 44368 10854 44398 10906
rect 44398 10854 44410 10906
rect 44410 10854 44424 10906
rect 44448 10854 44462 10906
rect 44462 10854 44474 10906
rect 44474 10854 44504 10906
rect 44528 10854 44538 10906
rect 44538 10854 44584 10906
rect 44288 10852 44344 10854
rect 44368 10852 44424 10854
rect 44448 10852 44504 10854
rect 44528 10852 44584 10854
rect 44288 9818 44344 9820
rect 44368 9818 44424 9820
rect 44448 9818 44504 9820
rect 44528 9818 44584 9820
rect 44288 9766 44334 9818
rect 44334 9766 44344 9818
rect 44368 9766 44398 9818
rect 44398 9766 44410 9818
rect 44410 9766 44424 9818
rect 44448 9766 44462 9818
rect 44462 9766 44474 9818
rect 44474 9766 44504 9818
rect 44528 9766 44538 9818
rect 44538 9766 44584 9818
rect 44288 9764 44344 9766
rect 44368 9764 44424 9766
rect 44448 9764 44504 9766
rect 44528 9764 44584 9766
rect 44288 8730 44344 8732
rect 44368 8730 44424 8732
rect 44448 8730 44504 8732
rect 44528 8730 44584 8732
rect 44288 8678 44334 8730
rect 44334 8678 44344 8730
rect 44368 8678 44398 8730
rect 44398 8678 44410 8730
rect 44410 8678 44424 8730
rect 44448 8678 44462 8730
rect 44462 8678 44474 8730
rect 44474 8678 44504 8730
rect 44528 8678 44538 8730
rect 44538 8678 44584 8730
rect 44288 8676 44344 8678
rect 44368 8676 44424 8678
rect 44448 8676 44504 8678
rect 44528 8676 44584 8678
rect 44288 7642 44344 7644
rect 44368 7642 44424 7644
rect 44448 7642 44504 7644
rect 44528 7642 44584 7644
rect 44288 7590 44334 7642
rect 44334 7590 44344 7642
rect 44368 7590 44398 7642
rect 44398 7590 44410 7642
rect 44410 7590 44424 7642
rect 44448 7590 44462 7642
rect 44462 7590 44474 7642
rect 44474 7590 44504 7642
rect 44528 7590 44538 7642
rect 44538 7590 44584 7642
rect 44288 7588 44344 7590
rect 44368 7588 44424 7590
rect 44448 7588 44504 7590
rect 44528 7588 44584 7590
rect 42246 3984 42302 4040
rect 44288 6554 44344 6556
rect 44368 6554 44424 6556
rect 44448 6554 44504 6556
rect 44528 6554 44584 6556
rect 44288 6502 44334 6554
rect 44334 6502 44344 6554
rect 44368 6502 44398 6554
rect 44398 6502 44410 6554
rect 44410 6502 44424 6554
rect 44448 6502 44462 6554
rect 44462 6502 44474 6554
rect 44474 6502 44504 6554
rect 44528 6502 44538 6554
rect 44538 6502 44584 6554
rect 44288 6500 44344 6502
rect 44368 6500 44424 6502
rect 44448 6500 44504 6502
rect 44528 6500 44584 6502
rect 44288 5466 44344 5468
rect 44368 5466 44424 5468
rect 44448 5466 44504 5468
rect 44528 5466 44584 5468
rect 44288 5414 44334 5466
rect 44334 5414 44344 5466
rect 44368 5414 44398 5466
rect 44398 5414 44410 5466
rect 44410 5414 44424 5466
rect 44448 5414 44462 5466
rect 44462 5414 44474 5466
rect 44474 5414 44504 5466
rect 44528 5414 44538 5466
rect 44538 5414 44584 5466
rect 44288 5412 44344 5414
rect 44368 5412 44424 5414
rect 44448 5412 44504 5414
rect 44528 5412 44584 5414
rect 44288 4378 44344 4380
rect 44368 4378 44424 4380
rect 44448 4378 44504 4380
rect 44528 4378 44584 4380
rect 44288 4326 44334 4378
rect 44334 4326 44344 4378
rect 44368 4326 44398 4378
rect 44398 4326 44410 4378
rect 44410 4326 44424 4378
rect 44448 4326 44462 4378
rect 44462 4326 44474 4378
rect 44474 4326 44504 4378
rect 44528 4326 44538 4378
rect 44538 4326 44584 4378
rect 44288 4324 44344 4326
rect 44368 4324 44424 4326
rect 44448 4324 44504 4326
rect 44528 4324 44584 4326
rect 44546 3984 44602 4040
rect 44288 3290 44344 3292
rect 44368 3290 44424 3292
rect 44448 3290 44504 3292
rect 44528 3290 44584 3292
rect 44288 3238 44334 3290
rect 44334 3238 44344 3290
rect 44368 3238 44398 3290
rect 44398 3238 44410 3290
rect 44410 3238 44424 3290
rect 44448 3238 44462 3290
rect 44462 3238 44474 3290
rect 44474 3238 44504 3290
rect 44528 3238 44538 3290
rect 44538 3238 44584 3290
rect 44288 3236 44344 3238
rect 44368 3236 44424 3238
rect 44448 3236 44504 3238
rect 44528 3236 44584 3238
rect 44288 2202 44344 2204
rect 44368 2202 44424 2204
rect 44448 2202 44504 2204
rect 44528 2202 44584 2204
rect 44288 2150 44334 2202
rect 44334 2150 44344 2202
rect 44368 2150 44398 2202
rect 44398 2150 44410 2202
rect 44410 2150 44424 2202
rect 44448 2150 44462 2202
rect 44462 2150 44474 2202
rect 44474 2150 44504 2202
rect 44528 2150 44538 2202
rect 44538 2150 44584 2202
rect 44288 2148 44344 2150
rect 44368 2148 44424 2150
rect 44448 2148 44504 2150
rect 44528 2148 44584 2150
rect 46570 9832 46626 9888
rect 45834 6704 45890 6760
rect 47030 9832 47086 9888
rect 46294 2760 46350 2816
rect 47582 6704 47638 6760
rect 47398 3984 47454 4040
rect 51510 23418 51566 23420
rect 51590 23418 51646 23420
rect 51670 23418 51726 23420
rect 51750 23418 51806 23420
rect 51510 23366 51556 23418
rect 51556 23366 51566 23418
rect 51590 23366 51620 23418
rect 51620 23366 51632 23418
rect 51632 23366 51646 23418
rect 51670 23366 51684 23418
rect 51684 23366 51696 23418
rect 51696 23366 51726 23418
rect 51750 23366 51760 23418
rect 51760 23366 51806 23418
rect 51510 23364 51566 23366
rect 51590 23364 51646 23366
rect 51670 23364 51726 23366
rect 51750 23364 51806 23366
rect 51510 22330 51566 22332
rect 51590 22330 51646 22332
rect 51670 22330 51726 22332
rect 51750 22330 51806 22332
rect 51510 22278 51556 22330
rect 51556 22278 51566 22330
rect 51590 22278 51620 22330
rect 51620 22278 51632 22330
rect 51632 22278 51646 22330
rect 51670 22278 51684 22330
rect 51684 22278 51696 22330
rect 51696 22278 51726 22330
rect 51750 22278 51760 22330
rect 51760 22278 51806 22330
rect 51510 22276 51566 22278
rect 51590 22276 51646 22278
rect 51670 22276 51726 22278
rect 51750 22276 51806 22278
rect 49146 6840 49202 6896
rect 51510 21242 51566 21244
rect 51590 21242 51646 21244
rect 51670 21242 51726 21244
rect 51750 21242 51806 21244
rect 51510 21190 51556 21242
rect 51556 21190 51566 21242
rect 51590 21190 51620 21242
rect 51620 21190 51632 21242
rect 51632 21190 51646 21242
rect 51670 21190 51684 21242
rect 51684 21190 51696 21242
rect 51696 21190 51726 21242
rect 51750 21190 51760 21242
rect 51760 21190 51806 21242
rect 51510 21188 51566 21190
rect 51590 21188 51646 21190
rect 51670 21188 51726 21190
rect 51750 21188 51806 21190
rect 51510 20154 51566 20156
rect 51590 20154 51646 20156
rect 51670 20154 51726 20156
rect 51750 20154 51806 20156
rect 51510 20102 51556 20154
rect 51556 20102 51566 20154
rect 51590 20102 51620 20154
rect 51620 20102 51632 20154
rect 51632 20102 51646 20154
rect 51670 20102 51684 20154
rect 51684 20102 51696 20154
rect 51696 20102 51726 20154
rect 51750 20102 51760 20154
rect 51760 20102 51806 20154
rect 51510 20100 51566 20102
rect 51590 20100 51646 20102
rect 51670 20100 51726 20102
rect 51750 20100 51806 20102
rect 51510 19066 51566 19068
rect 51590 19066 51646 19068
rect 51670 19066 51726 19068
rect 51750 19066 51806 19068
rect 51510 19014 51556 19066
rect 51556 19014 51566 19066
rect 51590 19014 51620 19066
rect 51620 19014 51632 19066
rect 51632 19014 51646 19066
rect 51670 19014 51684 19066
rect 51684 19014 51696 19066
rect 51696 19014 51726 19066
rect 51750 19014 51760 19066
rect 51760 19014 51806 19066
rect 51510 19012 51566 19014
rect 51590 19012 51646 19014
rect 51670 19012 51726 19014
rect 51750 19012 51806 19014
rect 58732 22874 58788 22876
rect 58812 22874 58868 22876
rect 58892 22874 58948 22876
rect 58972 22874 59028 22876
rect 58732 22822 58778 22874
rect 58778 22822 58788 22874
rect 58812 22822 58842 22874
rect 58842 22822 58854 22874
rect 58854 22822 58868 22874
rect 58892 22822 58906 22874
rect 58906 22822 58918 22874
rect 58918 22822 58948 22874
rect 58972 22822 58982 22874
rect 58982 22822 59028 22874
rect 58732 22820 58788 22822
rect 58812 22820 58868 22822
rect 58892 22820 58948 22822
rect 58972 22820 59028 22822
rect 58732 21786 58788 21788
rect 58812 21786 58868 21788
rect 58892 21786 58948 21788
rect 58972 21786 59028 21788
rect 58732 21734 58778 21786
rect 58778 21734 58788 21786
rect 58812 21734 58842 21786
rect 58842 21734 58854 21786
rect 58854 21734 58868 21786
rect 58892 21734 58906 21786
rect 58906 21734 58918 21786
rect 58918 21734 58948 21786
rect 58972 21734 58982 21786
rect 58982 21734 59028 21786
rect 58732 21732 58788 21734
rect 58812 21732 58868 21734
rect 58892 21732 58948 21734
rect 58972 21732 59028 21734
rect 51510 17978 51566 17980
rect 51590 17978 51646 17980
rect 51670 17978 51726 17980
rect 51750 17978 51806 17980
rect 51510 17926 51556 17978
rect 51556 17926 51566 17978
rect 51590 17926 51620 17978
rect 51620 17926 51632 17978
rect 51632 17926 51646 17978
rect 51670 17926 51684 17978
rect 51684 17926 51696 17978
rect 51696 17926 51726 17978
rect 51750 17926 51760 17978
rect 51760 17926 51806 17978
rect 51510 17924 51566 17926
rect 51590 17924 51646 17926
rect 51670 17924 51726 17926
rect 51750 17924 51806 17926
rect 51510 16890 51566 16892
rect 51590 16890 51646 16892
rect 51670 16890 51726 16892
rect 51750 16890 51806 16892
rect 51510 16838 51556 16890
rect 51556 16838 51566 16890
rect 51590 16838 51620 16890
rect 51620 16838 51632 16890
rect 51632 16838 51646 16890
rect 51670 16838 51684 16890
rect 51684 16838 51696 16890
rect 51696 16838 51726 16890
rect 51750 16838 51760 16890
rect 51760 16838 51806 16890
rect 51510 16836 51566 16838
rect 51590 16836 51646 16838
rect 51670 16836 51726 16838
rect 51750 16836 51806 16838
rect 51510 15802 51566 15804
rect 51590 15802 51646 15804
rect 51670 15802 51726 15804
rect 51750 15802 51806 15804
rect 51510 15750 51556 15802
rect 51556 15750 51566 15802
rect 51590 15750 51620 15802
rect 51620 15750 51632 15802
rect 51632 15750 51646 15802
rect 51670 15750 51684 15802
rect 51684 15750 51696 15802
rect 51696 15750 51726 15802
rect 51750 15750 51760 15802
rect 51760 15750 51806 15802
rect 51510 15748 51566 15750
rect 51590 15748 51646 15750
rect 51670 15748 51726 15750
rect 51750 15748 51806 15750
rect 51510 14714 51566 14716
rect 51590 14714 51646 14716
rect 51670 14714 51726 14716
rect 51750 14714 51806 14716
rect 51510 14662 51556 14714
rect 51556 14662 51566 14714
rect 51590 14662 51620 14714
rect 51620 14662 51632 14714
rect 51632 14662 51646 14714
rect 51670 14662 51684 14714
rect 51684 14662 51696 14714
rect 51696 14662 51726 14714
rect 51750 14662 51760 14714
rect 51760 14662 51806 14714
rect 51510 14660 51566 14662
rect 51590 14660 51646 14662
rect 51670 14660 51726 14662
rect 51750 14660 51806 14662
rect 51510 13626 51566 13628
rect 51590 13626 51646 13628
rect 51670 13626 51726 13628
rect 51750 13626 51806 13628
rect 51510 13574 51556 13626
rect 51556 13574 51566 13626
rect 51590 13574 51620 13626
rect 51620 13574 51632 13626
rect 51632 13574 51646 13626
rect 51670 13574 51684 13626
rect 51684 13574 51696 13626
rect 51696 13574 51726 13626
rect 51750 13574 51760 13626
rect 51760 13574 51806 13626
rect 51510 13572 51566 13574
rect 51590 13572 51646 13574
rect 51670 13572 51726 13574
rect 51750 13572 51806 13574
rect 52182 13368 52238 13424
rect 51510 12538 51566 12540
rect 51590 12538 51646 12540
rect 51670 12538 51726 12540
rect 51750 12538 51806 12540
rect 51510 12486 51556 12538
rect 51556 12486 51566 12538
rect 51590 12486 51620 12538
rect 51620 12486 51632 12538
rect 51632 12486 51646 12538
rect 51670 12486 51684 12538
rect 51684 12486 51696 12538
rect 51696 12486 51726 12538
rect 51750 12486 51760 12538
rect 51760 12486 51806 12538
rect 51510 12484 51566 12486
rect 51590 12484 51646 12486
rect 51670 12484 51726 12486
rect 51750 12484 51806 12486
rect 52734 12824 52790 12880
rect 49698 9580 49754 9616
rect 49698 9560 49700 9580
rect 49700 9560 49752 9580
rect 49752 9560 49754 9580
rect 51510 11450 51566 11452
rect 51590 11450 51646 11452
rect 51670 11450 51726 11452
rect 51750 11450 51806 11452
rect 51510 11398 51556 11450
rect 51556 11398 51566 11450
rect 51590 11398 51620 11450
rect 51620 11398 51632 11450
rect 51632 11398 51646 11450
rect 51670 11398 51684 11450
rect 51684 11398 51696 11450
rect 51696 11398 51726 11450
rect 51750 11398 51760 11450
rect 51760 11398 51806 11450
rect 51510 11396 51566 11398
rect 51590 11396 51646 11398
rect 51670 11396 51726 11398
rect 51750 11396 51806 11398
rect 51510 10362 51566 10364
rect 51590 10362 51646 10364
rect 51670 10362 51726 10364
rect 51750 10362 51806 10364
rect 51510 10310 51556 10362
rect 51556 10310 51566 10362
rect 51590 10310 51620 10362
rect 51620 10310 51632 10362
rect 51632 10310 51646 10362
rect 51670 10310 51684 10362
rect 51684 10310 51696 10362
rect 51696 10310 51726 10362
rect 51750 10310 51760 10362
rect 51760 10310 51806 10362
rect 51510 10308 51566 10310
rect 51590 10308 51646 10310
rect 51670 10308 51726 10310
rect 51750 10308 51806 10310
rect 51510 9274 51566 9276
rect 51590 9274 51646 9276
rect 51670 9274 51726 9276
rect 51750 9274 51806 9276
rect 51510 9222 51556 9274
rect 51556 9222 51566 9274
rect 51590 9222 51620 9274
rect 51620 9222 51632 9274
rect 51632 9222 51646 9274
rect 51670 9222 51684 9274
rect 51684 9222 51696 9274
rect 51696 9222 51726 9274
rect 51750 9222 51760 9274
rect 51760 9222 51806 9274
rect 51510 9220 51566 9222
rect 51590 9220 51646 9222
rect 51670 9220 51726 9222
rect 51750 9220 51806 9222
rect 51510 8186 51566 8188
rect 51590 8186 51646 8188
rect 51670 8186 51726 8188
rect 51750 8186 51806 8188
rect 51510 8134 51556 8186
rect 51556 8134 51566 8186
rect 51590 8134 51620 8186
rect 51620 8134 51632 8186
rect 51632 8134 51646 8186
rect 51670 8134 51684 8186
rect 51684 8134 51696 8186
rect 51696 8134 51726 8186
rect 51750 8134 51760 8186
rect 51760 8134 51806 8186
rect 51510 8132 51566 8134
rect 51590 8132 51646 8134
rect 51670 8132 51726 8134
rect 51750 8132 51806 8134
rect 51510 7098 51566 7100
rect 51590 7098 51646 7100
rect 51670 7098 51726 7100
rect 51750 7098 51806 7100
rect 51510 7046 51556 7098
rect 51556 7046 51566 7098
rect 51590 7046 51620 7098
rect 51620 7046 51632 7098
rect 51632 7046 51646 7098
rect 51670 7046 51684 7098
rect 51684 7046 51696 7098
rect 51696 7046 51726 7098
rect 51750 7046 51760 7098
rect 51760 7046 51806 7098
rect 51510 7044 51566 7046
rect 51590 7044 51646 7046
rect 51670 7044 51726 7046
rect 51750 7044 51806 7046
rect 49422 2896 49478 2952
rect 50342 3576 50398 3632
rect 51510 6010 51566 6012
rect 51590 6010 51646 6012
rect 51670 6010 51726 6012
rect 51750 6010 51806 6012
rect 51510 5958 51556 6010
rect 51556 5958 51566 6010
rect 51590 5958 51620 6010
rect 51620 5958 51632 6010
rect 51632 5958 51646 6010
rect 51670 5958 51684 6010
rect 51684 5958 51696 6010
rect 51696 5958 51726 6010
rect 51750 5958 51760 6010
rect 51760 5958 51806 6010
rect 51510 5956 51566 5958
rect 51590 5956 51646 5958
rect 51670 5956 51726 5958
rect 51750 5956 51806 5958
rect 52090 6840 52146 6896
rect 53746 13232 53802 13288
rect 50986 3984 51042 4040
rect 51510 4922 51566 4924
rect 51590 4922 51646 4924
rect 51670 4922 51726 4924
rect 51750 4922 51806 4924
rect 51510 4870 51556 4922
rect 51556 4870 51566 4922
rect 51590 4870 51620 4922
rect 51620 4870 51632 4922
rect 51632 4870 51646 4922
rect 51670 4870 51684 4922
rect 51684 4870 51696 4922
rect 51696 4870 51726 4922
rect 51750 4870 51760 4922
rect 51760 4870 51806 4922
rect 51510 4868 51566 4870
rect 51590 4868 51646 4870
rect 51670 4868 51726 4870
rect 51750 4868 51806 4870
rect 51510 3834 51566 3836
rect 51590 3834 51646 3836
rect 51670 3834 51726 3836
rect 51750 3834 51806 3836
rect 51510 3782 51556 3834
rect 51556 3782 51566 3834
rect 51590 3782 51620 3834
rect 51620 3782 51632 3834
rect 51632 3782 51646 3834
rect 51670 3782 51684 3834
rect 51684 3782 51696 3834
rect 51696 3782 51726 3834
rect 51750 3782 51760 3834
rect 51760 3782 51806 3834
rect 51510 3780 51566 3782
rect 51590 3780 51646 3782
rect 51670 3780 51726 3782
rect 51750 3780 51806 3782
rect 51170 2760 51226 2816
rect 51510 2746 51566 2748
rect 51590 2746 51646 2748
rect 51670 2746 51726 2748
rect 51750 2746 51806 2748
rect 51510 2694 51556 2746
rect 51556 2694 51566 2746
rect 51590 2694 51620 2746
rect 51620 2694 51632 2746
rect 51632 2694 51646 2746
rect 51670 2694 51684 2746
rect 51684 2694 51696 2746
rect 51696 2694 51726 2746
rect 51750 2694 51760 2746
rect 51760 2694 51806 2746
rect 51510 2692 51566 2694
rect 51590 2692 51646 2694
rect 51670 2692 51726 2694
rect 51750 2692 51806 2694
rect 52734 3576 52790 3632
rect 58732 20698 58788 20700
rect 58812 20698 58868 20700
rect 58892 20698 58948 20700
rect 58972 20698 59028 20700
rect 58732 20646 58778 20698
rect 58778 20646 58788 20698
rect 58812 20646 58842 20698
rect 58842 20646 58854 20698
rect 58854 20646 58868 20698
rect 58892 20646 58906 20698
rect 58906 20646 58918 20698
rect 58918 20646 58948 20698
rect 58972 20646 58982 20698
rect 58982 20646 59028 20698
rect 58732 20644 58788 20646
rect 58812 20644 58868 20646
rect 58892 20644 58948 20646
rect 58972 20644 59028 20646
rect 53102 3984 53158 4040
rect 53562 3304 53618 3360
rect 52734 2760 52790 2816
rect 56598 15000 56654 15056
rect 54758 2896 54814 2952
rect 58732 19610 58788 19612
rect 58812 19610 58868 19612
rect 58892 19610 58948 19612
rect 58972 19610 59028 19612
rect 58732 19558 58778 19610
rect 58778 19558 58788 19610
rect 58812 19558 58842 19610
rect 58842 19558 58854 19610
rect 58854 19558 58868 19610
rect 58892 19558 58906 19610
rect 58906 19558 58918 19610
rect 58918 19558 58948 19610
rect 58972 19558 58982 19610
rect 58982 19558 59028 19610
rect 58732 19556 58788 19558
rect 58812 19556 58868 19558
rect 58892 19556 58948 19558
rect 58972 19556 59028 19558
rect 58732 18522 58788 18524
rect 58812 18522 58868 18524
rect 58892 18522 58948 18524
rect 58972 18522 59028 18524
rect 58732 18470 58778 18522
rect 58778 18470 58788 18522
rect 58812 18470 58842 18522
rect 58842 18470 58854 18522
rect 58854 18470 58868 18522
rect 58892 18470 58906 18522
rect 58906 18470 58918 18522
rect 58918 18470 58948 18522
rect 58972 18470 58982 18522
rect 58982 18470 59028 18522
rect 58732 18468 58788 18470
rect 58812 18468 58868 18470
rect 58892 18468 58948 18470
rect 58972 18468 59028 18470
rect 58732 17434 58788 17436
rect 58812 17434 58868 17436
rect 58892 17434 58948 17436
rect 58972 17434 59028 17436
rect 58732 17382 58778 17434
rect 58778 17382 58788 17434
rect 58812 17382 58842 17434
rect 58842 17382 58854 17434
rect 58854 17382 58868 17434
rect 58892 17382 58906 17434
rect 58906 17382 58918 17434
rect 58918 17382 58948 17434
rect 58972 17382 58982 17434
rect 58982 17382 59028 17434
rect 58732 17380 58788 17382
rect 58812 17380 58868 17382
rect 58892 17380 58948 17382
rect 58972 17380 59028 17382
rect 58732 16346 58788 16348
rect 58812 16346 58868 16348
rect 58892 16346 58948 16348
rect 58972 16346 59028 16348
rect 58732 16294 58778 16346
rect 58778 16294 58788 16346
rect 58812 16294 58842 16346
rect 58842 16294 58854 16346
rect 58854 16294 58868 16346
rect 58892 16294 58906 16346
rect 58906 16294 58918 16346
rect 58918 16294 58948 16346
rect 58972 16294 58982 16346
rect 58982 16294 59028 16346
rect 58732 16292 58788 16294
rect 58812 16292 58868 16294
rect 58892 16292 58948 16294
rect 58972 16292 59028 16294
rect 58732 15258 58788 15260
rect 58812 15258 58868 15260
rect 58892 15258 58948 15260
rect 58972 15258 59028 15260
rect 58732 15206 58778 15258
rect 58778 15206 58788 15258
rect 58812 15206 58842 15258
rect 58842 15206 58854 15258
rect 58854 15206 58868 15258
rect 58892 15206 58906 15258
rect 58906 15206 58918 15258
rect 58918 15206 58948 15258
rect 58972 15206 58982 15258
rect 58982 15206 59028 15258
rect 58732 15204 58788 15206
rect 58812 15204 58868 15206
rect 58892 15204 58948 15206
rect 58972 15204 59028 15206
rect 58732 14170 58788 14172
rect 58812 14170 58868 14172
rect 58892 14170 58948 14172
rect 58972 14170 59028 14172
rect 58732 14118 58778 14170
rect 58778 14118 58788 14170
rect 58812 14118 58842 14170
rect 58842 14118 58854 14170
rect 58854 14118 58868 14170
rect 58892 14118 58906 14170
rect 58906 14118 58918 14170
rect 58918 14118 58948 14170
rect 58972 14118 58982 14170
rect 58982 14118 59028 14170
rect 58732 14116 58788 14118
rect 58812 14116 58868 14118
rect 58892 14116 58948 14118
rect 58972 14116 59028 14118
rect 58732 13082 58788 13084
rect 58812 13082 58868 13084
rect 58892 13082 58948 13084
rect 58972 13082 59028 13084
rect 58732 13030 58778 13082
rect 58778 13030 58788 13082
rect 58812 13030 58842 13082
rect 58842 13030 58854 13082
rect 58854 13030 58868 13082
rect 58892 13030 58906 13082
rect 58906 13030 58918 13082
rect 58918 13030 58948 13082
rect 58972 13030 58982 13082
rect 58982 13030 59028 13082
rect 58732 13028 58788 13030
rect 58812 13028 58868 13030
rect 58892 13028 58948 13030
rect 58972 13028 59028 13030
rect 57426 11736 57482 11792
rect 57426 3304 57482 3360
rect 58732 11994 58788 11996
rect 58812 11994 58868 11996
rect 58892 11994 58948 11996
rect 58972 11994 59028 11996
rect 58732 11942 58778 11994
rect 58778 11942 58788 11994
rect 58812 11942 58842 11994
rect 58842 11942 58854 11994
rect 58854 11942 58868 11994
rect 58892 11942 58906 11994
rect 58906 11942 58918 11994
rect 58918 11942 58948 11994
rect 58972 11942 58982 11994
rect 58982 11942 59028 11994
rect 58732 11940 58788 11942
rect 58812 11940 58868 11942
rect 58892 11940 58948 11942
rect 58972 11940 59028 11942
rect 58732 10906 58788 10908
rect 58812 10906 58868 10908
rect 58892 10906 58948 10908
rect 58972 10906 59028 10908
rect 58732 10854 58778 10906
rect 58778 10854 58788 10906
rect 58812 10854 58842 10906
rect 58842 10854 58854 10906
rect 58854 10854 58868 10906
rect 58892 10854 58906 10906
rect 58906 10854 58918 10906
rect 58918 10854 58948 10906
rect 58972 10854 58982 10906
rect 58982 10854 59028 10906
rect 58732 10852 58788 10854
rect 58812 10852 58868 10854
rect 58892 10852 58948 10854
rect 58972 10852 59028 10854
rect 58732 9818 58788 9820
rect 58812 9818 58868 9820
rect 58892 9818 58948 9820
rect 58972 9818 59028 9820
rect 58732 9766 58778 9818
rect 58778 9766 58788 9818
rect 58812 9766 58842 9818
rect 58842 9766 58854 9818
rect 58854 9766 58868 9818
rect 58892 9766 58906 9818
rect 58906 9766 58918 9818
rect 58918 9766 58948 9818
rect 58972 9766 58982 9818
rect 58982 9766 59028 9818
rect 58732 9764 58788 9766
rect 58812 9764 58868 9766
rect 58892 9764 58948 9766
rect 58972 9764 59028 9766
rect 58732 8730 58788 8732
rect 58812 8730 58868 8732
rect 58892 8730 58948 8732
rect 58972 8730 59028 8732
rect 58732 8678 58778 8730
rect 58778 8678 58788 8730
rect 58812 8678 58842 8730
rect 58842 8678 58854 8730
rect 58854 8678 58868 8730
rect 58892 8678 58906 8730
rect 58906 8678 58918 8730
rect 58918 8678 58948 8730
rect 58972 8678 58982 8730
rect 58982 8678 59028 8730
rect 58732 8676 58788 8678
rect 58812 8676 58868 8678
rect 58892 8676 58948 8678
rect 58972 8676 59028 8678
rect 58732 7642 58788 7644
rect 58812 7642 58868 7644
rect 58892 7642 58948 7644
rect 58972 7642 59028 7644
rect 58732 7590 58778 7642
rect 58778 7590 58788 7642
rect 58812 7590 58842 7642
rect 58842 7590 58854 7642
rect 58854 7590 58868 7642
rect 58892 7590 58906 7642
rect 58906 7590 58918 7642
rect 58918 7590 58948 7642
rect 58972 7590 58982 7642
rect 58982 7590 59028 7642
rect 58732 7588 58788 7590
rect 58812 7588 58868 7590
rect 58892 7588 58948 7590
rect 58972 7588 59028 7590
rect 58732 6554 58788 6556
rect 58812 6554 58868 6556
rect 58892 6554 58948 6556
rect 58972 6554 59028 6556
rect 58732 6502 58778 6554
rect 58778 6502 58788 6554
rect 58812 6502 58842 6554
rect 58842 6502 58854 6554
rect 58854 6502 58868 6554
rect 58892 6502 58906 6554
rect 58906 6502 58918 6554
rect 58918 6502 58948 6554
rect 58972 6502 58982 6554
rect 58982 6502 59028 6554
rect 58732 6500 58788 6502
rect 58812 6500 58868 6502
rect 58892 6500 58948 6502
rect 58972 6500 59028 6502
rect 58732 5466 58788 5468
rect 58812 5466 58868 5468
rect 58892 5466 58948 5468
rect 58972 5466 59028 5468
rect 58732 5414 58778 5466
rect 58778 5414 58788 5466
rect 58812 5414 58842 5466
rect 58842 5414 58854 5466
rect 58854 5414 58868 5466
rect 58892 5414 58906 5466
rect 58906 5414 58918 5466
rect 58918 5414 58948 5466
rect 58972 5414 58982 5466
rect 58982 5414 59028 5466
rect 58732 5412 58788 5414
rect 58812 5412 58868 5414
rect 58892 5412 58948 5414
rect 58972 5412 59028 5414
rect 58732 4378 58788 4380
rect 58812 4378 58868 4380
rect 58892 4378 58948 4380
rect 58972 4378 59028 4380
rect 58732 4326 58778 4378
rect 58778 4326 58788 4378
rect 58812 4326 58842 4378
rect 58842 4326 58854 4378
rect 58854 4326 58868 4378
rect 58892 4326 58906 4378
rect 58906 4326 58918 4378
rect 58918 4326 58948 4378
rect 58972 4326 58982 4378
rect 58982 4326 59028 4378
rect 58732 4324 58788 4326
rect 58812 4324 58868 4326
rect 58892 4324 58948 4326
rect 58972 4324 59028 4326
rect 58732 3290 58788 3292
rect 58812 3290 58868 3292
rect 58892 3290 58948 3292
rect 58972 3290 59028 3292
rect 58732 3238 58778 3290
rect 58778 3238 58788 3290
rect 58812 3238 58842 3290
rect 58842 3238 58854 3290
rect 58854 3238 58868 3290
rect 58892 3238 58906 3290
rect 58906 3238 58918 3290
rect 58918 3238 58948 3290
rect 58972 3238 58982 3290
rect 58982 3238 59028 3290
rect 58732 3236 58788 3238
rect 58812 3236 58868 3238
rect 58892 3236 58948 3238
rect 58972 3236 59028 3238
rect 58438 2760 58494 2816
rect 58732 2202 58788 2204
rect 58812 2202 58868 2204
rect 58892 2202 58948 2204
rect 58972 2202 59028 2204
rect 58732 2150 58778 2202
rect 58778 2150 58788 2202
rect 58812 2150 58842 2202
rect 58842 2150 58854 2202
rect 58854 2150 58868 2202
rect 58892 2150 58906 2202
rect 58906 2150 58918 2202
rect 58918 2150 58948 2202
rect 58972 2150 58982 2202
rect 58982 2150 59028 2202
rect 58732 2148 58788 2150
rect 58812 2148 58868 2150
rect 58892 2148 58948 2150
rect 58972 2148 59028 2150
<< metal3 >>
rect 8168 27776 8484 27777
rect 8168 27712 8174 27776
rect 8238 27712 8254 27776
rect 8318 27712 8334 27776
rect 8398 27712 8414 27776
rect 8478 27712 8484 27776
rect 8168 27711 8484 27712
rect 22612 27776 22928 27777
rect 22612 27712 22618 27776
rect 22682 27712 22698 27776
rect 22762 27712 22778 27776
rect 22842 27712 22858 27776
rect 22922 27712 22928 27776
rect 22612 27711 22928 27712
rect 37056 27776 37372 27777
rect 37056 27712 37062 27776
rect 37126 27712 37142 27776
rect 37206 27712 37222 27776
rect 37286 27712 37302 27776
rect 37366 27712 37372 27776
rect 37056 27711 37372 27712
rect 51500 27776 51816 27777
rect 51500 27712 51506 27776
rect 51570 27712 51586 27776
rect 51650 27712 51666 27776
rect 51730 27712 51746 27776
rect 51810 27712 51816 27776
rect 51500 27711 51816 27712
rect 15390 27232 15706 27233
rect 15390 27168 15396 27232
rect 15460 27168 15476 27232
rect 15540 27168 15556 27232
rect 15620 27168 15636 27232
rect 15700 27168 15706 27232
rect 15390 27167 15706 27168
rect 29834 27232 30150 27233
rect 29834 27168 29840 27232
rect 29904 27168 29920 27232
rect 29984 27168 30000 27232
rect 30064 27168 30080 27232
rect 30144 27168 30150 27232
rect 29834 27167 30150 27168
rect 44278 27232 44594 27233
rect 44278 27168 44284 27232
rect 44348 27168 44364 27232
rect 44428 27168 44444 27232
rect 44508 27168 44524 27232
rect 44588 27168 44594 27232
rect 44278 27167 44594 27168
rect 58722 27232 59038 27233
rect 58722 27168 58728 27232
rect 58792 27168 58808 27232
rect 58872 27168 58888 27232
rect 58952 27168 58968 27232
rect 59032 27168 59038 27232
rect 58722 27167 59038 27168
rect 8168 26688 8484 26689
rect 8168 26624 8174 26688
rect 8238 26624 8254 26688
rect 8318 26624 8334 26688
rect 8398 26624 8414 26688
rect 8478 26624 8484 26688
rect 8168 26623 8484 26624
rect 22612 26688 22928 26689
rect 22612 26624 22618 26688
rect 22682 26624 22698 26688
rect 22762 26624 22778 26688
rect 22842 26624 22858 26688
rect 22922 26624 22928 26688
rect 22612 26623 22928 26624
rect 37056 26688 37372 26689
rect 37056 26624 37062 26688
rect 37126 26624 37142 26688
rect 37206 26624 37222 26688
rect 37286 26624 37302 26688
rect 37366 26624 37372 26688
rect 37056 26623 37372 26624
rect 51500 26688 51816 26689
rect 51500 26624 51506 26688
rect 51570 26624 51586 26688
rect 51650 26624 51666 26688
rect 51730 26624 51746 26688
rect 51810 26624 51816 26688
rect 51500 26623 51816 26624
rect 15390 26144 15706 26145
rect 15390 26080 15396 26144
rect 15460 26080 15476 26144
rect 15540 26080 15556 26144
rect 15620 26080 15636 26144
rect 15700 26080 15706 26144
rect 15390 26079 15706 26080
rect 29834 26144 30150 26145
rect 29834 26080 29840 26144
rect 29904 26080 29920 26144
rect 29984 26080 30000 26144
rect 30064 26080 30080 26144
rect 30144 26080 30150 26144
rect 29834 26079 30150 26080
rect 44278 26144 44594 26145
rect 44278 26080 44284 26144
rect 44348 26080 44364 26144
rect 44428 26080 44444 26144
rect 44508 26080 44524 26144
rect 44588 26080 44594 26144
rect 44278 26079 44594 26080
rect 58722 26144 59038 26145
rect 58722 26080 58728 26144
rect 58792 26080 58808 26144
rect 58872 26080 58888 26144
rect 58952 26080 58968 26144
rect 59032 26080 59038 26144
rect 58722 26079 59038 26080
rect 8168 25600 8484 25601
rect 8168 25536 8174 25600
rect 8238 25536 8254 25600
rect 8318 25536 8334 25600
rect 8398 25536 8414 25600
rect 8478 25536 8484 25600
rect 8168 25535 8484 25536
rect 22612 25600 22928 25601
rect 22612 25536 22618 25600
rect 22682 25536 22698 25600
rect 22762 25536 22778 25600
rect 22842 25536 22858 25600
rect 22922 25536 22928 25600
rect 22612 25535 22928 25536
rect 37056 25600 37372 25601
rect 37056 25536 37062 25600
rect 37126 25536 37142 25600
rect 37206 25536 37222 25600
rect 37286 25536 37302 25600
rect 37366 25536 37372 25600
rect 37056 25535 37372 25536
rect 51500 25600 51816 25601
rect 51500 25536 51506 25600
rect 51570 25536 51586 25600
rect 51650 25536 51666 25600
rect 51730 25536 51746 25600
rect 51810 25536 51816 25600
rect 51500 25535 51816 25536
rect 15390 25056 15706 25057
rect 15390 24992 15396 25056
rect 15460 24992 15476 25056
rect 15540 24992 15556 25056
rect 15620 24992 15636 25056
rect 15700 24992 15706 25056
rect 15390 24991 15706 24992
rect 29834 25056 30150 25057
rect 29834 24992 29840 25056
rect 29904 24992 29920 25056
rect 29984 24992 30000 25056
rect 30064 24992 30080 25056
rect 30144 24992 30150 25056
rect 29834 24991 30150 24992
rect 44278 25056 44594 25057
rect 44278 24992 44284 25056
rect 44348 24992 44364 25056
rect 44428 24992 44444 25056
rect 44508 24992 44524 25056
rect 44588 24992 44594 25056
rect 44278 24991 44594 24992
rect 58722 25056 59038 25057
rect 58722 24992 58728 25056
rect 58792 24992 58808 25056
rect 58872 24992 58888 25056
rect 58952 24992 58968 25056
rect 59032 24992 59038 25056
rect 58722 24991 59038 24992
rect 8168 24512 8484 24513
rect 8168 24448 8174 24512
rect 8238 24448 8254 24512
rect 8318 24448 8334 24512
rect 8398 24448 8414 24512
rect 8478 24448 8484 24512
rect 8168 24447 8484 24448
rect 22612 24512 22928 24513
rect 22612 24448 22618 24512
rect 22682 24448 22698 24512
rect 22762 24448 22778 24512
rect 22842 24448 22858 24512
rect 22922 24448 22928 24512
rect 22612 24447 22928 24448
rect 37056 24512 37372 24513
rect 37056 24448 37062 24512
rect 37126 24448 37142 24512
rect 37206 24448 37222 24512
rect 37286 24448 37302 24512
rect 37366 24448 37372 24512
rect 37056 24447 37372 24448
rect 51500 24512 51816 24513
rect 51500 24448 51506 24512
rect 51570 24448 51586 24512
rect 51650 24448 51666 24512
rect 51730 24448 51746 24512
rect 51810 24448 51816 24512
rect 51500 24447 51816 24448
rect 15390 23968 15706 23969
rect 15390 23904 15396 23968
rect 15460 23904 15476 23968
rect 15540 23904 15556 23968
rect 15620 23904 15636 23968
rect 15700 23904 15706 23968
rect 15390 23903 15706 23904
rect 29834 23968 30150 23969
rect 29834 23904 29840 23968
rect 29904 23904 29920 23968
rect 29984 23904 30000 23968
rect 30064 23904 30080 23968
rect 30144 23904 30150 23968
rect 29834 23903 30150 23904
rect 44278 23968 44594 23969
rect 44278 23904 44284 23968
rect 44348 23904 44364 23968
rect 44428 23904 44444 23968
rect 44508 23904 44524 23968
rect 44588 23904 44594 23968
rect 44278 23903 44594 23904
rect 58722 23968 59038 23969
rect 58722 23904 58728 23968
rect 58792 23904 58808 23968
rect 58872 23904 58888 23968
rect 58952 23904 58968 23968
rect 59032 23904 59038 23968
rect 58722 23903 59038 23904
rect 8168 23424 8484 23425
rect 8168 23360 8174 23424
rect 8238 23360 8254 23424
rect 8318 23360 8334 23424
rect 8398 23360 8414 23424
rect 8478 23360 8484 23424
rect 8168 23359 8484 23360
rect 22612 23424 22928 23425
rect 22612 23360 22618 23424
rect 22682 23360 22698 23424
rect 22762 23360 22778 23424
rect 22842 23360 22858 23424
rect 22922 23360 22928 23424
rect 22612 23359 22928 23360
rect 37056 23424 37372 23425
rect 37056 23360 37062 23424
rect 37126 23360 37142 23424
rect 37206 23360 37222 23424
rect 37286 23360 37302 23424
rect 37366 23360 37372 23424
rect 37056 23359 37372 23360
rect 51500 23424 51816 23425
rect 51500 23360 51506 23424
rect 51570 23360 51586 23424
rect 51650 23360 51666 23424
rect 51730 23360 51746 23424
rect 51810 23360 51816 23424
rect 51500 23359 51816 23360
rect 15390 22880 15706 22881
rect 15390 22816 15396 22880
rect 15460 22816 15476 22880
rect 15540 22816 15556 22880
rect 15620 22816 15636 22880
rect 15700 22816 15706 22880
rect 15390 22815 15706 22816
rect 29834 22880 30150 22881
rect 29834 22816 29840 22880
rect 29904 22816 29920 22880
rect 29984 22816 30000 22880
rect 30064 22816 30080 22880
rect 30144 22816 30150 22880
rect 29834 22815 30150 22816
rect 44278 22880 44594 22881
rect 44278 22816 44284 22880
rect 44348 22816 44364 22880
rect 44428 22816 44444 22880
rect 44508 22816 44524 22880
rect 44588 22816 44594 22880
rect 44278 22815 44594 22816
rect 58722 22880 59038 22881
rect 58722 22816 58728 22880
rect 58792 22816 58808 22880
rect 58872 22816 58888 22880
rect 58952 22816 58968 22880
rect 59032 22816 59038 22880
rect 58722 22815 59038 22816
rect 8168 22336 8484 22337
rect 8168 22272 8174 22336
rect 8238 22272 8254 22336
rect 8318 22272 8334 22336
rect 8398 22272 8414 22336
rect 8478 22272 8484 22336
rect 8168 22271 8484 22272
rect 22612 22336 22928 22337
rect 22612 22272 22618 22336
rect 22682 22272 22698 22336
rect 22762 22272 22778 22336
rect 22842 22272 22858 22336
rect 22922 22272 22928 22336
rect 22612 22271 22928 22272
rect 37056 22336 37372 22337
rect 37056 22272 37062 22336
rect 37126 22272 37142 22336
rect 37206 22272 37222 22336
rect 37286 22272 37302 22336
rect 37366 22272 37372 22336
rect 37056 22271 37372 22272
rect 51500 22336 51816 22337
rect 51500 22272 51506 22336
rect 51570 22272 51586 22336
rect 51650 22272 51666 22336
rect 51730 22272 51746 22336
rect 51810 22272 51816 22336
rect 51500 22271 51816 22272
rect 15390 21792 15706 21793
rect 15390 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15706 21792
rect 15390 21727 15706 21728
rect 29834 21792 30150 21793
rect 29834 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30150 21792
rect 29834 21727 30150 21728
rect 44278 21792 44594 21793
rect 44278 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44594 21792
rect 44278 21727 44594 21728
rect 58722 21792 59038 21793
rect 58722 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59038 21792
rect 58722 21727 59038 21728
rect 27429 21722 27495 21725
rect 28073 21722 28139 21725
rect 27429 21720 28139 21722
rect 27429 21664 27434 21720
rect 27490 21664 28078 21720
rect 28134 21664 28139 21720
rect 27429 21662 28139 21664
rect 27429 21659 27495 21662
rect 28073 21659 28139 21662
rect 32213 21450 32279 21453
rect 32765 21450 32831 21453
rect 32213 21448 32831 21450
rect 32213 21392 32218 21448
rect 32274 21392 32770 21448
rect 32826 21392 32831 21448
rect 32213 21390 32831 21392
rect 32213 21387 32279 21390
rect 32765 21387 32831 21390
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 22612 21248 22928 21249
rect 22612 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22928 21248
rect 22612 21183 22928 21184
rect 37056 21248 37372 21249
rect 37056 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37372 21248
rect 37056 21183 37372 21184
rect 51500 21248 51816 21249
rect 51500 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51816 21248
rect 51500 21183 51816 21184
rect 16481 20772 16547 20773
rect 16430 20770 16436 20772
rect 16390 20710 16436 20770
rect 16500 20768 16547 20772
rect 16542 20712 16547 20768
rect 16430 20708 16436 20710
rect 16500 20708 16547 20712
rect 16481 20707 16547 20708
rect 15390 20704 15706 20705
rect 15390 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15706 20704
rect 15390 20639 15706 20640
rect 29834 20704 30150 20705
rect 29834 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30150 20704
rect 29834 20639 30150 20640
rect 44278 20704 44594 20705
rect 44278 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44594 20704
rect 44278 20639 44594 20640
rect 58722 20704 59038 20705
rect 58722 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59038 20704
rect 58722 20639 59038 20640
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 22612 20160 22928 20161
rect 22612 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22928 20160
rect 22612 20095 22928 20096
rect 37056 20160 37372 20161
rect 37056 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37372 20160
rect 37056 20095 37372 20096
rect 51500 20160 51816 20161
rect 51500 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51816 20160
rect 51500 20095 51816 20096
rect 15390 19616 15706 19617
rect 15390 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15706 19616
rect 15390 19551 15706 19552
rect 29834 19616 30150 19617
rect 29834 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30150 19616
rect 29834 19551 30150 19552
rect 44278 19616 44594 19617
rect 44278 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44594 19616
rect 44278 19551 44594 19552
rect 58722 19616 59038 19617
rect 58722 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59038 19616
rect 58722 19551 59038 19552
rect 6545 19410 6611 19413
rect 6678 19410 6684 19412
rect 6545 19408 6684 19410
rect 6545 19352 6550 19408
rect 6606 19352 6684 19408
rect 6545 19350 6684 19352
rect 6545 19347 6611 19350
rect 6678 19348 6684 19350
rect 6748 19348 6754 19412
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 22612 19072 22928 19073
rect 22612 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22928 19072
rect 22612 19007 22928 19008
rect 37056 19072 37372 19073
rect 37056 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37372 19072
rect 37056 19007 37372 19008
rect 51500 19072 51816 19073
rect 51500 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51816 19072
rect 51500 19007 51816 19008
rect 42885 18866 42951 18869
rect 43621 18866 43687 18869
rect 42885 18864 43687 18866
rect 42885 18808 42890 18864
rect 42946 18808 43626 18864
rect 43682 18808 43687 18864
rect 42885 18806 43687 18808
rect 42885 18803 42951 18806
rect 43621 18803 43687 18806
rect 31385 18730 31451 18733
rect 32489 18730 32555 18733
rect 31385 18728 32555 18730
rect 31385 18672 31390 18728
rect 31446 18672 32494 18728
rect 32550 18672 32555 18728
rect 31385 18670 32555 18672
rect 31385 18667 31451 18670
rect 32489 18667 32555 18670
rect 43345 18730 43411 18733
rect 45277 18730 45343 18733
rect 43345 18728 45343 18730
rect 43345 18672 43350 18728
rect 43406 18672 45282 18728
rect 45338 18672 45343 18728
rect 43345 18670 45343 18672
rect 43345 18667 43411 18670
rect 45277 18667 45343 18670
rect 15390 18528 15706 18529
rect 15390 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15706 18528
rect 15390 18463 15706 18464
rect 29834 18528 30150 18529
rect 29834 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30150 18528
rect 29834 18463 30150 18464
rect 44278 18528 44594 18529
rect 44278 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44594 18528
rect 44278 18463 44594 18464
rect 58722 18528 59038 18529
rect 58722 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59038 18528
rect 58722 18463 59038 18464
rect 27613 18186 27679 18189
rect 28349 18186 28415 18189
rect 27613 18184 28415 18186
rect 27613 18128 27618 18184
rect 27674 18128 28354 18184
rect 28410 18128 28415 18184
rect 27613 18126 28415 18128
rect 27613 18123 27679 18126
rect 28349 18123 28415 18126
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 22612 17984 22928 17985
rect 22612 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22928 17984
rect 22612 17919 22928 17920
rect 37056 17984 37372 17985
rect 37056 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37372 17984
rect 37056 17919 37372 17920
rect 51500 17984 51816 17985
rect 51500 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51816 17984
rect 51500 17919 51816 17920
rect 15390 17440 15706 17441
rect 15390 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15706 17440
rect 15390 17375 15706 17376
rect 29834 17440 30150 17441
rect 29834 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30150 17440
rect 29834 17375 30150 17376
rect 44278 17440 44594 17441
rect 44278 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44594 17440
rect 44278 17375 44594 17376
rect 58722 17440 59038 17441
rect 58722 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59038 17440
rect 58722 17375 59038 17376
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 22612 16896 22928 16897
rect 22612 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22928 16896
rect 22612 16831 22928 16832
rect 37056 16896 37372 16897
rect 37056 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37372 16896
rect 37056 16831 37372 16832
rect 51500 16896 51816 16897
rect 51500 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51816 16896
rect 51500 16831 51816 16832
rect 15390 16352 15706 16353
rect 15390 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15706 16352
rect 15390 16287 15706 16288
rect 29834 16352 30150 16353
rect 29834 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30150 16352
rect 29834 16287 30150 16288
rect 44278 16352 44594 16353
rect 44278 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44594 16352
rect 44278 16287 44594 16288
rect 58722 16352 59038 16353
rect 58722 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59038 16352
rect 58722 16287 59038 16288
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 22612 15808 22928 15809
rect 22612 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22928 15808
rect 22612 15743 22928 15744
rect 37056 15808 37372 15809
rect 37056 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37372 15808
rect 37056 15743 37372 15744
rect 51500 15808 51816 15809
rect 51500 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51816 15808
rect 51500 15743 51816 15744
rect 9581 15602 9647 15605
rect 26325 15602 26391 15605
rect 9581 15600 26391 15602
rect 9581 15544 9586 15600
rect 9642 15544 26330 15600
rect 26386 15544 26391 15600
rect 9581 15542 26391 15544
rect 9581 15539 9647 15542
rect 26325 15539 26391 15542
rect 15390 15264 15706 15265
rect 15390 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15706 15264
rect 15390 15199 15706 15200
rect 29834 15264 30150 15265
rect 29834 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30150 15264
rect 29834 15199 30150 15200
rect 44278 15264 44594 15265
rect 44278 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44594 15264
rect 44278 15199 44594 15200
rect 58722 15264 59038 15265
rect 58722 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59038 15264
rect 58722 15199 59038 15200
rect 7281 15058 7347 15061
rect 7925 15058 7991 15061
rect 56593 15058 56659 15061
rect 7281 15056 56659 15058
rect 7281 15000 7286 15056
rect 7342 15000 7930 15056
rect 7986 15000 56598 15056
rect 56654 15000 56659 15056
rect 7281 14998 56659 15000
rect 7281 14995 7347 14998
rect 7925 14995 7991 14998
rect 56593 14995 56659 14998
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 22612 14720 22928 14721
rect 22612 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22928 14720
rect 22612 14655 22928 14656
rect 37056 14720 37372 14721
rect 37056 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37372 14720
rect 37056 14655 37372 14656
rect 51500 14720 51816 14721
rect 51500 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51816 14720
rect 51500 14655 51816 14656
rect 15390 14176 15706 14177
rect 15390 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15706 14176
rect 15390 14111 15706 14112
rect 29834 14176 30150 14177
rect 29834 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30150 14176
rect 29834 14111 30150 14112
rect 44278 14176 44594 14177
rect 44278 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44594 14176
rect 44278 14111 44594 14112
rect 58722 14176 59038 14177
rect 58722 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59038 14176
rect 58722 14111 59038 14112
rect 42333 13836 42399 13837
rect 42333 13832 42380 13836
rect 42444 13834 42450 13836
rect 42333 13776 42338 13832
rect 42333 13772 42380 13776
rect 42444 13774 42490 13834
rect 42444 13772 42450 13774
rect 42333 13771 42399 13772
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 22612 13632 22928 13633
rect 22612 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22928 13632
rect 22612 13567 22928 13568
rect 37056 13632 37372 13633
rect 37056 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37372 13632
rect 37056 13567 37372 13568
rect 51500 13632 51816 13633
rect 51500 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51816 13632
rect 51500 13567 51816 13568
rect 23289 13562 23355 13565
rect 26233 13562 26299 13565
rect 23289 13560 26299 13562
rect 23289 13504 23294 13560
rect 23350 13504 26238 13560
rect 26294 13504 26299 13560
rect 23289 13502 26299 13504
rect 23289 13499 23355 13502
rect 26233 13499 26299 13502
rect 13721 13426 13787 13429
rect 52177 13426 52243 13429
rect 13721 13424 52243 13426
rect 13721 13368 13726 13424
rect 13782 13368 52182 13424
rect 52238 13368 52243 13424
rect 13721 13366 52243 13368
rect 13721 13363 13787 13366
rect 52177 13363 52243 13366
rect 12985 13290 13051 13293
rect 53741 13290 53807 13293
rect 12985 13288 53807 13290
rect 12985 13232 12990 13288
rect 13046 13232 53746 13288
rect 53802 13232 53807 13288
rect 12985 13230 53807 13232
rect 12985 13227 13051 13230
rect 53741 13227 53807 13230
rect 15390 13088 15706 13089
rect 15390 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15706 13088
rect 15390 13023 15706 13024
rect 29834 13088 30150 13089
rect 29834 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30150 13088
rect 29834 13023 30150 13024
rect 44278 13088 44594 13089
rect 44278 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44594 13088
rect 44278 13023 44594 13024
rect 58722 13088 59038 13089
rect 58722 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59038 13088
rect 58722 13023 59038 13024
rect 10409 12882 10475 12885
rect 52729 12882 52795 12885
rect 10409 12880 52795 12882
rect 10409 12824 10414 12880
rect 10470 12824 52734 12880
rect 52790 12824 52795 12880
rect 10409 12822 52795 12824
rect 10409 12819 10475 12822
rect 52729 12819 52795 12822
rect 9213 12746 9279 12749
rect 41873 12746 41939 12749
rect 9213 12744 41939 12746
rect 9213 12688 9218 12744
rect 9274 12688 41878 12744
rect 41934 12688 41939 12744
rect 9213 12686 41939 12688
rect 9213 12683 9279 12686
rect 41873 12683 41939 12686
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 22612 12544 22928 12545
rect 22612 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22928 12544
rect 22612 12479 22928 12480
rect 37056 12544 37372 12545
rect 37056 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37372 12544
rect 37056 12479 37372 12480
rect 51500 12544 51816 12545
rect 51500 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51816 12544
rect 51500 12479 51816 12480
rect 7557 12338 7623 12341
rect 12893 12338 12959 12341
rect 7557 12336 12959 12338
rect 7557 12280 7562 12336
rect 7618 12280 12898 12336
rect 12954 12280 12959 12336
rect 7557 12278 12959 12280
rect 7557 12275 7623 12278
rect 12893 12275 12959 12278
rect 30373 12202 30439 12205
rect 35065 12202 35131 12205
rect 30373 12200 35131 12202
rect 30373 12144 30378 12200
rect 30434 12144 35070 12200
rect 35126 12144 35131 12200
rect 30373 12142 35131 12144
rect 30373 12139 30439 12142
rect 35065 12139 35131 12142
rect 15390 12000 15706 12001
rect 15390 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15706 12000
rect 15390 11935 15706 11936
rect 29834 12000 30150 12001
rect 29834 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30150 12000
rect 29834 11935 30150 11936
rect 44278 12000 44594 12001
rect 44278 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44594 12000
rect 44278 11935 44594 11936
rect 58722 12000 59038 12001
rect 58722 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59038 12000
rect 58722 11935 59038 11936
rect 7005 11794 7071 11797
rect 57421 11794 57487 11797
rect 7005 11792 57487 11794
rect 7005 11736 7010 11792
rect 7066 11736 57426 11792
rect 57482 11736 57487 11792
rect 7005 11734 57487 11736
rect 7005 11731 7071 11734
rect 57421 11731 57487 11734
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 22612 11456 22928 11457
rect 22612 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22928 11456
rect 22612 11391 22928 11392
rect 37056 11456 37372 11457
rect 37056 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37372 11456
rect 37056 11391 37372 11392
rect 51500 11456 51816 11457
rect 51500 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51816 11456
rect 51500 11391 51816 11392
rect 10133 11250 10199 11253
rect 40033 11250 40099 11253
rect 10133 11248 40099 11250
rect 10133 11192 10138 11248
rect 10194 11192 40038 11248
rect 40094 11192 40099 11248
rect 10133 11190 40099 11192
rect 10133 11187 10199 11190
rect 40033 11187 40099 11190
rect 7097 11114 7163 11117
rect 35341 11114 35407 11117
rect 7097 11112 35407 11114
rect 7097 11056 7102 11112
rect 7158 11056 35346 11112
rect 35402 11056 35407 11112
rect 7097 11054 35407 11056
rect 7097 11051 7163 11054
rect 35341 11051 35407 11054
rect 15390 10912 15706 10913
rect 15390 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15706 10912
rect 15390 10847 15706 10848
rect 29834 10912 30150 10913
rect 29834 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30150 10912
rect 29834 10847 30150 10848
rect 44278 10912 44594 10913
rect 44278 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44594 10912
rect 44278 10847 44594 10848
rect 58722 10912 59038 10913
rect 58722 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59038 10912
rect 58722 10847 59038 10848
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 22612 10368 22928 10369
rect 22612 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22928 10368
rect 22612 10303 22928 10304
rect 37056 10368 37372 10369
rect 37056 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37372 10368
rect 37056 10303 37372 10304
rect 51500 10368 51816 10369
rect 51500 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51816 10368
rect 51500 10303 51816 10304
rect 46565 9890 46631 9893
rect 47025 9890 47091 9893
rect 46565 9888 47091 9890
rect 46565 9832 46570 9888
rect 46626 9832 47030 9888
rect 47086 9832 47091 9888
rect 46565 9830 47091 9832
rect 46565 9827 46631 9830
rect 47025 9827 47091 9830
rect 15390 9824 15706 9825
rect 15390 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15706 9824
rect 15390 9759 15706 9760
rect 29834 9824 30150 9825
rect 29834 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30150 9824
rect 29834 9759 30150 9760
rect 44278 9824 44594 9825
rect 44278 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44594 9824
rect 44278 9759 44594 9760
rect 58722 9824 59038 9825
rect 58722 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59038 9824
rect 58722 9759 59038 9760
rect 35934 9692 35940 9756
rect 36004 9754 36010 9756
rect 36353 9754 36419 9757
rect 36004 9752 36419 9754
rect 36004 9696 36358 9752
rect 36414 9696 36419 9752
rect 36004 9694 36419 9696
rect 36004 9692 36010 9694
rect 36353 9691 36419 9694
rect 40861 9618 40927 9621
rect 49693 9618 49759 9621
rect 40861 9616 49759 9618
rect 40861 9560 40866 9616
rect 40922 9560 49698 9616
rect 49754 9560 49759 9616
rect 40861 9558 49759 9560
rect 40861 9555 40927 9558
rect 49693 9555 49759 9558
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 22612 9280 22928 9281
rect 22612 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22928 9280
rect 22612 9215 22928 9216
rect 37056 9280 37372 9281
rect 37056 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37372 9280
rect 37056 9215 37372 9216
rect 51500 9280 51816 9281
rect 51500 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51816 9280
rect 51500 9215 51816 9216
rect 15390 8736 15706 8737
rect 15390 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15706 8736
rect 15390 8671 15706 8672
rect 29834 8736 30150 8737
rect 29834 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30150 8736
rect 29834 8671 30150 8672
rect 44278 8736 44594 8737
rect 44278 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44594 8736
rect 44278 8671 44594 8672
rect 58722 8736 59038 8737
rect 58722 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59038 8736
rect 58722 8671 59038 8672
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 22612 8192 22928 8193
rect 22612 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22928 8192
rect 22612 8127 22928 8128
rect 37056 8192 37372 8193
rect 37056 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37372 8192
rect 37056 8127 37372 8128
rect 51500 8192 51816 8193
rect 51500 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51816 8192
rect 51500 8127 51816 8128
rect 15390 7648 15706 7649
rect 15390 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15706 7648
rect 15390 7583 15706 7584
rect 29834 7648 30150 7649
rect 29834 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30150 7648
rect 29834 7583 30150 7584
rect 44278 7648 44594 7649
rect 44278 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44594 7648
rect 44278 7583 44594 7584
rect 58722 7648 59038 7649
rect 58722 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59038 7648
rect 58722 7583 59038 7584
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 22612 7104 22928 7105
rect 22612 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22928 7104
rect 22612 7039 22928 7040
rect 37056 7104 37372 7105
rect 37056 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37372 7104
rect 37056 7039 37372 7040
rect 51500 7104 51816 7105
rect 51500 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51816 7104
rect 51500 7039 51816 7040
rect 17493 7034 17559 7037
rect 19374 7034 19380 7036
rect 17493 7032 19380 7034
rect 17493 6976 17498 7032
rect 17554 6976 19380 7032
rect 17493 6974 19380 6976
rect 17493 6971 17559 6974
rect 19374 6972 19380 6974
rect 19444 6972 19450 7036
rect 12985 6898 13051 6901
rect 15377 6898 15443 6901
rect 12985 6896 15443 6898
rect 12985 6840 12990 6896
rect 13046 6840 15382 6896
rect 15438 6840 15443 6896
rect 12985 6838 15443 6840
rect 12985 6835 13051 6838
rect 15377 6835 15443 6838
rect 49141 6898 49207 6901
rect 52085 6898 52151 6901
rect 49141 6896 52151 6898
rect 49141 6840 49146 6896
rect 49202 6840 52090 6896
rect 52146 6840 52151 6896
rect 49141 6838 52151 6840
rect 49141 6835 49207 6838
rect 52085 6835 52151 6838
rect 45829 6762 45895 6765
rect 47577 6762 47643 6765
rect 45829 6760 47643 6762
rect 45829 6704 45834 6760
rect 45890 6704 47582 6760
rect 47638 6704 47643 6760
rect 45829 6702 47643 6704
rect 45829 6699 45895 6702
rect 47577 6699 47643 6702
rect 15390 6560 15706 6561
rect 15390 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15706 6560
rect 15390 6495 15706 6496
rect 29834 6560 30150 6561
rect 29834 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30150 6560
rect 29834 6495 30150 6496
rect 44278 6560 44594 6561
rect 44278 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44594 6560
rect 44278 6495 44594 6496
rect 58722 6560 59038 6561
rect 58722 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59038 6560
rect 58722 6495 59038 6496
rect 37457 6218 37523 6221
rect 38193 6218 38259 6221
rect 37457 6216 38259 6218
rect 37457 6160 37462 6216
rect 37518 6160 38198 6216
rect 38254 6160 38259 6216
rect 37457 6158 38259 6160
rect 37457 6155 37523 6158
rect 38193 6155 38259 6158
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 22612 6016 22928 6017
rect 22612 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22928 6016
rect 22612 5951 22928 5952
rect 37056 6016 37372 6017
rect 37056 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37372 6016
rect 37056 5951 37372 5952
rect 51500 6016 51816 6017
rect 51500 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51816 6016
rect 51500 5951 51816 5952
rect 34421 5538 34487 5541
rect 35934 5538 35940 5540
rect 34421 5536 35940 5538
rect 34421 5480 34426 5536
rect 34482 5480 35940 5536
rect 34421 5478 35940 5480
rect 34421 5475 34487 5478
rect 35934 5476 35940 5478
rect 36004 5476 36010 5540
rect 15390 5472 15706 5473
rect 15390 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15706 5472
rect 15390 5407 15706 5408
rect 29834 5472 30150 5473
rect 29834 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30150 5472
rect 29834 5407 30150 5408
rect 44278 5472 44594 5473
rect 44278 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44594 5472
rect 44278 5407 44594 5408
rect 58722 5472 59038 5473
rect 58722 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59038 5472
rect 58722 5407 59038 5408
rect 3969 4994 4035 4997
rect 7741 4994 7807 4997
rect 3969 4992 7807 4994
rect 3969 4936 3974 4992
rect 4030 4936 7746 4992
rect 7802 4936 7807 4992
rect 3969 4934 7807 4936
rect 3969 4931 4035 4934
rect 7741 4931 7807 4934
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 22612 4928 22928 4929
rect 22612 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22928 4928
rect 22612 4863 22928 4864
rect 37056 4928 37372 4929
rect 37056 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37372 4928
rect 37056 4863 37372 4864
rect 51500 4928 51816 4929
rect 51500 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51816 4928
rect 51500 4863 51816 4864
rect 30189 4722 30255 4725
rect 32397 4722 32463 4725
rect 30189 4720 32463 4722
rect 30189 4664 30194 4720
rect 30250 4664 32402 4720
rect 32458 4664 32463 4720
rect 30189 4662 32463 4664
rect 30189 4659 30255 4662
rect 32397 4659 32463 4662
rect 15390 4384 15706 4385
rect 15390 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15706 4384
rect 15390 4319 15706 4320
rect 29834 4384 30150 4385
rect 29834 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30150 4384
rect 29834 4319 30150 4320
rect 44278 4384 44594 4385
rect 44278 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44594 4384
rect 44278 4319 44594 4320
rect 58722 4384 59038 4385
rect 58722 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59038 4384
rect 58722 4319 59038 4320
rect 5901 4178 5967 4181
rect 6637 4178 6703 4181
rect 5901 4176 6703 4178
rect 5901 4120 5906 4176
rect 5962 4120 6642 4176
rect 6698 4120 6703 4176
rect 5901 4118 6703 4120
rect 5901 4115 5967 4118
rect 6637 4115 6703 4118
rect 5349 4042 5415 4045
rect 6678 4042 6684 4044
rect 5349 4040 6684 4042
rect 5349 3984 5354 4040
rect 5410 3984 6684 4040
rect 5349 3982 6684 3984
rect 5349 3979 5415 3982
rect 6678 3980 6684 3982
rect 6748 3980 6754 4044
rect 16430 3980 16436 4044
rect 16500 4042 16506 4044
rect 16849 4042 16915 4045
rect 16500 4040 16915 4042
rect 16500 3984 16854 4040
rect 16910 3984 16915 4040
rect 16500 3982 16915 3984
rect 16500 3980 16506 3982
rect 16849 3979 16915 3982
rect 19374 3980 19380 4044
rect 19444 4042 19450 4044
rect 19517 4042 19583 4045
rect 19444 4040 19583 4042
rect 19444 3984 19522 4040
rect 19578 3984 19583 4040
rect 19444 3982 19583 3984
rect 19444 3980 19450 3982
rect 19517 3979 19583 3982
rect 42241 4042 42307 4045
rect 42374 4042 42380 4044
rect 42241 4040 42380 4042
rect 42241 3984 42246 4040
rect 42302 3984 42380 4040
rect 42241 3982 42380 3984
rect 42241 3979 42307 3982
rect 42374 3980 42380 3982
rect 42444 3980 42450 4044
rect 44541 4042 44607 4045
rect 47393 4042 47459 4045
rect 44541 4040 47459 4042
rect 44541 3984 44546 4040
rect 44602 3984 47398 4040
rect 47454 3984 47459 4040
rect 44541 3982 47459 3984
rect 44541 3979 44607 3982
rect 47393 3979 47459 3982
rect 50981 4042 51047 4045
rect 53097 4042 53163 4045
rect 50981 4040 53163 4042
rect 50981 3984 50986 4040
rect 51042 3984 53102 4040
rect 53158 3984 53163 4040
rect 50981 3982 53163 3984
rect 50981 3979 51047 3982
rect 53097 3979 53163 3982
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 22612 3840 22928 3841
rect 22612 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22928 3840
rect 22612 3775 22928 3776
rect 37056 3840 37372 3841
rect 37056 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37372 3840
rect 37056 3775 37372 3776
rect 51500 3840 51816 3841
rect 51500 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51816 3840
rect 51500 3775 51816 3776
rect 50337 3634 50403 3637
rect 52729 3634 52795 3637
rect 50337 3632 52795 3634
rect 50337 3576 50342 3632
rect 50398 3576 52734 3632
rect 52790 3576 52795 3632
rect 50337 3574 52795 3576
rect 50337 3571 50403 3574
rect 52729 3571 52795 3574
rect 1393 3498 1459 3501
rect 29545 3498 29611 3501
rect 1393 3496 29611 3498
rect 1393 3440 1398 3496
rect 1454 3440 29550 3496
rect 29606 3440 29611 3496
rect 1393 3438 29611 3440
rect 1393 3435 1459 3438
rect 29545 3435 29611 3438
rect 53557 3362 53623 3365
rect 57421 3362 57487 3365
rect 53557 3360 57487 3362
rect 53557 3304 53562 3360
rect 53618 3304 57426 3360
rect 57482 3304 57487 3360
rect 53557 3302 57487 3304
rect 53557 3299 53623 3302
rect 57421 3299 57487 3302
rect 15390 3296 15706 3297
rect 15390 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15706 3296
rect 15390 3231 15706 3232
rect 29834 3296 30150 3297
rect 29834 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30150 3296
rect 29834 3231 30150 3232
rect 44278 3296 44594 3297
rect 44278 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44594 3296
rect 44278 3231 44594 3232
rect 58722 3296 59038 3297
rect 58722 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59038 3296
rect 58722 3231 59038 3232
rect 5993 2954 6059 2957
rect 7465 2954 7531 2957
rect 5993 2952 7531 2954
rect 5993 2896 5998 2952
rect 6054 2896 7470 2952
rect 7526 2896 7531 2952
rect 5993 2894 7531 2896
rect 5993 2891 6059 2894
rect 7465 2891 7531 2894
rect 49417 2954 49483 2957
rect 54753 2954 54819 2957
rect 49417 2952 54819 2954
rect 49417 2896 49422 2952
rect 49478 2896 54758 2952
rect 54814 2896 54819 2952
rect 49417 2894 54819 2896
rect 49417 2891 49483 2894
rect 54753 2891 54819 2894
rect 46289 2818 46355 2821
rect 51165 2818 51231 2821
rect 46289 2816 51231 2818
rect 46289 2760 46294 2816
rect 46350 2760 51170 2816
rect 51226 2760 51231 2816
rect 46289 2758 51231 2760
rect 46289 2755 46355 2758
rect 51165 2755 51231 2758
rect 52729 2818 52795 2821
rect 58433 2818 58499 2821
rect 52729 2816 58499 2818
rect 52729 2760 52734 2816
rect 52790 2760 58438 2816
rect 58494 2760 58499 2816
rect 52729 2758 58499 2760
rect 52729 2755 52795 2758
rect 58433 2755 58499 2758
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 22612 2752 22928 2753
rect 22612 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22928 2752
rect 22612 2687 22928 2688
rect 37056 2752 37372 2753
rect 37056 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37372 2752
rect 37056 2687 37372 2688
rect 51500 2752 51816 2753
rect 51500 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51816 2752
rect 51500 2687 51816 2688
rect 15390 2208 15706 2209
rect 15390 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15706 2208
rect 15390 2143 15706 2144
rect 29834 2208 30150 2209
rect 29834 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30150 2208
rect 29834 2143 30150 2144
rect 44278 2208 44594 2209
rect 44278 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44594 2208
rect 44278 2143 44594 2144
rect 58722 2208 59038 2209
rect 58722 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59038 2208
rect 58722 2143 59038 2144
<< via3 >>
rect 8174 27772 8238 27776
rect 8174 27716 8178 27772
rect 8178 27716 8234 27772
rect 8234 27716 8238 27772
rect 8174 27712 8238 27716
rect 8254 27772 8318 27776
rect 8254 27716 8258 27772
rect 8258 27716 8314 27772
rect 8314 27716 8318 27772
rect 8254 27712 8318 27716
rect 8334 27772 8398 27776
rect 8334 27716 8338 27772
rect 8338 27716 8394 27772
rect 8394 27716 8398 27772
rect 8334 27712 8398 27716
rect 8414 27772 8478 27776
rect 8414 27716 8418 27772
rect 8418 27716 8474 27772
rect 8474 27716 8478 27772
rect 8414 27712 8478 27716
rect 22618 27772 22682 27776
rect 22618 27716 22622 27772
rect 22622 27716 22678 27772
rect 22678 27716 22682 27772
rect 22618 27712 22682 27716
rect 22698 27772 22762 27776
rect 22698 27716 22702 27772
rect 22702 27716 22758 27772
rect 22758 27716 22762 27772
rect 22698 27712 22762 27716
rect 22778 27772 22842 27776
rect 22778 27716 22782 27772
rect 22782 27716 22838 27772
rect 22838 27716 22842 27772
rect 22778 27712 22842 27716
rect 22858 27772 22922 27776
rect 22858 27716 22862 27772
rect 22862 27716 22918 27772
rect 22918 27716 22922 27772
rect 22858 27712 22922 27716
rect 37062 27772 37126 27776
rect 37062 27716 37066 27772
rect 37066 27716 37122 27772
rect 37122 27716 37126 27772
rect 37062 27712 37126 27716
rect 37142 27772 37206 27776
rect 37142 27716 37146 27772
rect 37146 27716 37202 27772
rect 37202 27716 37206 27772
rect 37142 27712 37206 27716
rect 37222 27772 37286 27776
rect 37222 27716 37226 27772
rect 37226 27716 37282 27772
rect 37282 27716 37286 27772
rect 37222 27712 37286 27716
rect 37302 27772 37366 27776
rect 37302 27716 37306 27772
rect 37306 27716 37362 27772
rect 37362 27716 37366 27772
rect 37302 27712 37366 27716
rect 51506 27772 51570 27776
rect 51506 27716 51510 27772
rect 51510 27716 51566 27772
rect 51566 27716 51570 27772
rect 51506 27712 51570 27716
rect 51586 27772 51650 27776
rect 51586 27716 51590 27772
rect 51590 27716 51646 27772
rect 51646 27716 51650 27772
rect 51586 27712 51650 27716
rect 51666 27772 51730 27776
rect 51666 27716 51670 27772
rect 51670 27716 51726 27772
rect 51726 27716 51730 27772
rect 51666 27712 51730 27716
rect 51746 27772 51810 27776
rect 51746 27716 51750 27772
rect 51750 27716 51806 27772
rect 51806 27716 51810 27772
rect 51746 27712 51810 27716
rect 15396 27228 15460 27232
rect 15396 27172 15400 27228
rect 15400 27172 15456 27228
rect 15456 27172 15460 27228
rect 15396 27168 15460 27172
rect 15476 27228 15540 27232
rect 15476 27172 15480 27228
rect 15480 27172 15536 27228
rect 15536 27172 15540 27228
rect 15476 27168 15540 27172
rect 15556 27228 15620 27232
rect 15556 27172 15560 27228
rect 15560 27172 15616 27228
rect 15616 27172 15620 27228
rect 15556 27168 15620 27172
rect 15636 27228 15700 27232
rect 15636 27172 15640 27228
rect 15640 27172 15696 27228
rect 15696 27172 15700 27228
rect 15636 27168 15700 27172
rect 29840 27228 29904 27232
rect 29840 27172 29844 27228
rect 29844 27172 29900 27228
rect 29900 27172 29904 27228
rect 29840 27168 29904 27172
rect 29920 27228 29984 27232
rect 29920 27172 29924 27228
rect 29924 27172 29980 27228
rect 29980 27172 29984 27228
rect 29920 27168 29984 27172
rect 30000 27228 30064 27232
rect 30000 27172 30004 27228
rect 30004 27172 30060 27228
rect 30060 27172 30064 27228
rect 30000 27168 30064 27172
rect 30080 27228 30144 27232
rect 30080 27172 30084 27228
rect 30084 27172 30140 27228
rect 30140 27172 30144 27228
rect 30080 27168 30144 27172
rect 44284 27228 44348 27232
rect 44284 27172 44288 27228
rect 44288 27172 44344 27228
rect 44344 27172 44348 27228
rect 44284 27168 44348 27172
rect 44364 27228 44428 27232
rect 44364 27172 44368 27228
rect 44368 27172 44424 27228
rect 44424 27172 44428 27228
rect 44364 27168 44428 27172
rect 44444 27228 44508 27232
rect 44444 27172 44448 27228
rect 44448 27172 44504 27228
rect 44504 27172 44508 27228
rect 44444 27168 44508 27172
rect 44524 27228 44588 27232
rect 44524 27172 44528 27228
rect 44528 27172 44584 27228
rect 44584 27172 44588 27228
rect 44524 27168 44588 27172
rect 58728 27228 58792 27232
rect 58728 27172 58732 27228
rect 58732 27172 58788 27228
rect 58788 27172 58792 27228
rect 58728 27168 58792 27172
rect 58808 27228 58872 27232
rect 58808 27172 58812 27228
rect 58812 27172 58868 27228
rect 58868 27172 58872 27228
rect 58808 27168 58872 27172
rect 58888 27228 58952 27232
rect 58888 27172 58892 27228
rect 58892 27172 58948 27228
rect 58948 27172 58952 27228
rect 58888 27168 58952 27172
rect 58968 27228 59032 27232
rect 58968 27172 58972 27228
rect 58972 27172 59028 27228
rect 59028 27172 59032 27228
rect 58968 27168 59032 27172
rect 8174 26684 8238 26688
rect 8174 26628 8178 26684
rect 8178 26628 8234 26684
rect 8234 26628 8238 26684
rect 8174 26624 8238 26628
rect 8254 26684 8318 26688
rect 8254 26628 8258 26684
rect 8258 26628 8314 26684
rect 8314 26628 8318 26684
rect 8254 26624 8318 26628
rect 8334 26684 8398 26688
rect 8334 26628 8338 26684
rect 8338 26628 8394 26684
rect 8394 26628 8398 26684
rect 8334 26624 8398 26628
rect 8414 26684 8478 26688
rect 8414 26628 8418 26684
rect 8418 26628 8474 26684
rect 8474 26628 8478 26684
rect 8414 26624 8478 26628
rect 22618 26684 22682 26688
rect 22618 26628 22622 26684
rect 22622 26628 22678 26684
rect 22678 26628 22682 26684
rect 22618 26624 22682 26628
rect 22698 26684 22762 26688
rect 22698 26628 22702 26684
rect 22702 26628 22758 26684
rect 22758 26628 22762 26684
rect 22698 26624 22762 26628
rect 22778 26684 22842 26688
rect 22778 26628 22782 26684
rect 22782 26628 22838 26684
rect 22838 26628 22842 26684
rect 22778 26624 22842 26628
rect 22858 26684 22922 26688
rect 22858 26628 22862 26684
rect 22862 26628 22918 26684
rect 22918 26628 22922 26684
rect 22858 26624 22922 26628
rect 37062 26684 37126 26688
rect 37062 26628 37066 26684
rect 37066 26628 37122 26684
rect 37122 26628 37126 26684
rect 37062 26624 37126 26628
rect 37142 26684 37206 26688
rect 37142 26628 37146 26684
rect 37146 26628 37202 26684
rect 37202 26628 37206 26684
rect 37142 26624 37206 26628
rect 37222 26684 37286 26688
rect 37222 26628 37226 26684
rect 37226 26628 37282 26684
rect 37282 26628 37286 26684
rect 37222 26624 37286 26628
rect 37302 26684 37366 26688
rect 37302 26628 37306 26684
rect 37306 26628 37362 26684
rect 37362 26628 37366 26684
rect 37302 26624 37366 26628
rect 51506 26684 51570 26688
rect 51506 26628 51510 26684
rect 51510 26628 51566 26684
rect 51566 26628 51570 26684
rect 51506 26624 51570 26628
rect 51586 26684 51650 26688
rect 51586 26628 51590 26684
rect 51590 26628 51646 26684
rect 51646 26628 51650 26684
rect 51586 26624 51650 26628
rect 51666 26684 51730 26688
rect 51666 26628 51670 26684
rect 51670 26628 51726 26684
rect 51726 26628 51730 26684
rect 51666 26624 51730 26628
rect 51746 26684 51810 26688
rect 51746 26628 51750 26684
rect 51750 26628 51806 26684
rect 51806 26628 51810 26684
rect 51746 26624 51810 26628
rect 15396 26140 15460 26144
rect 15396 26084 15400 26140
rect 15400 26084 15456 26140
rect 15456 26084 15460 26140
rect 15396 26080 15460 26084
rect 15476 26140 15540 26144
rect 15476 26084 15480 26140
rect 15480 26084 15536 26140
rect 15536 26084 15540 26140
rect 15476 26080 15540 26084
rect 15556 26140 15620 26144
rect 15556 26084 15560 26140
rect 15560 26084 15616 26140
rect 15616 26084 15620 26140
rect 15556 26080 15620 26084
rect 15636 26140 15700 26144
rect 15636 26084 15640 26140
rect 15640 26084 15696 26140
rect 15696 26084 15700 26140
rect 15636 26080 15700 26084
rect 29840 26140 29904 26144
rect 29840 26084 29844 26140
rect 29844 26084 29900 26140
rect 29900 26084 29904 26140
rect 29840 26080 29904 26084
rect 29920 26140 29984 26144
rect 29920 26084 29924 26140
rect 29924 26084 29980 26140
rect 29980 26084 29984 26140
rect 29920 26080 29984 26084
rect 30000 26140 30064 26144
rect 30000 26084 30004 26140
rect 30004 26084 30060 26140
rect 30060 26084 30064 26140
rect 30000 26080 30064 26084
rect 30080 26140 30144 26144
rect 30080 26084 30084 26140
rect 30084 26084 30140 26140
rect 30140 26084 30144 26140
rect 30080 26080 30144 26084
rect 44284 26140 44348 26144
rect 44284 26084 44288 26140
rect 44288 26084 44344 26140
rect 44344 26084 44348 26140
rect 44284 26080 44348 26084
rect 44364 26140 44428 26144
rect 44364 26084 44368 26140
rect 44368 26084 44424 26140
rect 44424 26084 44428 26140
rect 44364 26080 44428 26084
rect 44444 26140 44508 26144
rect 44444 26084 44448 26140
rect 44448 26084 44504 26140
rect 44504 26084 44508 26140
rect 44444 26080 44508 26084
rect 44524 26140 44588 26144
rect 44524 26084 44528 26140
rect 44528 26084 44584 26140
rect 44584 26084 44588 26140
rect 44524 26080 44588 26084
rect 58728 26140 58792 26144
rect 58728 26084 58732 26140
rect 58732 26084 58788 26140
rect 58788 26084 58792 26140
rect 58728 26080 58792 26084
rect 58808 26140 58872 26144
rect 58808 26084 58812 26140
rect 58812 26084 58868 26140
rect 58868 26084 58872 26140
rect 58808 26080 58872 26084
rect 58888 26140 58952 26144
rect 58888 26084 58892 26140
rect 58892 26084 58948 26140
rect 58948 26084 58952 26140
rect 58888 26080 58952 26084
rect 58968 26140 59032 26144
rect 58968 26084 58972 26140
rect 58972 26084 59028 26140
rect 59028 26084 59032 26140
rect 58968 26080 59032 26084
rect 8174 25596 8238 25600
rect 8174 25540 8178 25596
rect 8178 25540 8234 25596
rect 8234 25540 8238 25596
rect 8174 25536 8238 25540
rect 8254 25596 8318 25600
rect 8254 25540 8258 25596
rect 8258 25540 8314 25596
rect 8314 25540 8318 25596
rect 8254 25536 8318 25540
rect 8334 25596 8398 25600
rect 8334 25540 8338 25596
rect 8338 25540 8394 25596
rect 8394 25540 8398 25596
rect 8334 25536 8398 25540
rect 8414 25596 8478 25600
rect 8414 25540 8418 25596
rect 8418 25540 8474 25596
rect 8474 25540 8478 25596
rect 8414 25536 8478 25540
rect 22618 25596 22682 25600
rect 22618 25540 22622 25596
rect 22622 25540 22678 25596
rect 22678 25540 22682 25596
rect 22618 25536 22682 25540
rect 22698 25596 22762 25600
rect 22698 25540 22702 25596
rect 22702 25540 22758 25596
rect 22758 25540 22762 25596
rect 22698 25536 22762 25540
rect 22778 25596 22842 25600
rect 22778 25540 22782 25596
rect 22782 25540 22838 25596
rect 22838 25540 22842 25596
rect 22778 25536 22842 25540
rect 22858 25596 22922 25600
rect 22858 25540 22862 25596
rect 22862 25540 22918 25596
rect 22918 25540 22922 25596
rect 22858 25536 22922 25540
rect 37062 25596 37126 25600
rect 37062 25540 37066 25596
rect 37066 25540 37122 25596
rect 37122 25540 37126 25596
rect 37062 25536 37126 25540
rect 37142 25596 37206 25600
rect 37142 25540 37146 25596
rect 37146 25540 37202 25596
rect 37202 25540 37206 25596
rect 37142 25536 37206 25540
rect 37222 25596 37286 25600
rect 37222 25540 37226 25596
rect 37226 25540 37282 25596
rect 37282 25540 37286 25596
rect 37222 25536 37286 25540
rect 37302 25596 37366 25600
rect 37302 25540 37306 25596
rect 37306 25540 37362 25596
rect 37362 25540 37366 25596
rect 37302 25536 37366 25540
rect 51506 25596 51570 25600
rect 51506 25540 51510 25596
rect 51510 25540 51566 25596
rect 51566 25540 51570 25596
rect 51506 25536 51570 25540
rect 51586 25596 51650 25600
rect 51586 25540 51590 25596
rect 51590 25540 51646 25596
rect 51646 25540 51650 25596
rect 51586 25536 51650 25540
rect 51666 25596 51730 25600
rect 51666 25540 51670 25596
rect 51670 25540 51726 25596
rect 51726 25540 51730 25596
rect 51666 25536 51730 25540
rect 51746 25596 51810 25600
rect 51746 25540 51750 25596
rect 51750 25540 51806 25596
rect 51806 25540 51810 25596
rect 51746 25536 51810 25540
rect 15396 25052 15460 25056
rect 15396 24996 15400 25052
rect 15400 24996 15456 25052
rect 15456 24996 15460 25052
rect 15396 24992 15460 24996
rect 15476 25052 15540 25056
rect 15476 24996 15480 25052
rect 15480 24996 15536 25052
rect 15536 24996 15540 25052
rect 15476 24992 15540 24996
rect 15556 25052 15620 25056
rect 15556 24996 15560 25052
rect 15560 24996 15616 25052
rect 15616 24996 15620 25052
rect 15556 24992 15620 24996
rect 15636 25052 15700 25056
rect 15636 24996 15640 25052
rect 15640 24996 15696 25052
rect 15696 24996 15700 25052
rect 15636 24992 15700 24996
rect 29840 25052 29904 25056
rect 29840 24996 29844 25052
rect 29844 24996 29900 25052
rect 29900 24996 29904 25052
rect 29840 24992 29904 24996
rect 29920 25052 29984 25056
rect 29920 24996 29924 25052
rect 29924 24996 29980 25052
rect 29980 24996 29984 25052
rect 29920 24992 29984 24996
rect 30000 25052 30064 25056
rect 30000 24996 30004 25052
rect 30004 24996 30060 25052
rect 30060 24996 30064 25052
rect 30000 24992 30064 24996
rect 30080 25052 30144 25056
rect 30080 24996 30084 25052
rect 30084 24996 30140 25052
rect 30140 24996 30144 25052
rect 30080 24992 30144 24996
rect 44284 25052 44348 25056
rect 44284 24996 44288 25052
rect 44288 24996 44344 25052
rect 44344 24996 44348 25052
rect 44284 24992 44348 24996
rect 44364 25052 44428 25056
rect 44364 24996 44368 25052
rect 44368 24996 44424 25052
rect 44424 24996 44428 25052
rect 44364 24992 44428 24996
rect 44444 25052 44508 25056
rect 44444 24996 44448 25052
rect 44448 24996 44504 25052
rect 44504 24996 44508 25052
rect 44444 24992 44508 24996
rect 44524 25052 44588 25056
rect 44524 24996 44528 25052
rect 44528 24996 44584 25052
rect 44584 24996 44588 25052
rect 44524 24992 44588 24996
rect 58728 25052 58792 25056
rect 58728 24996 58732 25052
rect 58732 24996 58788 25052
rect 58788 24996 58792 25052
rect 58728 24992 58792 24996
rect 58808 25052 58872 25056
rect 58808 24996 58812 25052
rect 58812 24996 58868 25052
rect 58868 24996 58872 25052
rect 58808 24992 58872 24996
rect 58888 25052 58952 25056
rect 58888 24996 58892 25052
rect 58892 24996 58948 25052
rect 58948 24996 58952 25052
rect 58888 24992 58952 24996
rect 58968 25052 59032 25056
rect 58968 24996 58972 25052
rect 58972 24996 59028 25052
rect 59028 24996 59032 25052
rect 58968 24992 59032 24996
rect 8174 24508 8238 24512
rect 8174 24452 8178 24508
rect 8178 24452 8234 24508
rect 8234 24452 8238 24508
rect 8174 24448 8238 24452
rect 8254 24508 8318 24512
rect 8254 24452 8258 24508
rect 8258 24452 8314 24508
rect 8314 24452 8318 24508
rect 8254 24448 8318 24452
rect 8334 24508 8398 24512
rect 8334 24452 8338 24508
rect 8338 24452 8394 24508
rect 8394 24452 8398 24508
rect 8334 24448 8398 24452
rect 8414 24508 8478 24512
rect 8414 24452 8418 24508
rect 8418 24452 8474 24508
rect 8474 24452 8478 24508
rect 8414 24448 8478 24452
rect 22618 24508 22682 24512
rect 22618 24452 22622 24508
rect 22622 24452 22678 24508
rect 22678 24452 22682 24508
rect 22618 24448 22682 24452
rect 22698 24508 22762 24512
rect 22698 24452 22702 24508
rect 22702 24452 22758 24508
rect 22758 24452 22762 24508
rect 22698 24448 22762 24452
rect 22778 24508 22842 24512
rect 22778 24452 22782 24508
rect 22782 24452 22838 24508
rect 22838 24452 22842 24508
rect 22778 24448 22842 24452
rect 22858 24508 22922 24512
rect 22858 24452 22862 24508
rect 22862 24452 22918 24508
rect 22918 24452 22922 24508
rect 22858 24448 22922 24452
rect 37062 24508 37126 24512
rect 37062 24452 37066 24508
rect 37066 24452 37122 24508
rect 37122 24452 37126 24508
rect 37062 24448 37126 24452
rect 37142 24508 37206 24512
rect 37142 24452 37146 24508
rect 37146 24452 37202 24508
rect 37202 24452 37206 24508
rect 37142 24448 37206 24452
rect 37222 24508 37286 24512
rect 37222 24452 37226 24508
rect 37226 24452 37282 24508
rect 37282 24452 37286 24508
rect 37222 24448 37286 24452
rect 37302 24508 37366 24512
rect 37302 24452 37306 24508
rect 37306 24452 37362 24508
rect 37362 24452 37366 24508
rect 37302 24448 37366 24452
rect 51506 24508 51570 24512
rect 51506 24452 51510 24508
rect 51510 24452 51566 24508
rect 51566 24452 51570 24508
rect 51506 24448 51570 24452
rect 51586 24508 51650 24512
rect 51586 24452 51590 24508
rect 51590 24452 51646 24508
rect 51646 24452 51650 24508
rect 51586 24448 51650 24452
rect 51666 24508 51730 24512
rect 51666 24452 51670 24508
rect 51670 24452 51726 24508
rect 51726 24452 51730 24508
rect 51666 24448 51730 24452
rect 51746 24508 51810 24512
rect 51746 24452 51750 24508
rect 51750 24452 51806 24508
rect 51806 24452 51810 24508
rect 51746 24448 51810 24452
rect 15396 23964 15460 23968
rect 15396 23908 15400 23964
rect 15400 23908 15456 23964
rect 15456 23908 15460 23964
rect 15396 23904 15460 23908
rect 15476 23964 15540 23968
rect 15476 23908 15480 23964
rect 15480 23908 15536 23964
rect 15536 23908 15540 23964
rect 15476 23904 15540 23908
rect 15556 23964 15620 23968
rect 15556 23908 15560 23964
rect 15560 23908 15616 23964
rect 15616 23908 15620 23964
rect 15556 23904 15620 23908
rect 15636 23964 15700 23968
rect 15636 23908 15640 23964
rect 15640 23908 15696 23964
rect 15696 23908 15700 23964
rect 15636 23904 15700 23908
rect 29840 23964 29904 23968
rect 29840 23908 29844 23964
rect 29844 23908 29900 23964
rect 29900 23908 29904 23964
rect 29840 23904 29904 23908
rect 29920 23964 29984 23968
rect 29920 23908 29924 23964
rect 29924 23908 29980 23964
rect 29980 23908 29984 23964
rect 29920 23904 29984 23908
rect 30000 23964 30064 23968
rect 30000 23908 30004 23964
rect 30004 23908 30060 23964
rect 30060 23908 30064 23964
rect 30000 23904 30064 23908
rect 30080 23964 30144 23968
rect 30080 23908 30084 23964
rect 30084 23908 30140 23964
rect 30140 23908 30144 23964
rect 30080 23904 30144 23908
rect 44284 23964 44348 23968
rect 44284 23908 44288 23964
rect 44288 23908 44344 23964
rect 44344 23908 44348 23964
rect 44284 23904 44348 23908
rect 44364 23964 44428 23968
rect 44364 23908 44368 23964
rect 44368 23908 44424 23964
rect 44424 23908 44428 23964
rect 44364 23904 44428 23908
rect 44444 23964 44508 23968
rect 44444 23908 44448 23964
rect 44448 23908 44504 23964
rect 44504 23908 44508 23964
rect 44444 23904 44508 23908
rect 44524 23964 44588 23968
rect 44524 23908 44528 23964
rect 44528 23908 44584 23964
rect 44584 23908 44588 23964
rect 44524 23904 44588 23908
rect 58728 23964 58792 23968
rect 58728 23908 58732 23964
rect 58732 23908 58788 23964
rect 58788 23908 58792 23964
rect 58728 23904 58792 23908
rect 58808 23964 58872 23968
rect 58808 23908 58812 23964
rect 58812 23908 58868 23964
rect 58868 23908 58872 23964
rect 58808 23904 58872 23908
rect 58888 23964 58952 23968
rect 58888 23908 58892 23964
rect 58892 23908 58948 23964
rect 58948 23908 58952 23964
rect 58888 23904 58952 23908
rect 58968 23964 59032 23968
rect 58968 23908 58972 23964
rect 58972 23908 59028 23964
rect 59028 23908 59032 23964
rect 58968 23904 59032 23908
rect 8174 23420 8238 23424
rect 8174 23364 8178 23420
rect 8178 23364 8234 23420
rect 8234 23364 8238 23420
rect 8174 23360 8238 23364
rect 8254 23420 8318 23424
rect 8254 23364 8258 23420
rect 8258 23364 8314 23420
rect 8314 23364 8318 23420
rect 8254 23360 8318 23364
rect 8334 23420 8398 23424
rect 8334 23364 8338 23420
rect 8338 23364 8394 23420
rect 8394 23364 8398 23420
rect 8334 23360 8398 23364
rect 8414 23420 8478 23424
rect 8414 23364 8418 23420
rect 8418 23364 8474 23420
rect 8474 23364 8478 23420
rect 8414 23360 8478 23364
rect 22618 23420 22682 23424
rect 22618 23364 22622 23420
rect 22622 23364 22678 23420
rect 22678 23364 22682 23420
rect 22618 23360 22682 23364
rect 22698 23420 22762 23424
rect 22698 23364 22702 23420
rect 22702 23364 22758 23420
rect 22758 23364 22762 23420
rect 22698 23360 22762 23364
rect 22778 23420 22842 23424
rect 22778 23364 22782 23420
rect 22782 23364 22838 23420
rect 22838 23364 22842 23420
rect 22778 23360 22842 23364
rect 22858 23420 22922 23424
rect 22858 23364 22862 23420
rect 22862 23364 22918 23420
rect 22918 23364 22922 23420
rect 22858 23360 22922 23364
rect 37062 23420 37126 23424
rect 37062 23364 37066 23420
rect 37066 23364 37122 23420
rect 37122 23364 37126 23420
rect 37062 23360 37126 23364
rect 37142 23420 37206 23424
rect 37142 23364 37146 23420
rect 37146 23364 37202 23420
rect 37202 23364 37206 23420
rect 37142 23360 37206 23364
rect 37222 23420 37286 23424
rect 37222 23364 37226 23420
rect 37226 23364 37282 23420
rect 37282 23364 37286 23420
rect 37222 23360 37286 23364
rect 37302 23420 37366 23424
rect 37302 23364 37306 23420
rect 37306 23364 37362 23420
rect 37362 23364 37366 23420
rect 37302 23360 37366 23364
rect 51506 23420 51570 23424
rect 51506 23364 51510 23420
rect 51510 23364 51566 23420
rect 51566 23364 51570 23420
rect 51506 23360 51570 23364
rect 51586 23420 51650 23424
rect 51586 23364 51590 23420
rect 51590 23364 51646 23420
rect 51646 23364 51650 23420
rect 51586 23360 51650 23364
rect 51666 23420 51730 23424
rect 51666 23364 51670 23420
rect 51670 23364 51726 23420
rect 51726 23364 51730 23420
rect 51666 23360 51730 23364
rect 51746 23420 51810 23424
rect 51746 23364 51750 23420
rect 51750 23364 51806 23420
rect 51806 23364 51810 23420
rect 51746 23360 51810 23364
rect 15396 22876 15460 22880
rect 15396 22820 15400 22876
rect 15400 22820 15456 22876
rect 15456 22820 15460 22876
rect 15396 22816 15460 22820
rect 15476 22876 15540 22880
rect 15476 22820 15480 22876
rect 15480 22820 15536 22876
rect 15536 22820 15540 22876
rect 15476 22816 15540 22820
rect 15556 22876 15620 22880
rect 15556 22820 15560 22876
rect 15560 22820 15616 22876
rect 15616 22820 15620 22876
rect 15556 22816 15620 22820
rect 15636 22876 15700 22880
rect 15636 22820 15640 22876
rect 15640 22820 15696 22876
rect 15696 22820 15700 22876
rect 15636 22816 15700 22820
rect 29840 22876 29904 22880
rect 29840 22820 29844 22876
rect 29844 22820 29900 22876
rect 29900 22820 29904 22876
rect 29840 22816 29904 22820
rect 29920 22876 29984 22880
rect 29920 22820 29924 22876
rect 29924 22820 29980 22876
rect 29980 22820 29984 22876
rect 29920 22816 29984 22820
rect 30000 22876 30064 22880
rect 30000 22820 30004 22876
rect 30004 22820 30060 22876
rect 30060 22820 30064 22876
rect 30000 22816 30064 22820
rect 30080 22876 30144 22880
rect 30080 22820 30084 22876
rect 30084 22820 30140 22876
rect 30140 22820 30144 22876
rect 30080 22816 30144 22820
rect 44284 22876 44348 22880
rect 44284 22820 44288 22876
rect 44288 22820 44344 22876
rect 44344 22820 44348 22876
rect 44284 22816 44348 22820
rect 44364 22876 44428 22880
rect 44364 22820 44368 22876
rect 44368 22820 44424 22876
rect 44424 22820 44428 22876
rect 44364 22816 44428 22820
rect 44444 22876 44508 22880
rect 44444 22820 44448 22876
rect 44448 22820 44504 22876
rect 44504 22820 44508 22876
rect 44444 22816 44508 22820
rect 44524 22876 44588 22880
rect 44524 22820 44528 22876
rect 44528 22820 44584 22876
rect 44584 22820 44588 22876
rect 44524 22816 44588 22820
rect 58728 22876 58792 22880
rect 58728 22820 58732 22876
rect 58732 22820 58788 22876
rect 58788 22820 58792 22876
rect 58728 22816 58792 22820
rect 58808 22876 58872 22880
rect 58808 22820 58812 22876
rect 58812 22820 58868 22876
rect 58868 22820 58872 22876
rect 58808 22816 58872 22820
rect 58888 22876 58952 22880
rect 58888 22820 58892 22876
rect 58892 22820 58948 22876
rect 58948 22820 58952 22876
rect 58888 22816 58952 22820
rect 58968 22876 59032 22880
rect 58968 22820 58972 22876
rect 58972 22820 59028 22876
rect 59028 22820 59032 22876
rect 58968 22816 59032 22820
rect 8174 22332 8238 22336
rect 8174 22276 8178 22332
rect 8178 22276 8234 22332
rect 8234 22276 8238 22332
rect 8174 22272 8238 22276
rect 8254 22332 8318 22336
rect 8254 22276 8258 22332
rect 8258 22276 8314 22332
rect 8314 22276 8318 22332
rect 8254 22272 8318 22276
rect 8334 22332 8398 22336
rect 8334 22276 8338 22332
rect 8338 22276 8394 22332
rect 8394 22276 8398 22332
rect 8334 22272 8398 22276
rect 8414 22332 8478 22336
rect 8414 22276 8418 22332
rect 8418 22276 8474 22332
rect 8474 22276 8478 22332
rect 8414 22272 8478 22276
rect 22618 22332 22682 22336
rect 22618 22276 22622 22332
rect 22622 22276 22678 22332
rect 22678 22276 22682 22332
rect 22618 22272 22682 22276
rect 22698 22332 22762 22336
rect 22698 22276 22702 22332
rect 22702 22276 22758 22332
rect 22758 22276 22762 22332
rect 22698 22272 22762 22276
rect 22778 22332 22842 22336
rect 22778 22276 22782 22332
rect 22782 22276 22838 22332
rect 22838 22276 22842 22332
rect 22778 22272 22842 22276
rect 22858 22332 22922 22336
rect 22858 22276 22862 22332
rect 22862 22276 22918 22332
rect 22918 22276 22922 22332
rect 22858 22272 22922 22276
rect 37062 22332 37126 22336
rect 37062 22276 37066 22332
rect 37066 22276 37122 22332
rect 37122 22276 37126 22332
rect 37062 22272 37126 22276
rect 37142 22332 37206 22336
rect 37142 22276 37146 22332
rect 37146 22276 37202 22332
rect 37202 22276 37206 22332
rect 37142 22272 37206 22276
rect 37222 22332 37286 22336
rect 37222 22276 37226 22332
rect 37226 22276 37282 22332
rect 37282 22276 37286 22332
rect 37222 22272 37286 22276
rect 37302 22332 37366 22336
rect 37302 22276 37306 22332
rect 37306 22276 37362 22332
rect 37362 22276 37366 22332
rect 37302 22272 37366 22276
rect 51506 22332 51570 22336
rect 51506 22276 51510 22332
rect 51510 22276 51566 22332
rect 51566 22276 51570 22332
rect 51506 22272 51570 22276
rect 51586 22332 51650 22336
rect 51586 22276 51590 22332
rect 51590 22276 51646 22332
rect 51646 22276 51650 22332
rect 51586 22272 51650 22276
rect 51666 22332 51730 22336
rect 51666 22276 51670 22332
rect 51670 22276 51726 22332
rect 51726 22276 51730 22332
rect 51666 22272 51730 22276
rect 51746 22332 51810 22336
rect 51746 22276 51750 22332
rect 51750 22276 51806 22332
rect 51806 22276 51810 22332
rect 51746 22272 51810 22276
rect 15396 21788 15460 21792
rect 15396 21732 15400 21788
rect 15400 21732 15456 21788
rect 15456 21732 15460 21788
rect 15396 21728 15460 21732
rect 15476 21788 15540 21792
rect 15476 21732 15480 21788
rect 15480 21732 15536 21788
rect 15536 21732 15540 21788
rect 15476 21728 15540 21732
rect 15556 21788 15620 21792
rect 15556 21732 15560 21788
rect 15560 21732 15616 21788
rect 15616 21732 15620 21788
rect 15556 21728 15620 21732
rect 15636 21788 15700 21792
rect 15636 21732 15640 21788
rect 15640 21732 15696 21788
rect 15696 21732 15700 21788
rect 15636 21728 15700 21732
rect 29840 21788 29904 21792
rect 29840 21732 29844 21788
rect 29844 21732 29900 21788
rect 29900 21732 29904 21788
rect 29840 21728 29904 21732
rect 29920 21788 29984 21792
rect 29920 21732 29924 21788
rect 29924 21732 29980 21788
rect 29980 21732 29984 21788
rect 29920 21728 29984 21732
rect 30000 21788 30064 21792
rect 30000 21732 30004 21788
rect 30004 21732 30060 21788
rect 30060 21732 30064 21788
rect 30000 21728 30064 21732
rect 30080 21788 30144 21792
rect 30080 21732 30084 21788
rect 30084 21732 30140 21788
rect 30140 21732 30144 21788
rect 30080 21728 30144 21732
rect 44284 21788 44348 21792
rect 44284 21732 44288 21788
rect 44288 21732 44344 21788
rect 44344 21732 44348 21788
rect 44284 21728 44348 21732
rect 44364 21788 44428 21792
rect 44364 21732 44368 21788
rect 44368 21732 44424 21788
rect 44424 21732 44428 21788
rect 44364 21728 44428 21732
rect 44444 21788 44508 21792
rect 44444 21732 44448 21788
rect 44448 21732 44504 21788
rect 44504 21732 44508 21788
rect 44444 21728 44508 21732
rect 44524 21788 44588 21792
rect 44524 21732 44528 21788
rect 44528 21732 44584 21788
rect 44584 21732 44588 21788
rect 44524 21728 44588 21732
rect 58728 21788 58792 21792
rect 58728 21732 58732 21788
rect 58732 21732 58788 21788
rect 58788 21732 58792 21788
rect 58728 21728 58792 21732
rect 58808 21788 58872 21792
rect 58808 21732 58812 21788
rect 58812 21732 58868 21788
rect 58868 21732 58872 21788
rect 58808 21728 58872 21732
rect 58888 21788 58952 21792
rect 58888 21732 58892 21788
rect 58892 21732 58948 21788
rect 58948 21732 58952 21788
rect 58888 21728 58952 21732
rect 58968 21788 59032 21792
rect 58968 21732 58972 21788
rect 58972 21732 59028 21788
rect 59028 21732 59032 21788
rect 58968 21728 59032 21732
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 22618 21244 22682 21248
rect 22618 21188 22622 21244
rect 22622 21188 22678 21244
rect 22678 21188 22682 21244
rect 22618 21184 22682 21188
rect 22698 21244 22762 21248
rect 22698 21188 22702 21244
rect 22702 21188 22758 21244
rect 22758 21188 22762 21244
rect 22698 21184 22762 21188
rect 22778 21244 22842 21248
rect 22778 21188 22782 21244
rect 22782 21188 22838 21244
rect 22838 21188 22842 21244
rect 22778 21184 22842 21188
rect 22858 21244 22922 21248
rect 22858 21188 22862 21244
rect 22862 21188 22918 21244
rect 22918 21188 22922 21244
rect 22858 21184 22922 21188
rect 37062 21244 37126 21248
rect 37062 21188 37066 21244
rect 37066 21188 37122 21244
rect 37122 21188 37126 21244
rect 37062 21184 37126 21188
rect 37142 21244 37206 21248
rect 37142 21188 37146 21244
rect 37146 21188 37202 21244
rect 37202 21188 37206 21244
rect 37142 21184 37206 21188
rect 37222 21244 37286 21248
rect 37222 21188 37226 21244
rect 37226 21188 37282 21244
rect 37282 21188 37286 21244
rect 37222 21184 37286 21188
rect 37302 21244 37366 21248
rect 37302 21188 37306 21244
rect 37306 21188 37362 21244
rect 37362 21188 37366 21244
rect 37302 21184 37366 21188
rect 51506 21244 51570 21248
rect 51506 21188 51510 21244
rect 51510 21188 51566 21244
rect 51566 21188 51570 21244
rect 51506 21184 51570 21188
rect 51586 21244 51650 21248
rect 51586 21188 51590 21244
rect 51590 21188 51646 21244
rect 51646 21188 51650 21244
rect 51586 21184 51650 21188
rect 51666 21244 51730 21248
rect 51666 21188 51670 21244
rect 51670 21188 51726 21244
rect 51726 21188 51730 21244
rect 51666 21184 51730 21188
rect 51746 21244 51810 21248
rect 51746 21188 51750 21244
rect 51750 21188 51806 21244
rect 51806 21188 51810 21244
rect 51746 21184 51810 21188
rect 16436 20768 16500 20772
rect 16436 20712 16486 20768
rect 16486 20712 16500 20768
rect 16436 20708 16500 20712
rect 15396 20700 15460 20704
rect 15396 20644 15400 20700
rect 15400 20644 15456 20700
rect 15456 20644 15460 20700
rect 15396 20640 15460 20644
rect 15476 20700 15540 20704
rect 15476 20644 15480 20700
rect 15480 20644 15536 20700
rect 15536 20644 15540 20700
rect 15476 20640 15540 20644
rect 15556 20700 15620 20704
rect 15556 20644 15560 20700
rect 15560 20644 15616 20700
rect 15616 20644 15620 20700
rect 15556 20640 15620 20644
rect 15636 20700 15700 20704
rect 15636 20644 15640 20700
rect 15640 20644 15696 20700
rect 15696 20644 15700 20700
rect 15636 20640 15700 20644
rect 29840 20700 29904 20704
rect 29840 20644 29844 20700
rect 29844 20644 29900 20700
rect 29900 20644 29904 20700
rect 29840 20640 29904 20644
rect 29920 20700 29984 20704
rect 29920 20644 29924 20700
rect 29924 20644 29980 20700
rect 29980 20644 29984 20700
rect 29920 20640 29984 20644
rect 30000 20700 30064 20704
rect 30000 20644 30004 20700
rect 30004 20644 30060 20700
rect 30060 20644 30064 20700
rect 30000 20640 30064 20644
rect 30080 20700 30144 20704
rect 30080 20644 30084 20700
rect 30084 20644 30140 20700
rect 30140 20644 30144 20700
rect 30080 20640 30144 20644
rect 44284 20700 44348 20704
rect 44284 20644 44288 20700
rect 44288 20644 44344 20700
rect 44344 20644 44348 20700
rect 44284 20640 44348 20644
rect 44364 20700 44428 20704
rect 44364 20644 44368 20700
rect 44368 20644 44424 20700
rect 44424 20644 44428 20700
rect 44364 20640 44428 20644
rect 44444 20700 44508 20704
rect 44444 20644 44448 20700
rect 44448 20644 44504 20700
rect 44504 20644 44508 20700
rect 44444 20640 44508 20644
rect 44524 20700 44588 20704
rect 44524 20644 44528 20700
rect 44528 20644 44584 20700
rect 44584 20644 44588 20700
rect 44524 20640 44588 20644
rect 58728 20700 58792 20704
rect 58728 20644 58732 20700
rect 58732 20644 58788 20700
rect 58788 20644 58792 20700
rect 58728 20640 58792 20644
rect 58808 20700 58872 20704
rect 58808 20644 58812 20700
rect 58812 20644 58868 20700
rect 58868 20644 58872 20700
rect 58808 20640 58872 20644
rect 58888 20700 58952 20704
rect 58888 20644 58892 20700
rect 58892 20644 58948 20700
rect 58948 20644 58952 20700
rect 58888 20640 58952 20644
rect 58968 20700 59032 20704
rect 58968 20644 58972 20700
rect 58972 20644 59028 20700
rect 59028 20644 59032 20700
rect 58968 20640 59032 20644
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 22618 20156 22682 20160
rect 22618 20100 22622 20156
rect 22622 20100 22678 20156
rect 22678 20100 22682 20156
rect 22618 20096 22682 20100
rect 22698 20156 22762 20160
rect 22698 20100 22702 20156
rect 22702 20100 22758 20156
rect 22758 20100 22762 20156
rect 22698 20096 22762 20100
rect 22778 20156 22842 20160
rect 22778 20100 22782 20156
rect 22782 20100 22838 20156
rect 22838 20100 22842 20156
rect 22778 20096 22842 20100
rect 22858 20156 22922 20160
rect 22858 20100 22862 20156
rect 22862 20100 22918 20156
rect 22918 20100 22922 20156
rect 22858 20096 22922 20100
rect 37062 20156 37126 20160
rect 37062 20100 37066 20156
rect 37066 20100 37122 20156
rect 37122 20100 37126 20156
rect 37062 20096 37126 20100
rect 37142 20156 37206 20160
rect 37142 20100 37146 20156
rect 37146 20100 37202 20156
rect 37202 20100 37206 20156
rect 37142 20096 37206 20100
rect 37222 20156 37286 20160
rect 37222 20100 37226 20156
rect 37226 20100 37282 20156
rect 37282 20100 37286 20156
rect 37222 20096 37286 20100
rect 37302 20156 37366 20160
rect 37302 20100 37306 20156
rect 37306 20100 37362 20156
rect 37362 20100 37366 20156
rect 37302 20096 37366 20100
rect 51506 20156 51570 20160
rect 51506 20100 51510 20156
rect 51510 20100 51566 20156
rect 51566 20100 51570 20156
rect 51506 20096 51570 20100
rect 51586 20156 51650 20160
rect 51586 20100 51590 20156
rect 51590 20100 51646 20156
rect 51646 20100 51650 20156
rect 51586 20096 51650 20100
rect 51666 20156 51730 20160
rect 51666 20100 51670 20156
rect 51670 20100 51726 20156
rect 51726 20100 51730 20156
rect 51666 20096 51730 20100
rect 51746 20156 51810 20160
rect 51746 20100 51750 20156
rect 51750 20100 51806 20156
rect 51806 20100 51810 20156
rect 51746 20096 51810 20100
rect 15396 19612 15460 19616
rect 15396 19556 15400 19612
rect 15400 19556 15456 19612
rect 15456 19556 15460 19612
rect 15396 19552 15460 19556
rect 15476 19612 15540 19616
rect 15476 19556 15480 19612
rect 15480 19556 15536 19612
rect 15536 19556 15540 19612
rect 15476 19552 15540 19556
rect 15556 19612 15620 19616
rect 15556 19556 15560 19612
rect 15560 19556 15616 19612
rect 15616 19556 15620 19612
rect 15556 19552 15620 19556
rect 15636 19612 15700 19616
rect 15636 19556 15640 19612
rect 15640 19556 15696 19612
rect 15696 19556 15700 19612
rect 15636 19552 15700 19556
rect 29840 19612 29904 19616
rect 29840 19556 29844 19612
rect 29844 19556 29900 19612
rect 29900 19556 29904 19612
rect 29840 19552 29904 19556
rect 29920 19612 29984 19616
rect 29920 19556 29924 19612
rect 29924 19556 29980 19612
rect 29980 19556 29984 19612
rect 29920 19552 29984 19556
rect 30000 19612 30064 19616
rect 30000 19556 30004 19612
rect 30004 19556 30060 19612
rect 30060 19556 30064 19612
rect 30000 19552 30064 19556
rect 30080 19612 30144 19616
rect 30080 19556 30084 19612
rect 30084 19556 30140 19612
rect 30140 19556 30144 19612
rect 30080 19552 30144 19556
rect 44284 19612 44348 19616
rect 44284 19556 44288 19612
rect 44288 19556 44344 19612
rect 44344 19556 44348 19612
rect 44284 19552 44348 19556
rect 44364 19612 44428 19616
rect 44364 19556 44368 19612
rect 44368 19556 44424 19612
rect 44424 19556 44428 19612
rect 44364 19552 44428 19556
rect 44444 19612 44508 19616
rect 44444 19556 44448 19612
rect 44448 19556 44504 19612
rect 44504 19556 44508 19612
rect 44444 19552 44508 19556
rect 44524 19612 44588 19616
rect 44524 19556 44528 19612
rect 44528 19556 44584 19612
rect 44584 19556 44588 19612
rect 44524 19552 44588 19556
rect 58728 19612 58792 19616
rect 58728 19556 58732 19612
rect 58732 19556 58788 19612
rect 58788 19556 58792 19612
rect 58728 19552 58792 19556
rect 58808 19612 58872 19616
rect 58808 19556 58812 19612
rect 58812 19556 58868 19612
rect 58868 19556 58872 19612
rect 58808 19552 58872 19556
rect 58888 19612 58952 19616
rect 58888 19556 58892 19612
rect 58892 19556 58948 19612
rect 58948 19556 58952 19612
rect 58888 19552 58952 19556
rect 58968 19612 59032 19616
rect 58968 19556 58972 19612
rect 58972 19556 59028 19612
rect 59028 19556 59032 19612
rect 58968 19552 59032 19556
rect 6684 19348 6748 19412
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 22618 19068 22682 19072
rect 22618 19012 22622 19068
rect 22622 19012 22678 19068
rect 22678 19012 22682 19068
rect 22618 19008 22682 19012
rect 22698 19068 22762 19072
rect 22698 19012 22702 19068
rect 22702 19012 22758 19068
rect 22758 19012 22762 19068
rect 22698 19008 22762 19012
rect 22778 19068 22842 19072
rect 22778 19012 22782 19068
rect 22782 19012 22838 19068
rect 22838 19012 22842 19068
rect 22778 19008 22842 19012
rect 22858 19068 22922 19072
rect 22858 19012 22862 19068
rect 22862 19012 22918 19068
rect 22918 19012 22922 19068
rect 22858 19008 22922 19012
rect 37062 19068 37126 19072
rect 37062 19012 37066 19068
rect 37066 19012 37122 19068
rect 37122 19012 37126 19068
rect 37062 19008 37126 19012
rect 37142 19068 37206 19072
rect 37142 19012 37146 19068
rect 37146 19012 37202 19068
rect 37202 19012 37206 19068
rect 37142 19008 37206 19012
rect 37222 19068 37286 19072
rect 37222 19012 37226 19068
rect 37226 19012 37282 19068
rect 37282 19012 37286 19068
rect 37222 19008 37286 19012
rect 37302 19068 37366 19072
rect 37302 19012 37306 19068
rect 37306 19012 37362 19068
rect 37362 19012 37366 19068
rect 37302 19008 37366 19012
rect 51506 19068 51570 19072
rect 51506 19012 51510 19068
rect 51510 19012 51566 19068
rect 51566 19012 51570 19068
rect 51506 19008 51570 19012
rect 51586 19068 51650 19072
rect 51586 19012 51590 19068
rect 51590 19012 51646 19068
rect 51646 19012 51650 19068
rect 51586 19008 51650 19012
rect 51666 19068 51730 19072
rect 51666 19012 51670 19068
rect 51670 19012 51726 19068
rect 51726 19012 51730 19068
rect 51666 19008 51730 19012
rect 51746 19068 51810 19072
rect 51746 19012 51750 19068
rect 51750 19012 51806 19068
rect 51806 19012 51810 19068
rect 51746 19008 51810 19012
rect 15396 18524 15460 18528
rect 15396 18468 15400 18524
rect 15400 18468 15456 18524
rect 15456 18468 15460 18524
rect 15396 18464 15460 18468
rect 15476 18524 15540 18528
rect 15476 18468 15480 18524
rect 15480 18468 15536 18524
rect 15536 18468 15540 18524
rect 15476 18464 15540 18468
rect 15556 18524 15620 18528
rect 15556 18468 15560 18524
rect 15560 18468 15616 18524
rect 15616 18468 15620 18524
rect 15556 18464 15620 18468
rect 15636 18524 15700 18528
rect 15636 18468 15640 18524
rect 15640 18468 15696 18524
rect 15696 18468 15700 18524
rect 15636 18464 15700 18468
rect 29840 18524 29904 18528
rect 29840 18468 29844 18524
rect 29844 18468 29900 18524
rect 29900 18468 29904 18524
rect 29840 18464 29904 18468
rect 29920 18524 29984 18528
rect 29920 18468 29924 18524
rect 29924 18468 29980 18524
rect 29980 18468 29984 18524
rect 29920 18464 29984 18468
rect 30000 18524 30064 18528
rect 30000 18468 30004 18524
rect 30004 18468 30060 18524
rect 30060 18468 30064 18524
rect 30000 18464 30064 18468
rect 30080 18524 30144 18528
rect 30080 18468 30084 18524
rect 30084 18468 30140 18524
rect 30140 18468 30144 18524
rect 30080 18464 30144 18468
rect 44284 18524 44348 18528
rect 44284 18468 44288 18524
rect 44288 18468 44344 18524
rect 44344 18468 44348 18524
rect 44284 18464 44348 18468
rect 44364 18524 44428 18528
rect 44364 18468 44368 18524
rect 44368 18468 44424 18524
rect 44424 18468 44428 18524
rect 44364 18464 44428 18468
rect 44444 18524 44508 18528
rect 44444 18468 44448 18524
rect 44448 18468 44504 18524
rect 44504 18468 44508 18524
rect 44444 18464 44508 18468
rect 44524 18524 44588 18528
rect 44524 18468 44528 18524
rect 44528 18468 44584 18524
rect 44584 18468 44588 18524
rect 44524 18464 44588 18468
rect 58728 18524 58792 18528
rect 58728 18468 58732 18524
rect 58732 18468 58788 18524
rect 58788 18468 58792 18524
rect 58728 18464 58792 18468
rect 58808 18524 58872 18528
rect 58808 18468 58812 18524
rect 58812 18468 58868 18524
rect 58868 18468 58872 18524
rect 58808 18464 58872 18468
rect 58888 18524 58952 18528
rect 58888 18468 58892 18524
rect 58892 18468 58948 18524
rect 58948 18468 58952 18524
rect 58888 18464 58952 18468
rect 58968 18524 59032 18528
rect 58968 18468 58972 18524
rect 58972 18468 59028 18524
rect 59028 18468 59032 18524
rect 58968 18464 59032 18468
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 22618 17980 22682 17984
rect 22618 17924 22622 17980
rect 22622 17924 22678 17980
rect 22678 17924 22682 17980
rect 22618 17920 22682 17924
rect 22698 17980 22762 17984
rect 22698 17924 22702 17980
rect 22702 17924 22758 17980
rect 22758 17924 22762 17980
rect 22698 17920 22762 17924
rect 22778 17980 22842 17984
rect 22778 17924 22782 17980
rect 22782 17924 22838 17980
rect 22838 17924 22842 17980
rect 22778 17920 22842 17924
rect 22858 17980 22922 17984
rect 22858 17924 22862 17980
rect 22862 17924 22918 17980
rect 22918 17924 22922 17980
rect 22858 17920 22922 17924
rect 37062 17980 37126 17984
rect 37062 17924 37066 17980
rect 37066 17924 37122 17980
rect 37122 17924 37126 17980
rect 37062 17920 37126 17924
rect 37142 17980 37206 17984
rect 37142 17924 37146 17980
rect 37146 17924 37202 17980
rect 37202 17924 37206 17980
rect 37142 17920 37206 17924
rect 37222 17980 37286 17984
rect 37222 17924 37226 17980
rect 37226 17924 37282 17980
rect 37282 17924 37286 17980
rect 37222 17920 37286 17924
rect 37302 17980 37366 17984
rect 37302 17924 37306 17980
rect 37306 17924 37362 17980
rect 37362 17924 37366 17980
rect 37302 17920 37366 17924
rect 51506 17980 51570 17984
rect 51506 17924 51510 17980
rect 51510 17924 51566 17980
rect 51566 17924 51570 17980
rect 51506 17920 51570 17924
rect 51586 17980 51650 17984
rect 51586 17924 51590 17980
rect 51590 17924 51646 17980
rect 51646 17924 51650 17980
rect 51586 17920 51650 17924
rect 51666 17980 51730 17984
rect 51666 17924 51670 17980
rect 51670 17924 51726 17980
rect 51726 17924 51730 17980
rect 51666 17920 51730 17924
rect 51746 17980 51810 17984
rect 51746 17924 51750 17980
rect 51750 17924 51806 17980
rect 51806 17924 51810 17980
rect 51746 17920 51810 17924
rect 15396 17436 15460 17440
rect 15396 17380 15400 17436
rect 15400 17380 15456 17436
rect 15456 17380 15460 17436
rect 15396 17376 15460 17380
rect 15476 17436 15540 17440
rect 15476 17380 15480 17436
rect 15480 17380 15536 17436
rect 15536 17380 15540 17436
rect 15476 17376 15540 17380
rect 15556 17436 15620 17440
rect 15556 17380 15560 17436
rect 15560 17380 15616 17436
rect 15616 17380 15620 17436
rect 15556 17376 15620 17380
rect 15636 17436 15700 17440
rect 15636 17380 15640 17436
rect 15640 17380 15696 17436
rect 15696 17380 15700 17436
rect 15636 17376 15700 17380
rect 29840 17436 29904 17440
rect 29840 17380 29844 17436
rect 29844 17380 29900 17436
rect 29900 17380 29904 17436
rect 29840 17376 29904 17380
rect 29920 17436 29984 17440
rect 29920 17380 29924 17436
rect 29924 17380 29980 17436
rect 29980 17380 29984 17436
rect 29920 17376 29984 17380
rect 30000 17436 30064 17440
rect 30000 17380 30004 17436
rect 30004 17380 30060 17436
rect 30060 17380 30064 17436
rect 30000 17376 30064 17380
rect 30080 17436 30144 17440
rect 30080 17380 30084 17436
rect 30084 17380 30140 17436
rect 30140 17380 30144 17436
rect 30080 17376 30144 17380
rect 44284 17436 44348 17440
rect 44284 17380 44288 17436
rect 44288 17380 44344 17436
rect 44344 17380 44348 17436
rect 44284 17376 44348 17380
rect 44364 17436 44428 17440
rect 44364 17380 44368 17436
rect 44368 17380 44424 17436
rect 44424 17380 44428 17436
rect 44364 17376 44428 17380
rect 44444 17436 44508 17440
rect 44444 17380 44448 17436
rect 44448 17380 44504 17436
rect 44504 17380 44508 17436
rect 44444 17376 44508 17380
rect 44524 17436 44588 17440
rect 44524 17380 44528 17436
rect 44528 17380 44584 17436
rect 44584 17380 44588 17436
rect 44524 17376 44588 17380
rect 58728 17436 58792 17440
rect 58728 17380 58732 17436
rect 58732 17380 58788 17436
rect 58788 17380 58792 17436
rect 58728 17376 58792 17380
rect 58808 17436 58872 17440
rect 58808 17380 58812 17436
rect 58812 17380 58868 17436
rect 58868 17380 58872 17436
rect 58808 17376 58872 17380
rect 58888 17436 58952 17440
rect 58888 17380 58892 17436
rect 58892 17380 58948 17436
rect 58948 17380 58952 17436
rect 58888 17376 58952 17380
rect 58968 17436 59032 17440
rect 58968 17380 58972 17436
rect 58972 17380 59028 17436
rect 59028 17380 59032 17436
rect 58968 17376 59032 17380
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 22618 16892 22682 16896
rect 22618 16836 22622 16892
rect 22622 16836 22678 16892
rect 22678 16836 22682 16892
rect 22618 16832 22682 16836
rect 22698 16892 22762 16896
rect 22698 16836 22702 16892
rect 22702 16836 22758 16892
rect 22758 16836 22762 16892
rect 22698 16832 22762 16836
rect 22778 16892 22842 16896
rect 22778 16836 22782 16892
rect 22782 16836 22838 16892
rect 22838 16836 22842 16892
rect 22778 16832 22842 16836
rect 22858 16892 22922 16896
rect 22858 16836 22862 16892
rect 22862 16836 22918 16892
rect 22918 16836 22922 16892
rect 22858 16832 22922 16836
rect 37062 16892 37126 16896
rect 37062 16836 37066 16892
rect 37066 16836 37122 16892
rect 37122 16836 37126 16892
rect 37062 16832 37126 16836
rect 37142 16892 37206 16896
rect 37142 16836 37146 16892
rect 37146 16836 37202 16892
rect 37202 16836 37206 16892
rect 37142 16832 37206 16836
rect 37222 16892 37286 16896
rect 37222 16836 37226 16892
rect 37226 16836 37282 16892
rect 37282 16836 37286 16892
rect 37222 16832 37286 16836
rect 37302 16892 37366 16896
rect 37302 16836 37306 16892
rect 37306 16836 37362 16892
rect 37362 16836 37366 16892
rect 37302 16832 37366 16836
rect 51506 16892 51570 16896
rect 51506 16836 51510 16892
rect 51510 16836 51566 16892
rect 51566 16836 51570 16892
rect 51506 16832 51570 16836
rect 51586 16892 51650 16896
rect 51586 16836 51590 16892
rect 51590 16836 51646 16892
rect 51646 16836 51650 16892
rect 51586 16832 51650 16836
rect 51666 16892 51730 16896
rect 51666 16836 51670 16892
rect 51670 16836 51726 16892
rect 51726 16836 51730 16892
rect 51666 16832 51730 16836
rect 51746 16892 51810 16896
rect 51746 16836 51750 16892
rect 51750 16836 51806 16892
rect 51806 16836 51810 16892
rect 51746 16832 51810 16836
rect 15396 16348 15460 16352
rect 15396 16292 15400 16348
rect 15400 16292 15456 16348
rect 15456 16292 15460 16348
rect 15396 16288 15460 16292
rect 15476 16348 15540 16352
rect 15476 16292 15480 16348
rect 15480 16292 15536 16348
rect 15536 16292 15540 16348
rect 15476 16288 15540 16292
rect 15556 16348 15620 16352
rect 15556 16292 15560 16348
rect 15560 16292 15616 16348
rect 15616 16292 15620 16348
rect 15556 16288 15620 16292
rect 15636 16348 15700 16352
rect 15636 16292 15640 16348
rect 15640 16292 15696 16348
rect 15696 16292 15700 16348
rect 15636 16288 15700 16292
rect 29840 16348 29904 16352
rect 29840 16292 29844 16348
rect 29844 16292 29900 16348
rect 29900 16292 29904 16348
rect 29840 16288 29904 16292
rect 29920 16348 29984 16352
rect 29920 16292 29924 16348
rect 29924 16292 29980 16348
rect 29980 16292 29984 16348
rect 29920 16288 29984 16292
rect 30000 16348 30064 16352
rect 30000 16292 30004 16348
rect 30004 16292 30060 16348
rect 30060 16292 30064 16348
rect 30000 16288 30064 16292
rect 30080 16348 30144 16352
rect 30080 16292 30084 16348
rect 30084 16292 30140 16348
rect 30140 16292 30144 16348
rect 30080 16288 30144 16292
rect 44284 16348 44348 16352
rect 44284 16292 44288 16348
rect 44288 16292 44344 16348
rect 44344 16292 44348 16348
rect 44284 16288 44348 16292
rect 44364 16348 44428 16352
rect 44364 16292 44368 16348
rect 44368 16292 44424 16348
rect 44424 16292 44428 16348
rect 44364 16288 44428 16292
rect 44444 16348 44508 16352
rect 44444 16292 44448 16348
rect 44448 16292 44504 16348
rect 44504 16292 44508 16348
rect 44444 16288 44508 16292
rect 44524 16348 44588 16352
rect 44524 16292 44528 16348
rect 44528 16292 44584 16348
rect 44584 16292 44588 16348
rect 44524 16288 44588 16292
rect 58728 16348 58792 16352
rect 58728 16292 58732 16348
rect 58732 16292 58788 16348
rect 58788 16292 58792 16348
rect 58728 16288 58792 16292
rect 58808 16348 58872 16352
rect 58808 16292 58812 16348
rect 58812 16292 58868 16348
rect 58868 16292 58872 16348
rect 58808 16288 58872 16292
rect 58888 16348 58952 16352
rect 58888 16292 58892 16348
rect 58892 16292 58948 16348
rect 58948 16292 58952 16348
rect 58888 16288 58952 16292
rect 58968 16348 59032 16352
rect 58968 16292 58972 16348
rect 58972 16292 59028 16348
rect 59028 16292 59032 16348
rect 58968 16288 59032 16292
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 22618 15804 22682 15808
rect 22618 15748 22622 15804
rect 22622 15748 22678 15804
rect 22678 15748 22682 15804
rect 22618 15744 22682 15748
rect 22698 15804 22762 15808
rect 22698 15748 22702 15804
rect 22702 15748 22758 15804
rect 22758 15748 22762 15804
rect 22698 15744 22762 15748
rect 22778 15804 22842 15808
rect 22778 15748 22782 15804
rect 22782 15748 22838 15804
rect 22838 15748 22842 15804
rect 22778 15744 22842 15748
rect 22858 15804 22922 15808
rect 22858 15748 22862 15804
rect 22862 15748 22918 15804
rect 22918 15748 22922 15804
rect 22858 15744 22922 15748
rect 37062 15804 37126 15808
rect 37062 15748 37066 15804
rect 37066 15748 37122 15804
rect 37122 15748 37126 15804
rect 37062 15744 37126 15748
rect 37142 15804 37206 15808
rect 37142 15748 37146 15804
rect 37146 15748 37202 15804
rect 37202 15748 37206 15804
rect 37142 15744 37206 15748
rect 37222 15804 37286 15808
rect 37222 15748 37226 15804
rect 37226 15748 37282 15804
rect 37282 15748 37286 15804
rect 37222 15744 37286 15748
rect 37302 15804 37366 15808
rect 37302 15748 37306 15804
rect 37306 15748 37362 15804
rect 37362 15748 37366 15804
rect 37302 15744 37366 15748
rect 51506 15804 51570 15808
rect 51506 15748 51510 15804
rect 51510 15748 51566 15804
rect 51566 15748 51570 15804
rect 51506 15744 51570 15748
rect 51586 15804 51650 15808
rect 51586 15748 51590 15804
rect 51590 15748 51646 15804
rect 51646 15748 51650 15804
rect 51586 15744 51650 15748
rect 51666 15804 51730 15808
rect 51666 15748 51670 15804
rect 51670 15748 51726 15804
rect 51726 15748 51730 15804
rect 51666 15744 51730 15748
rect 51746 15804 51810 15808
rect 51746 15748 51750 15804
rect 51750 15748 51806 15804
rect 51806 15748 51810 15804
rect 51746 15744 51810 15748
rect 15396 15260 15460 15264
rect 15396 15204 15400 15260
rect 15400 15204 15456 15260
rect 15456 15204 15460 15260
rect 15396 15200 15460 15204
rect 15476 15260 15540 15264
rect 15476 15204 15480 15260
rect 15480 15204 15536 15260
rect 15536 15204 15540 15260
rect 15476 15200 15540 15204
rect 15556 15260 15620 15264
rect 15556 15204 15560 15260
rect 15560 15204 15616 15260
rect 15616 15204 15620 15260
rect 15556 15200 15620 15204
rect 15636 15260 15700 15264
rect 15636 15204 15640 15260
rect 15640 15204 15696 15260
rect 15696 15204 15700 15260
rect 15636 15200 15700 15204
rect 29840 15260 29904 15264
rect 29840 15204 29844 15260
rect 29844 15204 29900 15260
rect 29900 15204 29904 15260
rect 29840 15200 29904 15204
rect 29920 15260 29984 15264
rect 29920 15204 29924 15260
rect 29924 15204 29980 15260
rect 29980 15204 29984 15260
rect 29920 15200 29984 15204
rect 30000 15260 30064 15264
rect 30000 15204 30004 15260
rect 30004 15204 30060 15260
rect 30060 15204 30064 15260
rect 30000 15200 30064 15204
rect 30080 15260 30144 15264
rect 30080 15204 30084 15260
rect 30084 15204 30140 15260
rect 30140 15204 30144 15260
rect 30080 15200 30144 15204
rect 44284 15260 44348 15264
rect 44284 15204 44288 15260
rect 44288 15204 44344 15260
rect 44344 15204 44348 15260
rect 44284 15200 44348 15204
rect 44364 15260 44428 15264
rect 44364 15204 44368 15260
rect 44368 15204 44424 15260
rect 44424 15204 44428 15260
rect 44364 15200 44428 15204
rect 44444 15260 44508 15264
rect 44444 15204 44448 15260
rect 44448 15204 44504 15260
rect 44504 15204 44508 15260
rect 44444 15200 44508 15204
rect 44524 15260 44588 15264
rect 44524 15204 44528 15260
rect 44528 15204 44584 15260
rect 44584 15204 44588 15260
rect 44524 15200 44588 15204
rect 58728 15260 58792 15264
rect 58728 15204 58732 15260
rect 58732 15204 58788 15260
rect 58788 15204 58792 15260
rect 58728 15200 58792 15204
rect 58808 15260 58872 15264
rect 58808 15204 58812 15260
rect 58812 15204 58868 15260
rect 58868 15204 58872 15260
rect 58808 15200 58872 15204
rect 58888 15260 58952 15264
rect 58888 15204 58892 15260
rect 58892 15204 58948 15260
rect 58948 15204 58952 15260
rect 58888 15200 58952 15204
rect 58968 15260 59032 15264
rect 58968 15204 58972 15260
rect 58972 15204 59028 15260
rect 59028 15204 59032 15260
rect 58968 15200 59032 15204
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 22618 14716 22682 14720
rect 22618 14660 22622 14716
rect 22622 14660 22678 14716
rect 22678 14660 22682 14716
rect 22618 14656 22682 14660
rect 22698 14716 22762 14720
rect 22698 14660 22702 14716
rect 22702 14660 22758 14716
rect 22758 14660 22762 14716
rect 22698 14656 22762 14660
rect 22778 14716 22842 14720
rect 22778 14660 22782 14716
rect 22782 14660 22838 14716
rect 22838 14660 22842 14716
rect 22778 14656 22842 14660
rect 22858 14716 22922 14720
rect 22858 14660 22862 14716
rect 22862 14660 22918 14716
rect 22918 14660 22922 14716
rect 22858 14656 22922 14660
rect 37062 14716 37126 14720
rect 37062 14660 37066 14716
rect 37066 14660 37122 14716
rect 37122 14660 37126 14716
rect 37062 14656 37126 14660
rect 37142 14716 37206 14720
rect 37142 14660 37146 14716
rect 37146 14660 37202 14716
rect 37202 14660 37206 14716
rect 37142 14656 37206 14660
rect 37222 14716 37286 14720
rect 37222 14660 37226 14716
rect 37226 14660 37282 14716
rect 37282 14660 37286 14716
rect 37222 14656 37286 14660
rect 37302 14716 37366 14720
rect 37302 14660 37306 14716
rect 37306 14660 37362 14716
rect 37362 14660 37366 14716
rect 37302 14656 37366 14660
rect 51506 14716 51570 14720
rect 51506 14660 51510 14716
rect 51510 14660 51566 14716
rect 51566 14660 51570 14716
rect 51506 14656 51570 14660
rect 51586 14716 51650 14720
rect 51586 14660 51590 14716
rect 51590 14660 51646 14716
rect 51646 14660 51650 14716
rect 51586 14656 51650 14660
rect 51666 14716 51730 14720
rect 51666 14660 51670 14716
rect 51670 14660 51726 14716
rect 51726 14660 51730 14716
rect 51666 14656 51730 14660
rect 51746 14716 51810 14720
rect 51746 14660 51750 14716
rect 51750 14660 51806 14716
rect 51806 14660 51810 14716
rect 51746 14656 51810 14660
rect 15396 14172 15460 14176
rect 15396 14116 15400 14172
rect 15400 14116 15456 14172
rect 15456 14116 15460 14172
rect 15396 14112 15460 14116
rect 15476 14172 15540 14176
rect 15476 14116 15480 14172
rect 15480 14116 15536 14172
rect 15536 14116 15540 14172
rect 15476 14112 15540 14116
rect 15556 14172 15620 14176
rect 15556 14116 15560 14172
rect 15560 14116 15616 14172
rect 15616 14116 15620 14172
rect 15556 14112 15620 14116
rect 15636 14172 15700 14176
rect 15636 14116 15640 14172
rect 15640 14116 15696 14172
rect 15696 14116 15700 14172
rect 15636 14112 15700 14116
rect 29840 14172 29904 14176
rect 29840 14116 29844 14172
rect 29844 14116 29900 14172
rect 29900 14116 29904 14172
rect 29840 14112 29904 14116
rect 29920 14172 29984 14176
rect 29920 14116 29924 14172
rect 29924 14116 29980 14172
rect 29980 14116 29984 14172
rect 29920 14112 29984 14116
rect 30000 14172 30064 14176
rect 30000 14116 30004 14172
rect 30004 14116 30060 14172
rect 30060 14116 30064 14172
rect 30000 14112 30064 14116
rect 30080 14172 30144 14176
rect 30080 14116 30084 14172
rect 30084 14116 30140 14172
rect 30140 14116 30144 14172
rect 30080 14112 30144 14116
rect 44284 14172 44348 14176
rect 44284 14116 44288 14172
rect 44288 14116 44344 14172
rect 44344 14116 44348 14172
rect 44284 14112 44348 14116
rect 44364 14172 44428 14176
rect 44364 14116 44368 14172
rect 44368 14116 44424 14172
rect 44424 14116 44428 14172
rect 44364 14112 44428 14116
rect 44444 14172 44508 14176
rect 44444 14116 44448 14172
rect 44448 14116 44504 14172
rect 44504 14116 44508 14172
rect 44444 14112 44508 14116
rect 44524 14172 44588 14176
rect 44524 14116 44528 14172
rect 44528 14116 44584 14172
rect 44584 14116 44588 14172
rect 44524 14112 44588 14116
rect 58728 14172 58792 14176
rect 58728 14116 58732 14172
rect 58732 14116 58788 14172
rect 58788 14116 58792 14172
rect 58728 14112 58792 14116
rect 58808 14172 58872 14176
rect 58808 14116 58812 14172
rect 58812 14116 58868 14172
rect 58868 14116 58872 14172
rect 58808 14112 58872 14116
rect 58888 14172 58952 14176
rect 58888 14116 58892 14172
rect 58892 14116 58948 14172
rect 58948 14116 58952 14172
rect 58888 14112 58952 14116
rect 58968 14172 59032 14176
rect 58968 14116 58972 14172
rect 58972 14116 59028 14172
rect 59028 14116 59032 14172
rect 58968 14112 59032 14116
rect 42380 13832 42444 13836
rect 42380 13776 42394 13832
rect 42394 13776 42444 13832
rect 42380 13772 42444 13776
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 22618 13628 22682 13632
rect 22618 13572 22622 13628
rect 22622 13572 22678 13628
rect 22678 13572 22682 13628
rect 22618 13568 22682 13572
rect 22698 13628 22762 13632
rect 22698 13572 22702 13628
rect 22702 13572 22758 13628
rect 22758 13572 22762 13628
rect 22698 13568 22762 13572
rect 22778 13628 22842 13632
rect 22778 13572 22782 13628
rect 22782 13572 22838 13628
rect 22838 13572 22842 13628
rect 22778 13568 22842 13572
rect 22858 13628 22922 13632
rect 22858 13572 22862 13628
rect 22862 13572 22918 13628
rect 22918 13572 22922 13628
rect 22858 13568 22922 13572
rect 37062 13628 37126 13632
rect 37062 13572 37066 13628
rect 37066 13572 37122 13628
rect 37122 13572 37126 13628
rect 37062 13568 37126 13572
rect 37142 13628 37206 13632
rect 37142 13572 37146 13628
rect 37146 13572 37202 13628
rect 37202 13572 37206 13628
rect 37142 13568 37206 13572
rect 37222 13628 37286 13632
rect 37222 13572 37226 13628
rect 37226 13572 37282 13628
rect 37282 13572 37286 13628
rect 37222 13568 37286 13572
rect 37302 13628 37366 13632
rect 37302 13572 37306 13628
rect 37306 13572 37362 13628
rect 37362 13572 37366 13628
rect 37302 13568 37366 13572
rect 51506 13628 51570 13632
rect 51506 13572 51510 13628
rect 51510 13572 51566 13628
rect 51566 13572 51570 13628
rect 51506 13568 51570 13572
rect 51586 13628 51650 13632
rect 51586 13572 51590 13628
rect 51590 13572 51646 13628
rect 51646 13572 51650 13628
rect 51586 13568 51650 13572
rect 51666 13628 51730 13632
rect 51666 13572 51670 13628
rect 51670 13572 51726 13628
rect 51726 13572 51730 13628
rect 51666 13568 51730 13572
rect 51746 13628 51810 13632
rect 51746 13572 51750 13628
rect 51750 13572 51806 13628
rect 51806 13572 51810 13628
rect 51746 13568 51810 13572
rect 15396 13084 15460 13088
rect 15396 13028 15400 13084
rect 15400 13028 15456 13084
rect 15456 13028 15460 13084
rect 15396 13024 15460 13028
rect 15476 13084 15540 13088
rect 15476 13028 15480 13084
rect 15480 13028 15536 13084
rect 15536 13028 15540 13084
rect 15476 13024 15540 13028
rect 15556 13084 15620 13088
rect 15556 13028 15560 13084
rect 15560 13028 15616 13084
rect 15616 13028 15620 13084
rect 15556 13024 15620 13028
rect 15636 13084 15700 13088
rect 15636 13028 15640 13084
rect 15640 13028 15696 13084
rect 15696 13028 15700 13084
rect 15636 13024 15700 13028
rect 29840 13084 29904 13088
rect 29840 13028 29844 13084
rect 29844 13028 29900 13084
rect 29900 13028 29904 13084
rect 29840 13024 29904 13028
rect 29920 13084 29984 13088
rect 29920 13028 29924 13084
rect 29924 13028 29980 13084
rect 29980 13028 29984 13084
rect 29920 13024 29984 13028
rect 30000 13084 30064 13088
rect 30000 13028 30004 13084
rect 30004 13028 30060 13084
rect 30060 13028 30064 13084
rect 30000 13024 30064 13028
rect 30080 13084 30144 13088
rect 30080 13028 30084 13084
rect 30084 13028 30140 13084
rect 30140 13028 30144 13084
rect 30080 13024 30144 13028
rect 44284 13084 44348 13088
rect 44284 13028 44288 13084
rect 44288 13028 44344 13084
rect 44344 13028 44348 13084
rect 44284 13024 44348 13028
rect 44364 13084 44428 13088
rect 44364 13028 44368 13084
rect 44368 13028 44424 13084
rect 44424 13028 44428 13084
rect 44364 13024 44428 13028
rect 44444 13084 44508 13088
rect 44444 13028 44448 13084
rect 44448 13028 44504 13084
rect 44504 13028 44508 13084
rect 44444 13024 44508 13028
rect 44524 13084 44588 13088
rect 44524 13028 44528 13084
rect 44528 13028 44584 13084
rect 44584 13028 44588 13084
rect 44524 13024 44588 13028
rect 58728 13084 58792 13088
rect 58728 13028 58732 13084
rect 58732 13028 58788 13084
rect 58788 13028 58792 13084
rect 58728 13024 58792 13028
rect 58808 13084 58872 13088
rect 58808 13028 58812 13084
rect 58812 13028 58868 13084
rect 58868 13028 58872 13084
rect 58808 13024 58872 13028
rect 58888 13084 58952 13088
rect 58888 13028 58892 13084
rect 58892 13028 58948 13084
rect 58948 13028 58952 13084
rect 58888 13024 58952 13028
rect 58968 13084 59032 13088
rect 58968 13028 58972 13084
rect 58972 13028 59028 13084
rect 59028 13028 59032 13084
rect 58968 13024 59032 13028
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 22618 12540 22682 12544
rect 22618 12484 22622 12540
rect 22622 12484 22678 12540
rect 22678 12484 22682 12540
rect 22618 12480 22682 12484
rect 22698 12540 22762 12544
rect 22698 12484 22702 12540
rect 22702 12484 22758 12540
rect 22758 12484 22762 12540
rect 22698 12480 22762 12484
rect 22778 12540 22842 12544
rect 22778 12484 22782 12540
rect 22782 12484 22838 12540
rect 22838 12484 22842 12540
rect 22778 12480 22842 12484
rect 22858 12540 22922 12544
rect 22858 12484 22862 12540
rect 22862 12484 22918 12540
rect 22918 12484 22922 12540
rect 22858 12480 22922 12484
rect 37062 12540 37126 12544
rect 37062 12484 37066 12540
rect 37066 12484 37122 12540
rect 37122 12484 37126 12540
rect 37062 12480 37126 12484
rect 37142 12540 37206 12544
rect 37142 12484 37146 12540
rect 37146 12484 37202 12540
rect 37202 12484 37206 12540
rect 37142 12480 37206 12484
rect 37222 12540 37286 12544
rect 37222 12484 37226 12540
rect 37226 12484 37282 12540
rect 37282 12484 37286 12540
rect 37222 12480 37286 12484
rect 37302 12540 37366 12544
rect 37302 12484 37306 12540
rect 37306 12484 37362 12540
rect 37362 12484 37366 12540
rect 37302 12480 37366 12484
rect 51506 12540 51570 12544
rect 51506 12484 51510 12540
rect 51510 12484 51566 12540
rect 51566 12484 51570 12540
rect 51506 12480 51570 12484
rect 51586 12540 51650 12544
rect 51586 12484 51590 12540
rect 51590 12484 51646 12540
rect 51646 12484 51650 12540
rect 51586 12480 51650 12484
rect 51666 12540 51730 12544
rect 51666 12484 51670 12540
rect 51670 12484 51726 12540
rect 51726 12484 51730 12540
rect 51666 12480 51730 12484
rect 51746 12540 51810 12544
rect 51746 12484 51750 12540
rect 51750 12484 51806 12540
rect 51806 12484 51810 12540
rect 51746 12480 51810 12484
rect 15396 11996 15460 12000
rect 15396 11940 15400 11996
rect 15400 11940 15456 11996
rect 15456 11940 15460 11996
rect 15396 11936 15460 11940
rect 15476 11996 15540 12000
rect 15476 11940 15480 11996
rect 15480 11940 15536 11996
rect 15536 11940 15540 11996
rect 15476 11936 15540 11940
rect 15556 11996 15620 12000
rect 15556 11940 15560 11996
rect 15560 11940 15616 11996
rect 15616 11940 15620 11996
rect 15556 11936 15620 11940
rect 15636 11996 15700 12000
rect 15636 11940 15640 11996
rect 15640 11940 15696 11996
rect 15696 11940 15700 11996
rect 15636 11936 15700 11940
rect 29840 11996 29904 12000
rect 29840 11940 29844 11996
rect 29844 11940 29900 11996
rect 29900 11940 29904 11996
rect 29840 11936 29904 11940
rect 29920 11996 29984 12000
rect 29920 11940 29924 11996
rect 29924 11940 29980 11996
rect 29980 11940 29984 11996
rect 29920 11936 29984 11940
rect 30000 11996 30064 12000
rect 30000 11940 30004 11996
rect 30004 11940 30060 11996
rect 30060 11940 30064 11996
rect 30000 11936 30064 11940
rect 30080 11996 30144 12000
rect 30080 11940 30084 11996
rect 30084 11940 30140 11996
rect 30140 11940 30144 11996
rect 30080 11936 30144 11940
rect 44284 11996 44348 12000
rect 44284 11940 44288 11996
rect 44288 11940 44344 11996
rect 44344 11940 44348 11996
rect 44284 11936 44348 11940
rect 44364 11996 44428 12000
rect 44364 11940 44368 11996
rect 44368 11940 44424 11996
rect 44424 11940 44428 11996
rect 44364 11936 44428 11940
rect 44444 11996 44508 12000
rect 44444 11940 44448 11996
rect 44448 11940 44504 11996
rect 44504 11940 44508 11996
rect 44444 11936 44508 11940
rect 44524 11996 44588 12000
rect 44524 11940 44528 11996
rect 44528 11940 44584 11996
rect 44584 11940 44588 11996
rect 44524 11936 44588 11940
rect 58728 11996 58792 12000
rect 58728 11940 58732 11996
rect 58732 11940 58788 11996
rect 58788 11940 58792 11996
rect 58728 11936 58792 11940
rect 58808 11996 58872 12000
rect 58808 11940 58812 11996
rect 58812 11940 58868 11996
rect 58868 11940 58872 11996
rect 58808 11936 58872 11940
rect 58888 11996 58952 12000
rect 58888 11940 58892 11996
rect 58892 11940 58948 11996
rect 58948 11940 58952 11996
rect 58888 11936 58952 11940
rect 58968 11996 59032 12000
rect 58968 11940 58972 11996
rect 58972 11940 59028 11996
rect 59028 11940 59032 11996
rect 58968 11936 59032 11940
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 22618 11452 22682 11456
rect 22618 11396 22622 11452
rect 22622 11396 22678 11452
rect 22678 11396 22682 11452
rect 22618 11392 22682 11396
rect 22698 11452 22762 11456
rect 22698 11396 22702 11452
rect 22702 11396 22758 11452
rect 22758 11396 22762 11452
rect 22698 11392 22762 11396
rect 22778 11452 22842 11456
rect 22778 11396 22782 11452
rect 22782 11396 22838 11452
rect 22838 11396 22842 11452
rect 22778 11392 22842 11396
rect 22858 11452 22922 11456
rect 22858 11396 22862 11452
rect 22862 11396 22918 11452
rect 22918 11396 22922 11452
rect 22858 11392 22922 11396
rect 37062 11452 37126 11456
rect 37062 11396 37066 11452
rect 37066 11396 37122 11452
rect 37122 11396 37126 11452
rect 37062 11392 37126 11396
rect 37142 11452 37206 11456
rect 37142 11396 37146 11452
rect 37146 11396 37202 11452
rect 37202 11396 37206 11452
rect 37142 11392 37206 11396
rect 37222 11452 37286 11456
rect 37222 11396 37226 11452
rect 37226 11396 37282 11452
rect 37282 11396 37286 11452
rect 37222 11392 37286 11396
rect 37302 11452 37366 11456
rect 37302 11396 37306 11452
rect 37306 11396 37362 11452
rect 37362 11396 37366 11452
rect 37302 11392 37366 11396
rect 51506 11452 51570 11456
rect 51506 11396 51510 11452
rect 51510 11396 51566 11452
rect 51566 11396 51570 11452
rect 51506 11392 51570 11396
rect 51586 11452 51650 11456
rect 51586 11396 51590 11452
rect 51590 11396 51646 11452
rect 51646 11396 51650 11452
rect 51586 11392 51650 11396
rect 51666 11452 51730 11456
rect 51666 11396 51670 11452
rect 51670 11396 51726 11452
rect 51726 11396 51730 11452
rect 51666 11392 51730 11396
rect 51746 11452 51810 11456
rect 51746 11396 51750 11452
rect 51750 11396 51806 11452
rect 51806 11396 51810 11452
rect 51746 11392 51810 11396
rect 15396 10908 15460 10912
rect 15396 10852 15400 10908
rect 15400 10852 15456 10908
rect 15456 10852 15460 10908
rect 15396 10848 15460 10852
rect 15476 10908 15540 10912
rect 15476 10852 15480 10908
rect 15480 10852 15536 10908
rect 15536 10852 15540 10908
rect 15476 10848 15540 10852
rect 15556 10908 15620 10912
rect 15556 10852 15560 10908
rect 15560 10852 15616 10908
rect 15616 10852 15620 10908
rect 15556 10848 15620 10852
rect 15636 10908 15700 10912
rect 15636 10852 15640 10908
rect 15640 10852 15696 10908
rect 15696 10852 15700 10908
rect 15636 10848 15700 10852
rect 29840 10908 29904 10912
rect 29840 10852 29844 10908
rect 29844 10852 29900 10908
rect 29900 10852 29904 10908
rect 29840 10848 29904 10852
rect 29920 10908 29984 10912
rect 29920 10852 29924 10908
rect 29924 10852 29980 10908
rect 29980 10852 29984 10908
rect 29920 10848 29984 10852
rect 30000 10908 30064 10912
rect 30000 10852 30004 10908
rect 30004 10852 30060 10908
rect 30060 10852 30064 10908
rect 30000 10848 30064 10852
rect 30080 10908 30144 10912
rect 30080 10852 30084 10908
rect 30084 10852 30140 10908
rect 30140 10852 30144 10908
rect 30080 10848 30144 10852
rect 44284 10908 44348 10912
rect 44284 10852 44288 10908
rect 44288 10852 44344 10908
rect 44344 10852 44348 10908
rect 44284 10848 44348 10852
rect 44364 10908 44428 10912
rect 44364 10852 44368 10908
rect 44368 10852 44424 10908
rect 44424 10852 44428 10908
rect 44364 10848 44428 10852
rect 44444 10908 44508 10912
rect 44444 10852 44448 10908
rect 44448 10852 44504 10908
rect 44504 10852 44508 10908
rect 44444 10848 44508 10852
rect 44524 10908 44588 10912
rect 44524 10852 44528 10908
rect 44528 10852 44584 10908
rect 44584 10852 44588 10908
rect 44524 10848 44588 10852
rect 58728 10908 58792 10912
rect 58728 10852 58732 10908
rect 58732 10852 58788 10908
rect 58788 10852 58792 10908
rect 58728 10848 58792 10852
rect 58808 10908 58872 10912
rect 58808 10852 58812 10908
rect 58812 10852 58868 10908
rect 58868 10852 58872 10908
rect 58808 10848 58872 10852
rect 58888 10908 58952 10912
rect 58888 10852 58892 10908
rect 58892 10852 58948 10908
rect 58948 10852 58952 10908
rect 58888 10848 58952 10852
rect 58968 10908 59032 10912
rect 58968 10852 58972 10908
rect 58972 10852 59028 10908
rect 59028 10852 59032 10908
rect 58968 10848 59032 10852
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 22618 10364 22682 10368
rect 22618 10308 22622 10364
rect 22622 10308 22678 10364
rect 22678 10308 22682 10364
rect 22618 10304 22682 10308
rect 22698 10364 22762 10368
rect 22698 10308 22702 10364
rect 22702 10308 22758 10364
rect 22758 10308 22762 10364
rect 22698 10304 22762 10308
rect 22778 10364 22842 10368
rect 22778 10308 22782 10364
rect 22782 10308 22838 10364
rect 22838 10308 22842 10364
rect 22778 10304 22842 10308
rect 22858 10364 22922 10368
rect 22858 10308 22862 10364
rect 22862 10308 22918 10364
rect 22918 10308 22922 10364
rect 22858 10304 22922 10308
rect 37062 10364 37126 10368
rect 37062 10308 37066 10364
rect 37066 10308 37122 10364
rect 37122 10308 37126 10364
rect 37062 10304 37126 10308
rect 37142 10364 37206 10368
rect 37142 10308 37146 10364
rect 37146 10308 37202 10364
rect 37202 10308 37206 10364
rect 37142 10304 37206 10308
rect 37222 10364 37286 10368
rect 37222 10308 37226 10364
rect 37226 10308 37282 10364
rect 37282 10308 37286 10364
rect 37222 10304 37286 10308
rect 37302 10364 37366 10368
rect 37302 10308 37306 10364
rect 37306 10308 37362 10364
rect 37362 10308 37366 10364
rect 37302 10304 37366 10308
rect 51506 10364 51570 10368
rect 51506 10308 51510 10364
rect 51510 10308 51566 10364
rect 51566 10308 51570 10364
rect 51506 10304 51570 10308
rect 51586 10364 51650 10368
rect 51586 10308 51590 10364
rect 51590 10308 51646 10364
rect 51646 10308 51650 10364
rect 51586 10304 51650 10308
rect 51666 10364 51730 10368
rect 51666 10308 51670 10364
rect 51670 10308 51726 10364
rect 51726 10308 51730 10364
rect 51666 10304 51730 10308
rect 51746 10364 51810 10368
rect 51746 10308 51750 10364
rect 51750 10308 51806 10364
rect 51806 10308 51810 10364
rect 51746 10304 51810 10308
rect 15396 9820 15460 9824
rect 15396 9764 15400 9820
rect 15400 9764 15456 9820
rect 15456 9764 15460 9820
rect 15396 9760 15460 9764
rect 15476 9820 15540 9824
rect 15476 9764 15480 9820
rect 15480 9764 15536 9820
rect 15536 9764 15540 9820
rect 15476 9760 15540 9764
rect 15556 9820 15620 9824
rect 15556 9764 15560 9820
rect 15560 9764 15616 9820
rect 15616 9764 15620 9820
rect 15556 9760 15620 9764
rect 15636 9820 15700 9824
rect 15636 9764 15640 9820
rect 15640 9764 15696 9820
rect 15696 9764 15700 9820
rect 15636 9760 15700 9764
rect 29840 9820 29904 9824
rect 29840 9764 29844 9820
rect 29844 9764 29900 9820
rect 29900 9764 29904 9820
rect 29840 9760 29904 9764
rect 29920 9820 29984 9824
rect 29920 9764 29924 9820
rect 29924 9764 29980 9820
rect 29980 9764 29984 9820
rect 29920 9760 29984 9764
rect 30000 9820 30064 9824
rect 30000 9764 30004 9820
rect 30004 9764 30060 9820
rect 30060 9764 30064 9820
rect 30000 9760 30064 9764
rect 30080 9820 30144 9824
rect 30080 9764 30084 9820
rect 30084 9764 30140 9820
rect 30140 9764 30144 9820
rect 30080 9760 30144 9764
rect 44284 9820 44348 9824
rect 44284 9764 44288 9820
rect 44288 9764 44344 9820
rect 44344 9764 44348 9820
rect 44284 9760 44348 9764
rect 44364 9820 44428 9824
rect 44364 9764 44368 9820
rect 44368 9764 44424 9820
rect 44424 9764 44428 9820
rect 44364 9760 44428 9764
rect 44444 9820 44508 9824
rect 44444 9764 44448 9820
rect 44448 9764 44504 9820
rect 44504 9764 44508 9820
rect 44444 9760 44508 9764
rect 44524 9820 44588 9824
rect 44524 9764 44528 9820
rect 44528 9764 44584 9820
rect 44584 9764 44588 9820
rect 44524 9760 44588 9764
rect 58728 9820 58792 9824
rect 58728 9764 58732 9820
rect 58732 9764 58788 9820
rect 58788 9764 58792 9820
rect 58728 9760 58792 9764
rect 58808 9820 58872 9824
rect 58808 9764 58812 9820
rect 58812 9764 58868 9820
rect 58868 9764 58872 9820
rect 58808 9760 58872 9764
rect 58888 9820 58952 9824
rect 58888 9764 58892 9820
rect 58892 9764 58948 9820
rect 58948 9764 58952 9820
rect 58888 9760 58952 9764
rect 58968 9820 59032 9824
rect 58968 9764 58972 9820
rect 58972 9764 59028 9820
rect 59028 9764 59032 9820
rect 58968 9760 59032 9764
rect 35940 9692 36004 9756
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 22618 9276 22682 9280
rect 22618 9220 22622 9276
rect 22622 9220 22678 9276
rect 22678 9220 22682 9276
rect 22618 9216 22682 9220
rect 22698 9276 22762 9280
rect 22698 9220 22702 9276
rect 22702 9220 22758 9276
rect 22758 9220 22762 9276
rect 22698 9216 22762 9220
rect 22778 9276 22842 9280
rect 22778 9220 22782 9276
rect 22782 9220 22838 9276
rect 22838 9220 22842 9276
rect 22778 9216 22842 9220
rect 22858 9276 22922 9280
rect 22858 9220 22862 9276
rect 22862 9220 22918 9276
rect 22918 9220 22922 9276
rect 22858 9216 22922 9220
rect 37062 9276 37126 9280
rect 37062 9220 37066 9276
rect 37066 9220 37122 9276
rect 37122 9220 37126 9276
rect 37062 9216 37126 9220
rect 37142 9276 37206 9280
rect 37142 9220 37146 9276
rect 37146 9220 37202 9276
rect 37202 9220 37206 9276
rect 37142 9216 37206 9220
rect 37222 9276 37286 9280
rect 37222 9220 37226 9276
rect 37226 9220 37282 9276
rect 37282 9220 37286 9276
rect 37222 9216 37286 9220
rect 37302 9276 37366 9280
rect 37302 9220 37306 9276
rect 37306 9220 37362 9276
rect 37362 9220 37366 9276
rect 37302 9216 37366 9220
rect 51506 9276 51570 9280
rect 51506 9220 51510 9276
rect 51510 9220 51566 9276
rect 51566 9220 51570 9276
rect 51506 9216 51570 9220
rect 51586 9276 51650 9280
rect 51586 9220 51590 9276
rect 51590 9220 51646 9276
rect 51646 9220 51650 9276
rect 51586 9216 51650 9220
rect 51666 9276 51730 9280
rect 51666 9220 51670 9276
rect 51670 9220 51726 9276
rect 51726 9220 51730 9276
rect 51666 9216 51730 9220
rect 51746 9276 51810 9280
rect 51746 9220 51750 9276
rect 51750 9220 51806 9276
rect 51806 9220 51810 9276
rect 51746 9216 51810 9220
rect 15396 8732 15460 8736
rect 15396 8676 15400 8732
rect 15400 8676 15456 8732
rect 15456 8676 15460 8732
rect 15396 8672 15460 8676
rect 15476 8732 15540 8736
rect 15476 8676 15480 8732
rect 15480 8676 15536 8732
rect 15536 8676 15540 8732
rect 15476 8672 15540 8676
rect 15556 8732 15620 8736
rect 15556 8676 15560 8732
rect 15560 8676 15616 8732
rect 15616 8676 15620 8732
rect 15556 8672 15620 8676
rect 15636 8732 15700 8736
rect 15636 8676 15640 8732
rect 15640 8676 15696 8732
rect 15696 8676 15700 8732
rect 15636 8672 15700 8676
rect 29840 8732 29904 8736
rect 29840 8676 29844 8732
rect 29844 8676 29900 8732
rect 29900 8676 29904 8732
rect 29840 8672 29904 8676
rect 29920 8732 29984 8736
rect 29920 8676 29924 8732
rect 29924 8676 29980 8732
rect 29980 8676 29984 8732
rect 29920 8672 29984 8676
rect 30000 8732 30064 8736
rect 30000 8676 30004 8732
rect 30004 8676 30060 8732
rect 30060 8676 30064 8732
rect 30000 8672 30064 8676
rect 30080 8732 30144 8736
rect 30080 8676 30084 8732
rect 30084 8676 30140 8732
rect 30140 8676 30144 8732
rect 30080 8672 30144 8676
rect 44284 8732 44348 8736
rect 44284 8676 44288 8732
rect 44288 8676 44344 8732
rect 44344 8676 44348 8732
rect 44284 8672 44348 8676
rect 44364 8732 44428 8736
rect 44364 8676 44368 8732
rect 44368 8676 44424 8732
rect 44424 8676 44428 8732
rect 44364 8672 44428 8676
rect 44444 8732 44508 8736
rect 44444 8676 44448 8732
rect 44448 8676 44504 8732
rect 44504 8676 44508 8732
rect 44444 8672 44508 8676
rect 44524 8732 44588 8736
rect 44524 8676 44528 8732
rect 44528 8676 44584 8732
rect 44584 8676 44588 8732
rect 44524 8672 44588 8676
rect 58728 8732 58792 8736
rect 58728 8676 58732 8732
rect 58732 8676 58788 8732
rect 58788 8676 58792 8732
rect 58728 8672 58792 8676
rect 58808 8732 58872 8736
rect 58808 8676 58812 8732
rect 58812 8676 58868 8732
rect 58868 8676 58872 8732
rect 58808 8672 58872 8676
rect 58888 8732 58952 8736
rect 58888 8676 58892 8732
rect 58892 8676 58948 8732
rect 58948 8676 58952 8732
rect 58888 8672 58952 8676
rect 58968 8732 59032 8736
rect 58968 8676 58972 8732
rect 58972 8676 59028 8732
rect 59028 8676 59032 8732
rect 58968 8672 59032 8676
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 22618 8188 22682 8192
rect 22618 8132 22622 8188
rect 22622 8132 22678 8188
rect 22678 8132 22682 8188
rect 22618 8128 22682 8132
rect 22698 8188 22762 8192
rect 22698 8132 22702 8188
rect 22702 8132 22758 8188
rect 22758 8132 22762 8188
rect 22698 8128 22762 8132
rect 22778 8188 22842 8192
rect 22778 8132 22782 8188
rect 22782 8132 22838 8188
rect 22838 8132 22842 8188
rect 22778 8128 22842 8132
rect 22858 8188 22922 8192
rect 22858 8132 22862 8188
rect 22862 8132 22918 8188
rect 22918 8132 22922 8188
rect 22858 8128 22922 8132
rect 37062 8188 37126 8192
rect 37062 8132 37066 8188
rect 37066 8132 37122 8188
rect 37122 8132 37126 8188
rect 37062 8128 37126 8132
rect 37142 8188 37206 8192
rect 37142 8132 37146 8188
rect 37146 8132 37202 8188
rect 37202 8132 37206 8188
rect 37142 8128 37206 8132
rect 37222 8188 37286 8192
rect 37222 8132 37226 8188
rect 37226 8132 37282 8188
rect 37282 8132 37286 8188
rect 37222 8128 37286 8132
rect 37302 8188 37366 8192
rect 37302 8132 37306 8188
rect 37306 8132 37362 8188
rect 37362 8132 37366 8188
rect 37302 8128 37366 8132
rect 51506 8188 51570 8192
rect 51506 8132 51510 8188
rect 51510 8132 51566 8188
rect 51566 8132 51570 8188
rect 51506 8128 51570 8132
rect 51586 8188 51650 8192
rect 51586 8132 51590 8188
rect 51590 8132 51646 8188
rect 51646 8132 51650 8188
rect 51586 8128 51650 8132
rect 51666 8188 51730 8192
rect 51666 8132 51670 8188
rect 51670 8132 51726 8188
rect 51726 8132 51730 8188
rect 51666 8128 51730 8132
rect 51746 8188 51810 8192
rect 51746 8132 51750 8188
rect 51750 8132 51806 8188
rect 51806 8132 51810 8188
rect 51746 8128 51810 8132
rect 15396 7644 15460 7648
rect 15396 7588 15400 7644
rect 15400 7588 15456 7644
rect 15456 7588 15460 7644
rect 15396 7584 15460 7588
rect 15476 7644 15540 7648
rect 15476 7588 15480 7644
rect 15480 7588 15536 7644
rect 15536 7588 15540 7644
rect 15476 7584 15540 7588
rect 15556 7644 15620 7648
rect 15556 7588 15560 7644
rect 15560 7588 15616 7644
rect 15616 7588 15620 7644
rect 15556 7584 15620 7588
rect 15636 7644 15700 7648
rect 15636 7588 15640 7644
rect 15640 7588 15696 7644
rect 15696 7588 15700 7644
rect 15636 7584 15700 7588
rect 29840 7644 29904 7648
rect 29840 7588 29844 7644
rect 29844 7588 29900 7644
rect 29900 7588 29904 7644
rect 29840 7584 29904 7588
rect 29920 7644 29984 7648
rect 29920 7588 29924 7644
rect 29924 7588 29980 7644
rect 29980 7588 29984 7644
rect 29920 7584 29984 7588
rect 30000 7644 30064 7648
rect 30000 7588 30004 7644
rect 30004 7588 30060 7644
rect 30060 7588 30064 7644
rect 30000 7584 30064 7588
rect 30080 7644 30144 7648
rect 30080 7588 30084 7644
rect 30084 7588 30140 7644
rect 30140 7588 30144 7644
rect 30080 7584 30144 7588
rect 44284 7644 44348 7648
rect 44284 7588 44288 7644
rect 44288 7588 44344 7644
rect 44344 7588 44348 7644
rect 44284 7584 44348 7588
rect 44364 7644 44428 7648
rect 44364 7588 44368 7644
rect 44368 7588 44424 7644
rect 44424 7588 44428 7644
rect 44364 7584 44428 7588
rect 44444 7644 44508 7648
rect 44444 7588 44448 7644
rect 44448 7588 44504 7644
rect 44504 7588 44508 7644
rect 44444 7584 44508 7588
rect 44524 7644 44588 7648
rect 44524 7588 44528 7644
rect 44528 7588 44584 7644
rect 44584 7588 44588 7644
rect 44524 7584 44588 7588
rect 58728 7644 58792 7648
rect 58728 7588 58732 7644
rect 58732 7588 58788 7644
rect 58788 7588 58792 7644
rect 58728 7584 58792 7588
rect 58808 7644 58872 7648
rect 58808 7588 58812 7644
rect 58812 7588 58868 7644
rect 58868 7588 58872 7644
rect 58808 7584 58872 7588
rect 58888 7644 58952 7648
rect 58888 7588 58892 7644
rect 58892 7588 58948 7644
rect 58948 7588 58952 7644
rect 58888 7584 58952 7588
rect 58968 7644 59032 7648
rect 58968 7588 58972 7644
rect 58972 7588 59028 7644
rect 59028 7588 59032 7644
rect 58968 7584 59032 7588
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 22618 7100 22682 7104
rect 22618 7044 22622 7100
rect 22622 7044 22678 7100
rect 22678 7044 22682 7100
rect 22618 7040 22682 7044
rect 22698 7100 22762 7104
rect 22698 7044 22702 7100
rect 22702 7044 22758 7100
rect 22758 7044 22762 7100
rect 22698 7040 22762 7044
rect 22778 7100 22842 7104
rect 22778 7044 22782 7100
rect 22782 7044 22838 7100
rect 22838 7044 22842 7100
rect 22778 7040 22842 7044
rect 22858 7100 22922 7104
rect 22858 7044 22862 7100
rect 22862 7044 22918 7100
rect 22918 7044 22922 7100
rect 22858 7040 22922 7044
rect 37062 7100 37126 7104
rect 37062 7044 37066 7100
rect 37066 7044 37122 7100
rect 37122 7044 37126 7100
rect 37062 7040 37126 7044
rect 37142 7100 37206 7104
rect 37142 7044 37146 7100
rect 37146 7044 37202 7100
rect 37202 7044 37206 7100
rect 37142 7040 37206 7044
rect 37222 7100 37286 7104
rect 37222 7044 37226 7100
rect 37226 7044 37282 7100
rect 37282 7044 37286 7100
rect 37222 7040 37286 7044
rect 37302 7100 37366 7104
rect 37302 7044 37306 7100
rect 37306 7044 37362 7100
rect 37362 7044 37366 7100
rect 37302 7040 37366 7044
rect 51506 7100 51570 7104
rect 51506 7044 51510 7100
rect 51510 7044 51566 7100
rect 51566 7044 51570 7100
rect 51506 7040 51570 7044
rect 51586 7100 51650 7104
rect 51586 7044 51590 7100
rect 51590 7044 51646 7100
rect 51646 7044 51650 7100
rect 51586 7040 51650 7044
rect 51666 7100 51730 7104
rect 51666 7044 51670 7100
rect 51670 7044 51726 7100
rect 51726 7044 51730 7100
rect 51666 7040 51730 7044
rect 51746 7100 51810 7104
rect 51746 7044 51750 7100
rect 51750 7044 51806 7100
rect 51806 7044 51810 7100
rect 51746 7040 51810 7044
rect 19380 6972 19444 7036
rect 15396 6556 15460 6560
rect 15396 6500 15400 6556
rect 15400 6500 15456 6556
rect 15456 6500 15460 6556
rect 15396 6496 15460 6500
rect 15476 6556 15540 6560
rect 15476 6500 15480 6556
rect 15480 6500 15536 6556
rect 15536 6500 15540 6556
rect 15476 6496 15540 6500
rect 15556 6556 15620 6560
rect 15556 6500 15560 6556
rect 15560 6500 15616 6556
rect 15616 6500 15620 6556
rect 15556 6496 15620 6500
rect 15636 6556 15700 6560
rect 15636 6500 15640 6556
rect 15640 6500 15696 6556
rect 15696 6500 15700 6556
rect 15636 6496 15700 6500
rect 29840 6556 29904 6560
rect 29840 6500 29844 6556
rect 29844 6500 29900 6556
rect 29900 6500 29904 6556
rect 29840 6496 29904 6500
rect 29920 6556 29984 6560
rect 29920 6500 29924 6556
rect 29924 6500 29980 6556
rect 29980 6500 29984 6556
rect 29920 6496 29984 6500
rect 30000 6556 30064 6560
rect 30000 6500 30004 6556
rect 30004 6500 30060 6556
rect 30060 6500 30064 6556
rect 30000 6496 30064 6500
rect 30080 6556 30144 6560
rect 30080 6500 30084 6556
rect 30084 6500 30140 6556
rect 30140 6500 30144 6556
rect 30080 6496 30144 6500
rect 44284 6556 44348 6560
rect 44284 6500 44288 6556
rect 44288 6500 44344 6556
rect 44344 6500 44348 6556
rect 44284 6496 44348 6500
rect 44364 6556 44428 6560
rect 44364 6500 44368 6556
rect 44368 6500 44424 6556
rect 44424 6500 44428 6556
rect 44364 6496 44428 6500
rect 44444 6556 44508 6560
rect 44444 6500 44448 6556
rect 44448 6500 44504 6556
rect 44504 6500 44508 6556
rect 44444 6496 44508 6500
rect 44524 6556 44588 6560
rect 44524 6500 44528 6556
rect 44528 6500 44584 6556
rect 44584 6500 44588 6556
rect 44524 6496 44588 6500
rect 58728 6556 58792 6560
rect 58728 6500 58732 6556
rect 58732 6500 58788 6556
rect 58788 6500 58792 6556
rect 58728 6496 58792 6500
rect 58808 6556 58872 6560
rect 58808 6500 58812 6556
rect 58812 6500 58868 6556
rect 58868 6500 58872 6556
rect 58808 6496 58872 6500
rect 58888 6556 58952 6560
rect 58888 6500 58892 6556
rect 58892 6500 58948 6556
rect 58948 6500 58952 6556
rect 58888 6496 58952 6500
rect 58968 6556 59032 6560
rect 58968 6500 58972 6556
rect 58972 6500 59028 6556
rect 59028 6500 59032 6556
rect 58968 6496 59032 6500
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 22618 6012 22682 6016
rect 22618 5956 22622 6012
rect 22622 5956 22678 6012
rect 22678 5956 22682 6012
rect 22618 5952 22682 5956
rect 22698 6012 22762 6016
rect 22698 5956 22702 6012
rect 22702 5956 22758 6012
rect 22758 5956 22762 6012
rect 22698 5952 22762 5956
rect 22778 6012 22842 6016
rect 22778 5956 22782 6012
rect 22782 5956 22838 6012
rect 22838 5956 22842 6012
rect 22778 5952 22842 5956
rect 22858 6012 22922 6016
rect 22858 5956 22862 6012
rect 22862 5956 22918 6012
rect 22918 5956 22922 6012
rect 22858 5952 22922 5956
rect 37062 6012 37126 6016
rect 37062 5956 37066 6012
rect 37066 5956 37122 6012
rect 37122 5956 37126 6012
rect 37062 5952 37126 5956
rect 37142 6012 37206 6016
rect 37142 5956 37146 6012
rect 37146 5956 37202 6012
rect 37202 5956 37206 6012
rect 37142 5952 37206 5956
rect 37222 6012 37286 6016
rect 37222 5956 37226 6012
rect 37226 5956 37282 6012
rect 37282 5956 37286 6012
rect 37222 5952 37286 5956
rect 37302 6012 37366 6016
rect 37302 5956 37306 6012
rect 37306 5956 37362 6012
rect 37362 5956 37366 6012
rect 37302 5952 37366 5956
rect 51506 6012 51570 6016
rect 51506 5956 51510 6012
rect 51510 5956 51566 6012
rect 51566 5956 51570 6012
rect 51506 5952 51570 5956
rect 51586 6012 51650 6016
rect 51586 5956 51590 6012
rect 51590 5956 51646 6012
rect 51646 5956 51650 6012
rect 51586 5952 51650 5956
rect 51666 6012 51730 6016
rect 51666 5956 51670 6012
rect 51670 5956 51726 6012
rect 51726 5956 51730 6012
rect 51666 5952 51730 5956
rect 51746 6012 51810 6016
rect 51746 5956 51750 6012
rect 51750 5956 51806 6012
rect 51806 5956 51810 6012
rect 51746 5952 51810 5956
rect 35940 5476 36004 5540
rect 15396 5468 15460 5472
rect 15396 5412 15400 5468
rect 15400 5412 15456 5468
rect 15456 5412 15460 5468
rect 15396 5408 15460 5412
rect 15476 5468 15540 5472
rect 15476 5412 15480 5468
rect 15480 5412 15536 5468
rect 15536 5412 15540 5468
rect 15476 5408 15540 5412
rect 15556 5468 15620 5472
rect 15556 5412 15560 5468
rect 15560 5412 15616 5468
rect 15616 5412 15620 5468
rect 15556 5408 15620 5412
rect 15636 5468 15700 5472
rect 15636 5412 15640 5468
rect 15640 5412 15696 5468
rect 15696 5412 15700 5468
rect 15636 5408 15700 5412
rect 29840 5468 29904 5472
rect 29840 5412 29844 5468
rect 29844 5412 29900 5468
rect 29900 5412 29904 5468
rect 29840 5408 29904 5412
rect 29920 5468 29984 5472
rect 29920 5412 29924 5468
rect 29924 5412 29980 5468
rect 29980 5412 29984 5468
rect 29920 5408 29984 5412
rect 30000 5468 30064 5472
rect 30000 5412 30004 5468
rect 30004 5412 30060 5468
rect 30060 5412 30064 5468
rect 30000 5408 30064 5412
rect 30080 5468 30144 5472
rect 30080 5412 30084 5468
rect 30084 5412 30140 5468
rect 30140 5412 30144 5468
rect 30080 5408 30144 5412
rect 44284 5468 44348 5472
rect 44284 5412 44288 5468
rect 44288 5412 44344 5468
rect 44344 5412 44348 5468
rect 44284 5408 44348 5412
rect 44364 5468 44428 5472
rect 44364 5412 44368 5468
rect 44368 5412 44424 5468
rect 44424 5412 44428 5468
rect 44364 5408 44428 5412
rect 44444 5468 44508 5472
rect 44444 5412 44448 5468
rect 44448 5412 44504 5468
rect 44504 5412 44508 5468
rect 44444 5408 44508 5412
rect 44524 5468 44588 5472
rect 44524 5412 44528 5468
rect 44528 5412 44584 5468
rect 44584 5412 44588 5468
rect 44524 5408 44588 5412
rect 58728 5468 58792 5472
rect 58728 5412 58732 5468
rect 58732 5412 58788 5468
rect 58788 5412 58792 5468
rect 58728 5408 58792 5412
rect 58808 5468 58872 5472
rect 58808 5412 58812 5468
rect 58812 5412 58868 5468
rect 58868 5412 58872 5468
rect 58808 5408 58872 5412
rect 58888 5468 58952 5472
rect 58888 5412 58892 5468
rect 58892 5412 58948 5468
rect 58948 5412 58952 5468
rect 58888 5408 58952 5412
rect 58968 5468 59032 5472
rect 58968 5412 58972 5468
rect 58972 5412 59028 5468
rect 59028 5412 59032 5468
rect 58968 5408 59032 5412
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 22618 4924 22682 4928
rect 22618 4868 22622 4924
rect 22622 4868 22678 4924
rect 22678 4868 22682 4924
rect 22618 4864 22682 4868
rect 22698 4924 22762 4928
rect 22698 4868 22702 4924
rect 22702 4868 22758 4924
rect 22758 4868 22762 4924
rect 22698 4864 22762 4868
rect 22778 4924 22842 4928
rect 22778 4868 22782 4924
rect 22782 4868 22838 4924
rect 22838 4868 22842 4924
rect 22778 4864 22842 4868
rect 22858 4924 22922 4928
rect 22858 4868 22862 4924
rect 22862 4868 22918 4924
rect 22918 4868 22922 4924
rect 22858 4864 22922 4868
rect 37062 4924 37126 4928
rect 37062 4868 37066 4924
rect 37066 4868 37122 4924
rect 37122 4868 37126 4924
rect 37062 4864 37126 4868
rect 37142 4924 37206 4928
rect 37142 4868 37146 4924
rect 37146 4868 37202 4924
rect 37202 4868 37206 4924
rect 37142 4864 37206 4868
rect 37222 4924 37286 4928
rect 37222 4868 37226 4924
rect 37226 4868 37282 4924
rect 37282 4868 37286 4924
rect 37222 4864 37286 4868
rect 37302 4924 37366 4928
rect 37302 4868 37306 4924
rect 37306 4868 37362 4924
rect 37362 4868 37366 4924
rect 37302 4864 37366 4868
rect 51506 4924 51570 4928
rect 51506 4868 51510 4924
rect 51510 4868 51566 4924
rect 51566 4868 51570 4924
rect 51506 4864 51570 4868
rect 51586 4924 51650 4928
rect 51586 4868 51590 4924
rect 51590 4868 51646 4924
rect 51646 4868 51650 4924
rect 51586 4864 51650 4868
rect 51666 4924 51730 4928
rect 51666 4868 51670 4924
rect 51670 4868 51726 4924
rect 51726 4868 51730 4924
rect 51666 4864 51730 4868
rect 51746 4924 51810 4928
rect 51746 4868 51750 4924
rect 51750 4868 51806 4924
rect 51806 4868 51810 4924
rect 51746 4864 51810 4868
rect 15396 4380 15460 4384
rect 15396 4324 15400 4380
rect 15400 4324 15456 4380
rect 15456 4324 15460 4380
rect 15396 4320 15460 4324
rect 15476 4380 15540 4384
rect 15476 4324 15480 4380
rect 15480 4324 15536 4380
rect 15536 4324 15540 4380
rect 15476 4320 15540 4324
rect 15556 4380 15620 4384
rect 15556 4324 15560 4380
rect 15560 4324 15616 4380
rect 15616 4324 15620 4380
rect 15556 4320 15620 4324
rect 15636 4380 15700 4384
rect 15636 4324 15640 4380
rect 15640 4324 15696 4380
rect 15696 4324 15700 4380
rect 15636 4320 15700 4324
rect 29840 4380 29904 4384
rect 29840 4324 29844 4380
rect 29844 4324 29900 4380
rect 29900 4324 29904 4380
rect 29840 4320 29904 4324
rect 29920 4380 29984 4384
rect 29920 4324 29924 4380
rect 29924 4324 29980 4380
rect 29980 4324 29984 4380
rect 29920 4320 29984 4324
rect 30000 4380 30064 4384
rect 30000 4324 30004 4380
rect 30004 4324 30060 4380
rect 30060 4324 30064 4380
rect 30000 4320 30064 4324
rect 30080 4380 30144 4384
rect 30080 4324 30084 4380
rect 30084 4324 30140 4380
rect 30140 4324 30144 4380
rect 30080 4320 30144 4324
rect 44284 4380 44348 4384
rect 44284 4324 44288 4380
rect 44288 4324 44344 4380
rect 44344 4324 44348 4380
rect 44284 4320 44348 4324
rect 44364 4380 44428 4384
rect 44364 4324 44368 4380
rect 44368 4324 44424 4380
rect 44424 4324 44428 4380
rect 44364 4320 44428 4324
rect 44444 4380 44508 4384
rect 44444 4324 44448 4380
rect 44448 4324 44504 4380
rect 44504 4324 44508 4380
rect 44444 4320 44508 4324
rect 44524 4380 44588 4384
rect 44524 4324 44528 4380
rect 44528 4324 44584 4380
rect 44584 4324 44588 4380
rect 44524 4320 44588 4324
rect 58728 4380 58792 4384
rect 58728 4324 58732 4380
rect 58732 4324 58788 4380
rect 58788 4324 58792 4380
rect 58728 4320 58792 4324
rect 58808 4380 58872 4384
rect 58808 4324 58812 4380
rect 58812 4324 58868 4380
rect 58868 4324 58872 4380
rect 58808 4320 58872 4324
rect 58888 4380 58952 4384
rect 58888 4324 58892 4380
rect 58892 4324 58948 4380
rect 58948 4324 58952 4380
rect 58888 4320 58952 4324
rect 58968 4380 59032 4384
rect 58968 4324 58972 4380
rect 58972 4324 59028 4380
rect 59028 4324 59032 4380
rect 58968 4320 59032 4324
rect 6684 3980 6748 4044
rect 16436 3980 16500 4044
rect 19380 3980 19444 4044
rect 42380 3980 42444 4044
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 22618 3836 22682 3840
rect 22618 3780 22622 3836
rect 22622 3780 22678 3836
rect 22678 3780 22682 3836
rect 22618 3776 22682 3780
rect 22698 3836 22762 3840
rect 22698 3780 22702 3836
rect 22702 3780 22758 3836
rect 22758 3780 22762 3836
rect 22698 3776 22762 3780
rect 22778 3836 22842 3840
rect 22778 3780 22782 3836
rect 22782 3780 22838 3836
rect 22838 3780 22842 3836
rect 22778 3776 22842 3780
rect 22858 3836 22922 3840
rect 22858 3780 22862 3836
rect 22862 3780 22918 3836
rect 22918 3780 22922 3836
rect 22858 3776 22922 3780
rect 37062 3836 37126 3840
rect 37062 3780 37066 3836
rect 37066 3780 37122 3836
rect 37122 3780 37126 3836
rect 37062 3776 37126 3780
rect 37142 3836 37206 3840
rect 37142 3780 37146 3836
rect 37146 3780 37202 3836
rect 37202 3780 37206 3836
rect 37142 3776 37206 3780
rect 37222 3836 37286 3840
rect 37222 3780 37226 3836
rect 37226 3780 37282 3836
rect 37282 3780 37286 3836
rect 37222 3776 37286 3780
rect 37302 3836 37366 3840
rect 37302 3780 37306 3836
rect 37306 3780 37362 3836
rect 37362 3780 37366 3836
rect 37302 3776 37366 3780
rect 51506 3836 51570 3840
rect 51506 3780 51510 3836
rect 51510 3780 51566 3836
rect 51566 3780 51570 3836
rect 51506 3776 51570 3780
rect 51586 3836 51650 3840
rect 51586 3780 51590 3836
rect 51590 3780 51646 3836
rect 51646 3780 51650 3836
rect 51586 3776 51650 3780
rect 51666 3836 51730 3840
rect 51666 3780 51670 3836
rect 51670 3780 51726 3836
rect 51726 3780 51730 3836
rect 51666 3776 51730 3780
rect 51746 3836 51810 3840
rect 51746 3780 51750 3836
rect 51750 3780 51806 3836
rect 51806 3780 51810 3836
rect 51746 3776 51810 3780
rect 15396 3292 15460 3296
rect 15396 3236 15400 3292
rect 15400 3236 15456 3292
rect 15456 3236 15460 3292
rect 15396 3232 15460 3236
rect 15476 3292 15540 3296
rect 15476 3236 15480 3292
rect 15480 3236 15536 3292
rect 15536 3236 15540 3292
rect 15476 3232 15540 3236
rect 15556 3292 15620 3296
rect 15556 3236 15560 3292
rect 15560 3236 15616 3292
rect 15616 3236 15620 3292
rect 15556 3232 15620 3236
rect 15636 3292 15700 3296
rect 15636 3236 15640 3292
rect 15640 3236 15696 3292
rect 15696 3236 15700 3292
rect 15636 3232 15700 3236
rect 29840 3292 29904 3296
rect 29840 3236 29844 3292
rect 29844 3236 29900 3292
rect 29900 3236 29904 3292
rect 29840 3232 29904 3236
rect 29920 3292 29984 3296
rect 29920 3236 29924 3292
rect 29924 3236 29980 3292
rect 29980 3236 29984 3292
rect 29920 3232 29984 3236
rect 30000 3292 30064 3296
rect 30000 3236 30004 3292
rect 30004 3236 30060 3292
rect 30060 3236 30064 3292
rect 30000 3232 30064 3236
rect 30080 3292 30144 3296
rect 30080 3236 30084 3292
rect 30084 3236 30140 3292
rect 30140 3236 30144 3292
rect 30080 3232 30144 3236
rect 44284 3292 44348 3296
rect 44284 3236 44288 3292
rect 44288 3236 44344 3292
rect 44344 3236 44348 3292
rect 44284 3232 44348 3236
rect 44364 3292 44428 3296
rect 44364 3236 44368 3292
rect 44368 3236 44424 3292
rect 44424 3236 44428 3292
rect 44364 3232 44428 3236
rect 44444 3292 44508 3296
rect 44444 3236 44448 3292
rect 44448 3236 44504 3292
rect 44504 3236 44508 3292
rect 44444 3232 44508 3236
rect 44524 3292 44588 3296
rect 44524 3236 44528 3292
rect 44528 3236 44584 3292
rect 44584 3236 44588 3292
rect 44524 3232 44588 3236
rect 58728 3292 58792 3296
rect 58728 3236 58732 3292
rect 58732 3236 58788 3292
rect 58788 3236 58792 3292
rect 58728 3232 58792 3236
rect 58808 3292 58872 3296
rect 58808 3236 58812 3292
rect 58812 3236 58868 3292
rect 58868 3236 58872 3292
rect 58808 3232 58872 3236
rect 58888 3292 58952 3296
rect 58888 3236 58892 3292
rect 58892 3236 58948 3292
rect 58948 3236 58952 3292
rect 58888 3232 58952 3236
rect 58968 3292 59032 3296
rect 58968 3236 58972 3292
rect 58972 3236 59028 3292
rect 59028 3236 59032 3292
rect 58968 3232 59032 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 22618 2748 22682 2752
rect 22618 2692 22622 2748
rect 22622 2692 22678 2748
rect 22678 2692 22682 2748
rect 22618 2688 22682 2692
rect 22698 2748 22762 2752
rect 22698 2692 22702 2748
rect 22702 2692 22758 2748
rect 22758 2692 22762 2748
rect 22698 2688 22762 2692
rect 22778 2748 22842 2752
rect 22778 2692 22782 2748
rect 22782 2692 22838 2748
rect 22838 2692 22842 2748
rect 22778 2688 22842 2692
rect 22858 2748 22922 2752
rect 22858 2692 22862 2748
rect 22862 2692 22918 2748
rect 22918 2692 22922 2748
rect 22858 2688 22922 2692
rect 37062 2748 37126 2752
rect 37062 2692 37066 2748
rect 37066 2692 37122 2748
rect 37122 2692 37126 2748
rect 37062 2688 37126 2692
rect 37142 2748 37206 2752
rect 37142 2692 37146 2748
rect 37146 2692 37202 2748
rect 37202 2692 37206 2748
rect 37142 2688 37206 2692
rect 37222 2748 37286 2752
rect 37222 2692 37226 2748
rect 37226 2692 37282 2748
rect 37282 2692 37286 2748
rect 37222 2688 37286 2692
rect 37302 2748 37366 2752
rect 37302 2692 37306 2748
rect 37306 2692 37362 2748
rect 37362 2692 37366 2748
rect 37302 2688 37366 2692
rect 51506 2748 51570 2752
rect 51506 2692 51510 2748
rect 51510 2692 51566 2748
rect 51566 2692 51570 2748
rect 51506 2688 51570 2692
rect 51586 2748 51650 2752
rect 51586 2692 51590 2748
rect 51590 2692 51646 2748
rect 51646 2692 51650 2748
rect 51586 2688 51650 2692
rect 51666 2748 51730 2752
rect 51666 2692 51670 2748
rect 51670 2692 51726 2748
rect 51726 2692 51730 2748
rect 51666 2688 51730 2692
rect 51746 2748 51810 2752
rect 51746 2692 51750 2748
rect 51750 2692 51806 2748
rect 51806 2692 51810 2748
rect 51746 2688 51810 2692
rect 15396 2204 15460 2208
rect 15396 2148 15400 2204
rect 15400 2148 15456 2204
rect 15456 2148 15460 2204
rect 15396 2144 15460 2148
rect 15476 2204 15540 2208
rect 15476 2148 15480 2204
rect 15480 2148 15536 2204
rect 15536 2148 15540 2204
rect 15476 2144 15540 2148
rect 15556 2204 15620 2208
rect 15556 2148 15560 2204
rect 15560 2148 15616 2204
rect 15616 2148 15620 2204
rect 15556 2144 15620 2148
rect 15636 2204 15700 2208
rect 15636 2148 15640 2204
rect 15640 2148 15696 2204
rect 15696 2148 15700 2204
rect 15636 2144 15700 2148
rect 29840 2204 29904 2208
rect 29840 2148 29844 2204
rect 29844 2148 29900 2204
rect 29900 2148 29904 2204
rect 29840 2144 29904 2148
rect 29920 2204 29984 2208
rect 29920 2148 29924 2204
rect 29924 2148 29980 2204
rect 29980 2148 29984 2204
rect 29920 2144 29984 2148
rect 30000 2204 30064 2208
rect 30000 2148 30004 2204
rect 30004 2148 30060 2204
rect 30060 2148 30064 2204
rect 30000 2144 30064 2148
rect 30080 2204 30144 2208
rect 30080 2148 30084 2204
rect 30084 2148 30140 2204
rect 30140 2148 30144 2204
rect 30080 2144 30144 2148
rect 44284 2204 44348 2208
rect 44284 2148 44288 2204
rect 44288 2148 44344 2204
rect 44344 2148 44348 2204
rect 44284 2144 44348 2148
rect 44364 2204 44428 2208
rect 44364 2148 44368 2204
rect 44368 2148 44424 2204
rect 44424 2148 44428 2204
rect 44364 2144 44428 2148
rect 44444 2204 44508 2208
rect 44444 2148 44448 2204
rect 44448 2148 44504 2204
rect 44504 2148 44508 2204
rect 44444 2144 44508 2148
rect 44524 2204 44588 2208
rect 44524 2148 44528 2204
rect 44528 2148 44584 2204
rect 44584 2148 44588 2204
rect 44524 2144 44588 2148
rect 58728 2204 58792 2208
rect 58728 2148 58732 2204
rect 58732 2148 58788 2204
rect 58788 2148 58792 2204
rect 58728 2144 58792 2148
rect 58808 2204 58872 2208
rect 58808 2148 58812 2204
rect 58812 2148 58868 2204
rect 58868 2148 58872 2204
rect 58808 2144 58872 2148
rect 58888 2204 58952 2208
rect 58888 2148 58892 2204
rect 58892 2148 58948 2204
rect 58948 2148 58952 2204
rect 58888 2144 58952 2148
rect 58968 2204 59032 2208
rect 58968 2148 58972 2204
rect 58972 2148 59028 2204
rect 59028 2148 59032 2204
rect 58968 2144 59032 2148
<< metal4 >>
rect 8166 27776 8486 27792
rect 8166 27712 8174 27776
rect 8238 27712 8254 27776
rect 8318 27712 8334 27776
rect 8398 27712 8414 27776
rect 8478 27712 8486 27776
rect 8166 26688 8486 27712
rect 8166 26624 8174 26688
rect 8238 26624 8254 26688
rect 8318 26624 8334 26688
rect 8398 26624 8414 26688
rect 8478 26624 8486 26688
rect 8166 25600 8486 26624
rect 8166 25536 8174 25600
rect 8238 25536 8254 25600
rect 8318 25536 8334 25600
rect 8398 25536 8414 25600
rect 8478 25536 8486 25600
rect 8166 24512 8486 25536
rect 8166 24448 8174 24512
rect 8238 24448 8254 24512
rect 8318 24448 8334 24512
rect 8398 24448 8414 24512
rect 8478 24448 8486 24512
rect 8166 23424 8486 24448
rect 8166 23360 8174 23424
rect 8238 23360 8254 23424
rect 8318 23360 8334 23424
rect 8398 23360 8414 23424
rect 8478 23360 8486 23424
rect 8166 22336 8486 23360
rect 8166 22272 8174 22336
rect 8238 22272 8254 22336
rect 8318 22272 8334 22336
rect 8398 22272 8414 22336
rect 8478 22272 8486 22336
rect 8166 21248 8486 22272
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 8166 20160 8486 21184
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 6683 19412 6749 19413
rect 6683 19348 6684 19412
rect 6748 19348 6749 19412
rect 6683 19347 6749 19348
rect 6686 4045 6746 19347
rect 8166 19072 8486 20096
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 8166 7104 8486 8128
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 8166 6016 8486 7040
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 8166 4928 8486 5952
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 6683 4044 6749 4045
rect 6683 3980 6684 4044
rect 6748 3980 6749 4044
rect 6683 3979 6749 3980
rect 8166 3840 8486 4864
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 2128 8486 2688
rect 15388 27232 15708 27792
rect 15388 27168 15396 27232
rect 15460 27168 15476 27232
rect 15540 27168 15556 27232
rect 15620 27168 15636 27232
rect 15700 27168 15708 27232
rect 15388 26144 15708 27168
rect 15388 26080 15396 26144
rect 15460 26080 15476 26144
rect 15540 26080 15556 26144
rect 15620 26080 15636 26144
rect 15700 26080 15708 26144
rect 15388 25056 15708 26080
rect 15388 24992 15396 25056
rect 15460 24992 15476 25056
rect 15540 24992 15556 25056
rect 15620 24992 15636 25056
rect 15700 24992 15708 25056
rect 15388 23968 15708 24992
rect 15388 23904 15396 23968
rect 15460 23904 15476 23968
rect 15540 23904 15556 23968
rect 15620 23904 15636 23968
rect 15700 23904 15708 23968
rect 15388 22880 15708 23904
rect 15388 22816 15396 22880
rect 15460 22816 15476 22880
rect 15540 22816 15556 22880
rect 15620 22816 15636 22880
rect 15700 22816 15708 22880
rect 15388 21792 15708 22816
rect 15388 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15708 21792
rect 15388 20704 15708 21728
rect 22610 27776 22930 27792
rect 22610 27712 22618 27776
rect 22682 27712 22698 27776
rect 22762 27712 22778 27776
rect 22842 27712 22858 27776
rect 22922 27712 22930 27776
rect 22610 26688 22930 27712
rect 22610 26624 22618 26688
rect 22682 26624 22698 26688
rect 22762 26624 22778 26688
rect 22842 26624 22858 26688
rect 22922 26624 22930 26688
rect 22610 25600 22930 26624
rect 22610 25536 22618 25600
rect 22682 25536 22698 25600
rect 22762 25536 22778 25600
rect 22842 25536 22858 25600
rect 22922 25536 22930 25600
rect 22610 24512 22930 25536
rect 22610 24448 22618 24512
rect 22682 24448 22698 24512
rect 22762 24448 22778 24512
rect 22842 24448 22858 24512
rect 22922 24448 22930 24512
rect 22610 23424 22930 24448
rect 22610 23360 22618 23424
rect 22682 23360 22698 23424
rect 22762 23360 22778 23424
rect 22842 23360 22858 23424
rect 22922 23360 22930 23424
rect 22610 22336 22930 23360
rect 22610 22272 22618 22336
rect 22682 22272 22698 22336
rect 22762 22272 22778 22336
rect 22842 22272 22858 22336
rect 22922 22272 22930 22336
rect 22610 21248 22930 22272
rect 22610 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22930 21248
rect 16435 20772 16501 20773
rect 16435 20708 16436 20772
rect 16500 20708 16501 20772
rect 16435 20707 16501 20708
rect 15388 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15708 20704
rect 15388 19616 15708 20640
rect 15388 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15708 19616
rect 15388 18528 15708 19552
rect 15388 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15708 18528
rect 15388 17440 15708 18464
rect 15388 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15708 17440
rect 15388 16352 15708 17376
rect 15388 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15708 16352
rect 15388 15264 15708 16288
rect 15388 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15708 15264
rect 15388 14176 15708 15200
rect 15388 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15708 14176
rect 15388 13088 15708 14112
rect 15388 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15708 13088
rect 15388 12000 15708 13024
rect 15388 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15708 12000
rect 15388 10912 15708 11936
rect 15388 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15708 10912
rect 15388 9824 15708 10848
rect 15388 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15708 9824
rect 15388 8736 15708 9760
rect 15388 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15708 8736
rect 15388 7648 15708 8672
rect 15388 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15708 7648
rect 15388 6560 15708 7584
rect 15388 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15708 6560
rect 15388 5472 15708 6496
rect 15388 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15708 5472
rect 15388 4384 15708 5408
rect 15388 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15708 4384
rect 15388 3296 15708 4320
rect 16438 4045 16498 20707
rect 22610 20160 22930 21184
rect 22610 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22930 20160
rect 22610 19072 22930 20096
rect 22610 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22930 19072
rect 22610 17984 22930 19008
rect 22610 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22930 17984
rect 22610 16896 22930 17920
rect 22610 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22930 16896
rect 22610 15808 22930 16832
rect 22610 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22930 15808
rect 22610 14720 22930 15744
rect 22610 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22930 14720
rect 22610 13632 22930 14656
rect 22610 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22930 13632
rect 22610 12544 22930 13568
rect 22610 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22930 12544
rect 22610 11456 22930 12480
rect 22610 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22930 11456
rect 22610 10368 22930 11392
rect 22610 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22930 10368
rect 22610 9280 22930 10304
rect 22610 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22930 9280
rect 22610 8192 22930 9216
rect 22610 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22930 8192
rect 22610 7104 22930 8128
rect 22610 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22930 7104
rect 19379 7036 19445 7037
rect 19379 6972 19380 7036
rect 19444 6972 19445 7036
rect 19379 6971 19445 6972
rect 19382 4045 19442 6971
rect 22610 6016 22930 7040
rect 22610 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22930 6016
rect 22610 4928 22930 5952
rect 22610 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22930 4928
rect 16435 4044 16501 4045
rect 16435 3980 16436 4044
rect 16500 3980 16501 4044
rect 16435 3979 16501 3980
rect 19379 4044 19445 4045
rect 19379 3980 19380 4044
rect 19444 3980 19445 4044
rect 19379 3979 19445 3980
rect 15388 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15708 3296
rect 15388 2208 15708 3232
rect 15388 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15708 2208
rect 15388 2128 15708 2144
rect 22610 3840 22930 4864
rect 22610 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22930 3840
rect 22610 2752 22930 3776
rect 22610 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22930 2752
rect 22610 2128 22930 2688
rect 29832 27232 30152 27792
rect 29832 27168 29840 27232
rect 29904 27168 29920 27232
rect 29984 27168 30000 27232
rect 30064 27168 30080 27232
rect 30144 27168 30152 27232
rect 29832 26144 30152 27168
rect 29832 26080 29840 26144
rect 29904 26080 29920 26144
rect 29984 26080 30000 26144
rect 30064 26080 30080 26144
rect 30144 26080 30152 26144
rect 29832 25056 30152 26080
rect 29832 24992 29840 25056
rect 29904 24992 29920 25056
rect 29984 24992 30000 25056
rect 30064 24992 30080 25056
rect 30144 24992 30152 25056
rect 29832 23968 30152 24992
rect 29832 23904 29840 23968
rect 29904 23904 29920 23968
rect 29984 23904 30000 23968
rect 30064 23904 30080 23968
rect 30144 23904 30152 23968
rect 29832 22880 30152 23904
rect 29832 22816 29840 22880
rect 29904 22816 29920 22880
rect 29984 22816 30000 22880
rect 30064 22816 30080 22880
rect 30144 22816 30152 22880
rect 29832 21792 30152 22816
rect 29832 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30152 21792
rect 29832 20704 30152 21728
rect 29832 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30152 20704
rect 29832 19616 30152 20640
rect 29832 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30152 19616
rect 29832 18528 30152 19552
rect 29832 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30152 18528
rect 29832 17440 30152 18464
rect 29832 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30152 17440
rect 29832 16352 30152 17376
rect 29832 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30152 16352
rect 29832 15264 30152 16288
rect 29832 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30152 15264
rect 29832 14176 30152 15200
rect 29832 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30152 14176
rect 29832 13088 30152 14112
rect 29832 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30152 13088
rect 29832 12000 30152 13024
rect 29832 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30152 12000
rect 29832 10912 30152 11936
rect 29832 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30152 10912
rect 29832 9824 30152 10848
rect 29832 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30152 9824
rect 29832 8736 30152 9760
rect 37054 27776 37374 27792
rect 37054 27712 37062 27776
rect 37126 27712 37142 27776
rect 37206 27712 37222 27776
rect 37286 27712 37302 27776
rect 37366 27712 37374 27776
rect 37054 26688 37374 27712
rect 37054 26624 37062 26688
rect 37126 26624 37142 26688
rect 37206 26624 37222 26688
rect 37286 26624 37302 26688
rect 37366 26624 37374 26688
rect 37054 25600 37374 26624
rect 37054 25536 37062 25600
rect 37126 25536 37142 25600
rect 37206 25536 37222 25600
rect 37286 25536 37302 25600
rect 37366 25536 37374 25600
rect 37054 24512 37374 25536
rect 37054 24448 37062 24512
rect 37126 24448 37142 24512
rect 37206 24448 37222 24512
rect 37286 24448 37302 24512
rect 37366 24448 37374 24512
rect 37054 23424 37374 24448
rect 37054 23360 37062 23424
rect 37126 23360 37142 23424
rect 37206 23360 37222 23424
rect 37286 23360 37302 23424
rect 37366 23360 37374 23424
rect 37054 22336 37374 23360
rect 37054 22272 37062 22336
rect 37126 22272 37142 22336
rect 37206 22272 37222 22336
rect 37286 22272 37302 22336
rect 37366 22272 37374 22336
rect 37054 21248 37374 22272
rect 37054 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37374 21248
rect 37054 20160 37374 21184
rect 37054 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37374 20160
rect 37054 19072 37374 20096
rect 37054 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37374 19072
rect 37054 17984 37374 19008
rect 37054 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37374 17984
rect 37054 16896 37374 17920
rect 37054 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37374 16896
rect 37054 15808 37374 16832
rect 37054 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37374 15808
rect 37054 14720 37374 15744
rect 37054 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37374 14720
rect 37054 13632 37374 14656
rect 44276 27232 44596 27792
rect 44276 27168 44284 27232
rect 44348 27168 44364 27232
rect 44428 27168 44444 27232
rect 44508 27168 44524 27232
rect 44588 27168 44596 27232
rect 44276 26144 44596 27168
rect 44276 26080 44284 26144
rect 44348 26080 44364 26144
rect 44428 26080 44444 26144
rect 44508 26080 44524 26144
rect 44588 26080 44596 26144
rect 44276 25056 44596 26080
rect 44276 24992 44284 25056
rect 44348 24992 44364 25056
rect 44428 24992 44444 25056
rect 44508 24992 44524 25056
rect 44588 24992 44596 25056
rect 44276 23968 44596 24992
rect 44276 23904 44284 23968
rect 44348 23904 44364 23968
rect 44428 23904 44444 23968
rect 44508 23904 44524 23968
rect 44588 23904 44596 23968
rect 44276 22880 44596 23904
rect 44276 22816 44284 22880
rect 44348 22816 44364 22880
rect 44428 22816 44444 22880
rect 44508 22816 44524 22880
rect 44588 22816 44596 22880
rect 44276 21792 44596 22816
rect 44276 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44596 21792
rect 44276 20704 44596 21728
rect 44276 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44596 20704
rect 44276 19616 44596 20640
rect 44276 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44596 19616
rect 44276 18528 44596 19552
rect 44276 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44596 18528
rect 44276 17440 44596 18464
rect 44276 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44596 17440
rect 44276 16352 44596 17376
rect 44276 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44596 16352
rect 44276 15264 44596 16288
rect 44276 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44596 15264
rect 44276 14176 44596 15200
rect 44276 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44596 14176
rect 42379 13836 42445 13837
rect 42379 13772 42380 13836
rect 42444 13772 42445 13836
rect 42379 13771 42445 13772
rect 37054 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37374 13632
rect 37054 12544 37374 13568
rect 37054 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37374 12544
rect 37054 11456 37374 12480
rect 37054 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37374 11456
rect 37054 10368 37374 11392
rect 37054 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37374 10368
rect 35939 9756 36005 9757
rect 35939 9692 35940 9756
rect 36004 9692 36005 9756
rect 35939 9691 36005 9692
rect 29832 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30152 8736
rect 29832 7648 30152 8672
rect 29832 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30152 7648
rect 29832 6560 30152 7584
rect 29832 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30152 6560
rect 29832 5472 30152 6496
rect 35942 5541 36002 9691
rect 37054 9280 37374 10304
rect 37054 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37374 9280
rect 37054 8192 37374 9216
rect 37054 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37374 8192
rect 37054 7104 37374 8128
rect 37054 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37374 7104
rect 37054 6016 37374 7040
rect 37054 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37374 6016
rect 35939 5540 36005 5541
rect 35939 5476 35940 5540
rect 36004 5476 36005 5540
rect 35939 5475 36005 5476
rect 29832 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30152 5472
rect 29832 4384 30152 5408
rect 29832 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30152 4384
rect 29832 3296 30152 4320
rect 29832 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30152 3296
rect 29832 2208 30152 3232
rect 29832 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30152 2208
rect 29832 2128 30152 2144
rect 37054 4928 37374 5952
rect 37054 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37374 4928
rect 37054 3840 37374 4864
rect 42382 4045 42442 13771
rect 44276 13088 44596 14112
rect 44276 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44596 13088
rect 44276 12000 44596 13024
rect 44276 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44596 12000
rect 44276 10912 44596 11936
rect 44276 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44596 10912
rect 44276 9824 44596 10848
rect 44276 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44596 9824
rect 44276 8736 44596 9760
rect 44276 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44596 8736
rect 44276 7648 44596 8672
rect 44276 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44596 7648
rect 44276 6560 44596 7584
rect 44276 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44596 6560
rect 44276 5472 44596 6496
rect 44276 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44596 5472
rect 44276 4384 44596 5408
rect 44276 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44596 4384
rect 42379 4044 42445 4045
rect 42379 3980 42380 4044
rect 42444 3980 42445 4044
rect 42379 3979 42445 3980
rect 37054 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37374 3840
rect 37054 2752 37374 3776
rect 37054 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37374 2752
rect 37054 2128 37374 2688
rect 44276 3296 44596 4320
rect 44276 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44596 3296
rect 44276 2208 44596 3232
rect 44276 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44596 2208
rect 44276 2128 44596 2144
rect 51498 27776 51818 27792
rect 51498 27712 51506 27776
rect 51570 27712 51586 27776
rect 51650 27712 51666 27776
rect 51730 27712 51746 27776
rect 51810 27712 51818 27776
rect 51498 26688 51818 27712
rect 51498 26624 51506 26688
rect 51570 26624 51586 26688
rect 51650 26624 51666 26688
rect 51730 26624 51746 26688
rect 51810 26624 51818 26688
rect 51498 25600 51818 26624
rect 51498 25536 51506 25600
rect 51570 25536 51586 25600
rect 51650 25536 51666 25600
rect 51730 25536 51746 25600
rect 51810 25536 51818 25600
rect 51498 24512 51818 25536
rect 51498 24448 51506 24512
rect 51570 24448 51586 24512
rect 51650 24448 51666 24512
rect 51730 24448 51746 24512
rect 51810 24448 51818 24512
rect 51498 23424 51818 24448
rect 51498 23360 51506 23424
rect 51570 23360 51586 23424
rect 51650 23360 51666 23424
rect 51730 23360 51746 23424
rect 51810 23360 51818 23424
rect 51498 22336 51818 23360
rect 51498 22272 51506 22336
rect 51570 22272 51586 22336
rect 51650 22272 51666 22336
rect 51730 22272 51746 22336
rect 51810 22272 51818 22336
rect 51498 21248 51818 22272
rect 51498 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51818 21248
rect 51498 20160 51818 21184
rect 51498 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51818 20160
rect 51498 19072 51818 20096
rect 51498 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51818 19072
rect 51498 17984 51818 19008
rect 51498 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51818 17984
rect 51498 16896 51818 17920
rect 51498 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51818 16896
rect 51498 15808 51818 16832
rect 51498 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51818 15808
rect 51498 14720 51818 15744
rect 51498 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51818 14720
rect 51498 13632 51818 14656
rect 51498 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51818 13632
rect 51498 12544 51818 13568
rect 51498 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51818 12544
rect 51498 11456 51818 12480
rect 51498 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51818 11456
rect 51498 10368 51818 11392
rect 51498 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51818 10368
rect 51498 9280 51818 10304
rect 51498 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51818 9280
rect 51498 8192 51818 9216
rect 51498 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51818 8192
rect 51498 7104 51818 8128
rect 51498 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51818 7104
rect 51498 6016 51818 7040
rect 51498 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51818 6016
rect 51498 4928 51818 5952
rect 51498 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51818 4928
rect 51498 3840 51818 4864
rect 51498 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51818 3840
rect 51498 2752 51818 3776
rect 51498 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51818 2752
rect 51498 2128 51818 2688
rect 58720 27232 59040 27792
rect 58720 27168 58728 27232
rect 58792 27168 58808 27232
rect 58872 27168 58888 27232
rect 58952 27168 58968 27232
rect 59032 27168 59040 27232
rect 58720 26144 59040 27168
rect 58720 26080 58728 26144
rect 58792 26080 58808 26144
rect 58872 26080 58888 26144
rect 58952 26080 58968 26144
rect 59032 26080 59040 26144
rect 58720 25056 59040 26080
rect 58720 24992 58728 25056
rect 58792 24992 58808 25056
rect 58872 24992 58888 25056
rect 58952 24992 58968 25056
rect 59032 24992 59040 25056
rect 58720 23968 59040 24992
rect 58720 23904 58728 23968
rect 58792 23904 58808 23968
rect 58872 23904 58888 23968
rect 58952 23904 58968 23968
rect 59032 23904 59040 23968
rect 58720 22880 59040 23904
rect 58720 22816 58728 22880
rect 58792 22816 58808 22880
rect 58872 22816 58888 22880
rect 58952 22816 58968 22880
rect 59032 22816 59040 22880
rect 58720 21792 59040 22816
rect 58720 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59040 21792
rect 58720 20704 59040 21728
rect 58720 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59040 20704
rect 58720 19616 59040 20640
rect 58720 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59040 19616
rect 58720 18528 59040 19552
rect 58720 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59040 18528
rect 58720 17440 59040 18464
rect 58720 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59040 17440
rect 58720 16352 59040 17376
rect 58720 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59040 16352
rect 58720 15264 59040 16288
rect 58720 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59040 15264
rect 58720 14176 59040 15200
rect 58720 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59040 14176
rect 58720 13088 59040 14112
rect 58720 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59040 13088
rect 58720 12000 59040 13024
rect 58720 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59040 12000
rect 58720 10912 59040 11936
rect 58720 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59040 10912
rect 58720 9824 59040 10848
rect 58720 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59040 9824
rect 58720 8736 59040 9760
rect 58720 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59040 8736
rect 58720 7648 59040 8672
rect 58720 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59040 7648
rect 58720 6560 59040 7584
rect 58720 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59040 6560
rect 58720 5472 59040 6496
rect 58720 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59040 5472
rect 58720 4384 59040 5408
rect 58720 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59040 4384
rect 58720 3296 59040 4320
rect 58720 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59040 3296
rect 58720 2208 59040 3232
rect 58720 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59040 2208
rect 58720 2128 59040 2144
use sky130_fd_sc_hd__inv_2  _0437_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0438_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0439_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0440_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0441_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0442_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0443_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0444_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0445_
timestamp 1688980957
transform 1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0446_
timestamp 1688980957
transform 1 0 8832 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0447_
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0448_
timestamp 1688980957
transform 1 0 9568 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0449_
timestamp 1688980957
transform 1 0 14536 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0450_
timestamp 1688980957
transform 1 0 12696 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0451_
timestamp 1688980957
transform 1 0 15272 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0452_
timestamp 1688980957
transform 1 0 17572 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0453_
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0454_
timestamp 1688980957
transform 1 0 19872 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0455_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0456_
timestamp 1688980957
transform 1 0 23644 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0457_
timestamp 1688980957
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0458_
timestamp 1688980957
transform 1 0 30544 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0459_
timestamp 1688980957
transform 1 0 28796 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0460_
timestamp 1688980957
transform 1 0 31464 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0461_
timestamp 1688980957
transform -1 0 35788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0462_
timestamp 1688980957
transform 1 0 32752 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0463_
timestamp 1688980957
transform -1 0 38732 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0464_
timestamp 1688980957
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0465_
timestamp 1688980957
transform 1 0 41676 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0466_
timestamp 1688980957
transform 1 0 42596 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0467_
timestamp 1688980957
transform -1 0 41952 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0468_
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0469_
timestamp 1688980957
transform 1 0 47748 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0470_
timestamp 1688980957
transform 1 0 47012 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0471_
timestamp 1688980957
transform -1 0 52624 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0472_
timestamp 1688980957
transform 1 0 50784 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0473_
timestamp 1688980957
transform -1 0 53636 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0474_
timestamp 1688980957
transform 1 0 52532 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0475_
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_4  _0476_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0477_
timestamp 1688980957
transform -1 0 4600 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0478_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0479_
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0480_
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0481_
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0482_
timestamp 1688980957
transform 1 0 15272 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0483_
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0484_
timestamp 1688980957
transform -1 0 16100 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0485_
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0486_
timestamp 1688980957
transform 1 0 20884 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0487_
timestamp 1688980957
transform 1 0 20608 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0488_
timestamp 1688980957
transform 1 0 23184 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0489_
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0490_
timestamp 1688980957
transform 1 0 25760 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0491_
timestamp 1688980957
transform 1 0 28612 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0492_
timestamp 1688980957
transform 1 0 28612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0494_
timestamp 1688980957
transform 1 0 35788 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0495_
timestamp 1688980957
transform 1 0 33580 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0496_
timestamp 1688980957
transform 1 0 38548 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0497_
timestamp 1688980957
transform 1 0 36892 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0498_
timestamp 1688980957
transform -1 0 42228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0499_
timestamp 1688980957
transform -1 0 43240 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0500_
timestamp 1688980957
transform 1 0 41676 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0501_
timestamp 1688980957
transform 1 0 44804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0502_
timestamp 1688980957
transform 1 0 48208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0503_
timestamp 1688980957
transform -1 0 47104 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0504_
timestamp 1688980957
transform -1 0 55752 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0505_
timestamp 1688980957
transform 1 0 50692 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0506_
timestamp 1688980957
transform -1 0 56120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0507_
timestamp 1688980957
transform -1 0 56028 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0508_
timestamp 1688980957
transform -1 0 55200 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0509_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0510_
timestamp 1688980957
transform -1 0 4232 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0511_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3588 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0512_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0513_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1688980957
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0515_
timestamp 1688980957
transform -1 0 6348 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0516_
timestamp 1688980957
transform -1 0 6808 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0517_
timestamp 1688980957
transform -1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0518_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0519_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0520_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0521_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0522_
timestamp 1688980957
transform -1 0 3680 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0523_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0524_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2944 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0525_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0526_
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0527_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0528_
timestamp 1688980957
transform 1 0 4692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0529_
timestamp 1688980957
transform -1 0 4324 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0530_
timestamp 1688980957
transform -1 0 5612 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0531_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_4  _0532_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0533_
timestamp 1688980957
transform -1 0 7912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0534_
timestamp 1688980957
transform -1 0 7728 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0535_
timestamp 1688980957
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0536_
timestamp 1688980957
transform 1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0537_
timestamp 1688980957
transform 1 0 12420 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0538_
timestamp 1688980957
transform -1 0 17756 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1688980957
transform -1 0 17480 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0540_
timestamp 1688980957
transform -1 0 18952 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0541_
timestamp 1688980957
transform -1 0 20976 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0542_
timestamp 1688980957
transform -1 0 23552 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0543_
timestamp 1688980957
transform -1 0 23644 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0544_
timestamp 1688980957
transform -1 0 26496 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0545_
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0546_
timestamp 1688980957
transform 1 0 26956 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0547_
timestamp 1688980957
transform -1 0 31004 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0548_
timestamp 1688980957
transform -1 0 33764 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0549_
timestamp 1688980957
transform -1 0 34408 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0550_
timestamp 1688980957
transform -1 0 38916 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1688980957
transform -1 0 36800 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0552_
timestamp 1688980957
transform -1 0 41400 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0553_
timestamp 1688980957
transform -1 0 40664 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0554_
timestamp 1688980957
transform -1 0 44252 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0555_
timestamp 1688980957
transform -1 0 45816 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0556_
timestamp 1688980957
transform 1 0 44344 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0557_
timestamp 1688980957
transform -1 0 48392 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1688980957
transform -1 0 50600 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1688980957
transform -1 0 49772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1688980957
transform 1 0 56764 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1688980957
transform -1 0 53544 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1688980957
transform 1 0 56856 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1688980957
transform 1 0 56856 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1688980957
transform 1 0 57592 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0565_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0568_
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1688980957
transform 1 0 9384 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0572_
timestamp 1688980957
transform 1 0 13064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0573_
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1688980957
transform 1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0575_
timestamp 1688980957
transform 1 0 20056 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0577_
timestamp 1688980957
transform 1 0 23460 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0578_
timestamp 1688980957
transform 1 0 22816 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 1688980957
transform 1 0 26496 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1688980957
transform 1 0 28888 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0581_
timestamp 1688980957
transform 1 0 28612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0582_
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0583_
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1688980957
transform 1 0 33488 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1688980957
transform -1 0 37904 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0587_
timestamp 1688980957
transform -1 0 40940 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1688980957
transform 1 0 41768 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1688980957
transform 1 0 41032 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1688980957
transform -1 0 45908 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 1688980957
transform 1 0 46920 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1688980957
transform 1 0 46184 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1688980957
transform 1 0 52992 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1688980957
transform -1 0 50876 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1688980957
transform -1 0 53544 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1688980957
transform 1 0 52072 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0598_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1688980957
transform -1 0 6256 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1688980957
transform 1 0 3864 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1688980957
transform 1 0 11040 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1688980957
transform -1 0 14996 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0606_
timestamp 1688980957
transform -1 0 17572 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1688980957
transform -1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1688980957
transform 1 0 22264 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 1688980957
transform 1 0 23920 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 1688980957
transform 1 0 27876 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1688980957
transform 1 0 29716 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1688980957
transform -1 0 33396 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0615_
timestamp 1688980957
transform 1 0 34040 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1688980957
transform -1 0 38088 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0617_
timestamp 1688980957
transform 1 0 36156 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1688980957
transform -1 0 39376 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1688980957
transform -1 0 42872 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1688980957
transform -1 0 45816 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1688980957
transform -1 0 43332 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1688980957
transform -1 0 48392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1688980957
transform 1 0 49220 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0625_
timestamp 1688980957
transform -1 0 49128 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1688980957
transform 1 0 54096 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1688980957
transform -1 0 52256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1688980957
transform -1 0 56120 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1688980957
transform 1 0 54464 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1688980957
transform 1 0 53176 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _0631_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6256 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1688980957
transform 1 0 7176 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1688980957
transform -1 0 7084 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1688980957
transform -1 0 11040 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform -1 0 12788 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1688980957
transform -1 0 18308 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1688980957
transform 1 0 18216 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1688980957
transform -1 0 20148 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1688980957
transform -1 0 22632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 23368 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0644_
timestamp 1688980957
transform -1 0 26864 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1688980957
transform 1 0 28888 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1688980957
transform 1 0 29992 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0647_
timestamp 1688980957
transform 1 0 33396 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0648_
timestamp 1688980957
transform -1 0 33856 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1688980957
transform -1 0 37996 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0650_
timestamp 1688980957
transform 1 0 35696 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0651_
timestamp 1688980957
transform -1 0 38824 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0652_
timestamp 1688980957
transform 1 0 39652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0653_
timestamp 1688980957
transform -1 0 44160 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0654_
timestamp 1688980957
transform -1 0 45632 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 1688980957
transform 1 0 43884 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0656_
timestamp 1688980957
transform -1 0 48024 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0657_
timestamp 1688980957
transform -1 0 50968 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1688980957
transform 1 0 50140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0659_
timestamp 1688980957
transform -1 0 56120 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0660_
timestamp 1688980957
transform -1 0 52624 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0661_
timestamp 1688980957
transform -1 0 55108 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0662_
timestamp 1688980957
transform 1 0 55936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0663_
timestamp 1688980957
transform -1 0 53544 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0664_
timestamp 1688980957
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0665_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5336 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0666_
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0667_
timestamp 1688980957
transform -1 0 3036 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0668_
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0669_
timestamp 1688980957
transform 1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_2  _0670_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1688980957
transform -1 0 6348 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0672_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0673_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7360 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0674_
timestamp 1688980957
transform 1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0675_
timestamp 1688980957
transform 1 0 6808 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0676_
timestamp 1688980957
transform 1 0 6348 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0677_
timestamp 1688980957
transform -1 0 9292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0678_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0679_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0681_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0682_
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1688980957
transform 1 0 10212 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0685_
timestamp 1688980957
transform 1 0 14444 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1688980957
transform 1 0 18400 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1688980957
transform 1 0 19780 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1688980957
transform 1 0 23828 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1688980957
transform 1 0 28704 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1688980957
transform -1 0 28612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1688980957
transform 1 0 31004 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1688980957
transform 1 0 34776 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1688980957
transform -1 0 33488 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1688980957
transform 1 0 37628 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1688980957
transform 1 0 36064 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1688980957
transform -1 0 41216 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1688980957
transform 1 0 41676 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1688980957
transform 1 0 40848 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1688980957
transform 1 0 44988 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1688980957
transform -1 0 48392 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1688980957
transform 1 0 46276 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1688980957
transform 1 0 54096 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1688980957
transform 1 0 50140 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1688980957
transform -1 0 54832 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1688980957
transform -1 0 55016 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1688980957
transform 1 0 54372 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _0712_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 1688980957
transform 1 0 7912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0717_
timestamp 1688980957
transform 1 0 11224 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1688980957
transform -1 0 17480 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1688980957
transform 1 0 15456 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0722_
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1688980957
transform 1 0 25392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1688980957
transform -1 0 26772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1688980957
transform -1 0 26864 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1688980957
transform 1 0 30084 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1688980957
transform -1 0 33304 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1688980957
transform -1 0 37996 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1688980957
transform -1 0 35788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1688980957
transform -1 0 39744 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0733_
timestamp 1688980957
transform 1 0 38548 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1688980957
transform 1 0 44068 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1688980957
transform 1 0 44068 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1688980957
transform 1 0 42964 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 1688980957
transform 1 0 46552 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1688980957
transform -1 0 50968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1688980957
transform -1 0 50968 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform -1 0 58052 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1688980957
transform 1 0 51520 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform -1 0 57500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1688980957
transform 1 0 56764 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1688980957
transform -1 0 57316 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0745_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7636 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__mux4_1  _0746_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0747_
timestamp 1688980957
transform -1 0 7176 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform 1 0 6532 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0749_
timestamp 1688980957
transform 1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0750_
timestamp 1688980957
transform -1 0 6256 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0751_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0754_
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0755_
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0757_
timestamp 1688980957
transform -1 0 11316 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0758_
timestamp 1688980957
transform -1 0 13432 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0759_
timestamp 1688980957
transform -1 0 12604 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1688980957
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1688980957
transform -1 0 12512 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0762_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0763_
timestamp 1688980957
transform 1 0 10580 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1688980957
transform -1 0 14260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0766_
timestamp 1688980957
transform -1 0 17480 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0767_
timestamp 1688980957
transform -1 0 17480 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1688980957
transform 1 0 16468 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1688980957
transform 1 0 16468 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0770_
timestamp 1688980957
transform -1 0 16468 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0771_
timestamp 1688980957
transform -1 0 16100 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0774_
timestamp 1688980957
transform -1 0 18308 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0775_
timestamp 1688980957
transform -1 0 18216 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1688980957
transform 1 0 18308 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1688980957
transform 1 0 18124 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0778_
timestamp 1688980957
transform -1 0 21160 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0779_
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1688980957
transform -1 0 20976 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 20240 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0782_
timestamp 1688980957
transform -1 0 23736 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0783_
timestamp 1688980957
transform 1 0 20884 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1688980957
transform 1 0 22080 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0786_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0787_
timestamp 1688980957
transform -1 0 23368 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1688980957
transform -1 0 24564 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0790_
timestamp 1688980957
transform 1 0 24472 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0791_
timestamp 1688980957
transform -1 0 27140 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1688980957
transform 1 0 26404 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1688980957
transform 1 0 25484 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0794_
timestamp 1688980957
transform -1 0 26864 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0795_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1688980957
transform -1 0 27784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1688980957
transform -1 0 27784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0798_
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0799_
timestamp 1688980957
transform -1 0 28888 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1688980957
transform 1 0 27784 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1688980957
transform 1 0 27232 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0802_
timestamp 1688980957
transform 1 0 29532 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0803_
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1688980957
transform 1 0 31464 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1688980957
transform 1 0 30360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0806_
timestamp 1688980957
transform -1 0 32568 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0807_
timestamp 1688980957
transform -1 0 32568 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1688980957
transform -1 0 32936 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0810_
timestamp 1688980957
transform -1 0 33580 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0811_
timestamp 1688980957
transform -1 0 34040 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1688980957
transform 1 0 33580 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1688980957
transform -1 0 33856 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0814_
timestamp 1688980957
transform -1 0 37720 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0815_
timestamp 1688980957
transform -1 0 37168 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1688980957
transform 1 0 35880 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0818_
timestamp 1688980957
transform -1 0 36616 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0819_
timestamp 1688980957
transform -1 0 35696 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1688980957
transform 1 0 35972 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1688980957
transform 1 0 35052 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0822_
timestamp 1688980957
transform -1 0 40572 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0823_
timestamp 1688980957
transform 1 0 37628 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1688980957
transform 1 0 39560 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1688980957
transform -1 0 39560 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0826_
timestamp 1688980957
transform -1 0 39652 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0827_
timestamp 1688980957
transform -1 0 39652 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 1688980957
transform -1 0 40664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform -1 0 40664 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0830_
timestamp 1688980957
transform -1 0 44344 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0831_
timestamp 1688980957
transform -1 0 43332 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp 1688980957
transform 1 0 42320 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1688980957
transform 1 0 41860 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0834_
timestamp 1688980957
transform -1 0 44804 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0835_
timestamp 1688980957
transform -1 0 44804 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp 1688980957
transform 1 0 43976 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 1688980957
transform 1 0 43424 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0838_
timestamp 1688980957
transform -1 0 44344 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0839_
timestamp 1688980957
transform 1 0 42596 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp 1688980957
transform -1 0 45632 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0842_
timestamp 1688980957
transform -1 0 47840 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0843_
timestamp 1688980957
transform 1 0 46552 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 1688980957
transform 1 0 48484 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1688980957
transform -1 0 47472 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0846_
timestamp 1688980957
transform -1 0 50324 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0847_
timestamp 1688980957
transform -1 0 50140 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1688980957
transform 1 0 49220 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1688980957
transform -1 0 49128 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0850_
timestamp 1688980957
transform -1 0 49496 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0851_
timestamp 1688980957
transform -1 0 49496 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1688980957
transform 1 0 49680 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1688980957
transform -1 0 49956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0854_
timestamp 1688980957
transform -1 0 57224 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0855_
timestamp 1688980957
transform -1 0 55200 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1688980957
transform 1 0 54372 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1688980957
transform 1 0 53268 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0858_
timestamp 1688980957
transform -1 0 52716 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0859_
timestamp 1688980957
transform 1 0 50600 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1688980957
transform -1 0 52348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0862_
timestamp 1688980957
transform -1 0 57500 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0863_
timestamp 1688980957
transform 1 0 54280 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1688980957
transform -1 0 56948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0865_
timestamp 1688980957
transform 1 0 57684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0866_
timestamp 1688980957
transform -1 0 57592 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0867_
timestamp 1688980957
transform -1 0 55936 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0868_
timestamp 1688980957
transform -1 0 57408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0869_
timestamp 1688980957
transform 1 0 56856 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0870_
timestamp 1688980957
transform -1 0 57592 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0871_
timestamp 1688980957
transform -1 0 53636 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0872_
timestamp 1688980957
transform -1 0 57592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1688980957
transform -1 0 57776 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _0874_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1688980957
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1688980957
transform 1 0 1840 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1688980957
transform -1 0 9660 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1688980957
transform 1 0 9016 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1688980957
transform 1 0 12512 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1688980957
transform 1 0 14536 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1688980957
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1688980957
transform 1 0 19688 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1688980957
transform 1 0 19320 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1688980957
transform 1 0 24104 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1688980957
transform 1 0 22816 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1688980957
transform 1 0 25300 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1688980957
transform 1 0 28244 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1688980957
transform 1 0 28520 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1688980957
transform 1 0 30176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1688980957
transform 1 0 32016 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1688980957
transform 1 0 37628 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1688980957
transform 1 0 39928 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1688980957
transform 1 0 41308 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1688980957
transform 1 0 40388 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1688980957
transform 1 0 46000 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1688980957
transform 1 0 46552 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1688980957
transform 1 0 45632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1688980957
transform 1 0 51888 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1688980957
transform 1 0 49312 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1688980957
transform 1 0 53268 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1688980957
transform 1 0 51796 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1688980957
transform -1 0 51888 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1688980957
transform -1 0 5428 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1688980957
transform 1 0 2024 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1688980957
transform 1 0 9200 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1688980957
transform 1 0 13800 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1688980957
transform 1 0 14628 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1688980957
transform 1 0 19412 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1688980957
transform 1 0 19136 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1688980957
transform 1 0 22448 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1688980957
transform 1 0 27968 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1688980957
transform 1 0 28704 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1688980957
transform 1 0 29532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1688980957
transform 1 0 34408 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1688980957
transform 1 0 32384 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1688980957
transform 1 0 37444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1688980957
transform 1 0 35420 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1688980957
transform 1 0 39928 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1688980957
transform 1 0 41308 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1688980957
transform 1 0 40296 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1688980957
transform 1 0 44068 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1688980957
transform 1 0 46736 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1688980957
transform 1 0 45724 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1688980957
transform 1 0 54556 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1688980957
transform 1 0 49220 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1688980957
transform 1 0 53728 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1688980957
transform 1 0 55292 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1688980957
transform 1 0 54556 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1688980957
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1688980957
transform 1 0 2392 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1688980957
transform -1 0 5336 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1688980957
transform 1 0 6348 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1688980957
transform 1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1688980957
transform -1 0 18952 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1688980957
transform -1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1688980957
transform -1 0 18768 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1688980957
transform -1 0 26680 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1688980957
transform 1 0 25944 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1688980957
transform 1 0 26956 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1688980957
transform -1 0 31188 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1688980957
transform 1 0 32568 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1688980957
transform 1 0 32660 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1688980957
transform 1 0 34776 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1688980957
transform 1 0 39744 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1688980957
transform 1 0 39652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1688980957
transform 1 0 43240 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1688980957
transform 1 0 44252 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1688980957
transform -1 0 49312 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1688980957
transform -1 0 51612 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1688980957
transform 1 0 48576 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1688980957
transform 1 0 56304 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1688980957
transform 1 0 52716 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1688980957
transform 1 0 56672 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1688980957
transform 1 0 56764 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1688980957
transform 1 0 56856 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1688980957
transform -1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1688980957
transform -1 0 10120 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1688980957
transform 1 0 13616 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1688980957
transform 1 0 14260 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1688980957
transform 1 0 16836 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1688980957
transform 1 0 19412 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1688980957
transform 1 0 23736 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1688980957
transform 1 0 22080 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1688980957
transform 1 0 25024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1688980957
transform 1 0 27968 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1688980957
transform 1 0 28520 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1688980957
transform 1 0 30084 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1688980957
transform 1 0 33764 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1688980957
transform 1 0 35420 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1688980957
transform 1 0 39836 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1688980957
transform 1 0 40848 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1688980957
transform 1 0 40388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1688980957
transform 1 0 46000 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1688980957
transform 1 0 45632 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1688980957
transform 1 0 51520 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1688980957
transform 1 0 50140 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1688980957
transform 1 0 51796 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1688980957
transform 1 0 51152 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1688980957
transform 1 0 50600 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1688980957
transform 1 0 5704 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1688980957
transform -1 0 11224 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1688980957
transform -1 0 11960 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1688980957
transform 1 0 16376 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1688980957
transform 1 0 13524 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1688980957
transform -1 0 18124 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1688980957
transform -1 0 19136 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1688980957
transform -1 0 22816 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1688980957
transform 1 0 25392 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1688980957
transform 1 0 22448 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1688980957
transform 1 0 27508 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1688980957
transform 1 0 28888 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1688980957
transform 1 0 30544 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1688980957
transform 1 0 32476 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1688980957
transform 1 0 36156 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1688980957
transform -1 0 38548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1688980957
transform 1 0 38180 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1688980957
transform 1 0 43424 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1688980957
transform -1 0 44344 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1688980957
transform -1 0 48392 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1688980957
transform 1 0 48576 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1688980957
transform 1 0 47840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1688980957
transform 1 0 53636 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1688980957
transform -1 0 51428 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1688980957
transform 1 0 53728 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1688980957
transform 1 0 53728 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1688980957
transform 1 0 51152 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1688980957
transform 1 0 6440 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1688980957
transform 1 0 11960 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1688980957
transform -1 0 12972 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1688980957
transform 1 0 16100 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1688980957
transform 1 0 17112 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1688980957
transform -1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1688980957
transform -1 0 22356 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1688980957
transform 1 0 22448 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1688980957
transform 1 0 26036 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1688980957
transform -1 0 26864 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1688980957
transform 1 0 27968 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1688980957
transform 1 0 32568 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1688980957
transform -1 0 39100 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1688980957
transform 1 0 34500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1688980957
transform 1 0 37536 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1688980957
transform 1 0 38548 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1688980957
transform 1 0 43056 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1688980957
transform 1 0 43792 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1688980957
transform 1 0 43332 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1688980957
transform -1 0 49036 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1688980957
transform 1 0 50140 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1688980957
transform 1 0 48116 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1688980957
transform 1 0 55200 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1688980957
transform -1 0 54004 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1688980957
transform -1 0 56580 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1688980957
transform 1 0 55292 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1688980957
transform 1 0 51704 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1071_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1072_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7912 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1688980957
transform -1 0 8280 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1688980957
transform 1 0 6624 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1075_
timestamp 1688980957
transform 1 0 8004 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1688980957
transform 1 0 9108 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1688980957
transform -1 0 13984 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1688980957
transform 1 0 14444 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1688980957
transform 1 0 17664 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1688980957
transform 1 0 22448 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1688980957
transform 1 0 28520 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1688980957
transform 1 0 29624 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1688980957
transform 1 0 32108 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1688980957
transform 1 0 37076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1688980957
transform 1 0 35512 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1688980957
transform 1 0 39836 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1688980957
transform 1 0 40848 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1688980957
transform 1 0 40296 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1688980957
transform 1 0 43424 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1688980957
transform -1 0 48116 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1688980957
transform 1 0 45632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1688980957
transform 1 0 52900 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1688980957
transform 1 0 48300 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1688980957
transform 1 0 53452 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1688980957
transform 1 0 53728 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1688980957
transform 1 0 54096 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1688980957
transform 1 0 9936 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1688980957
transform 1 0 10948 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1688980957
transform -1 0 18124 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1688980957
transform 1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1688980957
transform 1 0 19136 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1688980957
transform 1 0 21252 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1688980957
transform -1 0 22540 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1688980957
transform -1 0 26404 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1688980957
transform -1 0 26864 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1688980957
transform -1 0 31188 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1688980957
transform 1 0 30544 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1688980957
transform -1 0 39192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp 1688980957
transform 1 0 34500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp 1688980957
transform -1 0 41308 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1688980957
transform 1 0 38088 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1688980957
transform 1 0 42596 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1688980957
transform 1 0 43700 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1688980957
transform 1 0 42504 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1688980957
transform 1 0 46000 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1688980957
transform -1 0 51796 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1688980957
transform 1 0 48208 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1688980957
transform 1 0 56304 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1688980957
transform 1 0 50784 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1688980957
transform 1 0 56396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1688980957
transform 1 0 56672 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1688980957
transform 1 0 56028 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1688980957
transform 1 0 5796 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1688980957
transform -1 0 11408 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1688980957
transform -1 0 13616 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1688980957
transform -1 0 15824 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1688980957
transform 1 0 14996 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1688980957
transform 1 0 17664 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1688980957
transform 1 0 19596 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1688980957
transform -1 0 22540 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1688980957
transform 1 0 23368 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1688980957
transform 1 0 24748 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1688980957
transform 1 0 26220 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1688980957
transform 1 0 29900 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1688980957
transform 1 0 31556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1688980957
transform 1 0 33028 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1688980957
transform 1 0 34592 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1688980957
transform 1 0 37996 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1688980957
transform 1 0 38824 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1688980957
transform 1 0 40388 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1688980957
transform 1 0 42872 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1688980957
transform 1 0 46460 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1688980957
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1688980957
transform 1 0 48484 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1688980957
transform 1 0 51796 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1688980957
transform 1 0 51060 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1688980957
transform 1 0 56212 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1688980957
transform 1 0 56304 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1688980957
transform 1 0 56856 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__S asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0445__S
timestamp 1688980957
transform -1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__S
timestamp 1688980957
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__S
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__S
timestamp 1688980957
transform 1 0 9384 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__S
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__S
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__S
timestamp 1688980957
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__S
timestamp 1688980957
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__S
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__S
timestamp 1688980957
transform -1 0 19780 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__S
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__S
timestamp 1688980957
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0457__S
timestamp 1688980957
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__S
timestamp 1688980957
transform 1 0 31096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__S
timestamp 1688980957
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__S
timestamp 1688980957
transform 1 0 30452 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0461__S
timestamp 1688980957
transform 1 0 34776 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__S
timestamp 1688980957
transform 1 0 32568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__S
timestamp 1688980957
transform 1 0 40020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__S
timestamp 1688980957
transform 1 0 35880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__S
timestamp 1688980957
transform 1 0 40756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__S
timestamp 1688980957
transform 1 0 42596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__S
timestamp 1688980957
transform 1 0 40480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__S
timestamp 1688980957
transform 1 0 48208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__S
timestamp 1688980957
transform -1 0 47472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__S
timestamp 1688980957
transform 1 0 47012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__S
timestamp 1688980957
transform 1 0 52900 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__S
timestamp 1688980957
transform 1 0 51888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__S
timestamp 1688980957
transform 1 0 52900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__S
timestamp 1688980957
transform 1 0 52440 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__S
timestamp 1688980957
transform -1 0 53912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__S
timestamp 1688980957
transform 1 0 5704 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__S
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__S
timestamp 1688980957
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__S
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__S
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__S
timestamp 1688980957
transform 1 0 15640 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__S
timestamp 1688980957
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__S
timestamp 1688980957
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__S
timestamp 1688980957
transform -1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__S
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__S
timestamp 1688980957
transform 1 0 20976 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__S
timestamp 1688980957
transform 1 0 23000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__S
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__S
timestamp 1688980957
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__S
timestamp 1688980957
transform 1 0 28060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__S
timestamp 1688980957
transform -1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__S
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__S
timestamp 1688980957
transform 1 0 36432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__S
timestamp 1688980957
transform 1 0 36800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__S
timestamp 1688980957
transform 1 0 39192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__S
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__S
timestamp 1688980957
transform 1 0 42412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__S
timestamp 1688980957
transform 1 0 42688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__S
timestamp 1688980957
transform 1 0 41952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__S
timestamp 1688980957
transform 1 0 44620 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__S
timestamp 1688980957
transform -1 0 48208 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__S
timestamp 1688980957
transform 1 0 46092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__S
timestamp 1688980957
transform -1 0 54740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__S
timestamp 1688980957
transform 1 0 50508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__S
timestamp 1688980957
transform -1 0 56580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__S
timestamp 1688980957
transform 1 0 54648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__S
timestamp 1688980957
transform -1 0 55660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__B
timestamp 1688980957
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A_N
timestamp 1688980957
transform 1 0 4416 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A_N
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1688980957
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A_N
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__B
timestamp 1688980957
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__S
timestamp 1688980957
transform -1 0 6256 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__S
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__S
timestamp 1688980957
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__S
timestamp 1688980957
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__S
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__S
timestamp 1688980957
transform -1 0 16560 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__S
timestamp 1688980957
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__S
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__S
timestamp 1688980957
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__S
timestamp 1688980957
transform 1 0 22724 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__S
timestamp 1688980957
transform 1 0 22632 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__S
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__S
timestamp 1688980957
transform 1 0 27876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__S
timestamp 1688980957
transform 1 0 27324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__S
timestamp 1688980957
transform 1 0 31188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__S
timestamp 1688980957
transform 1 0 34040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__S
timestamp 1688980957
transform 1 0 33396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__S
timestamp 1688980957
transform 1 0 37720 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S
timestamp 1688980957
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__S
timestamp 1688980957
transform 1 0 40388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__S
timestamp 1688980957
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__S
timestamp 1688980957
transform 1 0 45172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__S
timestamp 1688980957
transform -1 0 44896 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__S
timestamp 1688980957
transform -1 0 44344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__S
timestamp 1688980957
transform 1 0 47380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__S
timestamp 1688980957
transform 1 0 49588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__S
timestamp 1688980957
transform 1 0 48760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__S
timestamp 1688980957
transform 1 0 56580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__S
timestamp 1688980957
transform 1 0 52900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__S
timestamp 1688980957
transform -1 0 58512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__S
timestamp 1688980957
transform 1 0 56488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__S
timestamp 1688980957
transform 1 0 57408 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__S
timestamp 1688980957
transform -1 0 4968 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__S
timestamp 1688980957
transform -1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__S
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__S
timestamp 1688980957
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__S
timestamp 1688980957
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__S
timestamp 1688980957
transform -1 0 16284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__S
timestamp 1688980957
transform 1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__S
timestamp 1688980957
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__S
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__S
timestamp 1688980957
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__S
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__S
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__S
timestamp 1688980957
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__S
timestamp 1688980957
transform 1 0 27508 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__S
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__S
timestamp 1688980957
transform 1 0 29716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__S
timestamp 1688980957
transform 1 0 30452 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__S
timestamp 1688980957
transform 1 0 34868 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__S
timestamp 1688980957
transform 1 0 33488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__S
timestamp 1688980957
transform 1 0 36892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__S
timestamp 1688980957
transform 1 0 36800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__S
timestamp 1688980957
transform 1 0 39928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__S
timestamp 1688980957
transform 1 0 41584 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__S
timestamp 1688980957
transform 1 0 40848 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__S
timestamp 1688980957
transform 1 0 44896 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__S
timestamp 1688980957
transform -1 0 46920 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__S
timestamp 1688980957
transform 1 0 45908 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__S
timestamp 1688980957
transform 1 0 52440 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__S
timestamp 1688980957
transform 1 0 52900 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__S
timestamp 1688980957
transform -1 0 56028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__S
timestamp 1688980957
transform 1 0 53728 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1688980957
transform 1 0 51888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1688980957
transform 1 0 5244 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__S
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__S
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__S
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__S
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__S
timestamp 1688980957
transform 1 0 21620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__S
timestamp 1688980957
transform 1 0 22080 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__S
timestamp 1688980957
transform 1 0 27232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__S
timestamp 1688980957
transform 1 0 24932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__S
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__S
timestamp 1688980957
transform 1 0 30728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__S
timestamp 1688980957
transform 1 0 34960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__S
timestamp 1688980957
transform 1 0 34132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__S
timestamp 1688980957
transform 1 0 36984 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__S
timestamp 1688980957
transform 1 0 36708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1688980957
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__S
timestamp 1688980957
transform 1 0 40388 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__S
timestamp 1688980957
transform 1 0 41952 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__S
timestamp 1688980957
transform 1 0 46552 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__S
timestamp 1688980957
transform -1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__S
timestamp 1688980957
transform 1 0 48576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__S
timestamp 1688980957
transform 1 0 49036 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__S
timestamp 1688980957
transform 1 0 48484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__S
timestamp 1688980957
transform 1 0 53912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__S
timestamp 1688980957
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__S
timestamp 1688980957
transform 1 0 49772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__S
timestamp 1688980957
transform 1 0 54096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__S
timestamp 1688980957
transform -1 0 54372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__S
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__S
timestamp 1688980957
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__S
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__S
timestamp 1688980957
transform -1 0 13064 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__S
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__S
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__S
timestamp 1688980957
transform 1 0 18032 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__S
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__S
timestamp 1688980957
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__S
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__S
timestamp 1688980957
transform 1 0 27140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__S
timestamp 1688980957
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__S
timestamp 1688980957
transform 1 0 29164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__S
timestamp 1688980957
transform 1 0 31004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__S
timestamp 1688980957
transform 1 0 34592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__S
timestamp 1688980957
transform -1 0 34500 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__S
timestamp 1688980957
transform 1 0 36616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__S
timestamp 1688980957
transform 1 0 35236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__S
timestamp 1688980957
transform 1 0 37536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__S
timestamp 1688980957
transform 1 0 40664 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__S
timestamp 1688980957
transform 1 0 43148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__S
timestamp 1688980957
transform 1 0 44620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__S
timestamp 1688980957
transform 1 0 44896 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__S
timestamp 1688980957
transform -1 0 47196 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__S
timestamp 1688980957
transform 1 0 49956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__S
timestamp 1688980957
transform 1 0 50324 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__S
timestamp 1688980957
transform 1 0 55108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__S
timestamp 1688980957
transform 1 0 53176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__S
timestamp 1688980957
transform -1 0 57868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__S
timestamp 1688980957
transform 1 0 55752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__S
timestamp 1688980957
transform -1 0 52348 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A1
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A1
timestamp 1688980957
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A1
timestamp 1688980957
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1688980957
transform 1 0 5336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A1
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B1
timestamp 1688980957
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__S
timestamp 1688980957
transform 1 0 4784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__S
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__S
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__S
timestamp 1688980957
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__S
timestamp 1688980957
transform 1 0 9568 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__S
timestamp 1688980957
transform -1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__S
timestamp 1688980957
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__S
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__S
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__S
timestamp 1688980957
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__S
timestamp 1688980957
transform 1 0 19596 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__S
timestamp 1688980957
transform 1 0 22724 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__S
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__S
timestamp 1688980957
transform 1 0 25760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__S
timestamp 1688980957
transform 1 0 28520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__S
timestamp 1688980957
transform 1 0 28612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__S
timestamp 1688980957
transform 1 0 30820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__S
timestamp 1688980957
transform 1 0 35236 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__S
timestamp 1688980957
transform 1 0 32476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__S
timestamp 1688980957
transform 1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__S
timestamp 1688980957
transform 1 0 35880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__S
timestamp 1688980957
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__S
timestamp 1688980957
transform -1 0 42228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__S
timestamp 1688980957
transform 1 0 40664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__S
timestamp 1688980957
transform 1 0 45172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__S
timestamp 1688980957
transform 1 0 47748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__S
timestamp 1688980957
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__S
timestamp 1688980957
transform 1 0 54372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__S
timestamp 1688980957
transform 1 0 49956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__S
timestamp 1688980957
transform -1 0 55200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__S
timestamp 1688980957
transform 1 0 54004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__S
timestamp 1688980957
transform 1 0 54188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__S
timestamp 1688980957
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__S
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__S
timestamp 1688980957
transform 1 0 10212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__S
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__S
timestamp 1688980957
transform 1 0 11040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__S
timestamp 1688980957
transform 1 0 16468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__S
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__S
timestamp 1688980957
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__S
timestamp 1688980957
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__S
timestamp 1688980957
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__S
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__S
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__S
timestamp 1688980957
transform 1 0 25760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__S
timestamp 1688980957
transform 1 0 25484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__S
timestamp 1688980957
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__S
timestamp 1688980957
transform 1 0 31280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__S
timestamp 1688980957
transform 1 0 33304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__S
timestamp 1688980957
transform 1 0 36984 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__S
timestamp 1688980957
transform 1 0 35788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__S
timestamp 1688980957
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__S
timestamp 1688980957
transform -1 0 38548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__S
timestamp 1688980957
transform 1 0 44436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__S
timestamp 1688980957
transform 1 0 43884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__S
timestamp 1688980957
transform 1 0 42780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S
timestamp 1688980957
transform 1 0 46368 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S
timestamp 1688980957
transform -1 0 50140 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__S
timestamp 1688980957
transform 1 0 50692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__S
timestamp 1688980957
transform -1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S
timestamp 1688980957
transform 1 0 51336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__S
timestamp 1688980957
transform 1 0 58052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__S
timestamp 1688980957
transform 1 0 56120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__S
timestamp 1688980957
transform 1 0 57500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S0
timestamp 1688980957
transform 1 0 7820 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S1
timestamp 1688980957
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S0
timestamp 1688980957
transform 1 0 7912 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S1
timestamp 1688980957
transform -1 0 8740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__S
timestamp 1688980957
transform 1 0 7544 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__S
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S0
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S1
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__S0
timestamp 1688980957
transform -1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__S1
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__S
timestamp 1688980957
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__S
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S0
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S1
timestamp 1688980957
transform 1 0 9292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__S0
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__S1
timestamp 1688980957
transform 1 0 6072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__S
timestamp 1688980957
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__S
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S0
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S1
timestamp 1688980957
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__S0
timestamp 1688980957
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__S1
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__S
timestamp 1688980957
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__S
timestamp 1688980957
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S0
timestamp 1688980957
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S1
timestamp 1688980957
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__S0
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__S1
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__S
timestamp 1688980957
transform 1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S
timestamp 1688980957
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S0
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S1
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__S0
timestamp 1688980957
transform 1 0 14352 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__S1
timestamp 1688980957
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__S
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S
timestamp 1688980957
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S0
timestamp 1688980957
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S1
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S0
timestamp 1688980957
transform 1 0 12880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S1
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__S
timestamp 1688980957
transform 1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S0
timestamp 1688980957
transform 1 0 15088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S1
timestamp 1688980957
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__S0
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__S1
timestamp 1688980957
transform 1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__S
timestamp 1688980957
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__S
timestamp 1688980957
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__S0
timestamp 1688980957
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__S1
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S0
timestamp 1688980957
transform 1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S1
timestamp 1688980957
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__S
timestamp 1688980957
transform 1 0 20792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__S
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S0
timestamp 1688980957
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S1
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S0
timestamp 1688980957
transform 1 0 19872 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S1
timestamp 1688980957
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__S
timestamp 1688980957
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__S
timestamp 1688980957
transform 1 0 17480 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S0
timestamp 1688980957
transform 1 0 21988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S1
timestamp 1688980957
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S0
timestamp 1688980957
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S1
timestamp 1688980957
transform -1 0 21436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp 1688980957
transform 1 0 23828 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__S
timestamp 1688980957
transform 1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S0
timestamp 1688980957
transform 1 0 24840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S1
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S0
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S1
timestamp 1688980957
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp 1688980957
transform 1 0 27416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__S
timestamp 1688980957
transform 1 0 20792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S0
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S1
timestamp 1688980957
transform 1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S0
timestamp 1688980957
transform 1 0 22264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S1
timestamp 1688980957
transform -1 0 24748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__S
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__S
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__S0
timestamp 1688980957
transform -1 0 29256 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__S1
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__S0
timestamp 1688980957
transform -1 0 26864 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__S1
timestamp 1688980957
transform 1 0 27140 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__S
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__S
timestamp 1688980957
transform -1 0 26956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__S0
timestamp 1688980957
transform 1 0 31832 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__S1
timestamp 1688980957
transform 1 0 31648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__S0
timestamp 1688980957
transform -1 0 32660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__S1
timestamp 1688980957
transform 1 0 31648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__S
timestamp 1688980957
transform 1 0 31280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__S
timestamp 1688980957
transform 1 0 29348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__S0
timestamp 1688980957
transform 1 0 34224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__S1
timestamp 1688980957
transform 1 0 33304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__S0
timestamp 1688980957
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__S1
timestamp 1688980957
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__S
timestamp 1688980957
transform 1 0 32476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__S
timestamp 1688980957
transform 1 0 32936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__S0
timestamp 1688980957
transform 1 0 32292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__S1
timestamp 1688980957
transform 1 0 33764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__S0
timestamp 1688980957
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__S1
timestamp 1688980957
transform 1 0 34224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__S
timestamp 1688980957
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__S
timestamp 1688980957
transform 1 0 33488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__S0
timestamp 1688980957
transform 1 0 36800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__S1
timestamp 1688980957
transform 1 0 36800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__S0
timestamp 1688980957
transform 1 0 35328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__S1
timestamp 1688980957
transform 1 0 35696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__S
timestamp 1688980957
transform 1 0 37076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__S
timestamp 1688980957
transform 1 0 35604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S0
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S1
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S0
timestamp 1688980957
transform 1 0 33396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S1
timestamp 1688980957
transform 1 0 33764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__S
timestamp 1688980957
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__S
timestamp 1688980957
transform 1 0 36616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S0
timestamp 1688980957
transform 1 0 38272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S1
timestamp 1688980957
transform 1 0 38640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__S0
timestamp 1688980957
transform 1 0 37444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__S1
timestamp 1688980957
transform 1 0 37444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__S
timestamp 1688980957
transform 1 0 40020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__S
timestamp 1688980957
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__S0
timestamp 1688980957
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__S1
timestamp 1688980957
transform 1 0 37536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__S0
timestamp 1688980957
transform -1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__S1
timestamp 1688980957
transform 1 0 37536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__S
timestamp 1688980957
transform -1 0 39836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__S
timestamp 1688980957
transform 1 0 42320 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__S0
timestamp 1688980957
transform 1 0 42044 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__S1
timestamp 1688980957
transform 1 0 41676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__S0
timestamp 1688980957
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__S1
timestamp 1688980957
transform 1 0 42596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__S
timestamp 1688980957
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__S
timestamp 1688980957
transform 1 0 42044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__S0
timestamp 1688980957
transform 1 0 43332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__S1
timestamp 1688980957
transform 1 0 45356 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__S0
timestamp 1688980957
transform 1 0 45540 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__S1
timestamp 1688980957
transform 1 0 45172 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__S
timestamp 1688980957
transform 1 0 43792 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__S
timestamp 1688980957
transform 1 0 42688 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__S0
timestamp 1688980957
transform 1 0 44528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__S1
timestamp 1688980957
transform 1 0 45172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S0
timestamp 1688980957
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S1
timestamp 1688980957
transform 1 0 44712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__S
timestamp 1688980957
transform 1 0 45172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__S
timestamp 1688980957
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__S0
timestamp 1688980957
transform 1 0 48484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__S1
timestamp 1688980957
transform 1 0 45724 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__S0
timestamp 1688980957
transform 1 0 49312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__S1
timestamp 1688980957
transform 1 0 46368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__S
timestamp 1688980957
transform 1 0 48576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__S
timestamp 1688980957
transform -1 0 47472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__S0
timestamp 1688980957
transform 1 0 48116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__S1
timestamp 1688980957
transform 1 0 49036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__S0
timestamp 1688980957
transform -1 0 48024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__S1
timestamp 1688980957
transform 1 0 48944 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__S
timestamp 1688980957
transform -1 0 49496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__S
timestamp 1688980957
transform 1 0 51060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__S0
timestamp 1688980957
transform 1 0 49680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__S1
timestamp 1688980957
transform 1 0 47380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__S0
timestamp 1688980957
transform 1 0 47288 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__S1
timestamp 1688980957
transform 1 0 48024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__S
timestamp 1688980957
transform 1 0 49496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__S
timestamp 1688980957
transform 1 0 46552 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__S0
timestamp 1688980957
transform 1 0 54924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__S1
timestamp 1688980957
transform 1 0 55936 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__S0
timestamp 1688980957
transform -1 0 52624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__S1
timestamp 1688980957
transform 1 0 53084 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__S
timestamp 1688980957
transform -1 0 54740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__S
timestamp 1688980957
transform 1 0 52440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__S0
timestamp 1688980957
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__S1
timestamp 1688980957
transform 1 0 49036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__S0
timestamp 1688980957
transform 1 0 50324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__S1
timestamp 1688980957
transform 1 0 50416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__S
timestamp 1688980957
transform 1 0 54464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__S
timestamp 1688980957
transform 1 0 53544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__S0
timestamp 1688980957
transform 1 0 55200 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__S1
timestamp 1688980957
transform 1 0 55568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__S0
timestamp 1688980957
transform 1 0 53728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__S1
timestamp 1688980957
transform 1 0 53360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__S
timestamp 1688980957
transform 1 0 51888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__S
timestamp 1688980957
transform 1 0 57592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__S0
timestamp 1688980957
transform 1 0 55476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__S1
timestamp 1688980957
transform 1 0 55844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__S0
timestamp 1688980957
transform 1 0 54188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__S1
timestamp 1688980957
transform 1 0 54556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__S
timestamp 1688980957
transform 1 0 56396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__S
timestamp 1688980957
transform 1 0 57960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__S0
timestamp 1688980957
transform 1 0 55752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__S1
timestamp 1688980957
transform 1 0 56212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__S0
timestamp 1688980957
transform 1 0 51336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__S1
timestamp 1688980957
transform -1 0 51704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__S
timestamp 1688980957
transform 1 0 56580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__S
timestamp 1688980957
transform 1 0 56764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__CLK
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__CLK
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__CLK
timestamp 1688980957
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__CLK
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__CLK
timestamp 1688980957
transform 1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__CLK
timestamp 1688980957
transform 1 0 19688 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__CLK
timestamp 1688980957
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__CLK
timestamp 1688980957
transform -1 0 28520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__CLK
timestamp 1688980957
transform 1 0 34408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__CLK
timestamp 1688980957
transform 1 0 42228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__CLK
timestamp 1688980957
transform -1 0 45632 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__CLK
timestamp 1688980957
transform 1 0 50784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__CLK
timestamp 1688980957
transform 1 0 51612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__CLK
timestamp 1688980957
transform 1 0 11684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__CLK
timestamp 1688980957
transform -1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__CLK
timestamp 1688980957
transform -1 0 17296 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__CLK
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__CLK
timestamp 1688980957
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__CLK
timestamp 1688980957
transform 1 0 23920 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__CLK
timestamp 1688980957
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__CLK
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__CLK
timestamp 1688980957
transform 1 0 27784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__CLK
timestamp 1688980957
transform 1 0 30544 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__CLK
timestamp 1688980957
transform 1 0 31280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__CLK
timestamp 1688980957
transform 1 0 35880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__CLK
timestamp 1688980957
transform 1 0 38916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__CLK
timestamp 1688980957
transform -1 0 35420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__CLK
timestamp 1688980957
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__CLK
timestamp 1688980957
transform 1 0 41124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__CLK
timestamp 1688980957
transform 1 0 45540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__CLK
timestamp 1688980957
transform 1 0 47748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__CLK
timestamp 1688980957
transform 1 0 50876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__CLK
timestamp 1688980957
transform 1 0 53544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__CLK
timestamp 1688980957
transform 1 0 55016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__CLK
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__CLK
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__CLK
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__CLK
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__CLK
timestamp 1688980957
transform 1 0 27416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__CLK
timestamp 1688980957
transform 1 0 27876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__CLK
timestamp 1688980957
transform 1 0 28980 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__CLK
timestamp 1688980957
transform 1 0 32384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__CLK
timestamp 1688980957
transform 1 0 38916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__CLK
timestamp 1688980957
transform -1 0 35052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__CLK
timestamp 1688980957
transform -1 0 42320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__CLK
timestamp 1688980957
transform -1 0 39744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__CLK
timestamp 1688980957
transform 1 0 45172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__CLK
timestamp 1688980957
transform 1 0 50324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__CLK
timestamp 1688980957
transform 1 0 48392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__CLK
timestamp 1688980957
transform 1 0 52532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__CLK
timestamp 1688980957
transform -1 0 58604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__CLK
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__CLK
timestamp 1688980957
transform 1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__CLK
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__CLK
timestamp 1688980957
transform 1 0 21988 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__CLK
timestamp 1688980957
transform 1 0 27784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__CLK
timestamp 1688980957
transform 1 0 28336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__CLK
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__CLK
timestamp 1688980957
transform 1 0 41860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__CLK
timestamp 1688980957
transform 1 0 45908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__CLK
timestamp 1688980957
transform 1 0 50968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__CLK
timestamp 1688980957
transform 1 0 50416 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__CLK
timestamp 1688980957
transform -1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__CLK
timestamp 1688980957
transform 1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__CLK
timestamp 1688980957
transform -1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__CLK
timestamp 1688980957
transform 1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__CLK
timestamp 1688980957
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__CLK
timestamp 1688980957
transform 1 0 21896 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__CLK
timestamp 1688980957
transform 1 0 28704 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__CLK
timestamp 1688980957
transform -1 0 30544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__CLK
timestamp 1688980957
transform 1 0 36708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__CLK
timestamp 1688980957
transform 1 0 43884 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__CLK
timestamp 1688980957
transform 1 0 48484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__CLK
timestamp 1688980957
transform 1 0 51428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__CLK
timestamp 1688980957
transform 1 0 53544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__CLK
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__CLK
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__CLK
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__CLK
timestamp 1688980957
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__CLK
timestamp 1688980957
transform 1 0 22172 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__CLK
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__CLK
timestamp 1688980957
transform 1 0 27968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__CLK
timestamp 1688980957
transform 1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__CLK
timestamp 1688980957
transform 1 0 33580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__CLK
timestamp 1688980957
transform 1 0 37444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__CLK
timestamp 1688980957
transform 1 0 45448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__CLK
timestamp 1688980957
transform 1 0 52624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__CLK
timestamp 1688980957
transform 1 0 55476 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__CLK
timestamp 1688980957
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__CLK
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__CLK
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__CLK
timestamp 1688980957
transform 1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__CLK
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__CLK
timestamp 1688980957
transform -1 0 19136 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__CLK
timestamp 1688980957
transform 1 0 23092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__CLK
timestamp 1688980957
transform 1 0 23920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1688980957
transform 1 0 25300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__CLK
timestamp 1688980957
transform 1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1688980957
transform 1 0 30452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__CLK
timestamp 1688980957
transform 1 0 35788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1688980957
transform 1 0 31924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1688980957
transform 1 0 41308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1688980957
transform 1 0 40664 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1688980957
transform 1 0 45724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1688980957
transform 1 0 45908 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1688980957
transform 1 0 50324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1688980957
transform 1 0 53176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1688980957
transform 1 0 53544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__CLK
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__CLK
timestamp 1688980957
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__CLK
timestamp 1688980957
transform 1 0 21068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__CLK
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__CLK
timestamp 1688980957
transform 1 0 26588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1688980957
transform 1 0 27876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__CLK
timestamp 1688980957
transform 1 0 29716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1688980957
transform 1 0 30360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__CLK
timestamp 1688980957
transform 1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__CLK
timestamp 1688980957
transform 1 0 41584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__CLK
timestamp 1688980957
transform 1 0 37904 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__CLK
timestamp 1688980957
transform 1 0 45172 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__CLK
timestamp 1688980957
transform 1 0 43976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__CLK
timestamp 1688980957
transform 1 0 47472 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__CLK
timestamp 1688980957
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__CLK
timestamp 1688980957
transform 1 0 52256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__CLK
timestamp 1688980957
transform 1 0 56488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__CLK
timestamp 1688980957
transform 1 0 2944 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__CLK
timestamp 1688980957
transform -1 0 1932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__CLK
timestamp 1688980957
transform -1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__CLK
timestamp 1688980957
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1688980957
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1688980957
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1688980957
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1688980957
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1688980957
transform 1 0 24840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1688980957
transform 1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1688980957
transform 1 0 25484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1688980957
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1688980957
transform -1 0 39744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1688980957
transform -1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1688980957
transform -1 0 57316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_wb_clk_i_A
timestamp 1688980957
transform -1 0 20608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 39652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1688980957
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1688980957
transform 1 0 19044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1688980957
transform 1 0 32016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1688980957
transform -1 0 40204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1688980957
transform 1 0 52440 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1688980957
transform 1 0 42596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1688980957
transform 1 0 49588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1688980957
transform -1 0 48392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1688980957
transform 1 0 37812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1688980957
transform 1 0 25208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1688980957
transform 1 0 15088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1688980957
transform 1 0 9476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout70_A
timestamp 1688980957
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout71_A
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_A
timestamp 1688980957
transform 1 0 39468 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout73_A
timestamp 1688980957
transform -1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_A
timestamp 1688980957
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_A
timestamp 1688980957
transform -1 0 35512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout76_A
timestamp 1688980957
transform -1 0 31280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout77_A
timestamp 1688980957
transform 1 0 9108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout78_A
timestamp 1688980957
transform -1 0 32936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout79_A
timestamp 1688980957
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout80_A
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout81_A
timestamp 1688980957
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout82_A
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_A
timestamp 1688980957
transform -1 0 9936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout84_A
timestamp 1688980957
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout85_A
timestamp 1688980957
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout86_A
timestamp 1688980957
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_A
timestamp 1688980957
transform -1 0 8556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout89_A
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_A
timestamp 1688980957
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_A
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_A
timestamp 1688980957
transform 1 0 46184 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout93_A
timestamp 1688980957
transform -1 0 32016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_A
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout96_A
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout97_A
timestamp 1688980957
transform 1 0 48024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout98_A
timestamp 1688980957
transform 1 0 30912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold625_A
timestamp 1688980957
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 20056 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1688980957
transform 1 0 15364 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1688980957
transform 1 0 6532 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1688980957
transform -1 0 21068 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1688980957
transform -1 0 31832 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1688980957
transform 1 0 37904 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1688980957
transform 1 0 49772 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1688980957
transform 1 0 49220 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1688980957
transform 1 0 35420 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1688980957
transform 1 0 25852 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1688980957
transform -1 0 17296 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1688980957
transform -1 0 8188 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout70 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29624 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout71
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout72 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout73
timestamp 1688980957
transform -1 0 7544 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout74
timestamp 1688980957
transform -1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout75
timestamp 1688980957
transform 1 0 35328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout76
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout77
timestamp 1688980957
transform -1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout78
timestamp 1688980957
transform 1 0 32384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout79
timestamp 1688980957
transform 1 0 12696 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout80
timestamp 1688980957
transform 1 0 31924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout81
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout82
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout83
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout84
timestamp 1688980957
transform 1 0 32476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout85
timestamp 1688980957
transform -1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout86
timestamp 1688980957
transform 1 0 33488 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout87
timestamp 1688980957
transform 1 0 8372 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout88
timestamp 1688980957
transform -1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout89
timestamp 1688980957
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout90 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8280 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout91
timestamp 1688980957
transform -1 0 8372 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout92
timestamp 1688980957
transform 1 0 44988 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout93
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout94 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout95
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout96
timestamp 1688980957
transform -1 0 8556 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout97
timestamp 1688980957
transform 1 0 48208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout98
timestamp 1688980957
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout99
timestamp 1688980957
transform 1 0 7636 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_66 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_85 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_173
timestamp 1688980957
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_191
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_480
timestamp 1688980957
transform 1 0 45264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_500
timestamp 1688980957
transform 1 0 47104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1688980957
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1688980957
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1688980957
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_605
timestamp 1688980957
transform 1 0 56764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_615
timestamp 1688980957
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_73
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_119
timestamp 1688980957
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_164
timestamp 1688980957
transform 1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_173
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_209 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_213
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_234
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_238
timestamp 1688980957
transform 1 0 23000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_263
timestamp 1688980957
transform 1 0 25300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_274
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_299
timestamp 1688980957
transform 1 0 28612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_346
timestamp 1688980957
transform 1 0 32936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_380
timestamp 1688980957
transform 1 0 36064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1688980957
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_425
timestamp 1688980957
transform 1 0 40204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1688980957
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_489
timestamp 1688980957
transform 1 0 46092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_494
timestamp 1688980957
transform 1 0 46552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_513
timestamp 1688980957
transform 1 0 48300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_539
timestamp 1688980957
transform 1 0 50692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1688980957
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_561
timestamp 1688980957
transform 1 0 52716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_595
timestamp 1688980957
transform 1 0 55844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_599
timestamp 1688980957
transform 1 0 56212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_21
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_39
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_110
timestamp 1688980957
transform 1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_150
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_299
timestamp 1688980957
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_312
timestamp 1688980957
transform 1 0 29808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_329
timestamp 1688980957
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_416
timestamp 1688980957
transform 1 0 39376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_424
timestamp 1688980957
transform 1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_452
timestamp 1688980957
transform 1 0 42688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_470
timestamp 1688980957
transform 1 0 44344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_474
timestamp 1688980957
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_525
timestamp 1688980957
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_530
timestamp 1688980957
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_533
timestamp 1688980957
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_586
timestamp 1688980957
transform 1 0 55016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_598
timestamp 1688980957
transform 1 0 56120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_624
timestamp 1688980957
transform 1 0 58512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_29
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_70
timestamp 1688980957
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_76
timestamp 1688980957
transform 1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_97
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_108
timestamp 1688980957
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_221
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_254
timestamp 1688980957
transform 1 0 24472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_263
timestamp 1688980957
transform 1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_290
timestamp 1688980957
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_294
timestamp 1688980957
transform 1 0 28152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_387
timestamp 1688980957
transform 1 0 36708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_434
timestamp 1688980957
transform 1 0 41032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_500
timestamp 1688980957
transform 1 0 47104 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_531
timestamp 1688980957
transform 1 0 49956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_541
timestamp 1688980957
transform 1 0 50876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_545
timestamp 1688980957
transform 1 0 51244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_557
timestamp 1688980957
transform 1 0 52348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_599
timestamp 1688980957
transform 1 0 56212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_50
timestamp 1688980957
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_119
timestamp 1688980957
transform 1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_145
timestamp 1688980957
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_148
timestamp 1688980957
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_176
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1688980957
transform 1 0 19596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_274
timestamp 1688980957
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_295
timestamp 1688980957
transform 1 0 28244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_299
timestamp 1688980957
transform 1 0 28612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_339
timestamp 1688980957
transform 1 0 32292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_343
timestamp 1688980957
transform 1 0 32660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_348
timestamp 1688980957
transform 1 0 33120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_384
timestamp 1688980957
transform 1 0 36432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_388
timestamp 1688980957
transform 1 0 36800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_417
timestamp 1688980957
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_425
timestamp 1688980957
transform 1 0 40204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_472
timestamp 1688980957
transform 1 0 44528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_494
timestamp 1688980957
transform 1 0 46552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_498
timestamp 1688980957
transform 1 0 46920 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_510
timestamp 1688980957
transform 1 0 48024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_530
timestamp 1688980957
transform 1 0 49864 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_568
timestamp 1688980957
transform 1 0 53360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_593
timestamp 1688980957
transform 1 0 55660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_597
timestamp 1688980957
transform 1 0 56028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_623
timestamp 1688980957
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_45
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_73
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_130
timestamp 1688980957
transform 1 0 13064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_135
timestamp 1688980957
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_139
timestamp 1688980957
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_151
timestamp 1688980957
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_156
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_196
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_229
timestamp 1688980957
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_257
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_290
timestamp 1688980957
transform 1 0 27784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_294
timestamp 1688980957
transform 1 0 28152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_298
timestamp 1688980957
transform 1 0 28520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_302
timestamp 1688980957
transform 1 0 28888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_306
timestamp 1688980957
transform 1 0 29256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_326
timestamp 1688980957
transform 1 0 31096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_330
timestamp 1688980957
transform 1 0 31464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_334
timestamp 1688980957
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_353
timestamp 1688980957
transform 1 0 33580 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_357
timestamp 1688980957
transform 1 0 33948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_369 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_406
timestamp 1688980957
transform 1 0 38456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_423
timestamp 1688980957
transform 1 0 40020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_427
timestamp 1688980957
transform 1 0 40388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_430
timestamp 1688980957
transform 1 0 40664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_443
timestamp 1688980957
transform 1 0 41860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_474
timestamp 1688980957
transform 1 0 44712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_490
timestamp 1688980957
transform 1 0 46184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_521
timestamp 1688980957
transform 1 0 49036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1688980957
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_561
timestamp 1688980957
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_577
timestamp 1688980957
transform 1 0 54188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_611
timestamp 1688980957
transform 1 0 57316 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_46
timestamp 1688980957
transform 1 0 5336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_52
timestamp 1688980957
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_94
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_116
timestamp 1688980957
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_122
timestamp 1688980957
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_126
timestamp 1688980957
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_149
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_154
timestamp 1688980957
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_166
timestamp 1688980957
transform 1 0 16376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_225
timestamp 1688980957
transform 1 0 21804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 1688980957
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_261
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_288
timestamp 1688980957
transform 1 0 27600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_300 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_313
timestamp 1688980957
transform 1 0 29900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_320
timestamp 1688980957
transform 1 0 30544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_324
timestamp 1688980957
transform 1 0 30912 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_328
timestamp 1688980957
transform 1 0 31280 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_340
timestamp 1688980957
transform 1 0 32384 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_354
timestamp 1688980957
transform 1 0 33672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_393
timestamp 1688980957
transform 1 0 37260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_397
timestamp 1688980957
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_418
timestamp 1688980957
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_425
timestamp 1688980957
transform 1 0 40204 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_431
timestamp 1688980957
transform 1 0 40756 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_440
timestamp 1688980957
transform 1 0 41584 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_463
timestamp 1688980957
transform 1 0 43700 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_472
timestamp 1688980957
transform 1 0 44528 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_481
timestamp 1688980957
transform 1 0 45356 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_489
timestamp 1688980957
transform 1 0 46092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_494
timestamp 1688980957
transform 1 0 46552 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_510
timestamp 1688980957
transform 1 0 48024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_514
timestamp 1688980957
transform 1 0 48392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_518
timestamp 1688980957
transform 1 0 48760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_529
timestamp 1688980957
transform 1 0 49772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_541
timestamp 1688980957
transform 1 0 50876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_550
timestamp 1688980957
transform 1 0 51704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_554
timestamp 1688980957
transform 1 0 52072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_564
timestamp 1688980957
transform 1 0 52992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_568
timestamp 1688980957
transform 1 0 53360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_586
timestamp 1688980957
transform 1 0 55016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_613
timestamp 1688980957
transform 1 0 57500 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_7
timestamp 1688980957
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_10
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_14
timestamp 1688980957
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_18
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_38
timestamp 1688980957
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_44
timestamp 1688980957
transform 1 0 5152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_48
timestamp 1688980957
transform 1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_52
timestamp 1688980957
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_80
timestamp 1688980957
transform 1 0 8464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_90
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_151
timestamp 1688980957
transform 1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_155
timestamp 1688980957
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_178
timestamp 1688980957
transform 1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_208
timestamp 1688980957
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_212
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_216
timestamp 1688980957
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_229
timestamp 1688980957
transform 1 0 22172 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_233
timestamp 1688980957
transform 1 0 22540 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_236
timestamp 1688980957
transform 1 0 22816 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_259
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_263
timestamp 1688980957
transform 1 0 25300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_266
timestamp 1688980957
transform 1 0 25576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_289
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_311
timestamp 1688980957
transform 1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_323
timestamp 1688980957
transform 1 0 30820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_327
timestamp 1688980957
transform 1 0 31188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_331
timestamp 1688980957
transform 1 0 31556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_353
timestamp 1688980957
transform 1 0 33580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_389
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_427
timestamp 1688980957
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_439
timestamp 1688980957
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_457
timestamp 1688980957
transform 1 0 43148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_465
timestamp 1688980957
transform 1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_470
timestamp 1688980957
transform 1 0 44344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_474
timestamp 1688980957
transform 1 0 44712 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_487
timestamp 1688980957
transform 1 0 45908 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_522
timestamp 1688980957
transform 1 0 49128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_549
timestamp 1688980957
transform 1 0 51612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_578
timestamp 1688980957
transform 1 0 54280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_590
timestamp 1688980957
transform 1 0 55384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_599
timestamp 1688980957
transform 1 0 56212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_603
timestamp 1688980957
transform 1 0 56580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_613
timestamp 1688980957
transform 1 0 57500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_38
timestamp 1688980957
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1688980957
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_89
timestamp 1688980957
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_114
timestamp 1688980957
transform 1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_187
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_201
timestamp 1688980957
transform 1 0 19596 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_205
timestamp 1688980957
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_228
timestamp 1688980957
transform 1 0 22080 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_248
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_261
timestamp 1688980957
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_266
timestamp 1688980957
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_286
timestamp 1688980957
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 1688980957
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_390
timestamp 1688980957
transform 1 0 36984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_416
timestamp 1688980957
transform 1 0 39376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_425
timestamp 1688980957
transform 1 0 40204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_450
timestamp 1688980957
transform 1 0 42504 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_456
timestamp 1688980957
transform 1 0 43056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_473
timestamp 1688980957
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_493
timestamp 1688980957
transform 1 0 46460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_537
timestamp 1688980957
transform 1 0 50508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_584
timestamp 1688980957
transform 1 0 54832 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_598
timestamp 1688980957
transform 1 0 56120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_77
timestamp 1688980957
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_103
timestamp 1688980957
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_107
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 1688980957
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_138
timestamp 1688980957
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_163
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_177
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_203
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_258
timestamp 1688980957
transform 1 0 24840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_298
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_325
timestamp 1688980957
transform 1 0 31004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_341
timestamp 1688980957
transform 1 0 32476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_388
timestamp 1688980957
transform 1 0 36800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_420
timestamp 1688980957
transform 1 0 39744 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_442
timestamp 1688980957
transform 1 0 41768 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_446
timestamp 1688980957
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 1688980957
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_514
timestamp 1688980957
transform 1 0 48392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_522
timestamp 1688980957
transform 1 0 49128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_526
timestamp 1688980957
transform 1 0 49496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_556
timestamp 1688980957
transform 1 0 52256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_585
timestamp 1688980957
transform 1 0 54924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_590
timestamp 1688980957
transform 1 0 55384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_613
timestamp 1688980957
transform 1 0 57500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_617
timestamp 1688980957
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_19
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_38
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_71
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_126
timestamp 1688980957
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_136
timestamp 1688980957
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_159
timestamp 1688980957
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_162
timestamp 1688980957
transform 1 0 16008 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_218
timestamp 1688980957
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_223
timestamp 1688980957
transform 1 0 21620 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_231
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_235
timestamp 1688980957
transform 1 0 22724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_248
timestamp 1688980957
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_293
timestamp 1688980957
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_305
timestamp 1688980957
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_335
timestamp 1688980957
transform 1 0 31924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_341
timestamp 1688980957
transform 1 0 32476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_350
timestamp 1688980957
transform 1 0 33304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_354
timestamp 1688980957
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_362
timestamp 1688980957
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_369
timestamp 1688980957
transform 1 0 35052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_398
timestamp 1688980957
transform 1 0 37720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_418
timestamp 1688980957
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_429
timestamp 1688980957
transform 1 0 40572 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_450
timestamp 1688980957
transform 1 0 42504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_464
timestamp 1688980957
transform 1 0 43792 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_473
timestamp 1688980957
transform 1 0 44620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_481
timestamp 1688980957
transform 1 0 45356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_493
timestamp 1688980957
transform 1 0 46460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_497
timestamp 1688980957
transform 1 0 46828 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_522
timestamp 1688980957
transform 1 0 49128 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_530
timestamp 1688980957
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_533
timestamp 1688980957
transform 1 0 50140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_538
timestamp 1688980957
transform 1 0 50600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_558
timestamp 1688980957
transform 1 0 52440 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_562
timestamp 1688980957
transform 1 0 52808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_568
timestamp 1688980957
transform 1 0 53360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_597
timestamp 1688980957
transform 1 0 56028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_601
timestamp 1688980957
transform 1 0 56396 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_620
timestamp 1688980957
transform 1 0 58144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_624
timestamp 1688980957
transform 1 0 58512 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_35
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_40
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_44
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_48
timestamp 1688980957
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_52
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_130
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_138
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_142
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_213
timestamp 1688980957
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_221
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_259
timestamp 1688980957
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_289
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_314
timestamp 1688980957
transform 1 0 29992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_331
timestamp 1688980957
transform 1 0 31556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_365
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_379
timestamp 1688980957
transform 1 0 35972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_388
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_401
timestamp 1688980957
transform 1 0 37996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_406
timestamp 1688980957
transform 1 0 38456 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_410
timestamp 1688980957
transform 1 0 38824 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_422
timestamp 1688980957
transform 1 0 39928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_430
timestamp 1688980957
transform 1 0 40664 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_474
timestamp 1688980957
transform 1 0 44712 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_486
timestamp 1688980957
transform 1 0 45816 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_498
timestamp 1688980957
transform 1 0 46920 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_513
timestamp 1688980957
transform 1 0 48300 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1688980957
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_529
timestamp 1688980957
transform 1 0 49772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_542
timestamp 1688980957
transform 1 0 50968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_546
timestamp 1688980957
transform 1 0 51336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_549
timestamp 1688980957
transform 1 0 51612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_554
timestamp 1688980957
transform 1 0 52072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_558
timestamp 1688980957
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_561
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_565
timestamp 1688980957
transform 1 0 53084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_570
timestamp 1688980957
transform 1 0 53544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_590
timestamp 1688980957
transform 1 0 55384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1688980957
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_39
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_51
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_57
timestamp 1688980957
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_60
timestamp 1688980957
transform 1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_64
timestamp 1688980957
transform 1 0 6992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_110
timestamp 1688980957
transform 1 0 11224 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_115
timestamp 1688980957
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_119
timestamp 1688980957
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_123
timestamp 1688980957
transform 1 0 12420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_135
timestamp 1688980957
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_192
timestamp 1688980957
transform 1 0 18768 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_210
timestamp 1688980957
transform 1 0 20424 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_222
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_234
timestamp 1688980957
transform 1 0 22632 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_237
timestamp 1688980957
transform 1 0 22908 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1688980957
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_284
timestamp 1688980957
transform 1 0 27232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_288
timestamp 1688980957
transform 1 0 27600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_292
timestamp 1688980957
transform 1 0 27968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_295
timestamp 1688980957
transform 1 0 28244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_313
timestamp 1688980957
transform 1 0 29900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_332
timestamp 1688980957
transform 1 0 31648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_336
timestamp 1688980957
transform 1 0 32016 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_385
timestamp 1688980957
transform 1 0 36524 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_393
timestamp 1688980957
transform 1 0 37260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_412
timestamp 1688980957
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_416
timestamp 1688980957
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_429
timestamp 1688980957
transform 1 0 40572 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_441
timestamp 1688980957
transform 1 0 41676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_449
timestamp 1688980957
transform 1 0 42412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_453
timestamp 1688980957
transform 1 0 42780 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_462
timestamp 1688980957
transform 1 0 43608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_468
timestamp 1688980957
transform 1 0 44160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_472
timestamp 1688980957
transform 1 0 44528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_481
timestamp 1688980957
transform 1 0 45356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_487
timestamp 1688980957
transform 1 0 45908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_491
timestamp 1688980957
transform 1 0 46276 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_494
timestamp 1688980957
transform 1 0 46552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_502
timestamp 1688980957
transform 1 0 47288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_514
timestamp 1688980957
transform 1 0 48392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_525
timestamp 1688980957
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_529
timestamp 1688980957
transform 1 0 49772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_533
timestamp 1688980957
transform 1 0 50140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_537
timestamp 1688980957
transform 1 0 50508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_556
timestamp 1688980957
transform 1 0 52256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_561
timestamp 1688980957
transform 1 0 52716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_565
timestamp 1688980957
transform 1 0 53084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_569
timestamp 1688980957
transform 1 0 53452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_572
timestamp 1688980957
transform 1 0 53728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_577
timestamp 1688980957
transform 1 0 54188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_581
timestamp 1688980957
transform 1 0 54556 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_584
timestamp 1688980957
transform 1 0 54832 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_597
timestamp 1688980957
transform 1 0 56028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_623
timestamp 1688980957
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_25
timestamp 1688980957
transform 1 0 3404 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_64
timestamp 1688980957
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_68
timestamp 1688980957
transform 1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_87
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_91
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_146
timestamp 1688980957
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_194
timestamp 1688980957
transform 1 0 18952 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_256
timestamp 1688980957
transform 1 0 24656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1688980957
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_286
timestamp 1688980957
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_290
timestamp 1688980957
transform 1 0 27784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_330
timestamp 1688980957
transform 1 0 31464 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_334
timestamp 1688980957
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_356
timestamp 1688980957
transform 1 0 33856 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_360
timestamp 1688980957
transform 1 0 34224 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_388
timestamp 1688980957
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_406
timestamp 1688980957
transform 1 0 38456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_438
timestamp 1688980957
transform 1 0 41400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_442
timestamp 1688980957
transform 1 0 41768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_446
timestamp 1688980957
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_492
timestamp 1688980957
transform 1 0 46368 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1688980957
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_557
timestamp 1688980957
transform 1 0 52348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_570
timestamp 1688980957
transform 1 0 53544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_605
timestamp 1688980957
transform 1 0 56764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 1688980957
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_46
timestamp 1688980957
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_64
timestamp 1688980957
transform 1 0 6992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1688980957
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_89
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_108
timestamp 1688980957
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_119
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_175
timestamp 1688980957
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_179
timestamp 1688980957
transform 1 0 17572 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_208
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_212
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_231
timestamp 1688980957
transform 1 0 22356 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_248
timestamp 1688980957
transform 1 0 23920 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_284
timestamp 1688980957
transform 1 0 27232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_288
timestamp 1688980957
transform 1 0 27600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_327
timestamp 1688980957
transform 1 0 31188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_362
timestamp 1688980957
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_386
timestamp 1688980957
transform 1 0 36616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_390
timestamp 1688980957
transform 1 0 36984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_416
timestamp 1688980957
transform 1 0 39376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_454
timestamp 1688980957
transform 1 0 42872 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_486
timestamp 1688980957
transform 1 0 45816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_533
timestamp 1688980957
transform 1 0 50140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_537
timestamp 1688980957
transform 1 0 50508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_586
timestamp 1688980957
transform 1 0 55016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_621
timestamp 1688980957
transform 1 0 58236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_11
timestamp 1688980957
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_37
timestamp 1688980957
transform 1 0 4508 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_74
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_86
timestamp 1688980957
transform 1 0 9016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_96
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1688980957
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_145
timestamp 1688980957
transform 1 0 14444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1688980957
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_173
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_185
timestamp 1688980957
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_214
timestamp 1688980957
transform 1 0 20792 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_234
timestamp 1688980957
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_257
timestamp 1688980957
transform 1 0 24748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_275
timestamp 1688980957
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_297
timestamp 1688980957
transform 1 0 28428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_325
timestamp 1688980957
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_333
timestamp 1688980957
transform 1 0 31740 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_364
timestamp 1688980957
transform 1 0 34592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_386
timestamp 1688980957
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_444
timestamp 1688980957
transform 1 0 41952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_465
timestamp 1688980957
transform 1 0 43884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_483
timestamp 1688980957
transform 1 0 45540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_487
timestamp 1688980957
transform 1 0 45908 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_513
timestamp 1688980957
transform 1 0 48300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_517
timestamp 1688980957
transform 1 0 48668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_557
timestamp 1688980957
transform 1 0 52348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_614
timestamp 1688980957
transform 1 0 57592 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_74
timestamp 1688980957
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_89
timestamp 1688980957
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_92
timestamp 1688980957
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_151
timestamp 1688980957
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_175
timestamp 1688980957
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_179
timestamp 1688980957
transform 1 0 17572 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_203
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_216
timestamp 1688980957
transform 1 0 20976 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_222
timestamp 1688980957
transform 1 0 21528 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_225
timestamp 1688980957
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_235
timestamp 1688980957
transform 1 0 22724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_243
timestamp 1688980957
transform 1 0 23460 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_247
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_281
timestamp 1688980957
transform 1 0 26956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_293
timestamp 1688980957
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_306
timestamp 1688980957
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_313
timestamp 1688980957
transform 1 0 29900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_325
timestamp 1688980957
transform 1 0 31004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_337
timestamp 1688980957
transform 1 0 32108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_369
timestamp 1688980957
transform 1 0 35052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_400
timestamp 1688980957
transform 1 0 37904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1688980957
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_445
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_453
timestamp 1688980957
transform 1 0 42780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_473
timestamp 1688980957
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_501
timestamp 1688980957
transform 1 0 47196 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_506
timestamp 1688980957
transform 1 0 47656 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_518
timestamp 1688980957
transform 1 0 48760 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 1688980957
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 1688980957
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 1688980957
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 1688980957
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_589
timestamp 1688980957
transform 1 0 55292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_593
timestamp 1688980957
transform 1 0 55660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_597
timestamp 1688980957
transform 1 0 56028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_612
timestamp 1688980957
transform 1 0 57408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_616
timestamp 1688980957
transform 1 0 57776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_620
timestamp 1688980957
transform 1 0 58144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_624
timestamp 1688980957
transform 1 0 58512 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_19
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_25
timestamp 1688980957
transform 1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_30
timestamp 1688980957
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_34
timestamp 1688980957
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_46
timestamp 1688980957
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 1688980957
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_67
timestamp 1688980957
transform 1 0 7268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_79
timestamp 1688980957
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_83
timestamp 1688980957
transform 1 0 8740 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_134
timestamp 1688980957
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_148
timestamp 1688980957
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_159
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_173
timestamp 1688980957
transform 1 0 17020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_185
timestamp 1688980957
transform 1 0 18124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_197
timestamp 1688980957
transform 1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_202
timestamp 1688980957
transform 1 0 19688 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_246
timestamp 1688980957
transform 1 0 23736 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_258
timestamp 1688980957
transform 1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_271
timestamp 1688980957
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_322
timestamp 1688980957
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_362
timestamp 1688980957
transform 1 0 34408 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_366
timestamp 1688980957
transform 1 0 34776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_370
timestamp 1688980957
transform 1 0 35144 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_374
timestamp 1688980957
transform 1 0 35512 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_379
timestamp 1688980957
transform 1 0 35972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_413
timestamp 1688980957
transform 1 0 39100 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_421
timestamp 1688980957
transform 1 0 39836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_441
timestamp 1688980957
transform 1 0 41676 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_445
timestamp 1688980957
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_449
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_453
timestamp 1688980957
transform 1 0 42780 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_459
timestamp 1688980957
transform 1 0 43332 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_471
timestamp 1688980957
transform 1 0 44436 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_485
timestamp 1688980957
transform 1 0 45724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_489
timestamp 1688980957
transform 1 0 46092 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_498
timestamp 1688980957
transform 1 0 46920 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 1688980957
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_517
timestamp 1688980957
transform 1 0 48668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_523
timestamp 1688980957
transform 1 0 49220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_528
timestamp 1688980957
transform 1 0 49680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_536
timestamp 1688980957
transform 1 0 50416 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_539
timestamp 1688980957
transform 1 0 50692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_543
timestamp 1688980957
transform 1 0 51060 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_548
timestamp 1688980957
transform 1 0 51520 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_565
timestamp 1688980957
transform 1 0 53084 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_577
timestamp 1688980957
transform 1 0 54188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_589
timestamp 1688980957
transform 1 0 55292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_593
timestamp 1688980957
transform 1 0 55660 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_596
timestamp 1688980957
transform 1 0 55936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_600
timestamp 1688980957
transform 1 0 56304 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_604
timestamp 1688980957
transform 1 0 56672 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_614
timestamp 1688980957
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_34
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_38
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_52
timestamp 1688980957
transform 1 0 5888 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_71
timestamp 1688980957
transform 1 0 7636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_102
timestamp 1688980957
transform 1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_134
timestamp 1688980957
transform 1 0 13432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_150
timestamp 1688980957
transform 1 0 14904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_170
timestamp 1688980957
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_181
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_236
timestamp 1688980957
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_262
timestamp 1688980957
transform 1 0 25208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_282
timestamp 1688980957
transform 1 0 27048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_286
timestamp 1688980957
transform 1 0 27416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_360
timestamp 1688980957
transform 1 0 34224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_373
timestamp 1688980957
transform 1 0 35420 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_382
timestamp 1688980957
transform 1 0 36248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_386
timestamp 1688980957
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_409
timestamp 1688980957
transform 1 0 38732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_413
timestamp 1688980957
transform 1 0 39100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_417
timestamp 1688980957
transform 1 0 39468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 1688980957
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_508
timestamp 1688980957
transform 1 0 47840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_524
timestamp 1688980957
transform 1 0 49312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_528
timestamp 1688980957
transform 1 0 49680 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_533
timestamp 1688980957
transform 1 0 50140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_541
timestamp 1688980957
transform 1 0 50876 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_544
timestamp 1688980957
transform 1 0 51152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_548
timestamp 1688980957
transform 1 0 51520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_575
timestamp 1688980957
transform 1 0 54004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_579
timestamp 1688980957
transform 1 0 54372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_583
timestamp 1688980957
transform 1 0 54740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 1688980957
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_589
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_593
timestamp 1688980957
transform 1 0 55660 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_620
timestamp 1688980957
transform 1 0 58144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_624
timestamp 1688980957
transform 1 0 58512 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_31
timestamp 1688980957
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_43
timestamp 1688980957
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_71
timestamp 1688980957
transform 1 0 7636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_98
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_138
timestamp 1688980957
transform 1 0 13800 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_144
timestamp 1688980957
transform 1 0 14352 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_173
timestamp 1688980957
transform 1 0 17020 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_192
timestamp 1688980957
transform 1 0 18768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_196
timestamp 1688980957
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_218
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_242
timestamp 1688980957
transform 1 0 23368 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_262
timestamp 1688980957
transform 1 0 25208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_290
timestamp 1688980957
transform 1 0 27784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_314
timestamp 1688980957
transform 1 0 29992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_386
timestamp 1688980957
transform 1 0 36616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_390
timestamp 1688980957
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_417
timestamp 1688980957
transform 1 0 39468 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_445
timestamp 1688980957
transform 1 0 42044 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_453
timestamp 1688980957
transform 1 0 42780 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_480
timestamp 1688980957
transform 1 0 45264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_484
timestamp 1688980957
transform 1 0 45632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_501
timestamp 1688980957
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_505
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_509
timestamp 1688980957
transform 1 0 47932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_537
timestamp 1688980957
transform 1 0 50508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_541
timestamp 1688980957
transform 1 0 50876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_570
timestamp 1688980957
transform 1 0 53544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_574
timestamp 1688980957
transform 1 0 53912 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_613
timestamp 1688980957
transform 1 0 57500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_617
timestamp 1688980957
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_20
timestamp 1688980957
transform 1 0 2944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_33
timestamp 1688980957
transform 1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_40
timestamp 1688980957
transform 1 0 4784 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_48
timestamp 1688980957
transform 1 0 5520 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_62
timestamp 1688980957
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_66
timestamp 1688980957
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_70
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_111
timestamp 1688980957
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_115
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_122
timestamp 1688980957
transform 1 0 12328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_126
timestamp 1688980957
transform 1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_130
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_134
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_163
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_205
timestamp 1688980957
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_218
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_236
timestamp 1688980957
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_240
timestamp 1688980957
transform 1 0 23184 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_300
timestamp 1688980957
transform 1 0 28704 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_329
timestamp 1688980957
transform 1 0 31372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_359
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_375
timestamp 1688980957
transform 1 0 35604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_414
timestamp 1688980957
transform 1 0 39192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_418
timestamp 1688980957
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_474
timestamp 1688980957
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_481
timestamp 1688980957
transform 1 0 45356 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_500
timestamp 1688980957
transform 1 0 47104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_526
timestamp 1688980957
transform 1 0 49496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_530
timestamp 1688980957
transform 1 0 49864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_550
timestamp 1688980957
transform 1 0 51704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_568
timestamp 1688980957
transform 1 0 53360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_605
timestamp 1688980957
transform 1 0 56764 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_622
timestamp 1688980957
transform 1 0 58328 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_26
timestamp 1688980957
transform 1 0 3496 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 1688980957
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_47
timestamp 1688980957
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_61
timestamp 1688980957
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_78
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_83
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_87
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_108
timestamp 1688980957
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_117
timestamp 1688980957
transform 1 0 11868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_140
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_150
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_163
timestamp 1688980957
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_202
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_215
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_266
timestamp 1688980957
transform 1 0 25576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_270
timestamp 1688980957
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_322
timestamp 1688980957
transform 1 0 30728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_360
timestamp 1688980957
transform 1 0 34224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_386
timestamp 1688980957
transform 1 0 36616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_390
timestamp 1688980957
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_419
timestamp 1688980957
transform 1 0 39652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_441
timestamp 1688980957
transform 1 0 41676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_445
timestamp 1688980957
transform 1 0 42044 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_485
timestamp 1688980957
transform 1 0 45724 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_489
timestamp 1688980957
transform 1 0 46092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_500
timestamp 1688980957
transform 1 0 47104 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_513
timestamp 1688980957
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_540
timestamp 1688980957
transform 1 0 50784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_556
timestamp 1688980957
transform 1 0 52256 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_577
timestamp 1688980957
transform 1 0 54188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_605
timestamp 1688980957
transform 1 0 56764 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_38
timestamp 1688980957
transform 1 0 4600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_50
timestamp 1688980957
transform 1 0 5704 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_56
timestamp 1688980957
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_59
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_68
timestamp 1688980957
transform 1 0 7360 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_89
timestamp 1688980957
transform 1 0 9292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_117
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_136
timestamp 1688980957
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_151
timestamp 1688980957
transform 1 0 14996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_160
timestamp 1688980957
transform 1 0 15824 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_169
timestamp 1688980957
transform 1 0 16652 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_180
timestamp 1688980957
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_191
timestamp 1688980957
transform 1 0 18676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_215
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_219
timestamp 1688980957
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_261
timestamp 1688980957
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_270
timestamp 1688980957
transform 1 0 25944 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_287
timestamp 1688980957
transform 1 0 27508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_291
timestamp 1688980957
transform 1 0 27876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_305
timestamp 1688980957
transform 1 0 29164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_318
timestamp 1688980957
transform 1 0 30360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_322
timestamp 1688980957
transform 1 0 30728 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_326
timestamp 1688980957
transform 1 0 31096 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_338
timestamp 1688980957
transform 1 0 32200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_342
timestamp 1688980957
transform 1 0 32568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_346
timestamp 1688980957
transform 1 0 32936 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_352
timestamp 1688980957
transform 1 0 33488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_355
timestamp 1688980957
transform 1 0 33764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_369
timestamp 1688980957
transform 1 0 35052 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_373
timestamp 1688980957
transform 1 0 35420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_388
timestamp 1688980957
transform 1 0 36800 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_393
timestamp 1688980957
transform 1 0 37260 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_397
timestamp 1688980957
transform 1 0 37628 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_408
timestamp 1688980957
transform 1 0 38640 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_439
timestamp 1688980957
transform 1 0 41492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_443
timestamp 1688980957
transform 1 0 41860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_447
timestamp 1688980957
transform 1 0 42228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_457
timestamp 1688980957
transform 1 0 43148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_469
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_473
timestamp 1688980957
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_477
timestamp 1688980957
transform 1 0 44988 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_481
timestamp 1688980957
transform 1 0 45356 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_497
timestamp 1688980957
transform 1 0 46828 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_509
timestamp 1688980957
transform 1 0 47932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_513
timestamp 1688980957
transform 1 0 48300 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_516
timestamp 1688980957
transform 1 0 48576 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_529
timestamp 1688980957
transform 1 0 49772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_533
timestamp 1688980957
transform 1 0 50140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_571
timestamp 1688980957
transform 1 0 53636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_575
timestamp 1688980957
transform 1 0 54004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_586
timestamp 1688980957
transform 1 0 55016 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 1688980957
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_601
timestamp 1688980957
transform 1 0 56396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_607
timestamp 1688980957
transform 1 0 56948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_611
timestamp 1688980957
transform 1 0 57316 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_40
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_48
timestamp 1688980957
transform 1 0 5520 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_52
timestamp 1688980957
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_94
timestamp 1688980957
transform 1 0 9752 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_151
timestamp 1688980957
transform 1 0 14996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_165
timestamp 1688980957
transform 1 0 16284 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_189
timestamp 1688980957
transform 1 0 18492 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_197
timestamp 1688980957
transform 1 0 19228 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_219
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_231
timestamp 1688980957
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_240
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_244
timestamp 1688980957
transform 1 0 23552 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_256
timestamp 1688980957
transform 1 0 24656 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_268
timestamp 1688980957
transform 1 0 25760 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_289
timestamp 1688980957
transform 1 0 27692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_324
timestamp 1688980957
transform 1 0 30912 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_328
timestamp 1688980957
transform 1 0 31280 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_348
timestamp 1688980957
transform 1 0 33120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_352
timestamp 1688980957
transform 1 0 33488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_370
timestamp 1688980957
transform 1 0 35144 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_374
timestamp 1688980957
transform 1 0 35512 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_378
timestamp 1688980957
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_390
timestamp 1688980957
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_417
timestamp 1688980957
transform 1 0 39468 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_445
timestamp 1688980957
transform 1 0 42044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_478
timestamp 1688980957
transform 1 0 45080 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_486
timestamp 1688980957
transform 1 0 45816 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_497
timestamp 1688980957
transform 1 0 46828 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_501
timestamp 1688980957
transform 1 0 47196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_513
timestamp 1688980957
transform 1 0 48300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_517
timestamp 1688980957
transform 1 0 48668 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_536
timestamp 1688980957
transform 1 0 50416 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_550
timestamp 1688980957
transform 1 0 51704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_554
timestamp 1688980957
transform 1 0 52072 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_561
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_573
timestamp 1688980957
transform 1 0 53820 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_587
timestamp 1688980957
transform 1 0 55108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_599
timestamp 1688980957
transform 1 0 56212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_611
timestamp 1688980957
transform 1 0 57316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_614
timestamp 1688980957
transform 1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_617
timestamp 1688980957
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_24
timestamp 1688980957
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_42
timestamp 1688980957
transform 1 0 4968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_93
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_96
timestamp 1688980957
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_118
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_135
timestamp 1688980957
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 1688980957
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_179
timestamp 1688980957
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_183
timestamp 1688980957
transform 1 0 17940 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_186
timestamp 1688980957
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_192
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_213
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_257
timestamp 1688980957
transform 1 0 24748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_269
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_286
timestamp 1688980957
transform 1 0 27416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_358
timestamp 1688980957
transform 1 0 34040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_362
timestamp 1688980957
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_382
timestamp 1688980957
transform 1 0 36248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_388
timestamp 1688980957
transform 1 0 36800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_413
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_417
timestamp 1688980957
transform 1 0 39468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_447
timestamp 1688980957
transform 1 0 42228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_485
timestamp 1688980957
transform 1 0 45724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_489
timestamp 1688980957
transform 1 0 46092 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_508
timestamp 1688980957
transform 1 0 47840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_512
timestamp 1688980957
transform 1 0 48208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_530
timestamp 1688980957
transform 1 0 49864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_537
timestamp 1688980957
transform 1 0 50508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_545
timestamp 1688980957
transform 1 0 51244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_548
timestamp 1688980957
transform 1 0 51520 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_571
timestamp 1688980957
transform 1 0 53636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_597
timestamp 1688980957
transform 1 0 56028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_614
timestamp 1688980957
transform 1 0 57592 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_31
timestamp 1688980957
transform 1 0 3956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_49
timestamp 1688980957
transform 1 0 5612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_87
timestamp 1688980957
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_91
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_95
timestamp 1688980957
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_99
timestamp 1688980957
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 1688980957
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_117
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_139
timestamp 1688980957
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_198
timestamp 1688980957
transform 1 0 19320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_254
timestamp 1688980957
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_260
timestamp 1688980957
transform 1 0 25024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_264
timestamp 1688980957
transform 1 0 25392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_267
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_297
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_314
timestamp 1688980957
transform 1 0 29992 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_426
timestamp 1688980957
transform 1 0 40296 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_444
timestamp 1688980957
transform 1 0 41952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_457
timestamp 1688980957
transform 1 0 43148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_477
timestamp 1688980957
transform 1 0 44988 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_481
timestamp 1688980957
transform 1 0 45356 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_500
timestamp 1688980957
transform 1 0 47104 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_534
timestamp 1688980957
transform 1 0 50232 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_570
timestamp 1688980957
transform 1 0 53544 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_574
timestamp 1688980957
transform 1 0 53912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_592
timestamp 1688980957
transform 1 0 55568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_596
timestamp 1688980957
transform 1 0 55936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_613
timestamp 1688980957
transform 1 0 57500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_46
timestamp 1688980957
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_58
timestamp 1688980957
transform 1 0 6440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_89
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_100
timestamp 1688980957
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_112
timestamp 1688980957
transform 1 0 11408 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_124
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1688980957
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_162
timestamp 1688980957
transform 1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_214
timestamp 1688980957
transform 1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_234
timestamp 1688980957
transform 1 0 22632 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_262
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_281
timestamp 1688980957
transform 1 0 26956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_293
timestamp 1688980957
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_299
timestamp 1688980957
transform 1 0 28612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_317
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_327
timestamp 1688980957
transform 1 0 31188 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_338
timestamp 1688980957
transform 1 0 32200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_361
timestamp 1688980957
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_413
timestamp 1688980957
transform 1 0 39100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_417
timestamp 1688980957
transform 1 0 39468 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_446
timestamp 1688980957
transform 1 0 42136 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_450
timestamp 1688980957
transform 1 0 42504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_470
timestamp 1688980957
transform 1 0 44344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_474
timestamp 1688980957
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_477
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_481
timestamp 1688980957
transform 1 0 45356 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_575
timestamp 1688980957
transform 1 0 54004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_589
timestamp 1688980957
transform 1 0 55292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_623
timestamp 1688980957
transform 1 0 58420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_11
timestamp 1688980957
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_38
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_82
timestamp 1688980957
transform 1 0 8648 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_117
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_131
timestamp 1688980957
transform 1 0 13156 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_143
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_147
timestamp 1688980957
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_150
timestamp 1688980957
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_163
timestamp 1688980957
transform 1 0 16100 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_185
timestamp 1688980957
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_195
timestamp 1688980957
transform 1 0 19044 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_221
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_233
timestamp 1688980957
transform 1 0 22540 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_241
timestamp 1688980957
transform 1 0 23276 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_266
timestamp 1688980957
transform 1 0 25576 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_270
timestamp 1688980957
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_292
timestamp 1688980957
transform 1 0 27968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_301
timestamp 1688980957
transform 1 0 28796 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_325
timestamp 1688980957
transform 1 0 31004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_333
timestamp 1688980957
transform 1 0 31740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_347
timestamp 1688980957
transform 1 0 33028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_352
timestamp 1688980957
transform 1 0 33488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_356
timestamp 1688980957
transform 1 0 33856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_360
timestamp 1688980957
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_364
timestamp 1688980957
transform 1 0 34592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_385
timestamp 1688980957
transform 1 0 36524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_389
timestamp 1688980957
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_409
timestamp 1688980957
transform 1 0 38732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_428
timestamp 1688980957
transform 1 0 40480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_438
timestamp 1688980957
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_446
timestamp 1688980957
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_469
timestamp 1688980957
transform 1 0 44252 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_481
timestamp 1688980957
transform 1 0 45356 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_493
timestamp 1688980957
transform 1 0 46460 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_501
timestamp 1688980957
transform 1 0 47196 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_505
timestamp 1688980957
transform 1 0 47564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_543
timestamp 1688980957
transform 1 0 51060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_578
timestamp 1688980957
transform 1 0 54280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_597
timestamp 1688980957
transform 1 0 56028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_601
timestamp 1688980957
transform 1 0 56396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_611
timestamp 1688980957
transform 1 0 57316 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 1688980957
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_37
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_49
timestamp 1688980957
transform 1 0 5612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_61
timestamp 1688980957
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_71
timestamp 1688980957
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_75
timestamp 1688980957
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_103
timestamp 1688980957
transform 1 0 10580 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_107
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_135
timestamp 1688980957
transform 1 0 13524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_149
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_168
timestamp 1688980957
transform 1 0 16560 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_180
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_184
timestamp 1688980957
transform 1 0 18032 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_187
timestamp 1688980957
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_205
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_214
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_218
timestamp 1688980957
transform 1 0 21160 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_231
timestamp 1688980957
transform 1 0 22356 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_235
timestamp 1688980957
transform 1 0 22724 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_247
timestamp 1688980957
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_261
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_274
timestamp 1688980957
transform 1 0 26312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_278
timestamp 1688980957
transform 1 0 26680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 1688980957
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_313
timestamp 1688980957
transform 1 0 29900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_334
timestamp 1688980957
transform 1 0 31832 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_338
timestamp 1688980957
transform 1 0 32200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_358
timestamp 1688980957
transform 1 0 34040 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_385
timestamp 1688980957
transform 1 0 36524 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_393
timestamp 1688980957
transform 1 0 37260 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_397
timestamp 1688980957
transform 1 0 37628 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_409
timestamp 1688980957
transform 1 0 38732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_417
timestamp 1688980957
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_461
timestamp 1688980957
transform 1 0 43516 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 1688980957
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_489
timestamp 1688980957
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_501
timestamp 1688980957
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_513
timestamp 1688980957
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_525
timestamp 1688980957
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 1688980957
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_533
timestamp 1688980957
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_545
timestamp 1688980957
transform 1 0 51244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_553
timestamp 1688980957
transform 1 0 51980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_581
timestamp 1688980957
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_587
timestamp 1688980957
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_605
timestamp 1688980957
transform 1 0 56764 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_622
timestamp 1688980957
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_85
timestamp 1688980957
transform 1 0 8924 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_143
timestamp 1688980957
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_155
timestamp 1688980957
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1688980957
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_242
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_248
timestamp 1688980957
transform 1 0 23920 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_251
timestamp 1688980957
transform 1 0 24196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_277
timestamp 1688980957
transform 1 0 26588 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_302
timestamp 1688980957
transform 1 0 28888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_306
timestamp 1688980957
transform 1 0 29256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_334
timestamp 1688980957
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_370
timestamp 1688980957
transform 1 0 35144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_378
timestamp 1688980957
transform 1 0 35880 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_387
timestamp 1688980957
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1688980957
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_401
timestamp 1688980957
transform 1 0 37996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_405
timestamp 1688980957
transform 1 0 38364 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_414
timestamp 1688980957
transform 1 0 39192 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_423
timestamp 1688980957
transform 1 0 40020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_427
timestamp 1688980957
transform 1 0 40388 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_458
timestamp 1688980957
transform 1 0 43240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_462
timestamp 1688980957
transform 1 0 43608 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_479
timestamp 1688980957
transform 1 0 45172 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_483
timestamp 1688980957
transform 1 0 45540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_495
timestamp 1688980957
transform 1 0 46644 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_503
timestamp 1688980957
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_505
timestamp 1688980957
transform 1 0 47564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_509
timestamp 1688980957
transform 1 0 47932 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_513
timestamp 1688980957
transform 1 0 48300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_525
timestamp 1688980957
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_538
timestamp 1688980957
transform 1 0 50600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_550
timestamp 1688980957
transform 1 0 51704 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_577
timestamp 1688980957
transform 1 0 54188 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_581
timestamp 1688980957
transform 1 0 54556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_593
timestamp 1688980957
transform 1 0 55660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_605
timestamp 1688980957
transform 1 0 56764 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_613
timestamp 1688980957
transform 1 0 57500 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_19
timestamp 1688980957
transform 1 0 2852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_38
timestamp 1688980957
transform 1 0 4600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_42
timestamp 1688980957
transform 1 0 4968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_89
timestamp 1688980957
transform 1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_104
timestamp 1688980957
transform 1 0 10672 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_147
timestamp 1688980957
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_156
timestamp 1688980957
transform 1 0 15456 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_160
timestamp 1688980957
transform 1 0 15824 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_166
timestamp 1688980957
transform 1 0 16376 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_186
timestamp 1688980957
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_213
timestamp 1688980957
transform 1 0 20700 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_249
timestamp 1688980957
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_257
timestamp 1688980957
transform 1 0 24748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_299
timestamp 1688980957
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_326
timestamp 1688980957
transform 1 0 31096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_330
timestamp 1688980957
transform 1 0 31464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_373
timestamp 1688980957
transform 1 0 35420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_377
timestamp 1688980957
transform 1 0 35788 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_398
timestamp 1688980957
transform 1 0 37720 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_418
timestamp 1688980957
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_438
timestamp 1688980957
transform 1 0 41400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_450
timestamp 1688980957
transform 1 0 42504 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 1688980957
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_488
timestamp 1688980957
transform 1 0 46000 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_492
timestamp 1688980957
transform 1 0 46368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_519
timestamp 1688980957
transform 1 0 48852 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_523
timestamp 1688980957
transform 1 0 49220 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_549
timestamp 1688980957
transform 1 0 51612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_585
timestamp 1688980957
transform 1 0 54924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_597
timestamp 1688980957
transform 1 0 56028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_614
timestamp 1688980957
transform 1 0 57592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_623
timestamp 1688980957
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_89
timestamp 1688980957
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_101
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_127
timestamp 1688980957
transform 1 0 12788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_131
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_163
timestamp 1688980957
transform 1 0 16100 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_212
timestamp 1688980957
transform 1 0 20608 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 1688980957
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_255
timestamp 1688980957
transform 1 0 24564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 1688980957
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_291
timestamp 1688980957
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_295
timestamp 1688980957
transform 1 0 28244 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_307
timestamp 1688980957
transform 1 0 29348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_326
timestamp 1688980957
transform 1 0 31096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_341
timestamp 1688980957
transform 1 0 32476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_367
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_373
timestamp 1688980957
transform 1 0 35420 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_390
timestamp 1688980957
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_397
timestamp 1688980957
transform 1 0 37628 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_443
timestamp 1688980957
transform 1 0 41860 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 1688980957
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_457
timestamp 1688980957
transform 1 0 43148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_493
timestamp 1688980957
transform 1 0 46460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_551
timestamp 1688980957
transform 1 0 51796 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_557
timestamp 1688980957
transform 1 0 52348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_597
timestamp 1688980957
transform 1 0 56028 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_38
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_48
timestamp 1688980957
transform 1 0 5520 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_52
timestamp 1688980957
transform 1 0 5888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_58
timestamp 1688980957
transform 1 0 6440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_79
timestamp 1688980957
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_101
timestamp 1688980957
transform 1 0 10396 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_117
timestamp 1688980957
transform 1 0 11868 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_129
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_137
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1688980957
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_218
timestamp 1688980957
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_222
timestamp 1688980957
transform 1 0 21528 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_225
timestamp 1688980957
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_229
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_249
timestamp 1688980957
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_261
timestamp 1688980957
transform 1 0 25116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_274
timestamp 1688980957
transform 1 0 26312 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_283
timestamp 1688980957
transform 1 0 27140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_287
timestamp 1688980957
transform 1 0 27508 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_291
timestamp 1688980957
transform 1 0 27876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_303
timestamp 1688980957
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_331
timestamp 1688980957
transform 1 0 31556 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_335
timestamp 1688980957
transform 1 0 31924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_347
timestamp 1688980957
transform 1 0 33028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_353
timestamp 1688980957
transform 1 0 33580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_405
timestamp 1688980957
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_416
timestamp 1688980957
transform 1 0 39376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_430
timestamp 1688980957
transform 1 0 40664 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_446
timestamp 1688980957
transform 1 0 42136 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_458
timestamp 1688980957
transform 1 0 43240 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_464
timestamp 1688980957
transform 1 0 43792 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_494
timestamp 1688980957
transform 1 0 46552 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_521
timestamp 1688980957
transform 1 0 49036 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_558
timestamp 1688980957
transform 1 0 52440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_562
timestamp 1688980957
transform 1 0 52808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_619
timestamp 1688980957
transform 1 0 58052 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_623
timestamp 1688980957
transform 1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_35
timestamp 1688980957
transform 1 0 4324 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_44
timestamp 1688980957
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_68
timestamp 1688980957
transform 1 0 7360 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_72
timestamp 1688980957
transform 1 0 7728 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_76
timestamp 1688980957
transform 1 0 8096 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_88
timestamp 1688980957
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_154
timestamp 1688980957
transform 1 0 15272 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_164
timestamp 1688980957
transform 1 0 16192 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_185
timestamp 1688980957
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_194
timestamp 1688980957
transform 1 0 18952 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_206
timestamp 1688980957
transform 1 0 20056 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_215
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_219
timestamp 1688980957
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_230
timestamp 1688980957
transform 1 0 22264 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_244
timestamp 1688980957
transform 1 0 23552 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_256
timestamp 1688980957
transform 1 0 24656 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_268
timestamp 1688980957
transform 1 0 25760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_289
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_308
timestamp 1688980957
transform 1 0 29440 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_328
timestamp 1688980957
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_398
timestamp 1688980957
transform 1 0 37720 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_404
timestamp 1688980957
transform 1 0 38272 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_407
timestamp 1688980957
transform 1 0 38548 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_421
timestamp 1688980957
transform 1 0 39836 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_433
timestamp 1688980957
transform 1 0 40940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_445
timestamp 1688980957
transform 1 0 42044 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 1688980957
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_473
timestamp 1688980957
transform 1 0 44620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_484
timestamp 1688980957
transform 1 0 45632 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_496
timestamp 1688980957
transform 1 0 46736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_505
timestamp 1688980957
transform 1 0 47564 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_522
timestamp 1688980957
transform 1 0 49128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_526
timestamp 1688980957
transform 1 0 49496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_530
timestamp 1688980957
transform 1 0 49864 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_533
timestamp 1688980957
transform 1 0 50140 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_545
timestamp 1688980957
transform 1 0 51244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_557
timestamp 1688980957
transform 1 0 52348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_561
timestamp 1688980957
transform 1 0 52716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_569
timestamp 1688980957
transform 1 0 53452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_579
timestamp 1688980957
transform 1 0 54372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_583
timestamp 1688980957
transform 1 0 54740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_594
timestamp 1688980957
transform 1 0 55752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_598
timestamp 1688980957
transform 1 0 56120 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_40
timestamp 1688980957
transform 1 0 4784 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_75
timestamp 1688980957
transform 1 0 8004 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_79
timestamp 1688980957
transform 1 0 8372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_101
timestamp 1688980957
transform 1 0 10396 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_124
timestamp 1688980957
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_136
timestamp 1688980957
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_161
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_176
timestamp 1688980957
transform 1 0 17296 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_185
timestamp 1688980957
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1688980957
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_239
timestamp 1688980957
transform 1 0 23092 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_243
timestamp 1688980957
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_259
timestamp 1688980957
transform 1 0 24932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_339
timestamp 1688980957
transform 1 0 32292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_358
timestamp 1688980957
transform 1 0 34040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_362
timestamp 1688980957
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_377
timestamp 1688980957
transform 1 0 35788 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_391
timestamp 1688980957
transform 1 0 37076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_395
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_398
timestamp 1688980957
transform 1 0 37720 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_425
timestamp 1688980957
transform 1 0 40204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_429
timestamp 1688980957
transform 1 0 40572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_469
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 1688980957
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_477
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_481
timestamp 1688980957
transform 1 0 45356 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_485
timestamp 1688980957
transform 1 0 45724 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_497
timestamp 1688980957
transform 1 0 46828 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_509
timestamp 1688980957
transform 1 0 47932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_512
timestamp 1688980957
transform 1 0 48208 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_520
timestamp 1688980957
transform 1 0 48944 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_523
timestamp 1688980957
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 1688980957
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_533
timestamp 1688980957
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_545
timestamp 1688980957
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_557
timestamp 1688980957
transform 1 0 52348 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_567
timestamp 1688980957
transform 1 0 53268 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_573
timestamp 1688980957
transform 1 0 53820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_576
timestamp 1688980957
transform 1 0 54096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_580
timestamp 1688980957
transform 1 0 54464 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_583
timestamp 1688980957
transform 1 0 54740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_587
timestamp 1688980957
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_613
timestamp 1688980957
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_82
timestamp 1688980957
transform 1 0 8648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_100
timestamp 1688980957
transform 1 0 10304 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_129
timestamp 1688980957
transform 1 0 12972 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_133
timestamp 1688980957
transform 1 0 13340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_153
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_157
timestamp 1688980957
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1688980957
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_178
timestamp 1688980957
transform 1 0 17480 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_190
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_194
timestamp 1688980957
transform 1 0 18952 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_221
timestamp 1688980957
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_231
timestamp 1688980957
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_248
timestamp 1688980957
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_260
timestamp 1688980957
transform 1 0 25024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_311
timestamp 1688980957
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_332
timestamp 1688980957
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_389
timestamp 1688980957
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_401
timestamp 1688980957
transform 1 0 37996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_428
timestamp 1688980957
transform 1 0 40480 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_453
timestamp 1688980957
transform 1 0 42780 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_492
timestamp 1688980957
transform 1 0 46368 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_496
timestamp 1688980957
transform 1 0 46736 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_505
timestamp 1688980957
transform 1 0 47564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_519
timestamp 1688980957
transform 1 0 48852 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_529
timestamp 1688980957
transform 1 0 49772 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_533
timestamp 1688980957
transform 1 0 50140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_541
timestamp 1688980957
transform 1 0 50876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_552
timestamp 1688980957
transform 1 0 51888 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_585
timestamp 1688980957
transform 1 0 54924 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_589
timestamp 1688980957
transform 1 0 55292 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_601
timestamp 1688980957
transform 1 0 56396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_613
timestamp 1688980957
transform 1 0 57500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_617
timestamp 1688980957
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_19
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_46
timestamp 1688980957
transform 1 0 5336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_74
timestamp 1688980957
transform 1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_82
timestamp 1688980957
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_101
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_135
timestamp 1688980957
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_155
timestamp 1688980957
transform 1 0 15364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_187
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_191
timestamp 1688980957
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_214
timestamp 1688980957
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_218
timestamp 1688980957
transform 1 0 21160 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_261
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_267
timestamp 1688980957
transform 1 0 25668 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_303
timestamp 1688980957
transform 1 0 28980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_317
timestamp 1688980957
transform 1 0 30268 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_339
timestamp 1688980957
transform 1 0 32292 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_361
timestamp 1688980957
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_438
timestamp 1688980957
transform 1 0 41400 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_518
timestamp 1688980957
transform 1 0 48760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_522
timestamp 1688980957
transform 1 0 49128 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_542
timestamp 1688980957
transform 1 0 50968 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_573
timestamp 1688980957
transform 1 0 53820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_585
timestamp 1688980957
transform 1 0 54924 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_598
timestamp 1688980957
transform 1 0 56120 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_610
timestamp 1688980957
transform 1 0 57224 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_622
timestamp 1688980957
transform 1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_29
timestamp 1688980957
transform 1 0 3772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_38
timestamp 1688980957
transform 1 0 4600 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_42
timestamp 1688980957
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1688980957
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_66
timestamp 1688980957
transform 1 0 7176 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_78
timestamp 1688980957
transform 1 0 8280 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_86
timestamp 1688980957
transform 1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_117
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_126
timestamp 1688980957
transform 1 0 12696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_130
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_165
timestamp 1688980957
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 1688980957
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_267
timestamp 1688980957
transform 1 0 25668 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_276
timestamp 1688980957
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_285
timestamp 1688980957
transform 1 0 27324 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_307
timestamp 1688980957
transform 1 0 29348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_321
timestamp 1688980957
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_333
timestamp 1688980957
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_345
timestamp 1688980957
transform 1 0 32844 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_372
timestamp 1688980957
transform 1 0 35328 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_389
timestamp 1688980957
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_401
timestamp 1688980957
transform 1 0 37996 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 1688980957
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_457
timestamp 1688980957
transform 1 0 43148 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_463
timestamp 1688980957
transform 1 0 43700 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_505
timestamp 1688980957
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_510
timestamp 1688980957
transform 1 0 48024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_549
timestamp 1688980957
transform 1 0 51612 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_561
timestamp 1688980957
transform 1 0 52716 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_565
timestamp 1688980957
transform 1 0 53084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_612
timestamp 1688980957
transform 1 0 57408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_617
timestamp 1688980957
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_62
timestamp 1688980957
transform 1 0 6808 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_74
timestamp 1688980957
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_182
timestamp 1688980957
transform 1 0 17848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_192
timestamp 1688980957
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_211
timestamp 1688980957
transform 1 0 20516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_223
timestamp 1688980957
transform 1 0 21620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_237
timestamp 1688980957
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_246
timestamp 1688980957
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_359
timestamp 1688980957
transform 1 0 34132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_386
timestamp 1688980957
transform 1 0 36616 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_390
timestamp 1688980957
transform 1 0 36984 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_402
timestamp 1688980957
transform 1 0 38088 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_414
timestamp 1688980957
transform 1 0 39192 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_429
timestamp 1688980957
transform 1 0 40572 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_441
timestamp 1688980957
transform 1 0 41676 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_453
timestamp 1688980957
transform 1 0 42780 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_465
timestamp 1688980957
transform 1 0 43884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_473
timestamp 1688980957
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_485
timestamp 1688980957
transform 1 0 45724 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_489
timestamp 1688980957
transform 1 0 46092 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_549
timestamp 1688980957
transform 1 0 51612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_568
timestamp 1688980957
transform 1 0 53360 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 1688980957
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_605
timestamp 1688980957
transform 1 0 56764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_617
timestamp 1688980957
transform 1 0 57868 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_145
timestamp 1688980957
transform 1 0 14444 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 1688980957
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_185
timestamp 1688980957
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_194
timestamp 1688980957
transform 1 0 18952 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_206
timestamp 1688980957
transform 1 0 20056 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_218
timestamp 1688980957
transform 1 0 21160 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 1688980957
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1688980957
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1688980957
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 1688980957
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 1688980957
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 1688980957
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 1688980957
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_485
timestamp 1688980957
transform 1 0 45724 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_493
timestamp 1688980957
transform 1 0 46460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_498
timestamp 1688980957
transform 1 0 46920 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_513
timestamp 1688980957
transform 1 0 48300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_525
timestamp 1688980957
transform 1 0 49404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_537
timestamp 1688980957
transform 1 0 50508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_549
timestamp 1688980957
transform 1 0 51612 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_557
timestamp 1688980957
transform 1 0 52348 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_577
timestamp 1688980957
transform 1 0 54188 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_589
timestamp 1688980957
transform 1 0 55292 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_601
timestamp 1688980957
transform 1 0 56396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_613
timestamp 1688980957
transform 1 0 57500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_617
timestamp 1688980957
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 1688980957
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 1688980957
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1688980957
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 1688980957
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 1688980957
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 1688980957
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 1688980957
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 1688980957
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 1688980957
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 1688980957
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 1688980957
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 1688980957
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 1688980957
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 1688980957
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 1688980957
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 1688980957
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 1688980957
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 1688980957
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 1688980957
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 1688980957
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 1688980957
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_613
timestamp 1688980957
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1688980957
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 1688980957
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_441
timestamp 1688980957
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 1688980957
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 1688980957
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 1688980957
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 1688980957
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 1688980957
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 1688980957
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 1688980957
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 1688980957
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 1688980957
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 1688980957
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 1688980957
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 1688980957
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 1688980957
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 1688980957
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 1688980957
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 1688980957
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 1688980957
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_617
timestamp 1688980957
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1688980957
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1688980957
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 1688980957
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 1688980957
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 1688980957
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 1688980957
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 1688980957
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 1688980957
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 1688980957
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 1688980957
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1688980957
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 1688980957
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 1688980957
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 1688980957
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 1688980957
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 1688980957
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 1688980957
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 1688980957
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 1688980957
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 1688980957
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 1688980957
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 1688980957
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 1688980957
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 1688980957
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 1688980957
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 1688980957
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 1688980957
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 1688980957
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 1688980957
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 1688980957
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 1688980957
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 1688980957
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 1688980957
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 1688980957
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 1688980957
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_617
timestamp 1688980957
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1688980957
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1688980957
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1688980957
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 1688980957
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 1688980957
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 1688980957
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 1688980957
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 1688980957
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 1688980957
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 1688980957
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 1688980957
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 1688980957
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 1688980957
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 1688980957
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 1688980957
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 1688980957
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 1688980957
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 1688980957
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1688980957
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1688980957
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 1688980957
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 1688980957
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 1688980957
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 1688980957
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 1688980957
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 1688980957
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 1688980957
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 1688980957
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 1688980957
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 1688980957
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 1688980957
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 1688980957
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 1688980957
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 1688980957
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 1688980957
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 1688980957
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 1688980957
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 1688980957
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_617
timestamp 1688980957
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_57
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 1688980957
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1688980957
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_281
timestamp 1688980957
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_293
timestamp 1688980957
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_337
timestamp 1688980957
transform 1 0 32108 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_349
timestamp 1688980957
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_393
timestamp 1688980957
transform 1 0 37260 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_405
timestamp 1688980957
transform 1 0 38364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_417
timestamp 1688980957
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_445
timestamp 1688980957
transform 1 0 42044 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_449
timestamp 1688980957
transform 1 0 42412 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_461
timestamp 1688980957
transform 1 0 43516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_473
timestamp 1688980957
transform 1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1688980957
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1688980957
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_501
timestamp 1688980957
transform 1 0 47196 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_505
timestamp 1688980957
transform 1 0 47564 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_517
timestamp 1688980957
transform 1 0 48668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_529
timestamp 1688980957
transform 1 0 49772 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1688980957
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 1688980957
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_557
timestamp 1688980957
transform 1 0 52348 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_561
timestamp 1688980957
transform 1 0 52716 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_573
timestamp 1688980957
transform 1 0 53820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_585
timestamp 1688980957
transform 1 0 54924 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1688980957
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1688980957
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_613
timestamp 1688980957
transform 1 0 57500 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_617
timestamp 1688980957
transform 1 0 57868 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 17664 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold7
timestamp 1688980957
transform -1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 9016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 20240 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 21436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 48300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold12
timestamp 1688980957
transform -1 0 45448 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 43608 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 27232 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold17
timestamp 1688980957
transform 1 0 30176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 30084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 19136 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 50692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold24
timestamp 1688980957
transform 1 0 47656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 49128 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 58604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold27
timestamp 1688980957
transform -1 0 53452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 52440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 21712 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 29164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 31740 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 30176 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 32844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 29440 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 11776 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold40
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 38916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 47196 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 58604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold45
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 54648 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 58604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 58604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 55016 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 54280 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold52
timestamp 1688980957
transform -1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 22172 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 45724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 45724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 25116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 24380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 30360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 29440 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 28888 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 50876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 50876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 50968 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 50048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 43884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 46368 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 29256 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 41952 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 40572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 55476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 56028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 45632 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 44804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 42044 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 42044 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 24196 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 58604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 56120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 58604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 57316 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 38088 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 39560 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 48300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 48668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 31556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 31924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 49128 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 47656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 46644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 46644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 22816 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 26036 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 27600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold101
timestamp 1688980957
transform -1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 11960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 53452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 52348 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 41584 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform 1 0 41676 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 42596 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 56028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 56764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 53452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 53544 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 53452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 54280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 54188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 54924 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 20240 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 41032 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 40296 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 42504 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 28520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 46184 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 44528 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 47472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 48392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 23644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 45908 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 44620 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 52532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 51796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 17388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform -1 0 39468 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 38456 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 38272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform -1 0 38272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 25116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform -1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform -1 0 37996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold148
timestamp 1688980957
transform -1 0 35512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform -1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 52348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 50048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold153
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 7728 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 54648 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold156
timestamp 1688980957
transform -1 0 58604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 55936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform 1 0 23092 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold159
timestamp 1688980957
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform 1 0 55292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform -1 0 55016 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 56948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform -1 0 56764 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform -1 0 35604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 23736 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform -1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 11040 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 39560 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 39744 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform 1 0 33580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform -1 0 33304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform -1 0 57500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform -1 0 56764 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 37904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform -1 0 37168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 37720 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 36984 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 58604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 56948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform 1 0 24932 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 27232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform -1 0 55660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 53268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 53452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform 1 0 33856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform -1 0 33856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 11592 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 10856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform -1 0 24012 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 27324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 26864 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 53452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 52532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform 1 0 29716 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold204
timestamp 1688980957
transform -1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform 1 0 27968 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform 1 0 25208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 25116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold209
timestamp 1688980957
transform -1 0 22080 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 22724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 13064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 12696 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 36892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold214
timestamp 1688980957
transform 1 0 36248 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform -1 0 36524 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 33764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform -1 0 54924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold219
timestamp 1688980957
transform -1 0 49128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform -1 0 46920 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform -1 0 44620 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold222
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 42044 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 45724 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 45080 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 32292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 32200 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform -1 0 36800 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 36248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 50416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 49680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 34316 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 33672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 33488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 34408 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 44896 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 45264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 34408 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 34316 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform 1 0 50048 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 51704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 43884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform -1 0 44620 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform -1 0 30268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform -1 0 38732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 37996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 22540 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform -1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform 1 0 35512 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform -1 0 46828 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform 1 0 12512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform -1 0 17204 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 15456 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform -1 0 46828 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform 1 0 40940 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform -1 0 42044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform -1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform -1 0 45724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform -1 0 44988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform 1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform -1 0 3036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform 1 0 27876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform -1 0 50232 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform -1 0 47840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform -1 0 16652 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform 1 0 41400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform -1 0 41952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform -1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform -1 0 39468 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform 1 0 21068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform -1 0 21068 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform -1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform -1 0 27048 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform 1 0 35512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 35144 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform 1 0 36064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform -1 0 36616 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform -1 0 38640 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform -1 0 39652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform -1 0 6992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform -1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform 1 0 22448 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform -1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform -1 0 43240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform -1 0 41676 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform -1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold297
timestamp 1688980957
transform 1 0 27048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform -1 0 26680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform 1 0 49128 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform -1 0 50048 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform -1 0 25208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform 1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform -1 0 8464 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform -1 0 8556 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 58604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold306
timestamp 1688980957
transform -1 0 56120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform -1 0 52256 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform 1 0 26404 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform -1 0 26312 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform -1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform -1 0 38824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform 1 0 38364 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform 1 0 56028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform -1 0 56028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform -1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform -1 0 24472 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform -1 0 24288 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform -1 0 3680 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform -1 0 58604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform -1 0 58604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 46092 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold325
timestamp 1688980957
transform 1 0 42412 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform -1 0 43516 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform -1 0 13064 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold328
timestamp 1688980957
transform 1 0 11316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform -1 0 11040 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform -1 0 20516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform 1 0 29624 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform -1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform 1 0 55292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform -1 0 55108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform -1 0 20608 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform -1 0 25760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform 1 0 49588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform -1 0 51060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform -1 0 42136 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform -1 0 29164 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform 1 0 27140 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform 1 0 50968 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform -1 0 52624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform -1 0 10212 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1688980957
transform -1 0 54556 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform -1 0 54280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1688980957
transform -1 0 13616 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold357
timestamp 1688980957
transform -1 0 40572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1688980957
transform -1 0 39192 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold359
timestamp 1688980957
transform -1 0 13892 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1688980957
transform -1 0 13156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold362
timestamp 1688980957
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1688980957
transform 1 0 21620 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1688980957
transform -1 0 55844 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold365
timestamp 1688980957
transform 1 0 52716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1688980957
transform -1 0 53452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1688980957
transform 1 0 53084 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1688980957
transform -1 0 53084 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 1688980957
transform -1 0 58604 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1688980957
transform -1 0 58604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1688980957
transform -1 0 41400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1688980957
transform -1 0 41860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 1688980957
transform 1 0 18768 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold374
timestamp 1688980957
transform -1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold375
timestamp 1688980957
transform -1 0 15824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold376
timestamp 1688980957
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold377
timestamp 1688980957
transform -1 0 20792 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 1688980957
transform 1 0 15824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 1688980957
transform -1 0 15824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 1688980957
transform -1 0 58420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 1688980957
transform -1 0 58604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold382
timestamp 1688980957
transform 1 0 56028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold383
timestamp 1688980957
transform -1 0 56028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 1688980957
transform -1 0 56028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 1688980957
transform -1 0 54924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 1688980957
transform -1 0 19320 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 1688980957
transform -1 0 19044 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold388
timestamp 1688980957
transform 1 0 20424 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold389
timestamp 1688980957
transform -1 0 20424 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 1688980957
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 1688980957
transform -1 0 9752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold392
timestamp 1688980957
transform -1 0 14996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold393
timestamp 1688980957
transform -1 0 13984 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold394
timestamp 1688980957
transform -1 0 52348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold395
timestamp 1688980957
transform 1 0 49312 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 1688980957
transform -1 0 52440 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold397
timestamp 1688980957
transform 1 0 11316 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 1688980957
transform -1 0 11224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold399
timestamp 1688980957
transform -1 0 46368 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold400
timestamp 1688980957
transform -1 0 46552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold401
timestamp 1688980957
transform -1 0 56764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold402
timestamp 1688980957
transform -1 0 57408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold403
timestamp 1688980957
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold404
timestamp 1688980957
transform -1 0 33028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 1688980957
transform -1 0 30820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold406
timestamp 1688980957
transform -1 0 25116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold407
timestamp 1688980957
transform -1 0 23552 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold408
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold409
timestamp 1688980957
transform -1 0 37628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold411
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold412
timestamp 1688980957
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold413
timestamp 1688980957
transform -1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold414
timestamp 1688980957
transform -1 0 17664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold415
timestamp 1688980957
transform 1 0 7912 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold416
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold417
timestamp 1688980957
transform 1 0 10488 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 1688980957
transform -1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 1688980957
transform -1 0 45632 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 1688980957
transform -1 0 46552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 1688980957
transform 1 0 53452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 1688980957
transform -1 0 53452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 1688980957
transform -1 0 50876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 1688980957
transform -1 0 49772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 1688980957
transform -1 0 46460 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 1688980957
transform -1 0 44252 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 1688980957
transform 1 0 16928 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 1688980957
transform -1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 1688980957
transform 1 0 9936 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 1688980957
transform -1 0 9936 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold432
timestamp 1688980957
transform -1 0 15916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 1688980957
transform 1 0 46736 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 1688980957
transform -1 0 48852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 1688980957
transform -1 0 12788 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 1688980957
transform -1 0 11408 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold437
timestamp 1688980957
transform 1 0 48392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 1688980957
transform -1 0 48392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 1688980957
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 1688980957
transform -1 0 14352 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 1688980957
transform -1 0 42228 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 1688980957
transform -1 0 51612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 1688980957
transform -1 0 51888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 1688980957
transform -1 0 46000 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 1688980957
transform -1 0 45724 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 1688980957
transform 1 0 43516 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 1688980957
transform -1 0 43516 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 1688980957
transform -1 0 35144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 1688980957
transform -1 0 34040 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 1688980957
transform -1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 1688980957
transform 1 0 49312 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 1688980957
transform 1 0 50968 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold456
timestamp 1688980957
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold457
timestamp 1688980957
transform -1 0 6808 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold458
timestamp 1688980957
transform -1 0 58604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold459
timestamp 1688980957
transform -1 0 57500 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold460
timestamp 1688980957
transform 1 0 4784 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 1688980957
transform 1 0 4416 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 1688980957
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 1688980957
transform -1 0 10304 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold464
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold465
timestamp 1688980957
transform -1 0 54372 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 1688980957
transform 1 0 26772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 1688980957
transform -1 0 26496 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 1688980957
transform 1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 1688980957
transform -1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold470
timestamp 1688980957
transform 1 0 4600 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 1688980957
transform -1 0 4600 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold473
timestamp 1688980957
transform -1 0 36616 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 1688980957
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold475
timestamp 1688980957
transform -1 0 46920 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold476
timestamp 1688980957
transform -1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 1688980957
transform -1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 1688980957
transform 1 0 48116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 1688980957
transform -1 0 48760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 1688980957
transform -1 0 13984 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold481
timestamp 1688980957
transform -1 0 13156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold482
timestamp 1688980957
transform 1 0 37628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold483
timestamp 1688980957
transform -1 0 36708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 1688980957
transform 1 0 17940 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 1688980957
transform -1 0 19688 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold486
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold487
timestamp 1688980957
transform -1 0 31740 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold488
timestamp 1688980957
transform -1 0 41400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 1688980957
transform -1 0 40756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold491
timestamp 1688980957
transform -1 0 37076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold492
timestamp 1688980957
transform -1 0 29348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold493
timestamp 1688980957
transform -1 0 28612 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold494
timestamp 1688980957
transform -1 0 35328 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold495
timestamp 1688980957
transform -1 0 34132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold496
timestamp 1688980957
transform -1 0 8556 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold497
timestamp 1688980957
transform -1 0 7636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold498
timestamp 1688980957
transform -1 0 8648 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold499
timestamp 1688980957
transform -1 0 7912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold500
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold501
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold502
timestamp 1688980957
transform 1 0 17480 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold503
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold504
timestamp 1688980957
transform -1 0 26680 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold505
timestamp 1688980957
transform -1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold506
timestamp 1688980957
transform -1 0 34868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold507
timestamp 1688980957
transform -1 0 30268 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold508
timestamp 1688980957
transform -1 0 29440 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold509
timestamp 1688980957
transform 1 0 31556 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold510
timestamp 1688980957
transform -1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold511
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold512
timestamp 1688980957
transform -1 0 13524 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold513
timestamp 1688980957
transform -1 0 41492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold514
timestamp 1688980957
transform -1 0 40572 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold515
timestamp 1688980957
transform 1 0 15456 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold516
timestamp 1688980957
transform -1 0 15456 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold517
timestamp 1688980957
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold518
timestamp 1688980957
transform -1 0 30268 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold519
timestamp 1688980957
transform 1 0 15548 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold520
timestamp 1688980957
transform -1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold521
timestamp 1688980957
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold522
timestamp 1688980957
transform -1 0 3680 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold523
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold524
timestamp 1688980957
transform -1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold525
timestamp 1688980957
transform 1 0 20700 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold526
timestamp 1688980957
transform -1 0 20516 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold527
timestamp 1688980957
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold528
timestamp 1688980957
transform -1 0 3772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold529
timestamp 1688980957
transform 1 0 18216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold530
timestamp 1688980957
transform -1 0 18124 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 1688980957
transform -1 0 18768 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 1688980957
transform -1 0 19688 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold533
timestamp 1688980957
transform 1 0 15272 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold534
timestamp 1688980957
transform -1 0 15272 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold535
timestamp 1688980957
transform -1 0 34592 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold536
timestamp 1688980957
transform -1 0 35420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold537
timestamp 1688980957
transform -1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold538
timestamp 1688980957
transform 1 0 18216 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold539
timestamp 1688980957
transform -1 0 23736 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold540
timestamp 1688980957
transform -1 0 22908 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold541
timestamp 1688980957
transform -1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold542
timestamp 1688980957
transform -1 0 24012 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold543
timestamp 1688980957
transform 1 0 21528 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold544
timestamp 1688980957
transform -1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold545
timestamp 1688980957
transform 1 0 1472 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold546
timestamp 1688980957
transform -1 0 2208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold547
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold548
timestamp 1688980957
transform -1 0 3220 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold549
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold550
timestamp 1688980957
transform 1 0 4232 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold551
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold552
timestamp 1688980957
transform -1 0 3680 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold553
timestamp 1688980957
transform -1 0 36984 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold554
timestamp 1688980957
transform -1 0 36432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold555
timestamp 1688980957
transform -1 0 49772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold556
timestamp 1688980957
transform -1 0 48300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold557
timestamp 1688980957
transform -1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold558
timestamp 1688980957
transform -1 0 33580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold559
timestamp 1688980957
transform -1 0 31924 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold560
timestamp 1688980957
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold561
timestamp 1688980957
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold562
timestamp 1688980957
transform 1 0 21344 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold563
timestamp 1688980957
transform -1 0 43148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold564
timestamp 1688980957
transform -1 0 42044 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold565
timestamp 1688980957
transform -1 0 28244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold566
timestamp 1688980957
transform -1 0 27508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold567
timestamp 1688980957
transform -1 0 35052 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold568
timestamp 1688980957
transform -1 0 34592 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold569
timestamp 1688980957
transform -1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold570
timestamp 1688980957
transform 1 0 12512 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold571
timestamp 1688980957
transform -1 0 26772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold572
timestamp 1688980957
transform -1 0 25300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold573
timestamp 1688980957
transform -1 0 50876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold574
timestamp 1688980957
transform -1 0 52348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold575
timestamp 1688980957
transform 1 0 14260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold576
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold577
timestamp 1688980957
transform -1 0 58420 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold578
timestamp 1688980957
transform -1 0 57500 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold579
timestamp 1688980957
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold580
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold581
timestamp 1688980957
transform 1 0 57868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold582
timestamp 1688980957
transform -1 0 58604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold583
timestamp 1688980957
transform -1 0 40020 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold584
timestamp 1688980957
transform -1 0 39284 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold585
timestamp 1688980957
transform -1 0 21344 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold586
timestamp 1688980957
transform -1 0 20608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold587
timestamp 1688980957
transform -1 0 47104 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold588
timestamp 1688980957
transform -1 0 46552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold589
timestamp 1688980957
transform -1 0 49772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold590
timestamp 1688980957
transform -1 0 49864 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold591
timestamp 1688980957
transform -1 0 52992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold592
timestamp 1688980957
transform -1 0 53084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold593
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold594
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold595
timestamp 1688980957
transform -1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold596
timestamp 1688980957
transform 1 0 4048 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold597
timestamp 1688980957
transform -1 0 36524 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold598
timestamp 1688980957
transform -1 0 35696 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold599
timestamp 1688980957
transform 1 0 9016 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold600
timestamp 1688980957
transform -1 0 12052 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold601
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold602
timestamp 1688980957
transform -1 0 16560 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold603
timestamp 1688980957
transform -1 0 6164 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold604
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold605
timestamp 1688980957
transform 1 0 7176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold606
timestamp 1688980957
transform -1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold607
timestamp 1688980957
transform -1 0 18768 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold608
timestamp 1688980957
transform -1 0 58604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold609
timestamp 1688980957
transform -1 0 58604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold610
timestamp 1688980957
transform -1 0 44988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold611
timestamp 1688980957
transform -1 0 44252 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold612
timestamp 1688980957
transform -1 0 28796 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold613
timestamp 1688980957
transform -1 0 27968 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold614
timestamp 1688980957
transform -1 0 25576 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold615
timestamp 1688980957
transform -1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold616
timestamp 1688980957
transform 1 0 53452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold617
timestamp 1688980957
transform -1 0 53452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold618
timestamp 1688980957
transform -1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold619
timestamp 1688980957
transform -1 0 41400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold620 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold621
timestamp 1688980957
transform 1 0 3956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold622
timestamp 1688980957
transform -1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold623
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold624
timestamp 1688980957
transform 1 0 2116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold625
timestamp 1688980957
transform -1 0 9108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold626
timestamp 1688980957
transform -1 0 51704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold627
timestamp 1688980957
transform -1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold628
timestamp 1688980957
transform -1 0 12236 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold629
timestamp 1688980957
transform -1 0 7176 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold630
timestamp 1688980957
transform -1 0 53636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold631
timestamp 1688980957
transform -1 0 26956 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold632
timestamp 1688980957
transform -1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold633
timestamp 1688980957
transform -1 0 55384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold634
timestamp 1688980957
transform -1 0 34500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold635
timestamp 1688980957
transform 1 0 17296 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold636
timestamp 1688980957
transform -1 0 16652 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold637
timestamp 1688980957
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold638
timestamp 1688980957
transform -1 0 44712 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold639
timestamp 1688980957
transform -1 0 36524 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold640
timestamp 1688980957
transform -1 0 8464 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold641
timestamp 1688980957
transform -1 0 54188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold642
timestamp 1688980957
transform -1 0 23368 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold643
timestamp 1688980957
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold644
timestamp 1688980957
transform -1 0 40020 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold645
timestamp 1688980957
transform -1 0 58604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold646
timestamp 1688980957
transform 1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold647
timestamp 1688980957
transform 1 0 50968 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold648
timestamp 1688980957
transform -1 0 39652 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold649
timestamp 1688980957
transform 1 0 11776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold650
timestamp 1688980957
transform -1 0 31648 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold651
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold652
timestamp 1688980957
transform -1 0 27416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold653
timestamp 1688980957
transform -1 0 43516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold654
timestamp 1688980957
transform -1 0 47840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold655
timestamp 1688980957
transform -1 0 30912 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold656
timestamp 1688980957
transform -1 0 43148 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold657
timestamp 1688980957
transform -1 0 31556 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 24196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 26772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 31464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 33672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 34500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 39376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 42136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform -1 0 42228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform -1 0 47104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 46276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 49588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 50784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform -1 0 53360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 55016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 9752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 57500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 16744 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform -1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1688980957
transform -1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output37 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 1688980957
transform 1 0 7268 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output39
timestamp 1688980957
transform -1 0 25300 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output40
timestamp 1688980957
transform -1 0 26864 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output41
timestamp 1688980957
transform 1 0 27140 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 1688980957
transform 1 0 27968 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 1688980957
transform -1 0 31924 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 1688980957
transform -1 0 33580 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output45
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output46
timestamp 1688980957
transform 1 0 36156 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output47
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output48
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output49
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output50
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 1688980957
transform -1 0 45356 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1688980957
transform -1 0 46828 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1688980957
transform -1 0 49036 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1688980957
transform 1 0 50324 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1688980957
transform -1 0 54188 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1688980957
transform 1 0 53636 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1688980957
transform -1 0 56764 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1688980957
transform -1 0 11408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1688980957
transform -1 0 58420 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1688980957
transform -1 0 57776 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1688980957
transform -1 0 13708 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1688980957
transform -1 0 13984 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1688980957
transform -1 0 20332 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1688980957
transform -1 0 21712 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 52624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 57776 0 1 27200
box -38 -48 130 592
<< labels >>
flabel metal4 s 8166 2128 8486 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 22610 2128 22930 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 37054 2128 37374 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 51498 2128 51818 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 15388 2128 15708 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 29832 2128 30152 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 44276 2128 44596 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 58720 2128 59040 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 5 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 6 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 7 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 8 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 9 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 10 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 11 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 12 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 13 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 14 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 15 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 16 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 17 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 18 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 19 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 20 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 21 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 22 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 23 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 24 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 25 nsew signal input
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 26 nsew signal input
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 27 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 28 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 29 nsew signal input
flabel metal2 s 57702 0 57758 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 30 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 31 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 32 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 33 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 34 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 35 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 36 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 37 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 38 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 39 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 40 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 41 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 42 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 43 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 44 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 45 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 46 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 47 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 48 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 49 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 50 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 51 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 52 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 53 nsew signal tristate
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 54 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 55 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 56 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 57 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 58 nsew signal tristate
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 59 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 60 nsew signal tristate
flabel metal2 s 56874 0 56930 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 61 nsew signal tristate
flabel metal2 s 58530 0 58586 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 62 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 63 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 64 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 65 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 66 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 67 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 68 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 69 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 70 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wbs_we_i
port 71 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
<< end >>
