magic
tech sky130A
magscale 1 2
timestamp 1727690133
<< viali >>
rect 37013 32385 37047 32419
rect 14105 32317 14139 32351
rect 14933 32317 14967 32351
rect 24593 32317 24627 32351
rect 24777 32317 24811 32351
rect 28181 32317 28215 32351
rect 28825 32317 28859 32351
rect 37289 32317 37323 32351
rect 10333 32181 10367 32215
rect 13461 32181 13495 32215
rect 14289 32181 14323 32215
rect 24041 32181 24075 32215
rect 25421 32181 25455 32215
rect 26709 32181 26743 32215
rect 27353 32181 27387 32215
rect 27537 32181 27571 32215
rect 28273 32181 28307 32215
rect 36369 32181 36403 32215
rect 37933 32181 37967 32215
rect 14105 31977 14139 32011
rect 23949 31977 23983 32011
rect 28457 31977 28491 32011
rect 13093 31909 13127 31943
rect 26893 31909 26927 31943
rect 14565 31841 14599 31875
rect 14657 31841 14691 31875
rect 23397 31841 23431 31875
rect 23489 31841 23523 31875
rect 26801 31841 26835 31875
rect 27445 31841 27479 31875
rect 27813 31841 27847 31875
rect 27997 31841 28031 31875
rect 36001 31841 36035 31875
rect 10333 31773 10367 31807
rect 11253 31773 11287 31807
rect 13921 31773 13955 31807
rect 15577 31773 15611 31807
rect 19073 31773 19107 31807
rect 19717 31773 19751 31807
rect 23121 31773 23155 31807
rect 24961 31773 24995 31807
rect 25697 31773 25731 31807
rect 26157 31773 26191 31807
rect 29193 31773 29227 31807
rect 31953 31773 31987 31807
rect 32505 31773 32539 31807
rect 35817 31773 35851 31807
rect 36553 31773 36587 31807
rect 36737 31773 36771 31807
rect 37289 31773 37323 31807
rect 37473 31773 37507 31807
rect 38117 31773 38151 31807
rect 12817 31705 12851 31739
rect 14473 31705 14507 31739
rect 27261 31705 27295 31739
rect 9689 31637 9723 31671
rect 10609 31637 10643 31671
rect 13277 31637 13311 31671
rect 15025 31637 15059 31671
rect 18429 31637 18463 31671
rect 19533 31637 19567 31671
rect 20361 31637 20395 31671
rect 23581 31637 23615 31671
rect 24409 31637 24443 31671
rect 25145 31637 25179 31671
rect 27353 31637 27387 31671
rect 28089 31637 28123 31671
rect 28549 31637 28583 31671
rect 29745 31637 29779 31671
rect 35265 31637 35299 31671
rect 9965 31433 9999 31467
rect 13369 31433 13403 31467
rect 20085 31433 20119 31467
rect 23581 31433 23615 31467
rect 28365 31433 28399 31467
rect 29193 31433 29227 31467
rect 29285 31433 29319 31467
rect 13461 31365 13495 31399
rect 23940 31365 23974 31399
rect 27252 31365 27286 31399
rect 28733 31365 28767 31399
rect 30021 31365 30055 31399
rect 31861 31365 31895 31399
rect 35440 31365 35474 31399
rect 9873 31297 9907 31331
rect 14096 31297 14130 31331
rect 18512 31297 18546 31331
rect 22457 31297 22491 31331
rect 25697 31297 25731 31331
rect 26985 31297 27019 31331
rect 28825 31297 28859 31331
rect 32404 31297 32438 31331
rect 33609 31297 33643 31331
rect 9413 31229 9447 31263
rect 10057 31229 10091 31263
rect 10885 31229 10919 31263
rect 11529 31229 11563 31263
rect 12357 31229 12391 31263
rect 13645 31229 13679 31263
rect 13829 31229 13863 31263
rect 15853 31229 15887 31263
rect 18245 31229 18279 31263
rect 19809 31229 19843 31263
rect 19993 31229 20027 31263
rect 21097 31229 21131 31263
rect 22201 31229 22235 31263
rect 23673 31229 23707 31263
rect 25145 31229 25179 31263
rect 26433 31229 26467 31263
rect 28549 31229 28583 31263
rect 29837 31229 29871 31263
rect 30573 31229 30607 31263
rect 32137 31229 32171 31263
rect 34161 31229 34195 31263
rect 34897 31229 34931 31263
rect 35173 31229 35207 31263
rect 37289 31229 37323 31263
rect 9505 31161 9539 31195
rect 13001 31161 13035 31195
rect 15209 31161 15243 31195
rect 20453 31161 20487 31195
rect 25053 31161 25087 31195
rect 33517 31161 33551 31195
rect 8769 31093 8803 31127
rect 10333 31093 10367 31127
rect 11345 31093 11379 31127
rect 12173 31093 12207 31127
rect 12909 31093 12943 31127
rect 15301 31093 15335 31127
rect 19625 31093 19659 31127
rect 20545 31093 20579 31127
rect 25881 31093 25915 31127
rect 34345 31093 34379 31127
rect 36553 31093 36587 31127
rect 37933 31093 37967 31127
rect 10793 30889 10827 30923
rect 13921 30889 13955 30923
rect 15577 30889 15611 30923
rect 19257 30889 19291 30923
rect 23305 30889 23339 30923
rect 24409 30889 24443 30923
rect 27629 30889 27663 30923
rect 29101 30889 29135 30923
rect 36369 30889 36403 30923
rect 10701 30821 10735 30855
rect 15485 30821 15519 30855
rect 33793 30821 33827 30855
rect 11345 30753 11379 30787
rect 14105 30753 14139 30787
rect 16129 30753 16163 30787
rect 16957 30753 16991 30787
rect 20637 30753 20671 30787
rect 21925 30753 21959 30787
rect 23581 30753 23615 30787
rect 30021 30753 30055 30787
rect 30113 30753 30147 30787
rect 34437 30753 34471 30787
rect 9321 30685 9355 30719
rect 9588 30685 9622 30719
rect 12173 30685 12207 30719
rect 12541 30685 12575 30719
rect 14372 30685 14406 30719
rect 16037 30685 16071 30719
rect 17693 30685 17727 30719
rect 20381 30685 20415 30719
rect 21281 30685 21315 30719
rect 21833 30685 21867 30719
rect 23765 30685 23799 30719
rect 25789 30685 25823 30719
rect 26249 30685 26283 30719
rect 27721 30685 27755 30719
rect 27988 30685 28022 30719
rect 30573 30685 30607 30719
rect 30941 30685 30975 30719
rect 32413 30685 32447 30719
rect 34989 30685 35023 30719
rect 37841 30685 37875 30719
rect 11161 30617 11195 30651
rect 11621 30617 11655 30651
rect 12808 30617 12842 30651
rect 15945 30617 15979 30651
rect 16405 30617 16439 30651
rect 17960 30617 17994 30651
rect 22192 30617 22226 30651
rect 25522 30617 25556 30651
rect 26494 30617 26528 30651
rect 29929 30617 29963 30651
rect 31208 30617 31242 30651
rect 32680 30617 32714 30651
rect 35256 30617 35290 30651
rect 37596 30617 37630 30651
rect 9229 30549 9263 30583
rect 11253 30549 11287 30583
rect 17601 30549 17635 30583
rect 19073 30549 19107 30583
rect 20729 30549 20763 30583
rect 23673 30549 23707 30583
rect 24133 30549 24167 30583
rect 29561 30549 29595 30583
rect 32321 30549 32355 30583
rect 33885 30549 33919 30583
rect 36461 30549 36495 30583
rect 11989 30345 12023 30379
rect 14013 30345 14047 30379
rect 16221 30345 16255 30379
rect 22201 30345 22235 30379
rect 30481 30345 30515 30379
rect 8300 30277 8334 30311
rect 12900 30277 12934 30311
rect 25053 30277 25087 30311
rect 34805 30277 34839 30311
rect 37749 30277 37783 30311
rect 10425 30209 10459 30243
rect 11161 30209 11195 30243
rect 11345 30209 11379 30243
rect 11897 30209 11931 30243
rect 12633 30209 12667 30243
rect 14908 30209 14942 30243
rect 15025 30209 15059 30243
rect 15761 30209 15795 30243
rect 15945 30209 15979 30243
rect 17141 30209 17175 30243
rect 17408 30209 17442 30243
rect 18797 30209 18831 30243
rect 19809 30209 19843 30243
rect 21097 30209 21131 30243
rect 23740 30209 23774 30243
rect 23857 30209 23891 30243
rect 24777 30209 24811 30243
rect 26801 30209 26835 30243
rect 27813 30209 27847 30243
rect 27972 30209 28006 30243
rect 28089 30209 28123 30243
rect 28825 30209 28859 30243
rect 29653 30209 29687 30243
rect 30573 30209 30607 30243
rect 30829 30209 30863 30243
rect 32940 30209 32974 30243
rect 33057 30209 33091 30243
rect 33793 30209 33827 30243
rect 33977 30209 34011 30243
rect 36185 30209 36219 30243
rect 37105 30209 37139 30243
rect 37657 30209 37691 30243
rect 8033 30141 8067 30175
rect 10149 30141 10183 30175
rect 10308 30141 10342 30175
rect 12173 30141 12207 30175
rect 14739 30141 14773 30175
rect 18613 30141 18647 30175
rect 19533 30141 19567 30175
rect 19650 30141 19684 30175
rect 22753 30141 22787 30175
rect 23581 30141 23615 30175
rect 24593 30141 24627 30175
rect 28365 30141 28399 30175
rect 29009 30141 29043 30175
rect 29837 30141 29871 30175
rect 32781 30141 32815 30175
rect 34253 30141 34287 30175
rect 34621 30141 34655 30175
rect 34713 30141 34747 30175
rect 35909 30141 35943 30175
rect 36068 30141 36102 30175
rect 36921 30141 36955 30175
rect 37841 30141 37875 30175
rect 38301 30141 38335 30175
rect 9413 30073 9447 30107
rect 10701 30073 10735 30107
rect 11529 30073 11563 30107
rect 15301 30073 15335 30107
rect 16957 30073 16991 30107
rect 19257 30073 19291 30107
rect 20453 30073 20487 30107
rect 24133 30073 24167 30107
rect 33333 30073 33367 30107
rect 35173 30073 35207 30107
rect 36461 30073 36495 30107
rect 37289 30073 37323 30107
rect 9505 30005 9539 30039
rect 14105 30005 14139 30039
rect 18521 30005 18555 30039
rect 20545 30005 20579 30039
rect 22937 30005 22971 30039
rect 27169 30005 27203 30039
rect 29101 30005 29135 30039
rect 31953 30005 31987 30039
rect 32137 30005 32171 30039
rect 35265 30005 35299 30039
rect 10977 29801 11011 29835
rect 13553 29801 13587 29835
rect 17601 29801 17635 29835
rect 19257 29801 19291 29835
rect 22753 29801 22787 29835
rect 23581 29801 23615 29835
rect 24869 29801 24903 29835
rect 28549 29801 28583 29835
rect 30665 29801 30699 29835
rect 33793 29801 33827 29835
rect 37289 29801 37323 29835
rect 31401 29733 31435 29767
rect 33885 29733 33919 29767
rect 37197 29733 37231 29767
rect 11621 29665 11655 29699
rect 12449 29665 12483 29699
rect 12909 29665 12943 29699
rect 13921 29665 13955 29699
rect 14565 29665 14599 29699
rect 14657 29665 14691 29699
rect 18797 29665 18831 29699
rect 18889 29665 18923 29699
rect 19901 29665 19935 29699
rect 20269 29665 20303 29699
rect 23397 29665 23431 29699
rect 24133 29665 24167 29699
rect 25421 29665 25455 29699
rect 27169 29665 27203 29699
rect 31309 29665 31343 29699
rect 32045 29665 32079 29699
rect 32781 29665 32815 29699
rect 33149 29665 33183 29699
rect 35173 29665 35207 29699
rect 37841 29665 37875 29699
rect 38301 29665 38335 29699
rect 6009 29597 6043 29631
rect 6745 29597 6779 29631
rect 9597 29597 9631 29631
rect 9864 29597 9898 29631
rect 18153 29597 18187 29631
rect 19717 29597 19751 29631
rect 23213 29597 23247 29631
rect 25237 29597 25271 29631
rect 27436 29597 27470 29631
rect 31769 29597 31803 29631
rect 33425 29597 33459 29631
rect 34437 29597 34471 29631
rect 35817 29597 35851 29631
rect 37657 29597 37691 29631
rect 9505 29529 9539 29563
rect 11437 29529 11471 29563
rect 11897 29529 11931 29563
rect 17509 29529 17543 29563
rect 23121 29529 23155 29563
rect 26801 29529 26835 29563
rect 30573 29529 30607 29563
rect 31861 29529 31895 29563
rect 33333 29529 33367 29563
rect 35725 29529 35759 29563
rect 36062 29529 36096 29563
rect 5365 29461 5399 29495
rect 6193 29461 6227 29495
rect 8769 29461 8803 29495
rect 11069 29461 11103 29495
rect 11529 29461 11563 29495
rect 14749 29461 14783 29495
rect 15117 29461 15151 29495
rect 18337 29461 18371 29495
rect 18705 29461 18739 29495
rect 19625 29461 19659 29495
rect 24685 29461 24719 29495
rect 25329 29461 25363 29495
rect 25973 29461 26007 29495
rect 26433 29461 26467 29495
rect 32229 29461 32263 29495
rect 32597 29461 32631 29495
rect 32689 29461 32723 29495
rect 34897 29461 34931 29495
rect 37749 29461 37783 29495
rect 5917 29257 5951 29291
rect 10149 29257 10183 29291
rect 14289 29257 14323 29291
rect 17509 29257 17543 29291
rect 18245 29257 18279 29291
rect 18705 29257 18739 29291
rect 31309 29257 31343 29291
rect 32965 29257 32999 29291
rect 34897 29257 34931 29291
rect 36369 29257 36403 29291
rect 36829 29257 36863 29291
rect 6377 29189 6411 29223
rect 11529 29189 11563 29223
rect 32413 29189 32447 29223
rect 5825 29121 5859 29155
rect 9036 29121 9070 29155
rect 10241 29121 10275 29155
rect 10885 29121 10919 29155
rect 11345 29121 11379 29155
rect 13277 29121 13311 29155
rect 18153 29121 18187 29155
rect 18613 29121 18647 29155
rect 19073 29121 19107 29155
rect 19625 29121 19659 29155
rect 31953 29121 31987 29155
rect 32505 29121 32539 29155
rect 33517 29121 33551 29155
rect 35265 29121 35299 29155
rect 36461 29121 36495 29155
rect 5365 29053 5399 29087
rect 6101 29053 6135 29087
rect 6929 29053 6963 29087
rect 8769 29053 8803 29087
rect 14933 29053 14967 29087
rect 17417 29053 17451 29087
rect 18797 29053 18831 29087
rect 32229 29053 32263 29087
rect 33885 29053 33919 29087
rect 36185 29053 36219 29087
rect 37841 29053 37875 29087
rect 5457 28985 5491 29019
rect 7389 28985 7423 29019
rect 23673 28985 23707 29019
rect 24869 28985 24903 29019
rect 27169 28985 27203 29019
rect 30757 28985 30791 29019
rect 31125 28985 31159 29019
rect 32873 28985 32907 29019
rect 35909 28985 35943 29019
rect 37289 28985 37323 29019
rect 4629 28917 4663 28951
rect 4721 28917 4755 28951
rect 13737 28917 13771 28951
rect 3801 28509 3835 28543
rect 4997 28509 5031 28543
rect 6469 28509 6503 28543
rect 7205 28509 7239 28543
rect 9781 28509 9815 28543
rect 11069 28509 11103 28543
rect 14473 28509 14507 28543
rect 18061 28509 18095 28543
rect 19901 28509 19935 28543
rect 23489 28509 23523 28543
rect 24409 28509 24443 28543
rect 25053 28509 25087 28543
rect 27353 28509 27387 28543
rect 28089 28509 28123 28543
rect 28825 28509 28859 28543
rect 33517 28509 33551 28543
rect 34253 28509 34287 28543
rect 37933 28509 37967 28543
rect 5242 28441 5276 28475
rect 13645 28441 13679 28475
rect 31125 28441 31159 28475
rect 35357 28441 35391 28475
rect 35541 28441 35575 28475
rect 4445 28373 4479 28407
rect 4721 28373 4755 28407
rect 6377 28373 6411 28407
rect 7113 28373 7147 28407
rect 7849 28373 7883 28407
rect 10333 28373 10367 28407
rect 10517 28373 10551 28407
rect 14381 28373 14415 28407
rect 15117 28373 15151 28407
rect 18613 28373 18647 28407
rect 18981 28373 19015 28407
rect 19349 28373 19383 28407
rect 22845 28373 22879 28407
rect 23765 28373 23799 28407
rect 26801 28373 26835 28407
rect 27537 28373 27571 28407
rect 28273 28373 28307 28407
rect 29193 28373 29227 28407
rect 31033 28373 31067 28407
rect 32413 28373 32447 28407
rect 32965 28373 32999 28407
rect 33701 28373 33735 28407
rect 36829 28373 36863 28407
rect 37381 28373 37415 28407
rect 4261 28169 4295 28203
rect 6377 28169 6411 28203
rect 8125 28169 8159 28203
rect 9781 28169 9815 28203
rect 10241 28169 10275 28203
rect 14473 28169 14507 28203
rect 16865 28169 16899 28203
rect 18337 28169 18371 28203
rect 19257 28169 19291 28203
rect 22477 28169 22511 28203
rect 28825 28169 28859 28203
rect 32597 28169 32631 28203
rect 36277 28169 36311 28203
rect 7512 28101 7546 28135
rect 14933 28101 14967 28135
rect 17049 28101 17083 28135
rect 27252 28101 27286 28135
rect 35081 28101 35115 28135
rect 4353 28033 4387 28067
rect 5937 28033 5971 28067
rect 10149 28033 10183 28067
rect 14841 28033 14875 28067
rect 15301 28033 15335 28067
rect 19349 28033 19383 28067
rect 23590 28033 23624 28067
rect 24685 28033 24719 28067
rect 26985 28033 27019 28067
rect 28917 28033 28951 28067
rect 31125 28033 31159 28067
rect 32505 28033 32539 28067
rect 36369 28033 36403 28067
rect 2421 27965 2455 27999
rect 3617 27965 3651 27999
rect 4169 27965 4203 27999
rect 6193 27965 6227 27999
rect 7757 27965 7791 27999
rect 9689 27965 9723 27999
rect 10425 27965 10459 27999
rect 11161 27965 11195 27999
rect 11529 27965 11563 27999
rect 13645 27965 13679 27999
rect 14381 27965 14415 27999
rect 15025 27965 15059 27999
rect 15853 27965 15887 27999
rect 19073 27965 19107 27999
rect 20085 27965 20119 27999
rect 23857 27965 23891 27999
rect 24501 27965 24535 27999
rect 26617 27965 26651 27999
rect 28641 27965 28675 27999
rect 29929 27965 29963 27999
rect 31953 27965 31987 27999
rect 32689 27965 32723 27999
rect 33517 27965 33551 27999
rect 33793 27965 33827 27999
rect 34529 27965 34563 27999
rect 35265 27965 35299 27999
rect 36185 27965 36219 27999
rect 37013 27965 37047 27999
rect 37841 27965 37875 27999
rect 4721 27897 4755 27931
rect 8953 27897 8987 27931
rect 19717 27897 19751 27931
rect 25605 27897 25639 27931
rect 28365 27897 28399 27931
rect 29377 27897 29411 27931
rect 32137 27897 32171 27931
rect 36737 27897 36771 27931
rect 2973 27829 3007 27863
rect 3065 27829 3099 27863
rect 4813 27829 4847 27863
rect 9045 27829 9079 27863
rect 10609 27829 10643 27863
rect 12173 27829 12207 27863
rect 12817 27829 12851 27863
rect 13001 27829 13035 27863
rect 13737 27829 13771 27863
rect 20729 27829 20763 27863
rect 22385 27829 22419 27863
rect 23949 27829 23983 27863
rect 25329 27829 25363 27863
rect 26065 27829 26099 27863
rect 29285 27829 29319 27863
rect 31309 27829 31343 27863
rect 32965 27829 32999 27863
rect 34345 27829 34379 27863
rect 35817 27829 35851 27863
rect 37289 27829 37323 27863
rect 2789 27625 2823 27659
rect 18337 27625 18371 27659
rect 24225 27625 24259 27659
rect 27077 27625 27111 27659
rect 29009 27625 29043 27659
rect 29377 27625 29411 27659
rect 5089 27557 5123 27591
rect 7849 27557 7883 27591
rect 9321 27557 9355 27591
rect 17509 27557 17543 27591
rect 19257 27557 19291 27591
rect 32689 27557 32723 27591
rect 33517 27557 33551 27591
rect 34989 27557 35023 27591
rect 1961 27489 1995 27523
rect 3341 27489 3375 27523
rect 4261 27489 4295 27523
rect 4445 27489 4479 27523
rect 5365 27489 5399 27523
rect 5825 27489 5859 27523
rect 6239 27489 6273 27523
rect 7113 27489 7147 27523
rect 10701 27489 10735 27523
rect 11253 27489 11287 27523
rect 11345 27489 11379 27523
rect 13737 27489 13771 27523
rect 16037 27489 16071 27523
rect 16129 27489 16163 27523
rect 18889 27489 18923 27523
rect 20637 27489 20671 27523
rect 22017 27489 22051 27523
rect 23673 27489 23707 27523
rect 24869 27489 24903 27523
rect 25053 27489 25087 27523
rect 25513 27489 25547 27523
rect 27169 27489 27203 27523
rect 27813 27489 27847 27523
rect 28206 27489 28240 27523
rect 28365 27489 28399 27523
rect 31309 27489 31343 27523
rect 32873 27489 32907 27523
rect 33057 27489 33091 27523
rect 34161 27489 34195 27523
rect 2053 27421 2087 27455
rect 4721 27421 4755 27455
rect 5181 27421 5215 27455
rect 6101 27421 6135 27455
rect 6377 27421 6411 27455
rect 8401 27421 8435 27455
rect 10434 27421 10468 27455
rect 12265 27421 12299 27455
rect 13093 27421 13127 27455
rect 13553 27421 13587 27455
rect 15485 27421 15519 27455
rect 16589 27421 16623 27455
rect 17693 27421 17727 27455
rect 20381 27421 20415 27455
rect 21373 27421 21407 27455
rect 22284 27421 22318 27455
rect 25697 27421 25731 27455
rect 27353 27421 27387 27455
rect 28089 27421 28123 27455
rect 30113 27421 30147 27455
rect 31217 27421 31251 27455
rect 36645 27421 36679 27455
rect 38117 27421 38151 27455
rect 2697 27353 2731 27387
rect 3157 27353 3191 27387
rect 9229 27353 9263 27387
rect 13645 27353 13679 27387
rect 15240 27353 15274 27387
rect 18245 27353 18279 27387
rect 18797 27353 18831 27387
rect 20913 27353 20947 27387
rect 23857 27353 23891 27387
rect 25964 27353 25998 27387
rect 31576 27353 31610 27387
rect 33609 27353 33643 27387
rect 36400 27353 36434 27387
rect 37872 27353 37906 27387
rect 3249 27285 3283 27319
rect 4629 27285 4663 27319
rect 7021 27285 7055 27319
rect 7757 27285 7791 27319
rect 10793 27285 10827 27319
rect 11161 27285 11195 27319
rect 11621 27285 11655 27319
rect 12449 27285 12483 27319
rect 13185 27285 13219 27319
rect 14105 27285 14139 27319
rect 15577 27285 15611 27319
rect 15945 27285 15979 27319
rect 18705 27285 18739 27319
rect 21925 27285 21959 27319
rect 23397 27285 23431 27319
rect 23765 27285 23799 27319
rect 24409 27285 24443 27319
rect 24777 27285 24811 27319
rect 29561 27285 29595 27319
rect 30573 27285 30607 27319
rect 33149 27285 33183 27319
rect 35265 27285 35299 27319
rect 36737 27285 36771 27319
rect 3525 27081 3559 27115
rect 3985 27081 4019 27115
rect 6377 27081 6411 27115
rect 9413 27081 9447 27115
rect 11345 27081 11379 27115
rect 11897 27081 11931 27115
rect 12265 27081 12299 27115
rect 13829 27081 13863 27115
rect 15761 27081 15795 27115
rect 17049 27081 17083 27115
rect 21097 27081 21131 27115
rect 21833 27081 21867 27115
rect 22293 27081 22327 27115
rect 24501 27081 24535 27115
rect 24961 27081 24995 27115
rect 26065 27081 26099 27115
rect 26433 27081 26467 27115
rect 28365 27081 28399 27115
rect 28733 27081 28767 27115
rect 29193 27081 29227 27115
rect 31953 27081 31987 27115
rect 34437 27081 34471 27115
rect 37289 27081 37323 27115
rect 3166 27013 3200 27047
rect 6193 27013 6227 27047
rect 8300 27013 8334 27047
rect 15853 27013 15887 27047
rect 26525 27013 26559 27047
rect 27252 27013 27286 27047
rect 30818 27013 30852 27047
rect 35348 27013 35382 27047
rect 37749 27013 37783 27047
rect 3433 26945 3467 26979
rect 3893 26945 3927 26979
rect 4445 26945 4479 26979
rect 7501 26945 7535 26979
rect 7757 26945 7791 26979
rect 8033 26945 8067 26979
rect 9505 26945 9539 26979
rect 10425 26945 10459 26979
rect 10542 26945 10576 26979
rect 12449 26945 12483 26979
rect 12716 26945 12750 26979
rect 14105 26945 14139 26979
rect 14841 26945 14875 26979
rect 14958 26945 14992 26979
rect 18357 26945 18391 26979
rect 18613 26945 18647 26979
rect 18705 26945 18739 26979
rect 18889 26945 18923 26979
rect 20545 26945 20579 26979
rect 21005 26945 21039 26979
rect 22201 26945 22235 26979
rect 22845 26945 22879 26979
rect 25605 26945 25639 26979
rect 26985 26945 27019 26979
rect 28825 26945 28859 26979
rect 29561 26945 29595 26979
rect 29653 26945 29687 26979
rect 32781 26945 32815 26979
rect 32940 26945 32974 26979
rect 33057 26945 33091 26979
rect 33977 26945 34011 26979
rect 37657 26945 37691 26979
rect 4077 26877 4111 26911
rect 9689 26877 9723 26911
rect 10701 26877 10735 26911
rect 11713 26877 11747 26911
rect 11805 26877 11839 26911
rect 13921 26877 13955 26911
rect 15117 26877 15151 26911
rect 16405 26877 16439 26911
rect 19625 26877 19659 26911
rect 19742 26877 19776 26911
rect 19901 26877 19935 26911
rect 21281 26877 21315 26911
rect 22385 26877 22419 26911
rect 22661 26877 22695 26911
rect 23305 26877 23339 26911
rect 23581 26877 23615 26911
rect 23698 26877 23732 26911
rect 23857 26877 23891 26911
rect 24685 26877 24719 26911
rect 24869 26877 24903 26911
rect 26617 26877 26651 26911
rect 28641 26877 28675 26911
rect 29377 26877 29411 26911
rect 30297 26877 30331 26911
rect 30573 26877 30607 26911
rect 33793 26877 33827 26911
rect 34529 26877 34563 26911
rect 34713 26877 34747 26911
rect 35081 26877 35115 26911
rect 37841 26877 37875 26911
rect 38301 26877 38335 26911
rect 10149 26809 10183 26843
rect 14565 26809 14599 26843
rect 19349 26809 19383 26843
rect 25329 26809 25363 26843
rect 33333 26809 33367 26843
rect 36461 26809 36495 26843
rect 2053 26741 2087 26775
rect 17233 26741 17267 26775
rect 20637 26741 20671 26775
rect 30021 26741 30055 26775
rect 32137 26741 32171 26775
rect 34069 26741 34103 26775
rect 36737 26741 36771 26775
rect 7113 26537 7147 26571
rect 9505 26537 9539 26571
rect 13185 26537 13219 26571
rect 14105 26537 14139 26571
rect 17601 26537 17635 26571
rect 24409 26537 24443 26571
rect 26525 26537 26559 26571
rect 29193 26537 29227 26571
rect 32597 26537 32631 26571
rect 34989 26537 35023 26571
rect 3617 26469 3651 26503
rect 4445 26469 4479 26503
rect 6009 26469 6043 26503
rect 8769 26469 8803 26503
rect 19073 26469 19107 26503
rect 23305 26469 23339 26503
rect 27077 26469 27111 26503
rect 32505 26469 32539 26503
rect 3801 26401 3835 26435
rect 4838 26401 4872 26435
rect 4997 26401 5031 26435
rect 6561 26401 6595 26435
rect 11529 26401 11563 26435
rect 13645 26401 13679 26435
rect 13737 26401 13771 26435
rect 15485 26401 15519 26435
rect 20637 26401 20671 26435
rect 21833 26401 21867 26435
rect 23949 26401 23983 26435
rect 25697 26401 25731 26435
rect 28457 26401 28491 26435
rect 31125 26401 31159 26435
rect 33977 26401 34011 26435
rect 35541 26401 35575 26435
rect 36461 26401 36495 26435
rect 36620 26401 36654 26435
rect 37013 26401 37047 26435
rect 37473 26401 37507 26435
rect 37657 26401 37691 26435
rect 38301 26401 38335 26435
rect 2237 26333 2271 26367
rect 2504 26333 2538 26367
rect 3985 26333 4019 26367
rect 4721 26333 4755 26367
rect 6745 26333 6779 26367
rect 7481 26333 7515 26367
rect 10885 26333 10919 26367
rect 12541 26333 12575 26367
rect 15218 26333 15252 26367
rect 16129 26333 16163 26367
rect 17693 26333 17727 26367
rect 21281 26333 21315 26367
rect 22089 26333 22123 26367
rect 24961 26333 24995 26367
rect 28549 26333 28583 26367
rect 30113 26333 30147 26367
rect 31392 26333 31426 26367
rect 34253 26333 34287 26367
rect 36737 26333 36771 26367
rect 6653 26265 6687 26299
rect 9321 26265 9355 26299
rect 10640 26265 10674 26299
rect 12265 26265 12299 26299
rect 17960 26265 17994 26299
rect 20392 26265 20426 26299
rect 20729 26265 20763 26299
rect 23765 26265 23799 26299
rect 25145 26265 25179 26299
rect 26065 26265 26099 26299
rect 26801 26265 26835 26299
rect 28212 26265 28246 26299
rect 29561 26265 29595 26299
rect 30941 26265 30975 26299
rect 33732 26265 33766 26299
rect 35357 26265 35391 26299
rect 35817 26265 35851 26299
rect 38117 26265 38151 26299
rect 38209 26265 38243 26299
rect 5641 26197 5675 26231
rect 7757 26197 7791 26231
rect 10977 26197 11011 26231
rect 11345 26197 11379 26231
rect 11437 26197 11471 26231
rect 13093 26197 13127 26231
rect 13553 26197 13587 26231
rect 15577 26197 15611 26231
rect 19257 26197 19291 26231
rect 23213 26197 23247 26231
rect 23673 26197 23707 26231
rect 35449 26197 35483 26231
rect 37749 26197 37783 26231
rect 3433 25993 3467 26027
rect 6745 25993 6779 26027
rect 6837 25993 6871 26027
rect 7481 25993 7515 26027
rect 10241 25993 10275 26027
rect 10701 25993 10735 26027
rect 11529 25993 11563 26027
rect 14841 25993 14875 26027
rect 17601 25993 17635 26027
rect 20085 25993 20119 26027
rect 27169 25993 27203 26027
rect 27353 25993 27387 26027
rect 27813 25993 27847 26027
rect 28457 25993 28491 26027
rect 31585 25993 31619 26027
rect 32137 25993 32171 26027
rect 32505 25993 32539 26027
rect 33333 25993 33367 26027
rect 33977 25993 34011 26027
rect 37289 25993 37323 26027
rect 38209 25993 38243 26027
rect 11253 25925 11287 25959
rect 13338 25925 13372 25959
rect 22968 25925 23002 25959
rect 32597 25925 32631 25959
rect 35449 25925 35483 25959
rect 35900 25925 35934 25959
rect 1961 25857 1995 25891
rect 2217 25857 2251 25891
rect 4557 25857 4591 25891
rect 4813 25857 4847 25891
rect 5457 25857 5491 25891
rect 8769 25857 8803 25891
rect 9036 25857 9070 25891
rect 10609 25857 10643 25891
rect 13093 25857 13127 25891
rect 14933 25857 14967 25891
rect 18705 25857 18739 25891
rect 18797 25857 18831 25891
rect 19717 25857 19751 25891
rect 20177 25857 20211 25891
rect 20729 25857 20763 25891
rect 23305 25857 23339 25891
rect 27721 25857 27755 25891
rect 34529 25857 34563 25891
rect 35633 25857 35667 25891
rect 37841 25857 37875 25891
rect 7021 25789 7055 25823
rect 10885 25789 10919 25823
rect 12081 25789 12115 25823
rect 14749 25789 14783 25823
rect 18245 25789 18279 25823
rect 18889 25789 18923 25823
rect 19441 25789 19475 25823
rect 19625 25789 19659 25823
rect 23213 25789 23247 25823
rect 27905 25789 27939 25823
rect 32689 25789 32723 25823
rect 33057 25789 33091 25823
rect 33241 25789 33275 25823
rect 10149 25721 10183 25755
rect 14473 25721 14507 25755
rect 15301 25721 15335 25755
rect 18337 25721 18371 25755
rect 34897 25721 34931 25755
rect 37013 25721 37047 25755
rect 3341 25653 3375 25687
rect 4905 25653 4939 25687
rect 6101 25653 6135 25687
rect 6377 25653 6411 25687
rect 17417 25653 17451 25687
rect 21833 25653 21867 25687
rect 24777 25653 24811 25687
rect 25329 25653 25363 25687
rect 31953 25653 31987 25687
rect 33701 25653 33735 25687
rect 2053 25449 2087 25483
rect 5825 25449 5859 25483
rect 10057 25449 10091 25483
rect 14473 25449 14507 25483
rect 19257 25449 19291 25483
rect 23581 25449 23615 25483
rect 24225 25449 24259 25483
rect 24685 25449 24719 25483
rect 32873 25449 32907 25483
rect 35081 25449 35115 25483
rect 35449 25449 35483 25483
rect 36277 25449 36311 25483
rect 38025 25449 38059 25483
rect 2789 25381 2823 25415
rect 3985 25381 4019 25415
rect 13829 25381 13863 25415
rect 18981 25381 19015 25415
rect 2697 25313 2731 25347
rect 3433 25313 3467 25347
rect 4629 25313 4663 25347
rect 5365 25313 5399 25347
rect 10701 25313 10735 25347
rect 19809 25313 19843 25347
rect 22937 25313 22971 25347
rect 29377 25313 29411 25347
rect 35725 25313 35759 25347
rect 36461 25313 36495 25347
rect 37473 25313 37507 25347
rect 4353 25245 4387 25279
rect 7021 25245 7055 25279
rect 8401 25245 8435 25279
rect 13277 25245 13311 25279
rect 16957 25245 16991 25279
rect 18061 25245 18095 25279
rect 26433 25245 26467 25279
rect 29009 25245 29043 25279
rect 30205 25245 30239 25279
rect 36737 25245 36771 25279
rect 3249 25177 3283 25211
rect 4813 25177 4847 25211
rect 9965 25177 9999 25211
rect 36645 25177 36679 25211
rect 3157 25109 3191 25143
rect 4445 25109 4479 25143
rect 7573 25109 7607 25143
rect 7757 25109 7791 25143
rect 11069 25109 11103 25143
rect 12725 25109 12759 25143
rect 16405 25109 16439 25143
rect 18613 25109 18647 25143
rect 25789 25109 25823 25143
rect 29561 25109 29595 25143
rect 37105 25109 37139 25143
rect 4537 24905 4571 24939
rect 4905 24905 4939 24939
rect 7021 24905 7055 24939
rect 12541 24905 12575 24939
rect 29561 24905 29595 24939
rect 8033 24837 8067 24871
rect 24961 24837 24995 24871
rect 28733 24837 28767 24871
rect 30021 24837 30055 24871
rect 3985 24769 4019 24803
rect 7389 24769 7423 24803
rect 11897 24769 11931 24803
rect 12449 24769 12483 24803
rect 17805 24769 17839 24803
rect 18061 24769 18095 24803
rect 25053 24769 25087 24803
rect 25421 24769 25455 24803
rect 28825 24769 28859 24803
rect 30573 24769 30607 24803
rect 7481 24701 7515 24735
rect 7573 24701 7607 24735
rect 8861 24701 8895 24735
rect 8953 24701 8987 24735
rect 12725 24701 12759 24735
rect 13001 24701 13035 24735
rect 13737 24701 13771 24735
rect 16129 24701 16163 24735
rect 18337 24701 18371 24735
rect 18889 24701 18923 24735
rect 24501 24701 24535 24735
rect 25237 24701 25271 24735
rect 25973 24701 26007 24735
rect 26157 24701 26191 24735
rect 28917 24701 28951 24735
rect 29285 24701 29319 24735
rect 29469 24701 29503 24735
rect 31309 24701 31343 24735
rect 35081 24701 35115 24735
rect 35909 24701 35943 24735
rect 37013 24701 37047 24735
rect 37841 24701 37875 24735
rect 24593 24633 24627 24667
rect 27813 24633 27847 24667
rect 28273 24633 28307 24667
rect 3709 24565 3743 24599
rect 8217 24565 8251 24599
rect 9597 24565 9631 24599
rect 12081 24565 12115 24599
rect 13553 24565 13587 24599
rect 14289 24565 14323 24599
rect 15577 24565 15611 24599
rect 16681 24565 16715 24599
rect 23857 24565 23891 24599
rect 26801 24565 26835 24599
rect 28365 24565 28399 24599
rect 29929 24565 29963 24599
rect 30757 24565 30791 24599
rect 34529 24565 34563 24599
rect 35357 24565 35391 24599
rect 36369 24565 36403 24599
rect 37289 24565 37323 24599
rect 4813 24361 4847 24395
rect 6929 24361 6963 24395
rect 11897 24361 11931 24395
rect 15761 24361 15795 24395
rect 24133 24361 24167 24395
rect 24409 24361 24443 24395
rect 26617 24361 26651 24395
rect 27629 24361 27663 24395
rect 29377 24361 29411 24395
rect 30297 24361 30331 24395
rect 31125 24361 31159 24395
rect 34529 24361 34563 24395
rect 37749 24361 37783 24395
rect 15669 24293 15703 24327
rect 11253 24225 11287 24259
rect 15209 24225 15243 24259
rect 16313 24225 16347 24259
rect 25973 24225 26007 24259
rect 27997 24225 28031 24259
rect 29653 24225 29687 24259
rect 32413 24225 32447 24259
rect 36369 24225 36403 24259
rect 38393 24225 38427 24259
rect 3433 24157 3467 24191
rect 4445 24157 4479 24191
rect 6377 24157 6411 24191
rect 7021 24157 7055 24191
rect 9045 24157 9079 24191
rect 13277 24157 13311 24191
rect 14657 24157 14691 24191
rect 16129 24157 16163 24191
rect 17969 24157 18003 24191
rect 18613 24157 18647 24191
rect 25789 24157 25823 24191
rect 26157 24157 26191 24191
rect 26709 24157 26743 24191
rect 28264 24157 28298 24191
rect 29837 24157 29871 24191
rect 30941 24157 30975 24191
rect 31677 24157 31711 24191
rect 34897 24157 34931 24191
rect 35541 24157 35575 24191
rect 36185 24157 36219 24191
rect 36636 24157 36670 24191
rect 7266 24089 7300 24123
rect 13032 24089 13066 24123
rect 14105 24089 14139 24123
rect 16221 24089 16255 24123
rect 17724 24089 17758 24123
rect 18061 24089 18095 24123
rect 25544 24089 25578 24123
rect 29929 24089 29963 24123
rect 2881 24021 2915 24055
rect 3801 24021 3835 24055
rect 5181 24021 5215 24055
rect 8401 24021 8435 24055
rect 9689 24021 9723 24055
rect 11805 24021 11839 24055
rect 13645 24021 13679 24055
rect 16589 24021 16623 24055
rect 26249 24021 26283 24055
rect 27353 24021 27387 24055
rect 30389 24021 30423 24055
rect 31861 24021 31895 24055
rect 35633 24021 35667 24055
rect 37841 24021 37875 24055
rect 3249 23817 3283 23851
rect 6101 23817 6135 23851
rect 6653 23817 6687 23851
rect 8585 23817 8619 23851
rect 13921 23817 13955 23851
rect 14381 23817 14415 23851
rect 16497 23817 16531 23851
rect 18797 23817 18831 23851
rect 22109 23817 22143 23851
rect 27353 23817 27387 23851
rect 30481 23817 30515 23851
rect 36921 23817 36955 23851
rect 3617 23749 3651 23783
rect 5825 23749 5859 23783
rect 7472 23749 7506 23783
rect 9790 23749 9824 23783
rect 11345 23749 11379 23783
rect 13308 23749 13342 23783
rect 19257 23749 19291 23783
rect 23664 23749 23698 23783
rect 27445 23749 27479 23783
rect 30849 23749 30883 23783
rect 3709 23681 3743 23715
rect 6745 23681 6779 23715
rect 11989 23681 12023 23715
rect 14013 23681 14047 23715
rect 14933 23681 14967 23715
rect 15117 23681 15151 23715
rect 15384 23681 15418 23715
rect 16865 23681 16899 23715
rect 17902 23681 17936 23715
rect 18061 23681 18095 23715
rect 19165 23681 19199 23715
rect 24869 23681 24903 23715
rect 25789 23681 25823 23715
rect 26065 23681 26099 23715
rect 28365 23681 28399 23715
rect 29352 23681 29386 23715
rect 30205 23681 30239 23715
rect 30941 23681 30975 23715
rect 31309 23681 31343 23715
rect 34069 23681 34103 23715
rect 34336 23681 34370 23715
rect 35541 23681 35575 23715
rect 35808 23681 35842 23715
rect 37289 23681 37323 23715
rect 3065 23613 3099 23647
rect 3893 23613 3927 23647
rect 4629 23613 4663 23647
rect 4813 23613 4847 23647
rect 6469 23613 6503 23647
rect 7205 23613 7239 23647
rect 10057 23613 10091 23647
rect 13553 23613 13587 23647
rect 13737 23613 13771 23647
rect 17049 23613 17083 23647
rect 17785 23613 17819 23647
rect 19349 23613 19383 23647
rect 20177 23613 20211 23647
rect 23397 23613 23431 23647
rect 25053 23613 25087 23647
rect 25906 23613 25940 23647
rect 27537 23613 27571 23647
rect 29193 23613 29227 23647
rect 29469 23613 29503 23647
rect 30389 23613 30423 23647
rect 31033 23613 31067 23647
rect 31861 23613 31895 23647
rect 33885 23613 33919 23647
rect 37841 23613 37875 23647
rect 8677 23545 8711 23579
rect 17509 23545 17543 23579
rect 24777 23545 24811 23579
rect 25513 23545 25547 23579
rect 26709 23545 26743 23579
rect 29745 23545 29779 23579
rect 2513 23477 2547 23511
rect 4077 23477 4111 23511
rect 5457 23477 5491 23511
rect 7113 23477 7147 23511
rect 12173 23477 12207 23511
rect 18705 23477 18739 23511
rect 19625 23477 19659 23511
rect 22477 23477 22511 23511
rect 26985 23477 27019 23511
rect 27813 23477 27847 23511
rect 28549 23477 28583 23511
rect 33333 23477 33367 23511
rect 35449 23477 35483 23511
rect 38209 23477 38243 23511
rect 4629 23273 4663 23307
rect 5457 23273 5491 23307
rect 6837 23273 6871 23307
rect 8953 23273 8987 23307
rect 9965 23273 9999 23307
rect 10425 23273 10459 23307
rect 15485 23273 15519 23307
rect 16957 23273 16991 23307
rect 18429 23273 18463 23307
rect 27721 23273 27755 23307
rect 29285 23273 29319 23307
rect 29561 23273 29595 23307
rect 32597 23273 32631 23307
rect 34713 23273 34747 23307
rect 11989 23205 12023 23239
rect 18705 23205 18739 23239
rect 3985 23137 4019 23171
rect 4077 23137 4111 23171
rect 5181 23137 5215 23171
rect 6009 23137 6043 23171
rect 6285 23137 6319 23171
rect 7849 23137 7883 23171
rect 8125 23137 8159 23171
rect 8585 23137 8619 23171
rect 8769 23137 8803 23171
rect 9597 23137 9631 23171
rect 13001 23137 13035 23171
rect 13277 23137 13311 23171
rect 13737 23137 13771 23171
rect 14657 23137 14691 23171
rect 17877 23137 17911 23171
rect 19441 23137 19475 23171
rect 21833 23137 21867 23171
rect 23765 23137 23799 23171
rect 24133 23137 24167 23171
rect 25973 23137 26007 23171
rect 26157 23137 26191 23171
rect 27261 23137 27295 23171
rect 34069 23137 34103 23171
rect 35265 23137 35299 23171
rect 36599 23137 36633 23171
rect 36737 23137 36771 23171
rect 37013 23137 37047 23171
rect 37657 23137 37691 23171
rect 2237 23069 2271 23103
rect 2504 23069 2538 23103
rect 4169 23069 4203 23103
rect 4997 23069 5031 23103
rect 7573 23069 7607 23103
rect 7711 23069 7745 23103
rect 9321 23069 9355 23103
rect 10609 23069 10643 23103
rect 12725 23069 12759 23103
rect 12884 23069 12918 23103
rect 13921 23069 13955 23103
rect 15669 23069 15703 23103
rect 18061 23069 18095 23103
rect 21281 23069 21315 23103
rect 23029 23069 23063 23103
rect 24409 23069 24443 23103
rect 27905 23069 27939 23103
rect 28161 23069 28195 23103
rect 30941 23069 30975 23103
rect 33241 23069 33275 23103
rect 35081 23069 35115 23103
rect 36461 23069 36495 23103
rect 37473 23069 37507 23103
rect 38393 23069 38427 23103
rect 5089 23001 5123 23035
rect 10854 23001 10888 23035
rect 22017 23001 22051 23035
rect 24676 23001 24710 23035
rect 26709 23001 26743 23035
rect 30696 23001 30730 23035
rect 33885 23001 33919 23035
rect 3617 22933 3651 22967
rect 4537 22933 4571 22967
rect 6929 22933 6963 22967
rect 9413 22933 9447 22967
rect 12081 22933 12115 22967
rect 14105 22933 14139 22967
rect 17969 22933 18003 22967
rect 20729 22933 20763 22967
rect 21925 22933 21959 22967
rect 22385 22933 22419 22967
rect 22477 22933 22511 22967
rect 23489 22933 23523 22967
rect 25789 22933 25823 22967
rect 26249 22933 26283 22967
rect 26617 22933 26651 22967
rect 32689 22933 32723 22967
rect 33517 22933 33551 22967
rect 33977 22933 34011 22967
rect 35173 22933 35207 22967
rect 35817 22933 35851 22967
rect 37749 22933 37783 22967
rect 6561 22729 6595 22763
rect 8493 22729 8527 22763
rect 9873 22729 9907 22763
rect 10701 22729 10735 22763
rect 13001 22729 13035 22763
rect 13369 22729 13403 22763
rect 18061 22729 18095 22763
rect 20913 22729 20947 22763
rect 22201 22729 22235 22763
rect 22293 22729 22327 22763
rect 25973 22729 26007 22763
rect 26065 22729 26099 22763
rect 28089 22729 28123 22763
rect 28641 22729 28675 22763
rect 33793 22729 33827 22763
rect 36093 22729 36127 22763
rect 36645 22729 36679 22763
rect 37105 22729 37139 22763
rect 38025 22729 38059 22763
rect 2228 22661 2262 22695
rect 7674 22661 7708 22695
rect 8401 22661 8435 22695
rect 11796 22661 11830 22695
rect 13461 22661 13495 22695
rect 14013 22661 14047 22695
rect 24860 22661 24894 22695
rect 35725 22661 35759 22695
rect 36737 22661 36771 22695
rect 1961 22593 1995 22627
rect 4353 22593 4387 22627
rect 4470 22593 4504 22627
rect 5917 22593 5951 22627
rect 7941 22593 7975 22627
rect 9413 22593 9447 22627
rect 11529 22593 11563 22627
rect 16681 22593 16715 22627
rect 16948 22593 16982 22627
rect 18705 22593 18739 22627
rect 21281 22593 21315 22627
rect 22661 22593 22695 22627
rect 24593 22593 24627 22627
rect 26617 22593 26651 22627
rect 28181 22593 28215 22627
rect 29765 22593 29799 22627
rect 30021 22593 30055 22627
rect 32321 22593 32355 22627
rect 32588 22593 32622 22627
rect 34917 22593 34951 22627
rect 35173 22593 35207 22627
rect 37657 22593 37691 22627
rect 3433 22525 3467 22559
rect 3617 22525 3651 22559
rect 4629 22525 4663 22559
rect 5273 22525 5307 22559
rect 8585 22525 8619 22559
rect 11345 22525 11379 22559
rect 13645 22525 13679 22559
rect 20821 22525 20855 22559
rect 21373 22525 21407 22559
rect 21557 22525 21591 22559
rect 22477 22525 22511 22559
rect 23213 22525 23247 22559
rect 23949 22525 23983 22559
rect 27721 22525 27755 22559
rect 27997 22525 28031 22559
rect 35449 22525 35483 22559
rect 35633 22525 35667 22559
rect 36461 22525 36495 22559
rect 37381 22525 37415 22559
rect 37565 22525 37599 22559
rect 4077 22457 4111 22491
rect 12909 22457 12943 22491
rect 21833 22457 21867 22491
rect 3341 22389 3375 22423
rect 5365 22389 5399 22423
rect 8033 22389 8067 22423
rect 8861 22389 8895 22423
rect 18153 22389 18187 22423
rect 20177 22389 20211 22423
rect 23397 22389 23431 22423
rect 28549 22389 28583 22423
rect 30389 22389 30423 22423
rect 33701 22389 33735 22423
rect 38301 22389 38335 22423
rect 3801 22185 3835 22219
rect 5641 22185 5675 22219
rect 7389 22185 7423 22219
rect 11805 22185 11839 22219
rect 16773 22185 16807 22219
rect 17693 22185 17727 22219
rect 25697 22185 25731 22219
rect 26709 22185 26743 22219
rect 34253 22185 34287 22219
rect 35449 22185 35483 22219
rect 37841 22185 37875 22219
rect 33885 22117 33919 22151
rect 37749 22117 37783 22151
rect 5181 22049 5215 22083
rect 8033 22049 8067 22083
rect 8493 22049 8527 22083
rect 12357 22049 12391 22083
rect 13185 22049 13219 22083
rect 16957 22049 16991 22083
rect 17141 22049 17175 22083
rect 19717 22049 19751 22083
rect 22405 22049 22439 22083
rect 22845 22049 22879 22083
rect 23765 22049 23799 22083
rect 26065 22049 26099 22083
rect 28365 22049 28399 22083
rect 32505 22049 32539 22083
rect 34805 22049 34839 22083
rect 35725 22049 35759 22083
rect 38393 22049 38427 22083
rect 2237 21981 2271 22015
rect 7757 21981 7791 22015
rect 11621 21981 11655 22015
rect 18245 21981 18279 22015
rect 19984 21981 20018 22015
rect 21833 21981 21867 22015
rect 21992 21981 22026 22015
rect 22109 21981 22143 22015
rect 23029 21981 23063 22015
rect 24409 21981 24443 22015
rect 24961 21981 24995 22015
rect 31861 21981 31895 22015
rect 36369 21981 36403 22015
rect 36636 21981 36670 22015
rect 2504 21913 2538 21947
rect 4936 21913 4970 21947
rect 12173 21913 12207 21947
rect 12633 21913 12667 21947
rect 32772 21913 32806 21947
rect 35081 21913 35115 21947
rect 35909 21913 35943 21947
rect 3617 21845 3651 21879
rect 6009 21845 6043 21879
rect 7849 21845 7883 21879
rect 10885 21845 10919 21879
rect 11069 21845 11103 21879
rect 12265 21845 12299 21879
rect 17233 21845 17267 21879
rect 17601 21845 17635 21879
rect 18705 21845 18739 21879
rect 21097 21845 21131 21879
rect 21189 21845 21223 21879
rect 23121 21845 23155 21879
rect 23489 21845 23523 21879
rect 23581 21845 23615 21879
rect 24225 21845 24259 21879
rect 32413 21845 32447 21879
rect 34989 21845 35023 21879
rect 35817 21845 35851 21879
rect 36277 21845 36311 21879
rect 2973 21641 3007 21675
rect 4261 21641 4295 21675
rect 7941 21641 7975 21675
rect 13829 21641 13863 21675
rect 21649 21641 21683 21675
rect 22569 21641 22603 21675
rect 24133 21641 24167 21675
rect 32781 21641 32815 21675
rect 33149 21641 33183 21675
rect 35449 21641 35483 21675
rect 37565 21641 37599 21675
rect 3341 21573 3375 21607
rect 20536 21573 20570 21607
rect 33241 21573 33275 21607
rect 37657 21573 37691 21607
rect 5549 21505 5583 21539
rect 12173 21505 12207 21539
rect 13461 21505 13495 21539
rect 16497 21505 16531 21539
rect 17141 21505 17175 21539
rect 17233 21505 17267 21539
rect 18521 21505 18555 21539
rect 23857 21505 23891 21539
rect 29929 21505 29963 21539
rect 32689 21505 32723 21539
rect 33793 21505 33827 21539
rect 34805 21505 34839 21539
rect 36093 21505 36127 21539
rect 3433 21437 3467 21471
rect 3617 21437 3651 21471
rect 10609 21437 10643 21471
rect 11345 21437 11379 21471
rect 12265 21437 12299 21471
rect 12357 21437 12391 21471
rect 15853 21437 15887 21471
rect 17325 21437 17359 21471
rect 17877 21437 17911 21471
rect 19165 21437 19199 21471
rect 20269 21437 20303 21471
rect 29653 21437 29687 21471
rect 29837 21437 29871 21471
rect 30389 21437 30423 21471
rect 30941 21437 30975 21471
rect 31769 21437 31803 21471
rect 33333 21437 33367 21471
rect 33609 21437 33643 21471
rect 34529 21437 34563 21471
rect 34646 21437 34680 21471
rect 36277 21437 36311 21471
rect 36829 21437 36863 21471
rect 37473 21437 37507 21471
rect 11805 21369 11839 21403
rect 15761 21369 15795 21403
rect 18613 21369 18647 21403
rect 30297 21369 30331 21403
rect 34253 21369 34287 21403
rect 35541 21369 35575 21403
rect 5825 21301 5859 21335
rect 9965 21301 9999 21335
rect 10701 21301 10735 21335
rect 12909 21301 12943 21335
rect 16773 21301 16807 21335
rect 19625 21301 19659 21335
rect 24593 21301 24627 21335
rect 29377 21301 29411 21335
rect 31125 21301 31159 21335
rect 38025 21301 38059 21335
rect 3801 21097 3835 21131
rect 10885 21097 10919 21131
rect 11713 21097 11747 21131
rect 16865 21097 16899 21131
rect 21741 21097 21775 21131
rect 23949 21097 23983 21131
rect 29377 21097 29411 21131
rect 30113 21097 30147 21131
rect 34161 21097 34195 21131
rect 36185 21097 36219 21131
rect 36737 21097 36771 21131
rect 37197 21097 37231 21131
rect 3617 21029 3651 21063
rect 19073 21029 19107 21063
rect 23213 21029 23247 21063
rect 37473 21029 37507 21063
rect 4445 20961 4479 20995
rect 11437 20961 11471 20995
rect 13645 20961 13679 20995
rect 13737 20961 13771 20995
rect 16773 20961 16807 20995
rect 18521 20961 18555 20995
rect 19717 20961 19751 20995
rect 19901 20961 19935 20995
rect 23305 20961 23339 20995
rect 27169 20961 27203 20995
rect 6653 20893 6687 20927
rect 7849 20893 7883 20927
rect 8309 20893 8343 20927
rect 11253 20893 11287 20927
rect 13093 20893 13127 20927
rect 14657 20893 14691 20927
rect 17989 20893 18023 20927
rect 18245 20893 18279 20927
rect 20361 20893 20395 20927
rect 21833 20893 21867 20927
rect 27261 20893 27295 20927
rect 31493 20893 31527 20927
rect 32781 20893 32815 20927
rect 33037 20893 33071 20927
rect 34437 20893 34471 20927
rect 7297 20825 7331 20859
rect 8953 20825 8987 20859
rect 11345 20825 11379 20859
rect 12826 20825 12860 20859
rect 14105 20825 14139 20859
rect 16037 20825 16071 20859
rect 20628 20825 20662 20859
rect 22100 20825 22134 20859
rect 25789 20825 25823 20859
rect 31226 20825 31260 20859
rect 34713 20825 34747 20859
rect 4813 20757 4847 20791
rect 7205 20757 7239 20791
rect 8677 20757 8711 20791
rect 10241 20757 10275 20791
rect 13185 20757 13219 20791
rect 13553 20757 13587 20791
rect 16129 20757 16163 20791
rect 18613 20757 18647 20791
rect 18705 20757 18739 20791
rect 19257 20757 19291 20791
rect 19625 20757 19659 20791
rect 26525 20757 26559 20791
rect 27905 20757 27939 20791
rect 29929 20757 29963 20791
rect 9781 20553 9815 20587
rect 11345 20553 11379 20587
rect 13737 20553 13771 20587
rect 15117 20553 15151 20587
rect 19073 20553 19107 20587
rect 19533 20553 19567 20587
rect 21925 20553 21959 20587
rect 26341 20553 26375 20587
rect 29837 20553 29871 20587
rect 31309 20553 31343 20587
rect 33333 20553 33367 20587
rect 34069 20553 34103 20587
rect 34989 20553 35023 20587
rect 3525 20485 3559 20519
rect 6920 20485 6954 20519
rect 10210 20485 10244 20519
rect 11805 20485 11839 20519
rect 16230 20485 16264 20519
rect 18981 20485 19015 20519
rect 30972 20485 31006 20519
rect 35357 20485 35391 20519
rect 3617 20417 3651 20451
rect 3985 20417 4019 20451
rect 8125 20417 8159 20451
rect 11897 20417 11931 20451
rect 12934 20417 12968 20451
rect 13093 20417 13127 20451
rect 14197 20417 14231 20451
rect 17141 20417 17175 20451
rect 18061 20417 18095 20451
rect 18178 20417 18212 20451
rect 18337 20417 18371 20451
rect 19441 20417 19475 20451
rect 22569 20417 22603 20451
rect 26249 20417 26283 20451
rect 27997 20417 28031 20451
rect 34621 20417 34655 20451
rect 3065 20349 3099 20383
rect 3801 20349 3835 20383
rect 4629 20349 4663 20383
rect 6653 20349 6687 20383
rect 8493 20349 8527 20383
rect 9965 20349 9999 20383
rect 12081 20349 12115 20383
rect 12541 20349 12575 20383
rect 12817 20349 12851 20383
rect 14013 20349 14047 20383
rect 14105 20349 14139 20383
rect 16497 20349 16531 20383
rect 17325 20349 17359 20383
rect 17785 20349 17819 20383
rect 19625 20349 19659 20383
rect 23305 20349 23339 20383
rect 23949 20349 23983 20383
rect 25789 20349 25823 20383
rect 26525 20349 26559 20383
rect 27629 20349 27663 20383
rect 31217 20349 31251 20383
rect 31861 20349 31895 20383
rect 3157 20281 3191 20315
rect 17049 20281 17083 20315
rect 24409 20281 24443 20315
rect 2421 20213 2455 20247
rect 4905 20213 4939 20247
rect 5549 20213 5583 20247
rect 8033 20213 8067 20247
rect 14565 20213 14599 20247
rect 22661 20213 22695 20247
rect 23397 20213 23431 20247
rect 25145 20213 25179 20247
rect 25881 20213 25915 20247
rect 26985 20213 27019 20247
rect 29285 20213 29319 20247
rect 3617 20009 3651 20043
rect 6837 20009 6871 20043
rect 9873 20009 9907 20043
rect 11989 20009 12023 20043
rect 17141 20009 17175 20043
rect 18981 20009 19015 20043
rect 23489 20009 23523 20043
rect 26893 20009 26927 20043
rect 27721 20009 27755 20043
rect 29377 20009 29411 20043
rect 22661 19941 22695 19975
rect 30757 19941 30791 19975
rect 2237 19873 2271 19907
rect 4445 19873 4479 19907
rect 6193 19873 6227 19907
rect 10609 19873 10643 19907
rect 13461 19873 13495 19907
rect 18613 19873 18647 19907
rect 19809 19873 19843 19907
rect 22109 19873 22143 19907
rect 22891 19873 22925 19907
rect 23029 19873 23063 19907
rect 24869 19873 24903 19907
rect 27077 19873 27111 19907
rect 27261 19873 27295 19907
rect 30205 19873 30239 19907
rect 30481 19873 30515 19907
rect 31401 19873 31435 19907
rect 33517 19873 33551 19907
rect 2504 19805 2538 19839
rect 4261 19805 4295 19839
rect 5181 19805 5215 19839
rect 6009 19805 6043 19839
rect 8309 19805 8343 19839
rect 9505 19805 9539 19839
rect 10865 19805 10899 19839
rect 14657 19805 14691 19839
rect 15761 19805 15795 19839
rect 21281 19805 21315 19839
rect 22293 19805 22327 19839
rect 24133 19805 24167 19839
rect 25513 19805 25547 19839
rect 27997 19805 28031 19839
rect 30364 19805 30398 19839
rect 31217 19805 31251 19839
rect 32045 19805 32079 19839
rect 32781 19805 32815 19839
rect 34529 19805 34563 19839
rect 35357 19805 35391 19839
rect 36093 19805 36127 19839
rect 36829 19805 36863 19839
rect 38485 19805 38519 19839
rect 4169 19737 4203 19771
rect 8064 19737 8098 19771
rect 8953 19737 8987 19771
rect 13216 19737 13250 19771
rect 14105 19737 14139 19771
rect 16028 19737 16062 19771
rect 18368 19737 18402 19771
rect 19257 19737 19291 19771
rect 23121 19737 23155 19771
rect 23581 19737 23615 19771
rect 24685 19737 24719 19771
rect 25780 19737 25814 19771
rect 28264 19737 28298 19771
rect 3801 19669 3835 19703
rect 4629 19669 4663 19703
rect 5365 19669 5399 19703
rect 6377 19669 6411 19703
rect 6469 19669 6503 19703
rect 6929 19669 6963 19703
rect 8677 19669 8711 19703
rect 12081 19669 12115 19703
rect 13829 19669 13863 19703
rect 17233 19669 17267 19703
rect 20729 19669 20763 19703
rect 21741 19669 21775 19703
rect 22201 19669 22235 19703
rect 25421 19669 25455 19703
rect 27353 19669 27387 19703
rect 29561 19669 29595 19703
rect 31493 19669 31527 19703
rect 32229 19669 32263 19703
rect 32965 19669 32999 19703
rect 33885 19669 33919 19703
rect 34713 19669 34747 19703
rect 35449 19669 35483 19703
rect 36185 19669 36219 19703
rect 37841 19669 37875 19703
rect 3249 19465 3283 19499
rect 5733 19465 5767 19499
rect 6193 19465 6227 19499
rect 12173 19465 12207 19499
rect 12725 19465 12759 19499
rect 13829 19465 13863 19499
rect 18705 19465 18739 19499
rect 20913 19465 20947 19499
rect 26709 19465 26743 19499
rect 30757 19465 30791 19499
rect 34437 19465 34471 19499
rect 34897 19465 34931 19499
rect 35357 19465 35391 19499
rect 36001 19465 36035 19499
rect 36461 19465 36495 19499
rect 5825 19397 5859 19431
rect 14381 19397 14415 19431
rect 14473 19397 14507 19431
rect 17325 19397 17359 19431
rect 22100 19397 22134 19431
rect 23305 19397 23339 19431
rect 24041 19397 24075 19431
rect 29276 19397 29310 19431
rect 37289 19397 37323 19431
rect 1869 19329 1903 19363
rect 2136 19329 2170 19363
rect 3341 19329 3375 19363
rect 4261 19329 4295 19363
rect 7732 19329 7766 19363
rect 8585 19329 8619 19363
rect 8769 19329 8803 19363
rect 9229 19329 9263 19363
rect 9689 19329 9723 19363
rect 12633 19329 12667 19363
rect 13185 19329 13219 19363
rect 18061 19329 18095 19363
rect 21281 19329 21315 19363
rect 21373 19329 21407 19363
rect 21833 19329 21867 19363
rect 25053 19329 25087 19363
rect 25309 19329 25343 19363
rect 26985 19329 27019 19363
rect 27169 19329 27203 19363
rect 27905 19329 27939 19363
rect 29009 19329 29043 19363
rect 30849 19329 30883 19363
rect 31861 19329 31895 19363
rect 34529 19329 34563 19363
rect 35265 19329 35299 19363
rect 36093 19329 36127 19363
rect 3525 19261 3559 19295
rect 4378 19261 4412 19295
rect 4537 19261 4571 19295
rect 5549 19261 5583 19295
rect 6929 19261 6963 19295
rect 7573 19261 7607 19295
rect 7849 19261 7883 19295
rect 9321 19261 9355 19295
rect 9505 19261 9539 19295
rect 10241 19261 10275 19295
rect 11345 19261 11379 19295
rect 12817 19261 12851 19295
rect 17417 19261 17451 19295
rect 17601 19261 17635 19295
rect 21465 19261 21499 19295
rect 23857 19261 23891 19295
rect 24593 19261 24627 19295
rect 28022 19261 28056 19295
rect 28181 19261 28215 19295
rect 30665 19261 30699 19295
rect 33977 19261 34011 19295
rect 34621 19261 34655 19295
rect 35449 19261 35483 19295
rect 35909 19261 35943 19295
rect 36737 19261 36771 19295
rect 37841 19261 37875 19295
rect 3985 19193 4019 19227
rect 8125 19193 8159 19227
rect 23213 19193 23247 19227
rect 26433 19193 26467 19227
rect 27629 19193 27663 19227
rect 30389 19193 30423 19227
rect 31217 19193 31251 19227
rect 33241 19193 33275 19227
rect 34069 19193 34103 19227
rect 5181 19125 5215 19159
rect 6653 19125 6687 19159
rect 8861 19125 8895 19159
rect 10701 19125 10735 19159
rect 11713 19125 11747 19159
rect 12265 19125 12299 19159
rect 15945 19125 15979 19159
rect 16957 19125 16991 19159
rect 28825 19125 28859 19159
rect 31309 19125 31343 19159
rect 33333 19125 33367 19159
rect 4629 18921 4663 18955
rect 8401 18921 8435 18955
rect 8769 18921 8803 18955
rect 12817 18921 12851 18955
rect 16497 18921 16531 18955
rect 17325 18921 17359 18955
rect 21373 18921 21407 18955
rect 23673 18921 23707 18955
rect 25145 18921 25179 18955
rect 26617 18921 26651 18955
rect 29285 18921 29319 18955
rect 31125 18921 31159 18955
rect 34529 18921 34563 18955
rect 38485 18921 38519 18955
rect 3617 18853 3651 18887
rect 2237 18785 2271 18819
rect 4445 18785 4479 18819
rect 5825 18785 5859 18819
rect 6009 18785 6043 18819
rect 6837 18785 6871 18819
rect 9505 18785 9539 18819
rect 12265 18785 12299 18819
rect 17049 18785 17083 18819
rect 17969 18785 18003 18819
rect 22268 18785 22302 18819
rect 22661 18785 22695 18819
rect 23121 18785 23155 18819
rect 25237 18785 25271 18819
rect 28089 18785 28123 18819
rect 30113 18785 30147 18819
rect 30573 18785 30607 18819
rect 31401 18785 31435 18819
rect 35817 18785 35851 18819
rect 35955 18785 35989 18819
rect 36369 18785 36403 18819
rect 37013 18785 37047 18819
rect 37105 18785 37139 18819
rect 1593 18717 1627 18751
rect 4169 18717 4203 18751
rect 5181 18717 5215 18751
rect 5733 18717 5767 18751
rect 7021 18717 7055 18751
rect 11529 18717 11563 18751
rect 19993 18717 20027 18751
rect 22109 18717 22143 18751
rect 22385 18717 22419 18751
rect 23305 18717 23339 18751
rect 25504 18717 25538 18751
rect 28733 18717 28767 18751
rect 30757 18717 30791 18751
rect 33149 18717 33183 18751
rect 33416 18717 33450 18751
rect 36093 18717 36127 18751
rect 36829 18717 36863 18751
rect 2145 18649 2179 18683
rect 2482 18649 2516 18683
rect 6561 18649 6595 18683
rect 7288 18649 7322 18683
rect 8953 18649 8987 18683
rect 20260 18649 20294 18683
rect 24041 18649 24075 18683
rect 27844 18649 27878 18683
rect 28181 18649 28215 18683
rect 29929 18649 29963 18683
rect 37372 18649 37406 18683
rect 3801 18581 3835 18615
rect 4261 18581 4295 18615
rect 5365 18581 5399 18615
rect 6193 18581 6227 18615
rect 6653 18581 6687 18615
rect 9873 18581 9907 18615
rect 10885 18581 10919 18615
rect 16405 18581 16439 18615
rect 21465 18581 21499 18615
rect 26709 18581 26743 18615
rect 29561 18581 29595 18615
rect 30021 18581 30055 18615
rect 30665 18581 30699 18615
rect 33057 18581 33091 18615
rect 34897 18581 34931 18615
rect 35173 18581 35207 18615
rect 5641 18377 5675 18411
rect 7757 18377 7791 18411
rect 10149 18377 10183 18411
rect 11529 18377 11563 18411
rect 11989 18377 12023 18411
rect 21649 18377 21683 18411
rect 25789 18377 25823 18411
rect 26249 18377 26283 18411
rect 27261 18377 27295 18411
rect 27721 18377 27755 18411
rect 28917 18377 28951 18411
rect 29929 18377 29963 18411
rect 30021 18377 30055 18411
rect 36461 18377 36495 18411
rect 37657 18377 37691 18411
rect 9597 18309 9631 18343
rect 22968 18309 23002 18343
rect 26157 18309 26191 18343
rect 2329 18241 2363 18275
rect 2596 18241 2630 18275
rect 4169 18241 4203 18275
rect 4629 18241 4663 18275
rect 6377 18241 6411 18275
rect 6644 18241 6678 18275
rect 11897 18241 11931 18275
rect 13093 18241 13127 18275
rect 20269 18241 20303 18275
rect 20536 18241 20570 18275
rect 24317 18241 24351 18275
rect 24593 18241 24627 18275
rect 27353 18241 27387 18275
rect 27813 18241 27847 18275
rect 29561 18241 29595 18275
rect 33517 18241 33551 18275
rect 33784 18241 33818 18275
rect 35081 18241 35115 18275
rect 35348 18241 35382 18275
rect 3893 18173 3927 18207
rect 4077 18173 4111 18207
rect 5181 18173 5215 18207
rect 11345 18173 11379 18207
rect 12081 18173 12115 18207
rect 12909 18173 12943 18207
rect 13645 18173 13679 18207
rect 15669 18173 15703 18207
rect 16497 18173 16531 18207
rect 17785 18173 17819 18207
rect 23213 18173 23247 18207
rect 23949 18173 23983 18207
rect 25697 18173 25731 18207
rect 26433 18173 26467 18207
rect 27169 18173 27203 18207
rect 28365 18173 28399 18207
rect 29745 18173 29779 18207
rect 37749 18173 37783 18207
rect 37841 18173 37875 18207
rect 38301 18173 38335 18207
rect 3709 18105 3743 18139
rect 4537 18105 4571 18139
rect 16957 18105 16991 18139
rect 6101 18037 6135 18071
rect 8309 18037 8343 18071
rect 10517 18037 10551 18071
rect 10701 18037 10735 18071
rect 12357 18037 12391 18071
rect 15117 18037 15151 18071
rect 15853 18037 15887 18071
rect 17233 18037 17267 18071
rect 21833 18037 21867 18071
rect 28733 18037 28767 18071
rect 30389 18037 30423 18071
rect 30757 18037 30791 18071
rect 34897 18037 34931 18071
rect 36737 18037 36771 18071
rect 37289 18037 37323 18071
rect 2973 17833 3007 17867
rect 3801 17833 3835 17867
rect 7113 17833 7147 17867
rect 15117 17833 15151 17867
rect 17417 17833 17451 17867
rect 20913 17833 20947 17867
rect 24685 17833 24719 17867
rect 26341 17833 26375 17867
rect 37381 17833 37415 17867
rect 7205 17765 7239 17799
rect 10241 17765 10275 17799
rect 17325 17765 17359 17799
rect 34713 17765 34747 17799
rect 36369 17765 36403 17799
rect 3617 17697 3651 17731
rect 4445 17697 4479 17731
rect 6469 17697 6503 17731
rect 7849 17697 7883 17731
rect 9597 17697 9631 17731
rect 10701 17697 10735 17731
rect 10793 17697 10827 17731
rect 12725 17697 12759 17731
rect 15669 17697 15703 17731
rect 18061 17697 18095 17731
rect 22109 17697 22143 17731
rect 22385 17697 22419 17731
rect 22569 17697 22603 17731
rect 23489 17697 23523 17731
rect 26893 17697 26927 17731
rect 27353 17697 27387 17731
rect 34529 17697 34563 17731
rect 35357 17697 35391 17731
rect 35633 17697 35667 17731
rect 37933 17697 37967 17731
rect 12193 17629 12227 17663
rect 12449 17629 12483 17663
rect 15945 17629 15979 17663
rect 27721 17629 27755 17663
rect 27997 17629 28031 17663
rect 35081 17629 35115 17663
rect 36921 17629 36955 17663
rect 4813 17561 4847 17595
rect 13645 17561 13679 17595
rect 16212 17561 16246 17595
rect 17785 17561 17819 17595
rect 19625 17561 19659 17595
rect 22661 17561 22695 17595
rect 24225 17561 24259 17595
rect 24961 17561 24995 17595
rect 35817 17561 35851 17595
rect 5089 17493 5123 17527
rect 10149 17493 10183 17527
rect 10609 17493 10643 17527
rect 11069 17493 11103 17527
rect 12817 17493 12851 17527
rect 12909 17493 12943 17527
rect 13277 17493 13311 17527
rect 14933 17493 14967 17527
rect 15485 17493 15519 17527
rect 15577 17493 15611 17527
rect 17877 17493 17911 17527
rect 18521 17493 18555 17527
rect 21465 17493 21499 17527
rect 21833 17493 21867 17527
rect 21925 17493 21959 17527
rect 23029 17493 23063 17527
rect 29745 17493 29779 17527
rect 33333 17493 33367 17527
rect 33793 17493 33827 17527
rect 33885 17493 33919 17527
rect 35173 17493 35207 17527
rect 35909 17493 35943 17527
rect 36277 17493 36311 17527
rect 4905 17289 4939 17323
rect 29193 17289 29227 17323
rect 34713 17289 34747 17323
rect 37657 17289 37691 17323
rect 4629 17221 4663 17255
rect 9505 17221 9539 17255
rect 15025 17221 15059 17255
rect 18613 17221 18647 17255
rect 20913 17221 20947 17255
rect 21833 17221 21867 17255
rect 33149 17221 33183 17255
rect 33600 17221 33634 17255
rect 4813 17153 4847 17187
rect 10221 17153 10255 17187
rect 14013 17153 14047 17187
rect 14473 17153 14507 17187
rect 15384 17153 15418 17187
rect 17315 17153 17349 17187
rect 18337 17153 18371 17187
rect 19165 17153 19199 17187
rect 21557 17153 21591 17187
rect 22385 17153 22419 17187
rect 29285 17153 29319 17187
rect 35081 17153 35115 17187
rect 36118 17153 36152 17187
rect 36921 17153 36955 17187
rect 37565 17153 37599 17187
rect 3433 17085 3467 17119
rect 4169 17085 4203 17119
rect 6193 17085 6227 17119
rect 7573 17085 7607 17119
rect 8309 17085 8343 17119
rect 9965 17085 9999 17119
rect 11529 17085 11563 17119
rect 11713 17085 11747 17119
rect 12449 17085 12483 17119
rect 12587 17085 12621 17119
rect 12725 17085 12759 17119
rect 15117 17085 15151 17119
rect 17463 17085 17497 17119
rect 17601 17085 17635 17119
rect 18521 17085 18555 17119
rect 23213 17085 23247 17119
rect 23857 17085 23891 17119
rect 26801 17085 26835 17119
rect 27629 17085 27663 17119
rect 28273 17085 28307 17119
rect 33333 17085 33367 17119
rect 35265 17085 35299 17119
rect 36001 17085 36035 17119
rect 36277 17085 36311 17119
rect 37473 17085 37507 17119
rect 38301 17085 38335 17119
rect 6653 17017 6687 17051
rect 8677 17017 8711 17051
rect 12173 17017 12207 17051
rect 13461 17017 13495 17051
rect 16497 17017 16531 17051
rect 17877 17017 17911 17051
rect 32781 17017 32815 17051
rect 35725 17017 35759 17051
rect 2789 16949 2823 16983
rect 3525 16949 3559 16983
rect 5273 16949 5307 16983
rect 5549 16949 5583 16983
rect 6929 16949 6963 16983
rect 7665 16949 7699 16983
rect 9781 16949 9815 16983
rect 11345 16949 11379 16983
rect 13369 16949 13403 16983
rect 16681 16949 16715 16983
rect 22569 16949 22603 16983
rect 23305 16949 23339 16983
rect 24317 16949 24351 16983
rect 26341 16949 26375 16983
rect 26985 16949 27019 16983
rect 27721 16949 27755 16983
rect 30389 16949 30423 16983
rect 38025 16949 38059 16983
rect 3617 16745 3651 16779
rect 7021 16745 7055 16779
rect 7849 16745 7883 16779
rect 12909 16745 12943 16779
rect 16221 16745 16255 16779
rect 16589 16745 16623 16779
rect 18061 16745 18095 16779
rect 21189 16745 21223 16779
rect 23121 16745 23155 16779
rect 24685 16745 24719 16779
rect 25973 16745 26007 16779
rect 26801 16745 26835 16779
rect 11437 16677 11471 16711
rect 37749 16677 37783 16711
rect 2053 16609 2087 16643
rect 2973 16609 3007 16643
rect 3157 16609 3191 16643
rect 4445 16609 4479 16643
rect 7297 16609 7331 16643
rect 9965 16609 9999 16643
rect 12817 16609 12851 16643
rect 14841 16609 14875 16643
rect 16681 16609 16715 16643
rect 22477 16609 22511 16643
rect 22661 16609 22695 16643
rect 24041 16609 24075 16643
rect 26157 16609 26191 16643
rect 26341 16609 26375 16643
rect 27353 16609 27387 16643
rect 27445 16609 27479 16643
rect 28181 16609 28215 16643
rect 28273 16609 28307 16643
rect 29101 16609 29135 16643
rect 30113 16609 30147 16643
rect 33149 16609 33183 16643
rect 36093 16609 36127 16643
rect 36369 16609 36403 16643
rect 2145 16541 2179 16575
rect 4997 16541 5031 16575
rect 5641 16541 5675 16575
rect 8493 16541 8527 16575
rect 10232 16541 10266 16575
rect 13461 16541 13495 16575
rect 15108 16541 15142 16575
rect 16948 16541 16982 16575
rect 18153 16541 18187 16575
rect 18705 16541 18739 16575
rect 22293 16541 22327 16575
rect 23213 16541 23247 16575
rect 25329 16541 25363 16575
rect 30481 16541 30515 16575
rect 32597 16541 32631 16575
rect 38393 16541 38427 16575
rect 3249 16473 3283 16507
rect 4169 16473 4203 16507
rect 5549 16473 5583 16507
rect 5886 16473 5920 16507
rect 7389 16473 7423 16507
rect 7941 16473 7975 16507
rect 12572 16473 12606 16507
rect 21281 16473 21315 16507
rect 27261 16473 27295 16507
rect 28549 16473 28583 16507
rect 30748 16473 30782 16507
rect 31953 16473 31987 16507
rect 33416 16473 33450 16507
rect 35848 16473 35882 16507
rect 36636 16473 36670 16507
rect 37841 16473 37875 16507
rect 2789 16405 2823 16439
rect 3801 16405 3835 16439
rect 4261 16405 4295 16439
rect 7481 16405 7515 16439
rect 11345 16405 11379 16439
rect 22753 16405 22787 16439
rect 25145 16405 25179 16439
rect 26433 16405 26467 16439
rect 26893 16405 26927 16439
rect 27721 16405 27755 16439
rect 28089 16405 28123 16439
rect 29561 16405 29595 16439
rect 31861 16405 31895 16439
rect 34529 16405 34563 16439
rect 34713 16405 34747 16439
rect 5457 16201 5491 16235
rect 5825 16201 5859 16235
rect 7849 16201 7883 16235
rect 7941 16201 7975 16235
rect 10517 16201 10551 16235
rect 12357 16201 12391 16235
rect 16221 16201 16255 16235
rect 17417 16201 17451 16235
rect 26341 16201 26375 16235
rect 29929 16201 29963 16235
rect 34713 16201 34747 16235
rect 36001 16201 36035 16235
rect 36093 16201 36127 16235
rect 37105 16201 37139 16235
rect 38025 16201 38059 16235
rect 2596 16133 2630 16167
rect 6736 16133 6770 16167
rect 16129 16133 16163 16167
rect 17049 16133 17083 16167
rect 18521 16133 18555 16167
rect 23060 16133 23094 16167
rect 28641 16133 28675 16167
rect 1685 16065 1719 16099
rect 4721 16065 4755 16099
rect 8309 16065 8343 16099
rect 8769 16065 8803 16099
rect 10793 16065 10827 16099
rect 11345 16065 11379 16099
rect 11897 16065 11931 16099
rect 11989 16065 12023 16099
rect 18153 16065 18187 16099
rect 23305 16065 23339 16099
rect 24521 16065 24555 16099
rect 24777 16065 24811 16099
rect 25053 16065 25087 16099
rect 26985 16065 27019 16099
rect 27252 16065 27286 16099
rect 30748 16065 30782 16099
rect 32137 16065 32171 16099
rect 34161 16065 34195 16099
rect 35357 16065 35391 16099
rect 36645 16065 36679 16099
rect 37657 16065 37691 16099
rect 2329 15997 2363 16031
rect 4537 15997 4571 16031
rect 5917 15997 5951 16031
rect 6101 15997 6135 16031
rect 6469 15997 6503 16031
rect 8401 15997 8435 16031
rect 8585 15997 8619 16031
rect 9321 15997 9355 16031
rect 11713 15997 11747 16031
rect 15301 15997 15335 16031
rect 16313 15997 16347 16031
rect 16773 15997 16807 16031
rect 16957 15997 16991 16031
rect 17509 15997 17543 16031
rect 30481 15997 30515 16031
rect 32689 15997 32723 16031
rect 33425 15997 33459 16031
rect 34805 15997 34839 16031
rect 34989 15997 35023 16031
rect 37381 15997 37415 16031
rect 37565 15997 37599 16031
rect 5365 15929 5399 15963
rect 15577 15929 15611 15963
rect 31861 15929 31895 15963
rect 2237 15861 2271 15895
rect 3709 15861 3743 15895
rect 15761 15861 15795 15895
rect 21925 15861 21959 15895
rect 23397 15861 23431 15895
rect 28365 15861 28399 15895
rect 32873 15861 32907 15895
rect 33609 15861 33643 15895
rect 34345 15861 34379 15895
rect 2145 15657 2179 15691
rect 5733 15657 5767 15691
rect 10057 15657 10091 15691
rect 15577 15657 15611 15691
rect 27445 15657 27479 15691
rect 33885 15657 33919 15691
rect 34713 15657 34747 15691
rect 35725 15657 35759 15691
rect 36369 15657 36403 15691
rect 37749 15657 37783 15691
rect 7665 15589 7699 15623
rect 12081 15589 12115 15623
rect 27537 15589 27571 15623
rect 32413 15589 32447 15623
rect 1593 15521 1627 15555
rect 4445 15521 4479 15555
rect 4838 15521 4872 15555
rect 4997 15521 5031 15555
rect 8125 15521 8159 15555
rect 8309 15521 8343 15555
rect 11989 15521 12023 15555
rect 12725 15521 12759 15555
rect 16129 15521 16163 15555
rect 16957 15521 16991 15555
rect 17049 15521 17083 15555
rect 17877 15521 17911 15555
rect 18337 15521 18371 15555
rect 23581 15521 23615 15555
rect 23765 15521 23799 15555
rect 25697 15521 25731 15555
rect 26065 15521 26099 15555
rect 29377 15521 29411 15555
rect 30297 15521 30331 15555
rect 31125 15521 31159 15555
rect 31401 15521 31435 15555
rect 31677 15521 31711 15555
rect 32137 15521 32171 15555
rect 32965 15521 32999 15555
rect 33425 15521 33459 15555
rect 34437 15521 34471 15555
rect 35357 15521 35391 15555
rect 38301 15521 38335 15555
rect 2237 15453 2271 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4721 15453 4755 15487
rect 6285 15453 6319 15487
rect 7113 15453 7147 15487
rect 7251 15453 7285 15487
rect 7389 15453 7423 15487
rect 11253 15453 11287 15487
rect 13461 15453 13495 15487
rect 17785 15453 17819 15487
rect 18521 15453 18555 15487
rect 19993 15453 20027 15487
rect 21649 15453 21683 15487
rect 23489 15453 23523 15487
rect 24869 15453 24903 15487
rect 26332 15453 26366 15487
rect 28661 15453 28695 15487
rect 28917 15453 28951 15487
rect 31263 15453 31297 15487
rect 32321 15453 32355 15487
rect 2504 15385 2538 15419
rect 8677 15385 8711 15419
rect 9965 15385 9999 15419
rect 12449 15385 12483 15419
rect 15485 15385 15519 15419
rect 21916 15385 21950 15419
rect 24685 15385 24719 15419
rect 30021 15385 30055 15419
rect 36461 15385 36495 15419
rect 1685 15317 1719 15351
rect 1777 15317 1811 15351
rect 3617 15317 3651 15351
rect 5641 15317 5675 15351
rect 6469 15317 6503 15351
rect 9229 15317 9263 15351
rect 11345 15317 11379 15351
rect 12541 15317 12575 15351
rect 12909 15317 12943 15351
rect 15025 15317 15059 15351
rect 16497 15317 16531 15351
rect 16865 15317 16899 15351
rect 17325 15317 17359 15351
rect 17693 15317 17727 15351
rect 18429 15317 18463 15351
rect 18889 15317 18923 15351
rect 20545 15317 20579 15351
rect 23029 15317 23063 15351
rect 23121 15317 23155 15351
rect 24225 15317 24259 15351
rect 29653 15317 29687 15351
rect 30113 15317 30147 15351
rect 30481 15317 30515 15351
rect 32781 15317 32815 15351
rect 32873 15317 32907 15351
rect 4169 15113 4203 15147
rect 5825 15113 5859 15147
rect 5917 15113 5951 15147
rect 6653 15113 6687 15147
rect 8125 15113 8159 15147
rect 8585 15113 8619 15147
rect 10977 15113 11011 15147
rect 12909 15113 12943 15147
rect 13277 15113 13311 15147
rect 14473 15113 14507 15147
rect 16681 15113 16715 15147
rect 17417 15113 17451 15147
rect 21833 15113 21867 15147
rect 26617 15113 26651 15147
rect 28917 15113 28951 15147
rect 32137 15113 32171 15147
rect 32597 15113 32631 15147
rect 33333 15113 33367 15147
rect 33977 15113 34011 15147
rect 34437 15113 34471 15147
rect 38301 15113 38335 15147
rect 2421 15045 2455 15079
rect 3034 15045 3068 15079
rect 7012 15045 7046 15079
rect 15761 15045 15795 15079
rect 30205 15045 30239 15079
rect 2329 14977 2363 15011
rect 4445 14977 4479 15011
rect 11785 14977 11819 15011
rect 13369 14977 13403 15011
rect 15945 14977 15979 15011
rect 18061 14977 18095 15011
rect 20473 14977 20507 15011
rect 20729 14977 20763 15011
rect 22477 14977 22511 15011
rect 23765 14977 23799 15011
rect 24501 14977 24535 15011
rect 25973 14977 26007 15011
rect 27788 14977 27822 15011
rect 29469 14977 29503 15011
rect 32505 14977 32539 15011
rect 33425 14977 33459 15011
rect 33885 14977 33919 15011
rect 2605 14909 2639 14943
rect 2789 14909 2823 14943
rect 5089 14909 5123 14943
rect 6101 14909 6135 14943
rect 6745 14909 6779 14943
rect 8401 14909 8435 14943
rect 8493 14909 8527 14943
rect 9597 14909 9631 14943
rect 11529 14909 11563 14943
rect 13185 14909 13219 14943
rect 17325 14909 17359 14943
rect 18199 14909 18233 14943
rect 18337 14909 18371 14943
rect 18613 14909 18647 14943
rect 19073 14909 19107 14943
rect 19257 14909 19291 14943
rect 22569 14909 22603 14943
rect 22753 14909 22787 14943
rect 23489 14909 23523 14943
rect 23627 14909 23661 14943
rect 25329 14909 25363 14943
rect 26065 14909 26099 14943
rect 26157 14909 26191 14943
rect 27629 14909 27663 14943
rect 27905 14909 27939 14943
rect 28641 14909 28675 14943
rect 28825 14909 28859 14943
rect 32689 14909 32723 14943
rect 33609 14909 33643 14943
rect 35081 14909 35115 14943
rect 35909 14909 35943 14943
rect 36553 14909 36587 14943
rect 37933 14909 37967 14943
rect 1869 14841 1903 14875
rect 8953 14841 8987 14875
rect 15301 14841 15335 14875
rect 23213 14841 23247 14875
rect 28181 14841 28215 14875
rect 1961 14773 1995 14807
rect 5457 14773 5491 14807
rect 9045 14773 9079 14807
rect 11345 14773 11379 14807
rect 13737 14773 13771 14807
rect 14105 14773 14139 14807
rect 16497 14773 16531 14807
rect 19349 14773 19383 14807
rect 24409 14773 24443 14807
rect 25605 14773 25639 14807
rect 26985 14773 27019 14807
rect 30113 14773 30147 14807
rect 31493 14773 31527 14807
rect 32965 14773 32999 14807
rect 34529 14773 34563 14807
rect 35265 14773 35299 14807
rect 37105 14773 37139 14807
rect 37289 14773 37323 14807
rect 3617 14569 3651 14603
rect 4169 14569 4203 14603
rect 7573 14569 7607 14603
rect 8769 14569 8803 14603
rect 11805 14569 11839 14603
rect 17693 14569 17727 14603
rect 19993 14569 20027 14603
rect 24133 14569 24167 14603
rect 24409 14569 24443 14603
rect 27905 14569 27939 14603
rect 28733 14569 28767 14603
rect 30941 14569 30975 14603
rect 32413 14569 32447 14603
rect 33241 14569 33275 14603
rect 34805 14569 34839 14603
rect 37013 14569 37047 14603
rect 15209 14501 15243 14535
rect 38117 14501 38151 14535
rect 1593 14433 1627 14467
rect 8125 14433 8159 14467
rect 12449 14433 12483 14467
rect 12725 14433 12759 14467
rect 13001 14433 13035 14467
rect 14749 14433 14783 14467
rect 19073 14433 19107 14467
rect 19441 14433 19475 14467
rect 19533 14433 19567 14467
rect 20637 14433 20671 14467
rect 24961 14433 24995 14467
rect 25789 14433 25823 14467
rect 26525 14433 26559 14467
rect 28549 14433 28583 14467
rect 29285 14433 29319 14467
rect 33149 14433 33183 14467
rect 33793 14433 33827 14467
rect 35357 14433 35391 14467
rect 37657 14433 37691 14467
rect 2237 14365 2271 14399
rect 5825 14365 5859 14399
rect 6193 14365 6227 14399
rect 6460 14365 6494 14399
rect 10333 14365 10367 14399
rect 12587 14365 12621 14399
rect 13461 14365 13495 14399
rect 13645 14365 13679 14399
rect 14565 14365 14599 14399
rect 16221 14365 16255 14399
rect 23673 14365 23707 14399
rect 29561 14365 29595 14399
rect 31033 14365 31067 14399
rect 35173 14365 35207 14399
rect 35633 14365 35667 14399
rect 37473 14365 37507 14399
rect 2145 14297 2179 14331
rect 2482 14297 2516 14331
rect 4261 14297 4295 14331
rect 9137 14297 9171 14331
rect 10600 14297 10634 14331
rect 15025 14297 15059 14331
rect 16488 14297 16522 14331
rect 18806 14297 18840 14331
rect 23428 14297 23462 14331
rect 25605 14297 25639 14331
rect 26792 14297 26826 14331
rect 27997 14297 28031 14331
rect 29828 14297 29862 14331
rect 31300 14297 31334 14331
rect 32505 14297 32539 14331
rect 35900 14297 35934 14331
rect 37565 14297 37599 14331
rect 11713 14229 11747 14263
rect 14105 14229 14139 14263
rect 14473 14229 14507 14263
rect 17601 14229 17635 14263
rect 19625 14229 19659 14263
rect 20085 14229 20119 14263
rect 22293 14229 22327 14263
rect 25237 14229 25271 14263
rect 25697 14229 25731 14263
rect 26341 14229 26375 14263
rect 34437 14229 34471 14263
rect 35265 14229 35299 14263
rect 37105 14229 37139 14263
rect 2697 14025 2731 14059
rect 6009 14025 6043 14059
rect 12909 14025 12943 14059
rect 18061 14025 18095 14059
rect 18889 14025 18923 14059
rect 24041 14025 24075 14059
rect 24961 14025 24995 14059
rect 25973 14025 26007 14059
rect 26341 14025 26375 14059
rect 26801 14025 26835 14059
rect 26985 14025 27019 14059
rect 27721 14025 27755 14059
rect 29561 14025 29595 14059
rect 30389 14025 30423 14059
rect 30573 14025 30607 14059
rect 32413 14025 32447 14059
rect 35173 14025 35207 14059
rect 37565 14025 37599 14059
rect 37657 14025 37691 14059
rect 38025 14025 38059 14059
rect 2237 13957 2271 13991
rect 7021 13957 7055 13991
rect 14749 13957 14783 13991
rect 16926 13957 16960 13991
rect 23489 13957 23523 13991
rect 3341 13889 3375 13923
rect 3709 13889 3743 13923
rect 3985 13889 4019 13923
rect 8217 13889 8251 13923
rect 9781 13889 9815 13923
rect 10517 13889 10551 13923
rect 10977 13889 11011 13923
rect 11069 13889 11103 13923
rect 11621 13889 11655 13923
rect 14197 13889 14231 13923
rect 14933 13889 14967 13923
rect 18153 13889 18187 13923
rect 19441 13889 19475 13923
rect 19901 13889 19935 13923
rect 22109 13889 22143 13923
rect 23581 13889 23615 13923
rect 24685 13889 24719 13923
rect 25513 13889 25547 13923
rect 26433 13889 26467 13923
rect 28273 13889 28307 13923
rect 29837 13889 29871 13923
rect 31217 13889 31251 13923
rect 33793 13889 33827 13923
rect 34060 13889 34094 13923
rect 36047 13889 36081 13923
rect 37105 13889 37139 13923
rect 4537 13821 4571 13855
rect 8401 13821 8435 13855
rect 9045 13821 9079 13855
rect 9965 13821 9999 13855
rect 11161 13821 11195 13855
rect 16681 13821 16715 13855
rect 18797 13821 18831 13855
rect 21557 13821 21591 13855
rect 22477 13821 22511 13855
rect 23397 13821 23431 13855
rect 26249 13821 26283 13855
rect 27537 13821 27571 13855
rect 35909 13821 35943 13855
rect 36185 13821 36219 13855
rect 36921 13821 36955 13855
rect 37473 13821 37507 13855
rect 23949 13753 23983 13787
rect 36461 13753 36495 13787
rect 6561 13685 6595 13719
rect 9413 13685 9447 13719
rect 10609 13685 10643 13719
rect 13645 13685 13679 13719
rect 33609 13685 33643 13719
rect 35265 13685 35299 13719
rect 38393 13685 38427 13719
rect 2973 13481 3007 13515
rect 10517 13481 10551 13515
rect 13369 13481 13403 13515
rect 14749 13481 14783 13515
rect 16405 13481 16439 13515
rect 23489 13481 23523 13515
rect 24593 13481 24627 13515
rect 25421 13481 25455 13515
rect 26617 13481 26651 13515
rect 27077 13481 27111 13515
rect 27997 13481 28031 13515
rect 36277 13481 36311 13515
rect 38209 13481 38243 13515
rect 17141 13413 17175 13447
rect 3617 13345 3651 13379
rect 9321 13345 9355 13379
rect 14105 13345 14139 13379
rect 17049 13345 17083 13379
rect 17693 13345 17727 13379
rect 18521 13345 18555 13379
rect 21557 13345 21591 13379
rect 24777 13345 24811 13379
rect 26065 13345 26099 13379
rect 36829 13345 36863 13379
rect 8769 13277 8803 13311
rect 9137 13277 9171 13311
rect 11897 13277 11931 13311
rect 11989 13277 12023 13311
rect 12256 13277 12290 13311
rect 13737 13277 13771 13311
rect 15761 13277 15795 13311
rect 16313 13277 16347 13311
rect 17509 13277 17543 13311
rect 22201 13277 22235 13311
rect 28457 13277 28491 13311
rect 30665 13277 30699 13311
rect 31953 13277 31987 13311
rect 32505 13277 32539 13311
rect 8033 13209 8067 13243
rect 11630 13209 11664 13243
rect 25697 13209 25731 13243
rect 28089 13209 28123 13243
rect 30481 13209 30515 13243
rect 34161 13209 34195 13243
rect 34989 13209 35023 13243
rect 37096 13209 37130 13243
rect 8125 13141 8159 13175
rect 10333 13141 10367 13175
rect 17601 13141 17635 13175
rect 17969 13141 18003 13175
rect 22109 13141 22143 13175
rect 27353 13141 27387 13175
rect 27721 13141 27755 13175
rect 31217 13141 31251 13175
rect 31309 13141 31343 13175
rect 34529 13141 34563 13175
rect 7941 12937 7975 12971
rect 11345 12937 11379 12971
rect 17049 12937 17083 12971
rect 24409 12937 24443 12971
rect 30665 12937 30699 12971
rect 31125 12937 31159 12971
rect 32413 12937 32447 12971
rect 36093 12937 36127 12971
rect 37289 12937 37323 12971
rect 38301 12937 38335 12971
rect 2789 12869 2823 12903
rect 4169 12869 4203 12903
rect 12541 12869 12575 12903
rect 17601 12869 17635 12903
rect 18705 12869 18739 12903
rect 22100 12869 22134 12903
rect 25145 12869 25179 12903
rect 27445 12869 27479 12903
rect 29837 12869 29871 12903
rect 34529 12869 34563 12903
rect 2697 12801 2731 12835
rect 2973 12801 3007 12835
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 9054 12801 9088 12835
rect 9413 12801 9447 12835
rect 10241 12801 10275 12835
rect 10701 12801 10735 12835
rect 12633 12801 12667 12835
rect 13001 12801 13035 12835
rect 13553 12801 13587 12835
rect 17509 12801 17543 12835
rect 18889 12801 18923 12835
rect 21833 12801 21867 12835
rect 23305 12801 23339 12835
rect 24133 12801 24167 12835
rect 25697 12801 25731 12835
rect 27353 12801 27387 12835
rect 31033 12801 31067 12835
rect 32505 12801 32539 12835
rect 34713 12801 34747 12835
rect 34980 12801 35014 12835
rect 36185 12801 36219 12835
rect 37841 12801 37875 12835
rect 3617 12733 3651 12767
rect 7297 12733 7331 12767
rect 9321 12733 9355 12767
rect 12817 12733 12851 12767
rect 14289 12733 14323 12767
rect 15945 12733 15979 12767
rect 17693 12733 17727 12767
rect 18153 12733 18187 12767
rect 20913 12733 20947 12767
rect 24961 12733 24995 12767
rect 26801 12733 26835 12767
rect 27537 12733 27571 12767
rect 28365 12733 28399 12767
rect 29101 12733 29135 12767
rect 30481 12733 30515 12767
rect 31217 12733 31251 12767
rect 31953 12733 31987 12767
rect 32229 12733 32263 12767
rect 33517 12733 33551 12767
rect 36737 12733 36771 12767
rect 2973 12665 3007 12699
rect 11805 12665 11839 12699
rect 17141 12665 17175 12699
rect 26985 12665 27019 12699
rect 3065 12597 3099 12631
rect 7849 12597 7883 12631
rect 12173 12597 12207 12631
rect 13737 12597 13771 12631
rect 16497 12597 16531 12631
rect 21557 12597 21591 12631
rect 23213 12597 23247 12631
rect 26157 12597 26191 12631
rect 27813 12597 27847 12631
rect 28549 12597 28583 12631
rect 29929 12597 29963 12631
rect 32873 12597 32907 12631
rect 32965 12597 32999 12631
rect 2881 12393 2915 12427
rect 2973 12393 3007 12427
rect 4261 12393 4295 12427
rect 6377 12393 6411 12427
rect 7297 12393 7331 12427
rect 8769 12393 8803 12427
rect 11437 12393 11471 12427
rect 12541 12393 12575 12427
rect 15945 12393 15979 12427
rect 18245 12393 18279 12427
rect 20545 12393 20579 12427
rect 28365 12393 28399 12427
rect 28457 12393 28491 12427
rect 30757 12393 30791 12427
rect 34897 12393 34931 12427
rect 35817 12393 35851 12427
rect 37473 12393 37507 12427
rect 37841 12393 37875 12427
rect 18153 12325 18187 12359
rect 27537 12325 27571 12359
rect 31953 12325 31987 12359
rect 33425 12325 33459 12359
rect 7389 12257 7423 12291
rect 9689 12257 9723 12291
rect 12081 12257 12115 12291
rect 13369 12257 13403 12291
rect 15117 12257 15151 12291
rect 16497 12257 16531 12291
rect 16773 12257 16807 12291
rect 18797 12257 18831 12291
rect 19901 12257 19935 12291
rect 22201 12257 22235 12291
rect 22661 12257 22695 12291
rect 23054 12257 23088 12291
rect 23213 12257 23247 12291
rect 25053 12257 25087 12291
rect 25421 12257 25455 12291
rect 26157 12257 26191 12291
rect 27721 12257 27755 12291
rect 27905 12257 27939 12291
rect 31401 12257 31435 12291
rect 31560 12257 31594 12291
rect 32781 12257 32815 12291
rect 32965 12257 32999 12291
rect 34069 12257 34103 12291
rect 35173 12257 35207 12291
rect 36461 12257 36495 12291
rect 38393 12257 38427 12291
rect 2329 12189 2363 12223
rect 3617 12189 3651 12223
rect 5365 12189 5399 12223
rect 6561 12189 6595 12223
rect 6745 12189 6779 12223
rect 7656 12189 7690 12223
rect 9137 12189 9171 12223
rect 10241 12189 10275 12223
rect 14657 12189 14691 12223
rect 15301 12189 15335 12223
rect 17029 12189 17063 12223
rect 21658 12189 21692 12223
rect 21925 12189 21959 12223
rect 22017 12189 22051 12223
rect 22937 12189 22971 12223
rect 25605 12189 25639 12223
rect 29009 12189 29043 12223
rect 30113 12189 30147 12223
rect 31677 12189 31711 12223
rect 32413 12189 32447 12223
rect 32597 12189 32631 12223
rect 4169 12121 4203 12155
rect 11069 12121 11103 12155
rect 15853 12121 15887 12155
rect 16313 12121 16347 12155
rect 23857 12121 23891 12155
rect 25513 12121 25547 12155
rect 26424 12121 26458 12155
rect 35357 12121 35391 12155
rect 35909 12121 35943 12155
rect 37565 12121 37599 12155
rect 4813 12053 4847 12087
rect 12725 12053 12759 12087
rect 13093 12053 13127 12087
rect 13185 12053 13219 12087
rect 13921 12053 13955 12087
rect 14105 12053 14139 12087
rect 16405 12053 16439 12087
rect 20453 12053 20487 12087
rect 24133 12053 24167 12087
rect 24409 12053 24443 12087
rect 24777 12053 24811 12087
rect 24869 12053 24903 12087
rect 25973 12053 26007 12087
rect 27997 12053 28031 12087
rect 29561 12053 29595 12087
rect 30573 12053 30607 12087
rect 33057 12053 33091 12087
rect 33517 12053 33551 12087
rect 34529 12053 34563 12087
rect 35449 12053 35483 12087
rect 37197 12053 37231 12087
rect 2421 11849 2455 11883
rect 3985 11849 4019 11883
rect 5374 11849 5408 11883
rect 7389 11849 7423 11883
rect 7849 11849 7883 11883
rect 11897 11849 11931 11883
rect 13461 11849 13495 11883
rect 13829 11849 13863 11883
rect 14289 11849 14323 11883
rect 20913 11849 20947 11883
rect 21373 11849 21407 11883
rect 26801 11849 26835 11883
rect 29193 11849 29227 11883
rect 29653 11849 29687 11883
rect 32137 11849 32171 11883
rect 38301 11849 38335 11883
rect 1777 11781 1811 11815
rect 1977 11781 2011 11815
rect 2872 11781 2906 11815
rect 4261 11781 4295 11815
rect 4675 11781 4709 11815
rect 12348 11781 12382 11815
rect 16252 11781 16286 11815
rect 21281 11781 21315 11815
rect 30196 11781 30230 11815
rect 34529 11781 34563 11815
rect 35786 11781 35820 11815
rect 37657 11781 37691 11815
rect 2329 11713 2363 11747
rect 2513 11713 2547 11747
rect 4997 11713 5031 11747
rect 5641 11713 5675 11747
rect 6929 11713 6963 11747
rect 7021 11713 7055 11747
rect 7757 11713 7791 11747
rect 8217 11713 8251 11747
rect 10517 11713 10551 11747
rect 11161 11713 11195 11747
rect 12081 11713 12115 11747
rect 13921 11713 13955 11747
rect 16497 11713 16531 11747
rect 17417 11713 17451 11747
rect 18613 11713 18647 11747
rect 19073 11713 19107 11747
rect 19533 11713 19567 11747
rect 22100 11713 22134 11747
rect 23397 11713 23431 11747
rect 24961 11713 24995 11747
rect 25688 11713 25722 11747
rect 27788 11713 27822 11747
rect 28825 11713 28859 11747
rect 29285 11713 29319 11747
rect 33250 11713 33284 11747
rect 33517 11713 33551 11747
rect 2605 11645 2639 11679
rect 7113 11645 7147 11679
rect 7941 11645 7975 11679
rect 8401 11645 8435 11679
rect 9137 11645 9171 11679
rect 9254 11645 9288 11679
rect 9413 11645 9447 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 13645 11645 13679 11679
rect 14933 11645 14967 11679
rect 17555 11645 17589 11679
rect 17693 11645 17727 11679
rect 18429 11645 18463 11679
rect 19165 11645 19199 11679
rect 19257 11645 19291 11679
rect 20085 11645 20119 11679
rect 21557 11645 21591 11679
rect 21833 11645 21867 11679
rect 24133 11645 24167 11679
rect 25421 11645 25455 11679
rect 27629 11645 27663 11679
rect 27905 11645 27939 11679
rect 28641 11645 28675 11679
rect 29009 11645 29043 11679
rect 29929 11645 29963 11679
rect 33977 11645 34011 11679
rect 34713 11645 34747 11679
rect 35541 11645 35575 11679
rect 37749 11645 37783 11679
rect 37841 11645 37875 11679
rect 6193 11577 6227 11611
rect 8861 11577 8895 11611
rect 10057 11577 10091 11611
rect 17969 11577 18003 11611
rect 28181 11577 28215 11611
rect 36921 11577 36955 11611
rect 1961 11509 1995 11543
rect 2145 11509 2179 11543
rect 4629 11509 4663 11543
rect 4813 11509 4847 11543
rect 5365 11509 5399 11543
rect 6561 11509 6595 11543
rect 10149 11509 10183 11543
rect 14381 11509 14415 11543
rect 15117 11509 15151 11543
rect 16773 11509 16807 11543
rect 18705 11509 18739 11543
rect 23213 11509 23247 11543
rect 24409 11509 24443 11543
rect 26985 11509 27019 11543
rect 31309 11509 31343 11543
rect 35265 11509 35299 11543
rect 37289 11509 37323 11543
rect 1501 11305 1535 11339
rect 5825 11305 5859 11339
rect 6193 11305 6227 11339
rect 8769 11305 8803 11339
rect 10609 11305 10643 11339
rect 12541 11305 12575 11339
rect 14841 11305 14875 11339
rect 15945 11305 15979 11339
rect 21741 11305 21775 11339
rect 21925 11305 21959 11339
rect 25053 11305 25087 11339
rect 27445 11305 27479 11339
rect 29101 11305 29135 11339
rect 30113 11305 30147 11339
rect 34713 11305 34747 11339
rect 35541 11305 35575 11339
rect 5365 11237 5399 11271
rect 5733 11237 5767 11271
rect 8953 11237 8987 11271
rect 19533 11237 19567 11271
rect 27353 11237 27387 11271
rect 36737 11237 36771 11271
rect 37473 11237 37507 11271
rect 5917 11169 5951 11203
rect 6653 11169 6687 11203
rect 10333 11169 10367 11203
rect 11069 11169 11103 11203
rect 14197 11169 14231 11203
rect 15485 11169 15519 11203
rect 17601 11169 17635 11203
rect 18061 11169 18095 11203
rect 23305 11169 23339 11203
rect 25973 11169 26007 11203
rect 28825 11169 28859 11203
rect 32965 11169 32999 11203
rect 33885 11169 33919 11203
rect 35265 11169 35299 11203
rect 36199 11169 36233 11203
rect 37381 11169 37415 11203
rect 38117 11169 38151 11203
rect 2053 11101 2087 11135
rect 2237 11101 2271 11135
rect 3801 11101 3835 11135
rect 7389 11101 7423 11135
rect 13665 11101 13699 11135
rect 13921 11101 13955 11135
rect 14473 11101 14507 11135
rect 18245 11101 18279 11135
rect 23038 11101 23072 11135
rect 24409 11101 24443 11135
rect 25789 11101 25823 11135
rect 26240 11101 26274 11135
rect 28569 11101 28603 11135
rect 31226 11101 31260 11135
rect 31493 11101 31527 11135
rect 33609 11101 33643 11135
rect 36323 11101 36357 11135
rect 36461 11101 36495 11135
rect 37197 11101 37231 11135
rect 2504 11033 2538 11067
rect 4046 11033 4080 11067
rect 7297 11033 7331 11067
rect 7634 11033 7668 11067
rect 10066 11033 10100 11067
rect 11336 11033 11370 11067
rect 14381 11033 14415 11067
rect 14933 11033 14967 11067
rect 16037 11033 16071 11067
rect 18889 11033 18923 11067
rect 23949 11033 23983 11067
rect 25329 11033 25363 11067
rect 32720 11033 32754 11067
rect 34529 11033 34563 11067
rect 35081 11033 35115 11067
rect 35173 11033 35207 11067
rect 37841 11033 37875 11067
rect 3617 10965 3651 10999
rect 5181 10965 5215 10999
rect 12449 10965 12483 10999
rect 18153 10965 18187 10999
rect 18613 10965 18647 10999
rect 23581 10965 23615 10999
rect 23857 10965 23891 10999
rect 31585 10965 31619 10999
rect 33057 10965 33091 10999
rect 37933 10965 37967 10999
rect 1685 10761 1719 10795
rect 2053 10761 2087 10795
rect 3341 10761 3375 10795
rect 4077 10761 4111 10795
rect 5365 10761 5399 10795
rect 6009 10761 6043 10795
rect 7757 10761 7791 10795
rect 8493 10761 8527 10795
rect 8953 10761 8987 10795
rect 10149 10761 10183 10795
rect 11529 10761 11563 10795
rect 12909 10761 12943 10795
rect 16957 10761 16991 10795
rect 18429 10761 18463 10795
rect 22201 10761 22235 10795
rect 23305 10761 23339 10795
rect 24225 10761 24259 10795
rect 26157 10761 26191 10795
rect 28181 10761 28215 10795
rect 28273 10761 28307 10795
rect 29285 10761 29319 10795
rect 29837 10761 29871 10795
rect 30481 10761 30515 10795
rect 30941 10761 30975 10795
rect 32505 10761 32539 10795
rect 34253 10761 34287 10795
rect 36093 10761 36127 10795
rect 36829 10761 36863 10795
rect 37565 10761 37599 10795
rect 37657 10761 37691 10795
rect 1961 10693 1995 10727
rect 3433 10693 3467 10727
rect 5641 10693 5675 10727
rect 5825 10693 5859 10727
rect 7665 10693 7699 10727
rect 22569 10693 22603 10727
rect 29929 10693 29963 10727
rect 32965 10693 32999 10727
rect 35366 10693 35400 10727
rect 1777 10625 1811 10659
rect 3580 10625 3614 10659
rect 4813 10625 4847 10659
rect 5089 10625 5123 10659
rect 5549 10625 5583 10659
rect 8401 10625 8435 10659
rect 8861 10625 8895 10659
rect 9413 10625 9447 10659
rect 10701 10625 10735 10659
rect 12357 10625 12391 10659
rect 15301 10625 15335 10659
rect 15761 10625 15795 10659
rect 16313 10625 16347 10659
rect 17049 10625 17083 10659
rect 17316 10625 17350 10659
rect 18521 10625 18555 10659
rect 19073 10625 19107 10659
rect 22661 10625 22695 10659
rect 23949 10625 23983 10659
rect 27353 10625 27387 10659
rect 27445 10625 27479 10659
rect 28733 10625 28767 10659
rect 30849 10625 30883 10659
rect 31309 10625 31343 10659
rect 31861 10625 31895 10659
rect 34069 10625 34103 10659
rect 35633 10625 35667 10659
rect 38117 10625 38151 10659
rect 2237 10557 2271 10591
rect 2329 10557 2363 10591
rect 2421 10557 2455 10591
rect 2513 10557 2547 10591
rect 2697 10557 2731 10591
rect 3801 10557 3835 10591
rect 9137 10557 9171 10591
rect 10057 10557 10091 10591
rect 12173 10557 12207 10591
rect 13001 10557 13035 10591
rect 13185 10557 13219 10591
rect 13921 10557 13955 10591
rect 14059 10557 14093 10591
rect 14197 10557 14231 10591
rect 15393 10557 15427 10591
rect 15577 10557 15611 10591
rect 22845 10557 22879 10591
rect 26801 10557 26835 10591
rect 27537 10557 27571 10591
rect 28365 10557 28399 10591
rect 31033 10557 31067 10591
rect 32229 10557 32263 10591
rect 32413 10557 32447 10591
rect 33517 10557 33551 10591
rect 36185 10557 36219 10591
rect 36277 10557 36311 10591
rect 37381 10557 37415 10591
rect 3709 10489 3743 10523
rect 13645 10489 13679 10523
rect 14841 10489 14875 10523
rect 26985 10489 27019 10523
rect 32873 10489 32907 10523
rect 5825 10421 5859 10455
rect 7205 10421 7239 10455
rect 14933 10421 14967 10455
rect 24685 10421 24719 10455
rect 25973 10421 26007 10455
rect 27813 10421 27847 10455
rect 30389 10421 30423 10455
rect 35725 10421 35759 10455
rect 38025 10421 38059 10455
rect 38301 10421 38335 10455
rect 2329 10217 2363 10251
rect 2605 10217 2639 10251
rect 5457 10217 5491 10251
rect 15853 10217 15887 10251
rect 18061 10217 18095 10251
rect 18245 10217 18279 10251
rect 27077 10217 27111 10251
rect 27169 10217 27203 10251
rect 30389 10217 30423 10251
rect 31309 10217 31343 10251
rect 34161 10217 34195 10251
rect 37657 10217 37691 10251
rect 38393 10217 38427 10251
rect 2513 10149 2547 10183
rect 5089 10149 5123 10183
rect 7481 10149 7515 10183
rect 7849 10149 7883 10183
rect 9873 10149 9907 10183
rect 12541 10149 12575 10183
rect 28181 10149 28215 10183
rect 30021 10149 30055 10183
rect 32413 10149 32447 10183
rect 3157 10081 3191 10115
rect 4629 10081 4663 10115
rect 5181 10081 5215 10115
rect 14933 10081 14967 10115
rect 16681 10081 16715 10115
rect 18797 10081 18831 10115
rect 27721 10081 27755 10115
rect 33057 10081 33091 10115
rect 33793 10081 33827 10115
rect 37749 10081 37783 10115
rect 4261 10013 4295 10047
rect 4721 10013 4755 10047
rect 8033 10013 8067 10047
rect 8953 10013 8987 10047
rect 12449 10013 12483 10047
rect 13921 10013 13955 10047
rect 31585 10013 31619 10047
rect 32045 10013 32079 10047
rect 34713 10013 34747 10047
rect 36277 10013 36311 10047
rect 2145 9945 2179 9979
rect 13676 9945 13710 9979
rect 14381 9945 14415 9979
rect 16948 9945 16982 9979
rect 34437 9945 34471 9979
rect 34980 9945 35014 9979
rect 36544 9945 36578 9979
rect 2355 9877 2389 9911
rect 4445 9877 4479 9911
rect 8585 9877 8619 9911
rect 9597 9877 9631 9911
rect 12081 9877 12115 9911
rect 15393 9877 15427 9911
rect 23029 9877 23063 9911
rect 26709 9877 26743 9911
rect 30757 9877 30791 9911
rect 32689 9877 32723 9911
rect 36093 9877 36127 9911
rect 2789 9673 2823 9707
rect 3065 9673 3099 9707
rect 4445 9673 4479 9707
rect 8125 9673 8159 9707
rect 17693 9673 17727 9707
rect 27629 9673 27663 9707
rect 36277 9673 36311 9707
rect 37289 9673 37323 9707
rect 4813 9605 4847 9639
rect 7757 9605 7791 9639
rect 8493 9605 8527 9639
rect 12817 9605 12851 9639
rect 17141 9605 17175 9639
rect 25421 9605 25455 9639
rect 34437 9605 34471 9639
rect 2605 9537 2639 9571
rect 2881 9537 2915 9571
rect 2973 9537 3007 9571
rect 3801 9537 3835 9571
rect 4286 9537 4320 9571
rect 4629 9537 4663 9571
rect 7665 9537 7699 9571
rect 8585 9537 8619 9571
rect 8953 9537 8987 9571
rect 12633 9537 12667 9571
rect 17233 9537 17267 9571
rect 18337 9537 18371 9571
rect 21649 9537 21683 9571
rect 22109 9537 22143 9571
rect 38485 9537 38519 9571
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 4169 9469 4203 9503
rect 6653 9469 6687 9503
rect 7849 9469 7883 9503
rect 8677 9469 8711 9503
rect 9505 9469 9539 9503
rect 16405 9469 16439 9503
rect 16957 9469 16991 9503
rect 18981 9469 19015 9503
rect 22937 9469 22971 9503
rect 23765 9469 23799 9503
rect 26157 9469 26191 9503
rect 29929 9469 29963 9503
rect 31217 9469 31251 9503
rect 32321 9469 32355 9503
rect 33793 9469 33827 9503
rect 34345 9469 34379 9503
rect 36829 9469 36863 9503
rect 37841 9469 37875 9503
rect 2881 9401 2915 9435
rect 7297 9401 7331 9435
rect 17601 9401 17635 9435
rect 29101 9401 29135 9435
rect 29837 9401 29871 9435
rect 38301 9401 38335 9435
rect 7205 9333 7239 9367
rect 9873 9333 9907 9367
rect 11989 9333 12023 9367
rect 18429 9333 18463 9367
rect 23213 9333 23247 9367
rect 25513 9333 25547 9367
rect 27169 9333 27203 9367
rect 29377 9333 29411 9367
rect 30573 9333 30607 9367
rect 30665 9333 30699 9367
rect 31585 9333 31619 9367
rect 32965 9333 32999 9367
rect 33333 9333 33367 9367
rect 35725 9333 35759 9367
rect 24685 9129 24719 9163
rect 31217 9129 31251 9163
rect 34345 9129 34379 9163
rect 35357 9129 35391 9163
rect 37749 9129 37783 9163
rect 3617 9061 3651 9095
rect 7297 9061 7331 9095
rect 9689 9061 9723 9095
rect 12081 9061 12115 9095
rect 26433 9061 26467 9095
rect 9045 8993 9079 9027
rect 10333 8993 10367 9027
rect 11989 8993 12023 9027
rect 12725 8993 12759 9027
rect 16773 8993 16807 9027
rect 35909 8993 35943 9027
rect 38301 8993 38335 9027
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 4537 8925 4571 8959
rect 6745 8925 6779 8959
rect 8502 8925 8536 8959
rect 8769 8925 8803 8959
rect 13461 8925 13495 8959
rect 15945 8925 15979 8959
rect 16865 8925 16899 8959
rect 18613 8925 18647 8959
rect 21097 8925 21131 8959
rect 22569 8925 22603 8959
rect 24041 8925 24075 8959
rect 25053 8925 25087 8959
rect 27077 8925 27111 8959
rect 27813 8925 27847 8959
rect 29745 8925 29779 8959
rect 30012 8925 30046 8959
rect 32597 8925 32631 8959
rect 33241 8925 33275 8959
rect 33977 8925 34011 8959
rect 36645 8925 36679 8959
rect 37381 8925 37415 8959
rect 4353 8857 4387 8891
rect 17132 8857 17166 8891
rect 18429 8857 18463 8891
rect 22324 8857 22358 8891
rect 23796 8857 23830 8891
rect 25320 8857 25354 8891
rect 28273 8857 28307 8891
rect 29009 8857 29043 8891
rect 32352 8857 32386 8891
rect 33425 8857 33459 8891
rect 3249 8789 3283 8823
rect 4629 8789 4663 8823
rect 7389 8789 7423 8823
rect 9229 8789 9263 8823
rect 9321 8789 9355 8823
rect 9781 8789 9815 8823
rect 11345 8789 11379 8823
rect 12449 8789 12483 8823
rect 12541 8789 12575 8823
rect 12909 8789 12943 8823
rect 15393 8789 15427 8823
rect 16129 8789 16163 8823
rect 18245 8789 18279 8823
rect 20453 8789 20487 8823
rect 21189 8789 21223 8823
rect 22661 8789 22695 8823
rect 26525 8789 26559 8823
rect 27261 8789 27295 8823
rect 28549 8789 28583 8823
rect 29377 8789 29411 8823
rect 31125 8789 31159 8823
rect 32689 8789 32723 8823
rect 34897 8789 34931 8823
rect 36093 8789 36127 8823
rect 36829 8789 36863 8823
rect 10333 8585 10367 8619
rect 13001 8585 13035 8619
rect 16865 8585 16899 8619
rect 26065 8585 26099 8619
rect 30849 8585 30883 8619
rect 30941 8585 30975 8619
rect 31309 8585 31343 8619
rect 33333 8585 33367 8619
rect 33701 8585 33735 8619
rect 35817 8585 35851 8619
rect 36737 8585 36771 8619
rect 38393 8585 38427 8619
rect 11866 8517 11900 8551
rect 13553 8517 13587 8551
rect 17408 8517 17442 8551
rect 29736 8517 29770 8551
rect 34069 8517 34103 8551
rect 36369 8517 36403 8551
rect 6469 8449 6503 8483
rect 6736 8449 6770 8483
rect 7941 8449 7975 8483
rect 8861 8449 8895 8483
rect 8978 8449 9012 8483
rect 9781 8449 9815 8483
rect 10241 8449 10275 8483
rect 11345 8449 11379 8483
rect 13461 8449 13495 8483
rect 13921 8449 13955 8483
rect 15117 8449 15151 8483
rect 15384 8449 15418 8483
rect 17141 8449 17175 8483
rect 20269 8449 20303 8483
rect 20525 8449 20559 8483
rect 22753 8449 22787 8483
rect 22870 8449 22904 8483
rect 24409 8449 24443 8483
rect 24685 8449 24719 8483
rect 24952 8449 24986 8483
rect 26157 8449 26191 8483
rect 27353 8449 27387 8483
rect 27813 8449 27847 8483
rect 31401 8449 31435 8483
rect 32505 8449 32539 8483
rect 33241 8449 33275 8483
rect 34345 8449 34379 8483
rect 34437 8449 34471 8483
rect 34704 8449 34738 8483
rect 37013 8449 37047 8483
rect 37289 8449 37323 8483
rect 38209 8449 38243 8483
rect 8125 8381 8159 8415
rect 9137 8381 9171 8415
rect 10425 8381 10459 8415
rect 11621 8381 11655 8415
rect 13737 8381 13771 8415
rect 14473 8381 14507 8415
rect 19165 8381 19199 8415
rect 19625 8381 19659 8415
rect 20177 8381 20211 8415
rect 21833 8381 21867 8415
rect 22017 8381 22051 8415
rect 23029 8381 23063 8415
rect 26709 8381 26743 8415
rect 27077 8381 27111 8415
rect 27261 8381 27295 8415
rect 28365 8381 28399 8415
rect 28549 8381 28583 8415
rect 29469 8381 29503 8415
rect 31585 8381 31619 8415
rect 32597 8381 32631 8415
rect 32781 8381 32815 8415
rect 33149 8381 33183 8415
rect 36093 8381 36127 8415
rect 36277 8381 36311 8415
rect 6193 8313 6227 8347
rect 7849 8313 7883 8347
rect 8585 8313 8619 8347
rect 13093 8313 13127 8347
rect 16497 8313 16531 8347
rect 18521 8313 18555 8347
rect 21649 8313 21683 8347
rect 22477 8313 22511 8347
rect 23673 8313 23707 8347
rect 27721 8313 27755 8347
rect 34161 8313 34195 8347
rect 37473 8313 37507 8347
rect 37749 8313 37783 8347
rect 9873 8245 9907 8279
rect 10701 8245 10735 8279
rect 18613 8245 18647 8279
rect 23765 8245 23799 8279
rect 29193 8245 29227 8279
rect 32137 8245 32171 8279
rect 36829 8245 36863 8279
rect 3893 8041 3927 8075
rect 4629 8041 4663 8075
rect 6653 8041 6687 8075
rect 13645 8041 13679 8075
rect 14841 8041 14875 8075
rect 15393 8041 15427 8075
rect 17049 8041 17083 8075
rect 20545 8041 20579 8075
rect 23581 8041 23615 8075
rect 24593 8041 24627 8075
rect 25605 8041 25639 8075
rect 27629 8041 27663 8075
rect 29837 8041 29871 8075
rect 32597 8041 32631 8075
rect 33609 8041 33643 8075
rect 36093 8041 36127 8075
rect 13277 7973 13311 8007
rect 15301 7973 15335 8007
rect 2881 7905 2915 7939
rect 4169 7905 4203 7939
rect 8769 7905 8803 7939
rect 15945 7905 15979 7939
rect 16313 7905 16347 7939
rect 17831 7905 17865 7939
rect 18245 7905 18279 7939
rect 18705 7905 18739 7939
rect 18889 7905 18923 7939
rect 19809 7905 19843 7939
rect 21189 7905 21223 7939
rect 23029 7905 23063 7939
rect 23121 7905 23155 7939
rect 25053 7905 25087 7939
rect 26341 7905 26375 7939
rect 26479 7905 26513 7939
rect 26617 7905 26651 7939
rect 26893 7905 26927 7939
rect 27353 7905 27387 7939
rect 27537 7905 27571 7939
rect 29377 7905 29411 7939
rect 30389 7905 30423 7939
rect 30665 7905 30699 7939
rect 30849 7905 30883 7939
rect 31309 7905 31343 7939
rect 31585 7905 31619 7939
rect 31702 7905 31736 7939
rect 31861 7905 31895 7939
rect 33149 7905 33183 7939
rect 33977 7905 34011 7939
rect 34713 7905 34747 7939
rect 38117 7905 38151 7939
rect 38301 7905 38335 7939
rect 2697 7837 2731 7871
rect 2789 7837 2823 7871
rect 4091 7837 4125 7871
rect 7297 7837 7331 7871
rect 8953 7837 8987 7871
rect 9781 7837 9815 7871
rect 10425 7837 10459 7871
rect 11897 7837 11931 7871
rect 15761 7837 15795 7871
rect 17693 7837 17727 7871
rect 17969 7837 18003 7871
rect 20913 7837 20947 7871
rect 21005 7837 21039 7871
rect 22753 7837 22787 7871
rect 29009 7837 29043 7871
rect 30205 7837 30239 7871
rect 33425 7837 33459 7871
rect 34069 7837 34103 7871
rect 36185 7837 36219 7871
rect 36452 7837 36486 7871
rect 3157 7769 3191 7803
rect 4813 7769 4847 7803
rect 8524 7769 8558 7803
rect 10692 7769 10726 7803
rect 12164 7769 12198 7803
rect 16497 7769 16531 7803
rect 22508 7769 22542 7803
rect 25237 7769 25271 7803
rect 28764 7769 28798 7803
rect 34980 7769 35014 7803
rect 3065 7701 3099 7735
rect 4445 7701 4479 7735
rect 4608 7701 4642 7735
rect 7389 7701 7423 7735
rect 10333 7701 10367 7735
rect 11805 7701 11839 7735
rect 15853 7701 15887 7735
rect 16589 7701 16623 7735
rect 16957 7701 16991 7735
rect 19257 7701 19291 7735
rect 21373 7701 21407 7735
rect 23213 7701 23247 7735
rect 23949 7701 23983 7735
rect 25145 7701 25179 7735
rect 25697 7701 25731 7735
rect 30297 7701 30331 7735
rect 32505 7701 32539 7735
rect 34161 7701 34195 7735
rect 34529 7701 34563 7735
rect 37565 7701 37599 7735
rect 37657 7701 37691 7735
rect 38025 7701 38059 7735
rect 8677 7497 8711 7531
rect 9137 7497 9171 7531
rect 14381 7497 14415 7531
rect 15761 7497 15795 7531
rect 18429 7497 18463 7531
rect 18521 7497 18555 7531
rect 18889 7497 18923 7531
rect 21373 7497 21407 7531
rect 24409 7497 24443 7531
rect 27261 7497 27295 7531
rect 28273 7497 28307 7531
rect 30297 7497 30331 7531
rect 33057 7497 33091 7531
rect 33793 7497 33827 7531
rect 35173 7497 35207 7531
rect 37289 7497 37323 7531
rect 5273 7429 5307 7463
rect 5457 7429 5491 7463
rect 10057 7429 10091 7463
rect 16405 7429 16439 7463
rect 30205 7429 30239 7463
rect 31432 7429 31466 7463
rect 32137 7429 32171 7463
rect 33425 7429 33459 7463
rect 3065 7361 3099 7395
rect 3801 7361 3835 7395
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 4169 7361 4203 7395
rect 5549 7361 5583 7395
rect 7472 7361 7506 7395
rect 9045 7361 9079 7395
rect 12792 7361 12826 7395
rect 12909 7361 12943 7395
rect 13829 7361 13863 7395
rect 14289 7361 14323 7395
rect 14749 7361 14783 7395
rect 15669 7361 15703 7395
rect 16681 7361 16715 7395
rect 16937 7361 16971 7395
rect 18981 7361 19015 7395
rect 22477 7361 22511 7395
rect 22569 7361 22603 7395
rect 25421 7361 25455 7395
rect 25688 7361 25722 7395
rect 27353 7361 27387 7395
rect 28365 7361 28399 7395
rect 32689 7361 32723 7395
rect 34345 7361 34379 7395
rect 34529 7361 34563 7395
rect 36068 7361 36102 7395
rect 36185 7361 36219 7395
rect 37105 7361 37139 7395
rect 37841 7361 37875 7395
rect 38209 7361 38243 7395
rect 2697 7293 2731 7327
rect 2973 7293 3007 7327
rect 4629 7293 4663 7327
rect 7205 7293 7239 7327
rect 9229 7293 9263 7327
rect 11897 7293 11931 7327
rect 12633 7293 12667 7327
rect 13185 7293 13219 7327
rect 13691 7293 13725 7327
rect 14473 7293 14507 7327
rect 15301 7293 15335 7327
rect 18245 7293 18279 7327
rect 19533 7293 19567 7327
rect 24961 7293 24995 7327
rect 27077 7293 27111 7327
rect 28733 7293 28767 7327
rect 31677 7293 31711 7327
rect 35909 7293 35943 7327
rect 36921 7293 36955 7327
rect 38393 7293 38427 7327
rect 5181 7225 5215 7259
rect 8585 7225 8619 7259
rect 23857 7225 23891 7259
rect 28089 7225 28123 7259
rect 29193 7225 29227 7259
rect 36461 7225 36495 7259
rect 3709 7157 3743 7191
rect 4445 7157 4479 7191
rect 5273 7157 5307 7191
rect 9689 7157 9723 7191
rect 11253 7157 11287 7191
rect 11989 7157 12023 7191
rect 13921 7157 13955 7191
rect 18061 7157 18095 7191
rect 21833 7157 21867 7191
rect 26801 7157 26835 7191
rect 27721 7157 27755 7191
rect 29469 7157 29503 7191
rect 33333 7157 33367 7191
rect 35265 7157 35299 7191
rect 38025 7157 38059 7191
rect 2237 6953 2271 6987
rect 5365 6953 5399 6987
rect 5917 6953 5951 6987
rect 10977 6953 11011 6987
rect 12081 6953 12115 6987
rect 13553 6953 13587 6987
rect 13921 6953 13955 6987
rect 16129 6953 16163 6987
rect 16589 6953 16623 6987
rect 18153 6953 18187 6987
rect 23489 6953 23523 6987
rect 25053 6953 25087 6987
rect 25329 6953 25363 6987
rect 27169 6953 27203 6987
rect 28825 6953 28859 6987
rect 34713 6953 34747 6987
rect 35909 6953 35943 6987
rect 28089 6885 28123 6919
rect 29193 6885 29227 6919
rect 3617 6817 3651 6851
rect 5549 6817 5583 6851
rect 8953 6817 8987 6851
rect 9597 6817 9631 6851
rect 11253 6817 11287 6851
rect 12173 6817 12207 6851
rect 14657 6817 14691 6851
rect 15669 6817 15703 6851
rect 17141 6817 17175 6851
rect 17509 6817 17543 6851
rect 17601 6817 17635 6851
rect 18705 6817 18739 6851
rect 21005 6817 21039 6851
rect 22017 6817 22051 6851
rect 22109 6817 22143 6851
rect 22845 6817 22879 6851
rect 22937 6817 22971 6851
rect 25697 6817 25731 6851
rect 26985 6817 27019 6851
rect 27721 6817 27755 6851
rect 30757 6817 30791 6851
rect 31309 6817 31343 6851
rect 32321 6817 32355 6851
rect 33793 6817 33827 6851
rect 35541 6817 35575 6851
rect 37933 6817 37967 6851
rect 3350 6749 3384 6783
rect 3801 6749 3835 6783
rect 5181 6749 5215 6783
rect 5641 6749 5675 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 7021 6749 7055 6783
rect 10425 6749 10459 6783
rect 11529 6749 11563 6783
rect 16405 6749 16439 6783
rect 22201 6749 22235 6783
rect 24041 6749 24075 6783
rect 25973 6749 26007 6783
rect 28457 6749 28491 6783
rect 29377 6749 29411 6783
rect 30113 6749 30147 6783
rect 30665 6749 30699 6783
rect 31769 6749 31803 6783
rect 32505 6749 32539 6783
rect 33241 6749 33275 6783
rect 33977 6749 34011 6783
rect 34529 6749 34563 6783
rect 34897 6749 34931 6783
rect 35449 6749 35483 6783
rect 36093 6749 36127 6783
rect 37565 6749 37599 6783
rect 37749 6749 37783 6783
rect 38301 6749 38335 6783
rect 12440 6681 12474 6715
rect 24593 6681 24627 6715
rect 25881 6681 25915 6715
rect 26433 6681 26467 6715
rect 37298 6681 37332 6715
rect 3985 6613 4019 6647
rect 4537 6613 4571 6647
rect 8309 6613 8343 6647
rect 14105 6613 14139 6647
rect 17693 6613 17727 6647
rect 18061 6613 18095 6647
rect 20637 6613 20671 6647
rect 21281 6613 21315 6647
rect 21649 6613 21683 6647
rect 22569 6613 22603 6647
rect 23029 6613 23063 6647
rect 23397 6613 23431 6647
rect 26341 6613 26375 6647
rect 29745 6613 29779 6647
rect 33057 6613 33091 6647
rect 34069 6613 34103 6647
rect 34989 6613 35023 6647
rect 35357 6613 35391 6647
rect 36185 6613 36219 6647
rect 2145 6409 2179 6443
rect 3157 6409 3191 6443
rect 5457 6409 5491 6443
rect 8861 6409 8895 6443
rect 9321 6409 9355 6443
rect 10517 6409 10551 6443
rect 12357 6409 12391 6443
rect 12725 6409 12759 6443
rect 13185 6409 13219 6443
rect 14841 6409 14875 6443
rect 22937 6409 22971 6443
rect 28549 6409 28583 6443
rect 30205 6409 30239 6443
rect 32965 6409 32999 6443
rect 34069 6409 34103 6443
rect 34897 6409 34931 6443
rect 37933 6409 37967 6443
rect 4292 6341 4326 6375
rect 7297 6341 7331 6375
rect 8585 6341 8619 6375
rect 12817 6341 12851 6375
rect 23397 6341 23431 6375
rect 24869 6341 24903 6375
rect 1961 6273 1995 6307
rect 2145 6273 2179 6307
rect 2605 6273 2639 6307
rect 3065 6273 3099 6307
rect 5273 6273 5307 6307
rect 5733 6273 5767 6307
rect 5825 6273 5859 6307
rect 5917 6273 5951 6307
rect 6101 6273 6135 6307
rect 9229 6273 9263 6307
rect 13829 6273 13863 6307
rect 15485 6273 15519 6307
rect 15577 6273 15611 6307
rect 22293 6273 22327 6307
rect 23581 6273 23615 6307
rect 23857 6273 23891 6307
rect 24685 6273 24719 6307
rect 25789 6273 25823 6307
rect 26249 6273 26283 6307
rect 27905 6273 27939 6307
rect 28365 6273 28399 6307
rect 28733 6273 28767 6307
rect 29193 6273 29227 6307
rect 31769 6273 31803 6307
rect 33149 6273 33183 6307
rect 35449 6273 35483 6307
rect 36369 6273 36403 6307
rect 37289 6273 37323 6307
rect 38209 6273 38243 6307
rect 2697 6205 2731 6239
rect 4537 6205 4571 6239
rect 11253 6205 11287 6239
rect 11529 6205 11563 6239
rect 12173 6205 12207 6239
rect 13001 6205 13035 6239
rect 15853 6205 15887 6239
rect 17601 6205 17635 6239
rect 18245 6205 18279 6239
rect 18705 6205 18739 6239
rect 20821 6205 20855 6239
rect 22017 6205 22051 6239
rect 24501 6205 24535 6239
rect 25973 6205 26007 6239
rect 26157 6205 26191 6239
rect 26985 6205 27019 6239
rect 27537 6205 27571 6239
rect 28089 6205 28123 6239
rect 29009 6205 29043 6239
rect 29653 6205 29687 6239
rect 30849 6205 30883 6239
rect 31585 6205 31619 6239
rect 32689 6205 32723 6239
rect 33517 6205 33551 6239
rect 34713 6205 34747 6239
rect 36185 6205 36219 6239
rect 36921 6205 36955 6239
rect 38393 6205 38427 6239
rect 8217 6137 8251 6171
rect 10241 6137 10275 6171
rect 14473 6137 14507 6171
rect 20269 6137 20303 6171
rect 24133 6137 24167 6171
rect 2329 6069 2363 6103
rect 2789 6069 2823 6103
rect 2881 6069 2915 6103
rect 4721 6069 4755 6103
rect 7757 6069 7791 6103
rect 9781 6069 9815 6103
rect 10701 6069 10735 6103
rect 15117 6069 15151 6103
rect 15301 6069 15335 6103
rect 16497 6069 16531 6103
rect 16957 6069 16991 6103
rect 17693 6069 17727 6103
rect 20545 6069 20579 6103
rect 21373 6069 21407 6103
rect 23213 6069 23247 6103
rect 25145 6069 25179 6103
rect 26617 6069 26651 6103
rect 27721 6069 27755 6103
rect 29377 6069 29411 6103
rect 30297 6069 30331 6103
rect 31033 6069 31067 6103
rect 31953 6069 31987 6103
rect 32137 6069 32171 6103
rect 34161 6069 34195 6103
rect 35633 6069 35667 6103
rect 38025 6069 38059 6103
rect 3617 5865 3651 5899
rect 5641 5865 5675 5899
rect 6377 5865 6411 5899
rect 8217 5865 8251 5899
rect 12633 5865 12667 5899
rect 13001 5865 13035 5899
rect 14473 5865 14507 5899
rect 15761 5865 15795 5899
rect 17693 5865 17727 5899
rect 20913 5865 20947 5899
rect 24225 5865 24259 5899
rect 24409 5865 24443 5899
rect 26341 5865 26375 5899
rect 36185 5865 36219 5899
rect 10517 5797 10551 5831
rect 12357 5797 12391 5831
rect 16773 5797 16807 5831
rect 3341 5729 3375 5763
rect 5181 5729 5215 5763
rect 10425 5729 10459 5763
rect 11161 5729 11195 5763
rect 11713 5729 11747 5763
rect 11897 5729 11931 5763
rect 16313 5729 16347 5763
rect 17049 5729 17083 5763
rect 20085 5729 20119 5763
rect 21465 5729 21499 5763
rect 24133 5729 24167 5763
rect 34161 5729 34195 5763
rect 35541 5729 35575 5763
rect 36369 5729 36403 5763
rect 2513 5661 2547 5695
rect 2667 5661 2701 5695
rect 3433 5661 3467 5695
rect 4914 5661 4948 5695
rect 6745 5661 6779 5695
rect 7573 5661 7607 5695
rect 7849 5661 7883 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 10977 5661 11011 5695
rect 11989 5661 12023 5695
rect 13461 5661 13495 5695
rect 13553 5661 13587 5695
rect 14657 5661 14691 5695
rect 14749 5661 14783 5695
rect 15669 5661 15703 5695
rect 16221 5661 16255 5695
rect 17233 5661 17267 5695
rect 18337 5661 18371 5695
rect 19625 5661 19659 5695
rect 20177 5661 20211 5695
rect 21833 5661 21867 5695
rect 22753 5661 22787 5695
rect 23397 5661 23431 5695
rect 23949 5661 23983 5695
rect 24593 5661 24627 5695
rect 24777 5661 24811 5695
rect 25697 5661 25731 5695
rect 25881 5661 25915 5695
rect 28457 5661 28491 5695
rect 29193 5661 29227 5695
rect 30205 5661 30239 5695
rect 31953 5661 31987 5695
rect 32045 5661 32079 5695
rect 34069 5661 34103 5695
rect 34345 5661 34379 5695
rect 35265 5661 35299 5695
rect 36553 5661 36587 5695
rect 37289 5661 37323 5695
rect 38301 5661 38335 5695
rect 2881 5593 2915 5627
rect 2973 5593 3007 5627
rect 9321 5593 9355 5627
rect 9689 5593 9723 5627
rect 12541 5593 12575 5627
rect 14933 5593 14967 5627
rect 17325 5593 17359 5627
rect 17785 5593 17819 5627
rect 20821 5593 20855 5627
rect 21281 5593 21315 5627
rect 22385 5593 22419 5627
rect 24225 5593 24259 5627
rect 27813 5593 27847 5627
rect 31708 5593 31742 5627
rect 34713 5593 34747 5627
rect 35725 5593 35759 5627
rect 3801 5525 3835 5559
rect 6009 5525 6043 5559
rect 7665 5525 7699 5559
rect 8769 5525 8803 5559
rect 9781 5525 9815 5559
rect 10885 5525 10919 5559
rect 13737 5525 13771 5559
rect 15025 5525 15059 5559
rect 16129 5525 16163 5559
rect 18705 5525 18739 5559
rect 21373 5525 21407 5559
rect 23765 5525 23799 5559
rect 25421 5525 25455 5559
rect 25513 5525 25547 5559
rect 27905 5525 27939 5559
rect 28641 5525 28675 5559
rect 29653 5525 29687 5559
rect 30573 5525 30607 5559
rect 32229 5525 32263 5559
rect 32781 5525 32815 5559
rect 34529 5525 34563 5559
rect 35817 5525 35851 5559
rect 36645 5525 36679 5559
rect 37013 5525 37047 5559
rect 3525 5321 3559 5355
rect 4537 5321 4571 5355
rect 5273 5321 5307 5355
rect 8033 5321 8067 5355
rect 8953 5321 8987 5355
rect 10517 5321 10551 5355
rect 11069 5321 11103 5355
rect 12357 5321 12391 5355
rect 12817 5321 12851 5355
rect 18061 5321 18095 5355
rect 21833 5321 21867 5355
rect 26249 5321 26283 5355
rect 27721 5321 27755 5355
rect 30849 5321 30883 5355
rect 31677 5321 31711 5355
rect 32413 5321 32447 5355
rect 32873 5321 32907 5355
rect 37565 5321 37599 5355
rect 14749 5253 14783 5287
rect 16497 5253 16531 5287
rect 21281 5253 21315 5287
rect 22385 5253 22419 5287
rect 29736 5253 29770 5287
rect 34406 5253 34440 5287
rect 2973 5185 3007 5219
rect 3164 5185 3198 5219
rect 3311 5185 3345 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 4721 5185 4755 5219
rect 5733 5185 5767 5219
rect 5917 5185 5951 5219
rect 6009 5185 6043 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6929 5185 6963 5219
rect 8677 5185 8711 5219
rect 8769 5185 8803 5219
rect 10977 5185 11011 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12449 5185 12483 5219
rect 13645 5185 13679 5219
rect 14381 5185 14415 5219
rect 16948 5185 16982 5219
rect 18705 5185 18739 5219
rect 19073 5185 19107 5219
rect 22017 5185 22051 5219
rect 23489 5185 23523 5219
rect 24685 5185 24719 5219
rect 24869 5185 24903 5219
rect 25136 5185 25170 5219
rect 26525 5185 26559 5219
rect 26709 5185 26743 5219
rect 27353 5185 27387 5219
rect 28549 5185 28583 5219
rect 29469 5185 29503 5219
rect 31309 5185 31343 5219
rect 31953 5185 31987 5219
rect 32505 5185 32539 5219
rect 33517 5185 33551 5219
rect 33885 5185 33919 5219
rect 33977 5185 34011 5219
rect 34161 5185 34195 5219
rect 37105 5185 37139 5219
rect 37289 5185 37323 5219
rect 38485 5185 38519 5219
rect 2697 5117 2731 5151
rect 2881 5117 2915 5151
rect 7481 5117 7515 5151
rect 9229 5117 9263 5151
rect 9873 5117 9907 5151
rect 11161 5117 11195 5151
rect 12173 5117 12207 5151
rect 13461 5117 13495 5151
rect 14197 5117 14231 5151
rect 16681 5117 16715 5151
rect 18521 5117 18555 5151
rect 19257 5117 19291 5151
rect 20085 5117 20119 5151
rect 20269 5117 20303 5151
rect 20821 5117 20855 5151
rect 21373 5117 21407 5151
rect 21557 5117 21591 5151
rect 23121 5117 23155 5151
rect 24225 5117 24259 5151
rect 27077 5117 27111 5151
rect 27261 5117 27295 5151
rect 28365 5117 28399 5151
rect 29101 5117 29135 5151
rect 31033 5117 31067 5151
rect 31217 5117 31251 5151
rect 32229 5117 32263 5151
rect 36645 5117 36679 5151
rect 38117 5117 38151 5151
rect 2789 5049 2823 5083
rect 5641 5049 5675 5083
rect 7941 5049 7975 5083
rect 10609 5049 10643 5083
rect 20913 5049 20947 5083
rect 31769 5049 31803 5083
rect 3617 4981 3651 5015
rect 3893 4981 3927 5015
rect 4445 4981 4479 5015
rect 6009 4981 6043 5015
rect 6561 4981 6595 5015
rect 9781 4981 9815 5015
rect 11989 4981 12023 5015
rect 12909 4981 12943 5015
rect 14565 4981 14599 5015
rect 18337 4981 18371 5015
rect 18889 4981 18923 5015
rect 19441 4981 19475 5015
rect 24501 4981 24535 5015
rect 26341 4981 26375 5015
rect 27813 4981 27847 5015
rect 32965 4981 32999 5015
rect 33701 4981 33735 5015
rect 35541 4981 35575 5015
rect 37473 4981 37507 5015
rect 38301 4981 38335 5015
rect 3249 4777 3283 4811
rect 8585 4777 8619 4811
rect 11069 4777 11103 4811
rect 16497 4777 16531 4811
rect 19349 4777 19383 4811
rect 21005 4777 21039 4811
rect 23121 4777 23155 4811
rect 24685 4777 24719 4811
rect 28917 4777 28951 4811
rect 29285 4777 29319 4811
rect 29653 4777 29687 4811
rect 32321 4777 32355 4811
rect 33701 4777 33735 4811
rect 34529 4777 34563 4811
rect 35173 4777 35207 4811
rect 4169 4709 4203 4743
rect 4997 4709 5031 4743
rect 26709 4709 26743 4743
rect 32413 4709 32447 4743
rect 36369 4709 36403 4743
rect 3617 4641 3651 4675
rect 4813 4641 4847 4675
rect 6193 4641 6227 4675
rect 7113 4641 7147 4675
rect 9689 4641 9723 4675
rect 11161 4641 11195 4675
rect 11805 4641 11839 4675
rect 12081 4641 12115 4675
rect 12198 4641 12232 4675
rect 13553 4641 13587 4675
rect 13737 4641 13771 4675
rect 14473 4641 14507 4675
rect 17233 4641 17267 4675
rect 17785 4641 17819 4675
rect 18245 4641 18279 4675
rect 18521 4641 18555 4675
rect 19625 4641 19659 4675
rect 21879 4641 21913 4675
rect 22017 4641 22051 4675
rect 22293 4641 22327 4675
rect 22753 4641 22787 4675
rect 23489 4641 23523 4675
rect 23673 4641 23707 4675
rect 25329 4641 25363 4675
rect 27169 4641 27203 4675
rect 29285 4641 29319 4675
rect 30113 4641 30147 4675
rect 30205 4641 30239 4675
rect 30665 4641 30699 4675
rect 31125 4641 31159 4675
rect 31539 4641 31573 4675
rect 32873 4641 32907 4675
rect 33057 4641 33091 4675
rect 33609 4641 33643 4675
rect 33885 4641 33919 4675
rect 34069 4641 34103 4675
rect 35081 4641 35115 4675
rect 35817 4641 35851 4675
rect 35976 4641 36010 4675
rect 37105 4641 37139 4675
rect 3985 4573 4019 4607
rect 4353 4573 4387 4607
rect 4629 4573 4663 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 5641 4573 5675 4607
rect 6377 4573 6411 4607
rect 7205 4573 7239 4607
rect 9137 4573 9171 4607
rect 9321 4573 9355 4607
rect 9945 4573 9979 4607
rect 11345 4573 11379 4607
rect 12357 4573 12391 4607
rect 13001 4573 13035 4607
rect 13461 4573 13495 4607
rect 14105 4573 14139 4607
rect 15117 4573 15151 4607
rect 17371 4573 17405 4607
rect 17509 4573 17543 4607
rect 18429 4573 18463 4607
rect 18705 4573 18739 4607
rect 19533 4573 19567 4607
rect 19881 4573 19915 4607
rect 21741 4573 21775 4607
rect 22937 4573 22971 4607
rect 23213 4573 23247 4607
rect 25145 4573 25179 4607
rect 26157 4573 26191 4607
rect 26295 4573 26329 4607
rect 26433 4573 26467 4607
rect 27353 4573 27387 4607
rect 28558 4573 28592 4607
rect 28825 4573 28859 4607
rect 29101 4573 29135 4607
rect 30481 4573 30515 4607
rect 31401 4573 31435 4607
rect 31677 4573 31711 4607
rect 32781 4573 32815 4607
rect 33425 4573 33459 4607
rect 33701 4573 33735 4607
rect 34161 4573 34195 4607
rect 34897 4573 34931 4607
rect 36093 4573 36127 4607
rect 36829 4573 36863 4607
rect 37013 4573 37047 4607
rect 4997 4505 5031 4539
rect 7450 4505 7484 4539
rect 15384 4505 15418 4539
rect 29377 4505 29411 4539
rect 37350 4505 37384 4539
rect 2881 4437 2915 4471
rect 3801 4437 3835 4471
rect 4445 4437 4479 4471
rect 5181 4437 5215 4471
rect 5457 4437 5491 4471
rect 5825 4437 5859 4471
rect 6469 4437 6503 4471
rect 9505 4437 9539 4471
rect 13093 4437 13127 4471
rect 14289 4437 14323 4471
rect 15025 4437 15059 4471
rect 16589 4437 16623 4471
rect 18889 4437 18923 4471
rect 21097 4437 21131 4471
rect 23765 4437 23799 4471
rect 24133 4437 24167 4471
rect 25053 4437 25087 4471
rect 25513 4437 25547 4471
rect 27445 4437 27479 4471
rect 30021 4437 30055 4471
rect 33241 4437 33275 4471
rect 34713 4437 34747 4471
rect 38485 4437 38519 4471
rect 6577 4233 6611 4267
rect 6837 4233 6871 4267
rect 11621 4233 11655 4267
rect 18061 4233 18095 4267
rect 18521 4233 18555 4267
rect 18889 4233 18923 4267
rect 19533 4233 19567 4267
rect 20269 4233 20303 4267
rect 23673 4233 23707 4267
rect 26985 4233 27019 4267
rect 27353 4233 27387 4267
rect 32137 4233 32171 4267
rect 33333 4233 33367 4267
rect 33609 4233 33643 4267
rect 37289 4233 37323 4267
rect 37657 4233 37691 4267
rect 3065 4165 3099 4199
rect 3525 4165 3559 4199
rect 6377 4165 6411 4199
rect 9229 4165 9263 4199
rect 10210 4165 10244 4199
rect 12734 4165 12768 4199
rect 19441 4165 19475 4199
rect 23765 4165 23799 4199
rect 26433 4165 26467 4199
rect 28181 4165 28215 4199
rect 28365 4165 28399 4199
rect 2697 4097 2731 4131
rect 3433 4097 3467 4131
rect 3709 4097 3743 4131
rect 4537 4097 4571 4131
rect 4813 4097 4847 4131
rect 5181 4097 5215 4131
rect 6101 4097 6135 4131
rect 7950 4097 7984 4131
rect 8217 4097 8251 4131
rect 8493 4097 8527 4131
rect 9413 4097 9447 4131
rect 9682 4097 9716 4131
rect 9965 4097 9999 4131
rect 13001 4097 13035 4131
rect 13645 4097 13679 4131
rect 14657 4097 14691 4131
rect 15669 4097 15703 4131
rect 16129 4097 16163 4131
rect 16221 4097 16255 4131
rect 16681 4097 16715 4131
rect 16948 4097 16982 4131
rect 18429 4097 18463 4131
rect 19165 4097 19199 4131
rect 19717 4097 19751 4131
rect 19993 4097 20027 4131
rect 21382 4097 21416 4131
rect 22100 4097 22134 4131
rect 24317 4097 24351 4131
rect 24501 4097 24535 4131
rect 24593 4097 24627 4131
rect 24860 4097 24894 4131
rect 26525 4097 26559 4131
rect 27997 4097 28031 4131
rect 29552 4097 29586 4131
rect 31125 4097 31159 4131
rect 31217 4097 31251 4131
rect 31769 4097 31803 4131
rect 31953 4097 31987 4131
rect 32689 4097 32723 4131
rect 33425 4097 33459 4131
rect 33793 4097 33827 4131
rect 33885 4097 33919 4131
rect 34152 4097 34186 4131
rect 35357 4097 35391 4131
rect 35624 4097 35658 4131
rect 37105 4097 37139 4131
rect 38301 4097 38335 4131
rect 4261 4029 4295 4063
rect 4905 4029 4939 4063
rect 5549 4029 5583 4063
rect 9505 4029 9539 4063
rect 14473 4029 14507 4063
rect 15025 4029 15059 4063
rect 16313 4029 16347 4063
rect 18245 4029 18279 4063
rect 19349 4029 19383 4063
rect 19809 4029 19843 4063
rect 21649 4029 21683 4063
rect 21833 4029 21867 4063
rect 23857 4029 23891 4063
rect 26709 4029 26743 4063
rect 27445 4029 27479 4063
rect 27537 4029 27571 4063
rect 28549 4029 28583 4063
rect 29285 4029 29319 4063
rect 31401 4029 31435 4063
rect 37749 4029 37783 4063
rect 37933 4029 37967 4063
rect 38485 4029 38519 4063
rect 2237 3961 2271 3995
rect 4997 3961 5031 3995
rect 6745 3961 6779 3995
rect 9873 3961 9907 3995
rect 11345 3961 11379 3995
rect 15761 3961 15795 3995
rect 23213 3961 23247 3995
rect 25973 3961 26007 3995
rect 29193 3961 29227 3995
rect 31585 3961 31619 3995
rect 36737 3961 36771 3995
rect 2605 3893 2639 3927
rect 2789 3893 2823 3927
rect 3893 3893 3927 3927
rect 3985 3893 4019 3927
rect 4169 3893 4203 3927
rect 4629 3893 4663 3927
rect 5365 3893 5399 3927
rect 6561 3893 6595 3927
rect 9413 3893 9447 3927
rect 13093 3893 13127 3927
rect 13921 3893 13955 3927
rect 14841 3893 14875 3927
rect 18981 3893 19015 3927
rect 19349 3893 19383 3927
rect 20177 3893 20211 3927
rect 23305 3893 23339 3927
rect 24133 3893 24167 3927
rect 26065 3893 26099 3927
rect 30665 3893 30699 3927
rect 30757 3893 30791 3927
rect 33149 3893 33183 3927
rect 35265 3893 35299 3927
rect 36921 3893 36955 3927
rect 38117 3893 38151 3927
rect 2145 3689 2179 3723
rect 2881 3689 2915 3723
rect 3433 3689 3467 3723
rect 3617 3689 3651 3723
rect 9137 3689 9171 3723
rect 14381 3689 14415 3723
rect 17969 3689 18003 3723
rect 20729 3689 20763 3723
rect 22201 3689 22235 3723
rect 24409 3689 24443 3723
rect 25145 3689 25179 3723
rect 26893 3689 26927 3723
rect 29193 3689 29227 3723
rect 29653 3689 29687 3723
rect 31401 3689 31435 3723
rect 32873 3689 32907 3723
rect 34713 3689 34747 3723
rect 37749 3689 37783 3723
rect 2421 3621 2455 3655
rect 7389 3621 7423 3655
rect 8309 3621 8343 3655
rect 10057 3621 10091 3655
rect 11069 3621 11103 3655
rect 12633 3621 12667 3655
rect 17877 3621 17911 3655
rect 23029 3621 23063 3655
rect 26801 3621 26835 3655
rect 3065 3553 3099 3587
rect 3801 3553 3835 3587
rect 4997 3553 5031 3587
rect 6009 3553 6043 3587
rect 8401 3553 8435 3587
rect 12449 3553 12483 3587
rect 12909 3553 12943 3587
rect 14749 3553 14783 3587
rect 17233 3553 17267 3587
rect 17417 3553 17451 3587
rect 18521 3553 18555 3587
rect 18705 3553 18739 3587
rect 22385 3553 22419 3587
rect 23673 3553 23707 3587
rect 25421 3553 25455 3587
rect 27445 3553 27479 3587
rect 29009 3553 29043 3587
rect 32689 3553 32723 3587
rect 35265 3553 35299 3587
rect 35541 3553 35575 3587
rect 35909 3553 35943 3587
rect 38209 3553 38243 3587
rect 1869 3485 1903 3519
rect 1961 3485 1995 3519
rect 2237 3485 2271 3519
rect 2697 3485 2731 3519
rect 3893 3485 3927 3519
rect 4077 3485 4111 3519
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 5733 3485 5767 3519
rect 5917 3485 5951 3519
rect 6285 3485 6319 3519
rect 8033 3485 8067 3519
rect 8125 3485 8159 3519
rect 8585 3485 8619 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9781 3485 9815 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 12193 3485 12227 3519
rect 12817 3485 12851 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 14381 3485 14415 3519
rect 14473 3485 14507 3519
rect 15301 3485 15335 3519
rect 17049 3485 17083 3519
rect 17509 3485 17543 3519
rect 18889 3485 18923 3519
rect 19257 3485 19291 3519
rect 20085 3485 20119 3519
rect 20821 3485 20855 3519
rect 22569 3485 22603 3519
rect 24041 3485 24075 3519
rect 24225 3485 24259 3519
rect 24961 3485 24995 3519
rect 25329 3485 25363 3519
rect 27629 3485 27663 3519
rect 28365 3485 28399 3519
rect 29377 3485 29411 3519
rect 29837 3485 29871 3519
rect 31309 3485 31343 3519
rect 31953 3485 31987 3519
rect 33057 3485 33091 3519
rect 34437 3485 34471 3519
rect 35081 3485 35115 3519
rect 35725 3485 35759 3519
rect 37473 3485 37507 3519
rect 37749 3485 37783 3519
rect 38117 3485 38151 3519
rect 4721 3417 4755 3451
rect 5181 3417 5215 3451
rect 14657 3417 14691 3451
rect 16782 3417 16816 3451
rect 21088 3417 21122 3451
rect 25688 3417 25722 3451
rect 31064 3417 31098 3451
rect 32137 3417 32171 3451
rect 33609 3417 33643 3451
rect 36277 3417 36311 3451
rect 1685 3349 1719 3383
rect 3433 3349 3467 3383
rect 5089 3349 5123 3383
rect 5365 3349 5399 3383
rect 5549 3349 5583 3383
rect 8769 3349 8803 3383
rect 10977 3349 11011 3383
rect 13921 3349 13955 3383
rect 14197 3349 14231 3383
rect 15669 3349 15703 3383
rect 19073 3349 19107 3383
rect 19901 3349 19935 3383
rect 22661 3349 22695 3383
rect 23121 3349 23155 3383
rect 23857 3349 23891 3383
rect 28273 3349 28307 3383
rect 29929 3349 29963 3383
rect 35173 3349 35207 3383
rect 37565 3349 37599 3383
rect 1777 3145 1811 3179
rect 2421 3145 2455 3179
rect 5549 3145 5583 3179
rect 6377 3145 6411 3179
rect 7113 3145 7147 3179
rect 11253 3145 11287 3179
rect 11713 3145 11747 3179
rect 17141 3145 17175 3179
rect 19441 3145 19475 3179
rect 21833 3145 21867 3179
rect 22109 3145 22143 3179
rect 24961 3145 24995 3179
rect 26617 3145 26651 3179
rect 26985 3145 27019 3179
rect 30205 3145 30239 3179
rect 36461 3145 36495 3179
rect 2329 3077 2363 3111
rect 3617 3077 3651 3111
rect 16681 3077 16715 3111
rect 37289 3077 37323 3111
rect 1501 3009 1535 3043
rect 2053 3009 2087 3043
rect 2605 3009 2639 3043
rect 2697 3009 2731 3043
rect 3157 3009 3191 3043
rect 3433 3009 3467 3043
rect 4905 3009 4939 3043
rect 5273 3009 5307 3043
rect 7297 3009 7331 3043
rect 7481 3009 7515 3043
rect 7573 3009 7607 3043
rect 7849 3009 7883 3043
rect 8033 3009 8067 3043
rect 8125 3009 8159 3043
rect 9689 3009 9723 3043
rect 11069 3009 11103 3043
rect 11529 3009 11563 3043
rect 11805 3009 11839 3043
rect 13277 3009 13311 3043
rect 13737 3009 13771 3043
rect 15301 3009 15335 3043
rect 16957 3009 16991 3043
rect 18705 3009 18739 3043
rect 19533 3009 19567 3043
rect 22017 3009 22051 3043
rect 22661 3009 22695 3043
rect 24133 3009 24167 3043
rect 26341 3009 26375 3043
rect 26801 3009 26835 3043
rect 27169 3009 27203 3043
rect 27445 3009 27479 3043
rect 30113 3009 30147 3043
rect 30389 3009 30423 3043
rect 31769 3009 31803 3043
rect 32597 3009 32631 3043
rect 34161 3009 34195 3043
rect 34897 3009 34931 3043
rect 36369 3009 36403 3043
rect 38025 3009 38059 3043
rect 38209 3009 38243 3043
rect 38393 3009 38427 3043
rect 3065 2941 3099 2975
rect 3249 2941 3283 2975
rect 3893 2941 3927 2975
rect 6193 2941 6227 2975
rect 6929 2941 6963 2975
rect 7665 2941 7699 2975
rect 8585 2941 8619 2975
rect 10057 2941 10091 2975
rect 12265 2941 12299 2975
rect 14105 2941 14139 2975
rect 15577 2941 15611 2975
rect 16773 2941 16807 2975
rect 17509 2941 17543 2975
rect 18889 2941 18923 2975
rect 20085 2941 20119 2975
rect 21097 2941 21131 2975
rect 23029 2941 23063 2975
rect 24409 2941 24443 2975
rect 25237 2941 25271 2975
rect 27721 2941 27755 2975
rect 28917 2941 28951 2975
rect 30757 2941 30791 2975
rect 32505 2941 32539 2975
rect 32965 2941 32999 2975
rect 34253 2941 34287 2975
rect 35173 2941 35207 2975
rect 37013 2941 37047 2975
rect 37933 2941 37967 2975
rect 2513 2873 2547 2907
rect 2789 2873 2823 2907
rect 21649 2873 21683 2907
rect 32229 2873 32263 2907
rect 2237 2805 2271 2839
rect 3157 2805 3191 2839
rect 5457 2805 5491 2839
rect 13461 2805 13495 2839
rect 16681 2805 16715 2839
rect 32597 2805 32631 2839
rect 2973 2601 3007 2635
rect 3801 2601 3835 2635
rect 8769 2601 8803 2635
rect 9137 2601 9171 2635
rect 11713 2601 11747 2635
rect 14381 2601 14415 2635
rect 16957 2601 16991 2635
rect 19257 2601 19291 2635
rect 20177 2601 20211 2635
rect 23305 2601 23339 2635
rect 24225 2601 24259 2635
rect 25881 2601 25915 2635
rect 26617 2601 26651 2635
rect 29101 2601 29135 2635
rect 31033 2601 31067 2635
rect 33609 2601 33643 2635
rect 34345 2601 34379 2635
rect 36185 2601 36219 2635
rect 36921 2601 36955 2635
rect 37289 2601 37323 2635
rect 38025 2601 38059 2635
rect 4077 2533 4111 2567
rect 6561 2533 6595 2567
rect 12449 2533 12483 2567
rect 16865 2533 16899 2567
rect 19809 2533 19843 2567
rect 31769 2533 31803 2567
rect 1961 2465 1995 2499
rect 7113 2465 7147 2499
rect 10609 2465 10643 2499
rect 13001 2465 13035 2499
rect 18337 2465 18371 2499
rect 20729 2465 20763 2499
rect 23857 2465 23891 2499
rect 27629 2465 27663 2499
rect 30021 2465 30055 2499
rect 35173 2465 35207 2499
rect 36737 2465 36771 2499
rect 37841 2465 37875 2499
rect 1685 2397 1719 2431
rect 3525 2397 3559 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 8125 2397 8159 2431
rect 8953 2397 8987 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 11529 2397 11563 2431
rect 12081 2397 12115 2431
rect 12541 2397 12575 2431
rect 14105 2397 14139 2431
rect 15025 2397 15059 2431
rect 15301 2397 15335 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 20269 2397 20303 2431
rect 23213 2397 23247 2431
rect 24041 2397 24075 2431
rect 25605 2397 25639 2431
rect 26433 2397 26467 2431
rect 26801 2397 26835 2431
rect 26985 2397 27019 2431
rect 28457 2397 28491 2431
rect 29193 2397 29227 2431
rect 29745 2397 29779 2431
rect 31585 2397 31619 2431
rect 31953 2397 31987 2431
rect 33517 2397 33551 2431
rect 34161 2397 34195 2431
rect 34529 2397 34563 2431
rect 34713 2397 34747 2431
rect 37105 2397 37139 2431
rect 38209 2397 38243 2431
rect 38393 2397 38427 2431
rect 5089 2329 5123 2363
rect 9873 2329 9907 2363
rect 16129 2329 16163 2363
rect 22109 2329 22143 2363
rect 24593 2329 24627 2363
rect 32321 2329 32355 2363
rect 14289 2261 14323 2295
rect 29377 2261 29411 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 37001 32419 37059 32425
rect 37001 32385 37013 32419
rect 37047 32416 37059 32419
rect 37366 32416 37372 32428
rect 37047 32388 37372 32416
rect 37047 32385 37059 32388
rect 37001 32379 37059 32385
rect 37366 32376 37372 32388
rect 37424 32376 37430 32428
rect 14090 32308 14096 32360
rect 14148 32308 14154 32360
rect 14921 32351 14979 32357
rect 14921 32317 14933 32351
rect 14967 32348 14979 32351
rect 15010 32348 15016 32360
rect 14967 32320 15016 32348
rect 14967 32317 14979 32320
rect 14921 32311 14979 32317
rect 15010 32308 15016 32320
rect 15068 32308 15074 32360
rect 24578 32308 24584 32360
rect 24636 32308 24642 32360
rect 24765 32351 24823 32357
rect 24765 32317 24777 32351
rect 24811 32317 24823 32351
rect 24765 32311 24823 32317
rect 28169 32351 28227 32357
rect 28169 32317 28181 32351
rect 28215 32348 28227 32351
rect 28442 32348 28448 32360
rect 28215 32320 28448 32348
rect 28215 32317 28227 32320
rect 28169 32311 28227 32317
rect 23934 32240 23940 32292
rect 23992 32280 23998 32292
rect 24780 32280 24808 32311
rect 28442 32308 28448 32320
rect 28500 32308 28506 32360
rect 28810 32308 28816 32360
rect 28868 32308 28874 32360
rect 36630 32308 36636 32360
rect 36688 32348 36694 32360
rect 37277 32351 37335 32357
rect 37277 32348 37289 32351
rect 36688 32320 37289 32348
rect 36688 32308 36694 32320
rect 37277 32317 37289 32320
rect 37323 32317 37335 32351
rect 37277 32311 37335 32317
rect 23992 32252 24808 32280
rect 23992 32240 23998 32252
rect 10042 32172 10048 32224
rect 10100 32212 10106 32224
rect 10321 32215 10379 32221
rect 10321 32212 10333 32215
rect 10100 32184 10333 32212
rect 10100 32172 10106 32184
rect 10321 32181 10333 32184
rect 10367 32181 10379 32215
rect 10321 32175 10379 32181
rect 13446 32172 13452 32224
rect 13504 32172 13510 32224
rect 14274 32172 14280 32224
rect 14332 32172 14338 32224
rect 24026 32172 24032 32224
rect 24084 32172 24090 32224
rect 25406 32172 25412 32224
rect 25464 32172 25470 32224
rect 26602 32172 26608 32224
rect 26660 32212 26666 32224
rect 26697 32215 26755 32221
rect 26697 32212 26709 32215
rect 26660 32184 26709 32212
rect 26660 32172 26666 32184
rect 26697 32181 26709 32184
rect 26743 32181 26755 32215
rect 26697 32175 26755 32181
rect 27062 32172 27068 32224
rect 27120 32212 27126 32224
rect 27341 32215 27399 32221
rect 27341 32212 27353 32215
rect 27120 32184 27353 32212
rect 27120 32172 27126 32184
rect 27341 32181 27353 32184
rect 27387 32181 27399 32215
rect 27341 32175 27399 32181
rect 27522 32172 27528 32224
rect 27580 32172 27586 32224
rect 28258 32172 28264 32224
rect 28316 32172 28322 32224
rect 36354 32172 36360 32224
rect 36412 32172 36418 32224
rect 37734 32172 37740 32224
rect 37792 32212 37798 32224
rect 37921 32215 37979 32221
rect 37921 32212 37933 32215
rect 37792 32184 37933 32212
rect 37792 32172 37798 32184
rect 37921 32181 37933 32184
rect 37967 32181 37979 32215
rect 37921 32175 37979 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 14090 31968 14096 32020
rect 14148 31968 14154 32020
rect 14274 31968 14280 32020
rect 14332 31968 14338 32020
rect 23934 31968 23940 32020
rect 23992 31968 23998 32020
rect 24026 31968 24032 32020
rect 24084 31968 24090 32020
rect 28258 31968 28264 32020
rect 28316 31968 28322 32020
rect 28442 31968 28448 32020
rect 28500 31968 28506 32020
rect 10042 31900 10048 31952
rect 10100 31940 10106 31952
rect 13081 31943 13139 31949
rect 13081 31940 13093 31943
rect 10100 31912 13093 31940
rect 10100 31900 10106 31912
rect 13081 31909 13093 31912
rect 13127 31940 13139 31943
rect 13127 31912 14228 31940
rect 13127 31909 13139 31912
rect 13081 31903 13139 31909
rect 10321 31807 10379 31813
rect 10321 31773 10333 31807
rect 10367 31804 10379 31807
rect 10410 31804 10416 31816
rect 10367 31776 10416 31804
rect 10367 31773 10379 31776
rect 10321 31767 10379 31773
rect 10410 31764 10416 31776
rect 10468 31764 10474 31816
rect 11238 31764 11244 31816
rect 11296 31764 11302 31816
rect 13906 31764 13912 31816
rect 13964 31764 13970 31816
rect 14200 31804 14228 31912
rect 14292 31872 14320 31968
rect 14553 31875 14611 31881
rect 14553 31872 14565 31875
rect 14292 31844 14565 31872
rect 14553 31841 14565 31844
rect 14599 31841 14611 31875
rect 14553 31835 14611 31841
rect 14645 31875 14703 31881
rect 14645 31841 14657 31875
rect 14691 31841 14703 31875
rect 14645 31835 14703 31841
rect 23385 31875 23443 31881
rect 23385 31841 23397 31875
rect 23431 31841 23443 31875
rect 23385 31835 23443 31841
rect 23477 31875 23535 31881
rect 23477 31841 23489 31875
rect 23523 31872 23535 31875
rect 24044 31872 24072 31968
rect 26881 31943 26939 31949
rect 26881 31909 26893 31943
rect 26927 31909 26939 31943
rect 26881 31903 26939 31909
rect 27080 31912 27844 31940
rect 23523 31844 24072 31872
rect 23523 31841 23535 31844
rect 23477 31835 23535 31841
rect 14660 31804 14688 31835
rect 14200 31776 14688 31804
rect 15562 31764 15568 31816
rect 15620 31764 15626 31816
rect 19058 31764 19064 31816
rect 19116 31764 19122 31816
rect 19242 31764 19248 31816
rect 19300 31804 19306 31816
rect 19705 31807 19763 31813
rect 19705 31804 19717 31807
rect 19300 31776 19717 31804
rect 19300 31764 19306 31776
rect 19705 31773 19717 31776
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31804 23167 31807
rect 23400 31804 23428 31835
rect 24762 31832 24768 31884
rect 24820 31832 24826 31884
rect 26602 31832 26608 31884
rect 26660 31832 26666 31884
rect 26789 31875 26847 31881
rect 26789 31841 26801 31875
rect 26835 31872 26847 31875
rect 26896 31872 26924 31903
rect 27080 31884 27108 31912
rect 26835 31844 26924 31872
rect 26835 31841 26847 31844
rect 26789 31835 26847 31841
rect 27062 31832 27068 31884
rect 27120 31832 27126 31884
rect 27816 31881 27844 31912
rect 27433 31875 27491 31881
rect 27433 31841 27445 31875
rect 27479 31841 27491 31875
rect 27433 31835 27491 31841
rect 27801 31875 27859 31881
rect 27801 31841 27813 31875
rect 27847 31841 27859 31875
rect 27801 31835 27859 31841
rect 27985 31875 28043 31881
rect 27985 31841 27997 31875
rect 28031 31872 28043 31875
rect 28276 31872 28304 31968
rect 28031 31844 28304 31872
rect 28031 31841 28043 31844
rect 27985 31835 28043 31841
rect 24780 31804 24808 31832
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 23155 31776 24808 31804
rect 24872 31776 24961 31804
rect 23155 31773 23167 31776
rect 23109 31767 23167 31773
rect 12805 31739 12863 31745
rect 12805 31705 12817 31739
rect 12851 31736 12863 31739
rect 14461 31739 14519 31745
rect 12851 31708 13676 31736
rect 12851 31705 12863 31708
rect 12805 31699 12863 31705
rect 13648 31680 13676 31708
rect 14461 31705 14473 31739
rect 14507 31736 14519 31739
rect 14734 31736 14740 31748
rect 14507 31708 14740 31736
rect 14507 31705 14519 31708
rect 14461 31699 14519 31705
rect 14734 31696 14740 31708
rect 14792 31696 14798 31748
rect 23934 31696 23940 31748
rect 23992 31736 23998 31748
rect 24872 31736 24900 31776
rect 24949 31773 24961 31776
rect 24995 31773 25007 31807
rect 24949 31767 25007 31773
rect 25222 31764 25228 31816
rect 25280 31804 25286 31816
rect 25685 31807 25743 31813
rect 25685 31804 25697 31807
rect 25280 31776 25697 31804
rect 25280 31764 25286 31776
rect 25685 31773 25697 31776
rect 25731 31773 25743 31807
rect 25685 31767 25743 31773
rect 26145 31807 26203 31813
rect 26145 31773 26157 31807
rect 26191 31804 26203 31807
rect 26326 31804 26332 31816
rect 26191 31776 26332 31804
rect 26191 31773 26203 31776
rect 26145 31767 26203 31773
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 26620 31804 26648 31832
rect 27448 31804 27476 31835
rect 34698 31832 34704 31884
rect 34756 31872 34762 31884
rect 35989 31875 36047 31881
rect 35989 31872 36001 31875
rect 34756 31844 36001 31872
rect 34756 31832 34762 31844
rect 35989 31841 36001 31844
rect 36035 31841 36047 31875
rect 35989 31835 36047 31841
rect 26620 31776 27476 31804
rect 29178 31764 29184 31816
rect 29236 31764 29242 31816
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 31941 31807 31999 31813
rect 31941 31804 31953 31807
rect 31812 31776 31953 31804
rect 31812 31764 31818 31776
rect 31941 31773 31953 31776
rect 31987 31773 31999 31807
rect 31941 31767 31999 31773
rect 32030 31764 32036 31816
rect 32088 31804 32094 31816
rect 32493 31807 32551 31813
rect 32493 31804 32505 31807
rect 32088 31776 32505 31804
rect 32088 31764 32094 31776
rect 32493 31773 32505 31776
rect 32539 31773 32551 31807
rect 32493 31767 32551 31773
rect 35434 31764 35440 31816
rect 35492 31804 35498 31816
rect 35805 31807 35863 31813
rect 35805 31804 35817 31807
rect 35492 31776 35817 31804
rect 35492 31764 35498 31776
rect 35805 31773 35817 31776
rect 35851 31773 35863 31807
rect 35805 31767 35863 31773
rect 36446 31764 36452 31816
rect 36504 31804 36510 31816
rect 36541 31807 36599 31813
rect 36541 31804 36553 31807
rect 36504 31776 36553 31804
rect 36504 31764 36510 31776
rect 36541 31773 36553 31776
rect 36587 31773 36599 31807
rect 36541 31767 36599 31773
rect 36722 31764 36728 31816
rect 36780 31764 36786 31816
rect 36906 31764 36912 31816
rect 36964 31804 36970 31816
rect 37277 31807 37335 31813
rect 37277 31804 37289 31807
rect 36964 31776 37289 31804
rect 36964 31764 36970 31776
rect 37277 31773 37289 31776
rect 37323 31773 37335 31807
rect 37277 31767 37335 31773
rect 37458 31764 37464 31816
rect 37516 31764 37522 31816
rect 38102 31764 38108 31816
rect 38160 31764 38166 31816
rect 23992 31708 24900 31736
rect 27249 31739 27307 31745
rect 23992 31696 23998 31708
rect 27249 31705 27261 31739
rect 27295 31736 27307 31739
rect 29270 31736 29276 31748
rect 27295 31708 29276 31736
rect 27295 31705 27307 31708
rect 27249 31699 27307 31705
rect 29270 31696 29276 31708
rect 29328 31696 29334 31748
rect 9674 31628 9680 31680
rect 9732 31628 9738 31680
rect 10594 31628 10600 31680
rect 10652 31628 10658 31680
rect 13262 31628 13268 31680
rect 13320 31628 13326 31680
rect 13630 31628 13636 31680
rect 13688 31628 13694 31680
rect 14642 31628 14648 31680
rect 14700 31668 14706 31680
rect 15013 31671 15071 31677
rect 15013 31668 15025 31671
rect 14700 31640 15025 31668
rect 14700 31628 14706 31640
rect 15013 31637 15025 31640
rect 15059 31637 15071 31671
rect 15013 31631 15071 31637
rect 18417 31671 18475 31677
rect 18417 31637 18429 31671
rect 18463 31668 18475 31671
rect 18506 31668 18512 31680
rect 18463 31640 18512 31668
rect 18463 31637 18475 31640
rect 18417 31631 18475 31637
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 19334 31628 19340 31680
rect 19392 31668 19398 31680
rect 19521 31671 19579 31677
rect 19521 31668 19533 31671
rect 19392 31640 19533 31668
rect 19392 31628 19398 31640
rect 19521 31637 19533 31640
rect 19567 31637 19579 31671
rect 19521 31631 19579 31637
rect 20346 31628 20352 31680
rect 20404 31628 20410 31680
rect 23569 31671 23627 31677
rect 23569 31637 23581 31671
rect 23615 31668 23627 31671
rect 23658 31668 23664 31680
rect 23615 31640 23664 31668
rect 23615 31637 23627 31640
rect 23569 31631 23627 31637
rect 23658 31628 23664 31640
rect 23716 31628 23722 31680
rect 24394 31628 24400 31680
rect 24452 31628 24458 31680
rect 25130 31628 25136 31680
rect 25188 31628 25194 31680
rect 27341 31671 27399 31677
rect 27341 31637 27353 31671
rect 27387 31668 27399 31671
rect 28077 31671 28135 31677
rect 28077 31668 28089 31671
rect 27387 31640 28089 31668
rect 27387 31637 27399 31640
rect 27341 31631 27399 31637
rect 28077 31637 28089 31640
rect 28123 31668 28135 31671
rect 28442 31668 28448 31680
rect 28123 31640 28448 31668
rect 28123 31637 28135 31640
rect 28077 31631 28135 31637
rect 28442 31628 28448 31640
rect 28500 31628 28506 31680
rect 28534 31628 28540 31680
rect 28592 31628 28598 31680
rect 29730 31628 29736 31680
rect 29788 31628 29794 31680
rect 35253 31671 35311 31677
rect 35253 31637 35265 31671
rect 35299 31668 35311 31671
rect 35342 31668 35348 31680
rect 35299 31640 35348 31668
rect 35299 31637 35311 31640
rect 35253 31631 35311 31637
rect 35342 31628 35348 31640
rect 35400 31628 35406 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 9953 31467 10011 31473
rect 9953 31464 9965 31467
rect 9732 31436 9965 31464
rect 9732 31424 9738 31436
rect 9953 31433 9965 31436
rect 9999 31433 10011 31467
rect 9953 31427 10011 31433
rect 13262 31424 13268 31476
rect 13320 31464 13326 31476
rect 13357 31467 13415 31473
rect 13357 31464 13369 31467
rect 13320 31436 13369 31464
rect 13320 31424 13326 31436
rect 13357 31433 13369 31436
rect 13403 31433 13415 31467
rect 13357 31427 13415 31433
rect 16114 31424 16120 31476
rect 16172 31464 16178 31476
rect 19334 31464 19340 31476
rect 16172 31436 19340 31464
rect 16172 31424 16178 31436
rect 13449 31399 13507 31405
rect 13449 31365 13461 31399
rect 13495 31396 13507 31399
rect 14734 31396 14740 31408
rect 13495 31368 14740 31396
rect 13495 31365 13507 31368
rect 13449 31359 13507 31365
rect 14734 31356 14740 31368
rect 14792 31356 14798 31408
rect 9861 31331 9919 31337
rect 9861 31297 9873 31331
rect 9907 31328 9919 31331
rect 11054 31328 11060 31340
rect 9907 31300 11060 31328
rect 9907 31297 9919 31300
rect 9861 31291 9919 31297
rect 11054 31288 11060 31300
rect 11112 31288 11118 31340
rect 14090 31337 14096 31340
rect 14084 31291 14096 31337
rect 14090 31288 14096 31291
rect 14148 31288 14154 31340
rect 18506 31337 18512 31340
rect 18500 31291 18512 31337
rect 18564 31328 18570 31340
rect 18564 31300 18600 31328
rect 18506 31288 18512 31291
rect 18564 31288 18570 31300
rect 9401 31263 9459 31269
rect 9401 31229 9413 31263
rect 9447 31260 9459 31263
rect 9447 31232 9536 31260
rect 9447 31229 9459 31232
rect 9401 31223 9459 31229
rect 9508 31201 9536 31232
rect 10042 31220 10048 31272
rect 10100 31220 10106 31272
rect 10870 31220 10876 31272
rect 10928 31220 10934 31272
rect 11514 31220 11520 31272
rect 11572 31220 11578 31272
rect 12345 31263 12403 31269
rect 12345 31229 12357 31263
rect 12391 31229 12403 31263
rect 12345 31223 12403 31229
rect 9493 31195 9551 31201
rect 9493 31161 9505 31195
rect 9539 31161 9551 31195
rect 12360 31192 12388 31223
rect 13630 31220 13636 31272
rect 13688 31220 13694 31272
rect 13722 31220 13728 31272
rect 13780 31260 13786 31272
rect 13817 31263 13875 31269
rect 13817 31260 13829 31263
rect 13780 31232 13829 31260
rect 13780 31220 13786 31232
rect 13817 31229 13829 31232
rect 13863 31229 13875 31263
rect 15838 31260 15844 31272
rect 13817 31223 13875 31229
rect 15212 31232 15844 31260
rect 15212 31201 15240 31232
rect 15838 31220 15844 31232
rect 15896 31220 15902 31272
rect 18230 31220 18236 31272
rect 18288 31220 18294 31272
rect 19260 31260 19288 31436
rect 19334 31424 19340 31436
rect 19392 31424 19398 31476
rect 20073 31467 20131 31473
rect 20073 31433 20085 31467
rect 20119 31464 20131 31467
rect 20346 31464 20352 31476
rect 20119 31436 20352 31464
rect 20119 31433 20131 31436
rect 20073 31427 20131 31433
rect 20346 31424 20352 31436
rect 20404 31424 20410 31476
rect 23569 31467 23627 31473
rect 23569 31433 23581 31467
rect 23615 31464 23627 31467
rect 23842 31464 23848 31476
rect 23615 31436 23848 31464
rect 23615 31433 23627 31436
rect 23569 31427 23627 31433
rect 23842 31424 23848 31436
rect 23900 31464 23906 31476
rect 23900 31436 25728 31464
rect 23900 31424 23906 31436
rect 23928 31399 23986 31405
rect 23928 31365 23940 31399
rect 23974 31396 23986 31399
rect 25130 31396 25136 31408
rect 23974 31368 25136 31396
rect 23974 31365 23986 31368
rect 23928 31359 23986 31365
rect 25130 31356 25136 31368
rect 25188 31356 25194 31408
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22445 31331 22503 31337
rect 22445 31328 22457 31331
rect 22336 31300 22457 31328
rect 22336 31288 22342 31300
rect 22445 31297 22457 31300
rect 22491 31297 22503 31331
rect 22445 31291 22503 31297
rect 24762 31288 24768 31340
rect 24820 31328 24826 31340
rect 25700 31337 25728 31436
rect 28074 31424 28080 31476
rect 28132 31464 28138 31476
rect 28353 31467 28411 31473
rect 28353 31464 28365 31467
rect 28132 31436 28365 31464
rect 28132 31424 28138 31436
rect 28353 31433 28365 31436
rect 28399 31464 28411 31467
rect 28810 31464 28816 31476
rect 28399 31436 28816 31464
rect 28399 31433 28411 31436
rect 28353 31427 28411 31433
rect 28810 31424 28816 31436
rect 28868 31424 28874 31476
rect 29178 31424 29184 31476
rect 29236 31424 29242 31476
rect 29270 31424 29276 31476
rect 29328 31424 29334 31476
rect 27240 31399 27298 31405
rect 25884 31368 27200 31396
rect 25685 31331 25743 31337
rect 24820 31300 25452 31328
rect 24820 31288 24826 31300
rect 19797 31263 19855 31269
rect 19797 31260 19809 31263
rect 19260 31232 19809 31260
rect 19797 31229 19809 31232
rect 19843 31229 19855 31263
rect 19797 31223 19855 31229
rect 19978 31220 19984 31272
rect 20036 31220 20042 31272
rect 21085 31263 21143 31269
rect 21085 31260 21097 31263
rect 20456 31232 21097 31260
rect 20456 31201 20484 31232
rect 21085 31229 21097 31232
rect 21131 31229 21143 31263
rect 22189 31263 22247 31269
rect 22189 31260 22201 31263
rect 21085 31223 21143 31229
rect 22066 31232 22201 31260
rect 12989 31195 13047 31201
rect 12989 31192 13001 31195
rect 12360 31164 13001 31192
rect 9493 31155 9551 31161
rect 12989 31161 13001 31164
rect 13035 31161 13047 31195
rect 12989 31155 13047 31161
rect 15197 31195 15255 31201
rect 15197 31161 15209 31195
rect 15243 31161 15255 31195
rect 15197 31155 15255 31161
rect 20441 31195 20499 31201
rect 20441 31161 20453 31195
rect 20487 31161 20499 31195
rect 20441 31155 20499 31161
rect 8754 31084 8760 31136
rect 8812 31084 8818 31136
rect 10318 31084 10324 31136
rect 10376 31084 10382 31136
rect 11330 31084 11336 31136
rect 11388 31084 11394 31136
rect 12158 31084 12164 31136
rect 12216 31084 12222 31136
rect 12894 31084 12900 31136
rect 12952 31084 12958 31136
rect 15286 31084 15292 31136
rect 15344 31084 15350 31136
rect 19150 31084 19156 31136
rect 19208 31124 19214 31136
rect 19610 31124 19616 31136
rect 19208 31096 19616 31124
rect 19208 31084 19214 31096
rect 19610 31084 19616 31096
rect 19668 31084 19674 31136
rect 20530 31084 20536 31136
rect 20588 31084 20594 31136
rect 21910 31084 21916 31136
rect 21968 31124 21974 31136
rect 22066 31124 22094 31232
rect 22189 31229 22201 31232
rect 22235 31229 22247 31263
rect 23661 31263 23719 31269
rect 23661 31260 23673 31263
rect 22189 31223 22247 31229
rect 23492 31232 23673 31260
rect 23492 31192 23520 31232
rect 23661 31229 23673 31232
rect 23707 31229 23719 31263
rect 23661 31223 23719 31229
rect 24670 31220 24676 31272
rect 24728 31260 24734 31272
rect 25133 31263 25191 31269
rect 25133 31260 25145 31263
rect 24728 31232 25145 31260
rect 24728 31220 24734 31232
rect 25133 31229 25145 31232
rect 25179 31229 25191 31263
rect 25424 31260 25452 31300
rect 25685 31297 25697 31331
rect 25731 31297 25743 31331
rect 25685 31291 25743 31297
rect 25884 31260 25912 31368
rect 26142 31288 26148 31340
rect 26200 31328 26206 31340
rect 26973 31331 27031 31337
rect 26973 31328 26985 31331
rect 26200 31300 26985 31328
rect 26200 31288 26206 31300
rect 26973 31297 26985 31300
rect 27019 31297 27031 31331
rect 27172 31328 27200 31368
rect 27240 31365 27252 31399
rect 27286 31396 27298 31399
rect 27522 31396 27528 31408
rect 27286 31368 27528 31396
rect 27286 31365 27298 31368
rect 27240 31359 27298 31365
rect 27522 31356 27528 31368
rect 27580 31356 27586 31408
rect 28721 31399 28779 31405
rect 28721 31365 28733 31399
rect 28767 31396 28779 31399
rect 30009 31399 30067 31405
rect 30009 31396 30021 31399
rect 28767 31368 30021 31396
rect 28767 31365 28779 31368
rect 28721 31359 28779 31365
rect 30009 31365 30021 31368
rect 30055 31365 30067 31399
rect 30009 31359 30067 31365
rect 31849 31399 31907 31405
rect 31849 31365 31861 31399
rect 31895 31396 31907 31399
rect 33318 31396 33324 31408
rect 31895 31368 33324 31396
rect 31895 31365 31907 31368
rect 31849 31359 31907 31365
rect 33318 31356 33324 31368
rect 33376 31356 33382 31408
rect 35428 31399 35486 31405
rect 35428 31365 35440 31399
rect 35474 31396 35486 31399
rect 36354 31396 36360 31408
rect 35474 31368 36360 31396
rect 35474 31365 35486 31368
rect 35428 31359 35486 31365
rect 36354 31356 36360 31368
rect 36412 31356 36418 31408
rect 27172 31300 28028 31328
rect 26973 31291 27031 31297
rect 25424 31232 25912 31260
rect 26421 31263 26479 31269
rect 25133 31223 25191 31229
rect 26421 31229 26433 31263
rect 26467 31229 26479 31263
rect 28000 31260 28028 31300
rect 28442 31288 28448 31340
rect 28500 31328 28506 31340
rect 28813 31331 28871 31337
rect 28813 31328 28825 31331
rect 28500 31300 28825 31328
rect 28500 31288 28506 31300
rect 28813 31297 28825 31300
rect 28859 31328 28871 31331
rect 29454 31328 29460 31340
rect 28859 31300 29460 31328
rect 28859 31297 28871 31300
rect 28813 31291 28871 31297
rect 29454 31288 29460 31300
rect 29512 31288 29518 31340
rect 32392 31331 32450 31337
rect 32392 31297 32404 31331
rect 32438 31328 32450 31331
rect 33597 31331 33655 31337
rect 33597 31328 33609 31331
rect 32438 31300 33609 31328
rect 32438 31297 32450 31300
rect 32392 31291 32450 31297
rect 33597 31297 33609 31300
rect 33643 31297 33655 31331
rect 33597 31291 33655 31297
rect 28537 31263 28595 31269
rect 28537 31260 28549 31263
rect 28000 31232 28549 31260
rect 26421 31223 26479 31229
rect 28537 31229 28549 31232
rect 28583 31229 28595 31263
rect 28537 31223 28595 31229
rect 23492 31164 23704 31192
rect 23492 31124 23520 31164
rect 21968 31096 23520 31124
rect 23676 31124 23704 31164
rect 24854 31152 24860 31204
rect 24912 31192 24918 31204
rect 25041 31195 25099 31201
rect 25041 31192 25053 31195
rect 24912 31164 25053 31192
rect 24912 31152 24918 31164
rect 25041 31161 25053 31164
rect 25087 31192 25099 31195
rect 26436 31192 26464 31223
rect 25087 31164 26464 31192
rect 25087 31161 25099 31164
rect 25041 31155 25099 31161
rect 24946 31124 24952 31136
rect 23676 31096 24952 31124
rect 21968 31084 21974 31096
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 25866 31084 25872 31136
rect 25924 31084 25930 31136
rect 28552 31124 28580 31223
rect 28626 31220 28632 31272
rect 28684 31260 28690 31272
rect 29825 31263 29883 31269
rect 29825 31260 29837 31263
rect 28684 31232 29837 31260
rect 28684 31220 28690 31232
rect 29825 31229 29837 31232
rect 29871 31229 29883 31263
rect 29825 31223 29883 31229
rect 29914 31220 29920 31272
rect 29972 31260 29978 31272
rect 30561 31263 30619 31269
rect 30561 31260 30573 31263
rect 29972 31232 30573 31260
rect 29972 31220 29978 31232
rect 30561 31229 30573 31232
rect 30607 31229 30619 31263
rect 30561 31223 30619 31229
rect 32125 31263 32183 31269
rect 32125 31229 32137 31263
rect 32171 31229 32183 31263
rect 32125 31223 32183 31229
rect 29730 31124 29736 31136
rect 28552 31096 29736 31124
rect 29730 31084 29736 31096
rect 29788 31124 29794 31136
rect 31110 31124 31116 31136
rect 29788 31096 31116 31124
rect 29788 31084 29794 31096
rect 31110 31084 31116 31096
rect 31168 31084 31174 31136
rect 32140 31124 32168 31223
rect 34146 31220 34152 31272
rect 34204 31220 34210 31272
rect 34885 31263 34943 31269
rect 34885 31229 34897 31263
rect 34931 31229 34943 31263
rect 34885 31223 34943 31229
rect 35161 31263 35219 31269
rect 35161 31229 35173 31263
rect 35207 31229 35219 31263
rect 35161 31223 35219 31229
rect 33505 31195 33563 31201
rect 33505 31161 33517 31195
rect 33551 31192 33563 31195
rect 33778 31192 33784 31204
rect 33551 31164 33784 31192
rect 33551 31161 33563 31164
rect 33505 31155 33563 31161
rect 33778 31152 33784 31164
rect 33836 31192 33842 31204
rect 34900 31192 34928 31223
rect 33836 31164 34928 31192
rect 33836 31152 33842 31164
rect 32306 31124 32312 31136
rect 32140 31096 32312 31124
rect 32306 31084 32312 31096
rect 32364 31084 32370 31136
rect 34330 31084 34336 31136
rect 34388 31084 34394 31136
rect 35176 31124 35204 31223
rect 36814 31220 36820 31272
rect 36872 31260 36878 31272
rect 37277 31263 37335 31269
rect 37277 31260 37289 31263
rect 36872 31232 37289 31260
rect 36872 31220 36878 31232
rect 37277 31229 37289 31232
rect 37323 31229 37335 31263
rect 37277 31223 37335 31229
rect 35802 31124 35808 31136
rect 35176 31096 35808 31124
rect 35802 31084 35808 31096
rect 35860 31084 35866 31136
rect 36170 31084 36176 31136
rect 36228 31124 36234 31136
rect 36538 31124 36544 31136
rect 36228 31096 36544 31124
rect 36228 31084 36234 31096
rect 36538 31084 36544 31096
rect 36596 31084 36602 31136
rect 37918 31084 37924 31136
rect 37976 31084 37982 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 10781 30923 10839 30929
rect 10781 30889 10793 30923
rect 10827 30920 10839 30923
rect 10870 30920 10876 30932
rect 10827 30892 10876 30920
rect 10827 30889 10839 30892
rect 10781 30883 10839 30889
rect 10870 30880 10876 30892
rect 10928 30880 10934 30932
rect 11514 30880 11520 30932
rect 11572 30880 11578 30932
rect 13909 30923 13967 30929
rect 13909 30889 13921 30923
rect 13955 30920 13967 30923
rect 15010 30920 15016 30932
rect 13955 30892 15016 30920
rect 13955 30889 13967 30892
rect 13909 30883 13967 30889
rect 15010 30880 15016 30892
rect 15068 30880 15074 30932
rect 15562 30880 15568 30932
rect 15620 30880 15626 30932
rect 19242 30880 19248 30932
rect 19300 30880 19306 30932
rect 23293 30923 23351 30929
rect 23293 30889 23305 30923
rect 23339 30920 23351 30923
rect 23750 30920 23756 30932
rect 23339 30892 23756 30920
rect 23339 30889 23351 30892
rect 23293 30883 23351 30889
rect 23750 30880 23756 30892
rect 23808 30920 23814 30932
rect 23934 30920 23940 30932
rect 23808 30892 23940 30920
rect 23808 30880 23814 30892
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 24397 30923 24455 30929
rect 24397 30889 24409 30923
rect 24443 30920 24455 30923
rect 24578 30920 24584 30932
rect 24443 30892 24584 30920
rect 24443 30889 24455 30892
rect 24397 30883 24455 30889
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 26602 30920 26608 30932
rect 24688 30892 26608 30920
rect 10689 30855 10747 30861
rect 10689 30821 10701 30855
rect 10735 30852 10747 30855
rect 11532 30852 11560 30880
rect 10735 30824 11560 30852
rect 15473 30855 15531 30861
rect 10735 30821 10747 30824
rect 10689 30815 10747 30821
rect 15473 30821 15485 30855
rect 15519 30852 15531 30855
rect 15746 30852 15752 30864
rect 15519 30824 15752 30852
rect 15519 30821 15531 30824
rect 15473 30815 15531 30821
rect 15746 30812 15752 30824
rect 15804 30852 15810 30864
rect 15804 30824 16988 30852
rect 15804 30812 15810 30824
rect 11330 30744 11336 30796
rect 11388 30784 11394 30796
rect 11388 30756 12434 30784
rect 11388 30744 11394 30756
rect 9306 30676 9312 30728
rect 9364 30676 9370 30728
rect 9576 30719 9634 30725
rect 9576 30685 9588 30719
rect 9622 30716 9634 30719
rect 10594 30716 10600 30728
rect 9622 30688 10600 30716
rect 9622 30685 9634 30688
rect 9576 30679 9634 30685
rect 10594 30676 10600 30688
rect 10652 30676 10658 30728
rect 11422 30676 11428 30728
rect 11480 30716 11486 30728
rect 12161 30719 12219 30725
rect 12161 30716 12173 30719
rect 11480 30688 12173 30716
rect 11480 30676 11486 30688
rect 12161 30685 12173 30688
rect 12207 30685 12219 30719
rect 12161 30679 12219 30685
rect 11149 30651 11207 30657
rect 11149 30617 11161 30651
rect 11195 30648 11207 30651
rect 11609 30651 11667 30657
rect 11609 30648 11621 30651
rect 11195 30620 11621 30648
rect 11195 30617 11207 30620
rect 11149 30611 11207 30617
rect 11609 30617 11621 30620
rect 11655 30617 11667 30651
rect 11609 30611 11667 30617
rect 9217 30583 9275 30589
rect 9217 30549 9229 30583
rect 9263 30580 9275 30583
rect 10134 30580 10140 30592
rect 9263 30552 10140 30580
rect 9263 30549 9275 30552
rect 9217 30543 9275 30549
rect 10134 30540 10140 30552
rect 10192 30540 10198 30592
rect 11054 30540 11060 30592
rect 11112 30580 11118 30592
rect 11241 30583 11299 30589
rect 11241 30580 11253 30583
rect 11112 30552 11253 30580
rect 11112 30540 11118 30552
rect 11241 30549 11253 30552
rect 11287 30580 11299 30583
rect 11698 30580 11704 30592
rect 11287 30552 11704 30580
rect 11287 30549 11299 30552
rect 11241 30543 11299 30549
rect 11698 30540 11704 30552
rect 11756 30540 11762 30592
rect 12406 30580 12434 30756
rect 13722 30744 13728 30796
rect 13780 30784 13786 30796
rect 14093 30787 14151 30793
rect 14093 30784 14105 30787
rect 13780 30756 14105 30784
rect 13780 30744 13786 30756
rect 14093 30753 14105 30756
rect 14139 30753 14151 30787
rect 14093 30747 14151 30753
rect 15764 30756 16068 30784
rect 12529 30719 12587 30725
rect 12529 30685 12541 30719
rect 12575 30716 12587 30719
rect 12618 30716 12624 30728
rect 12575 30688 12624 30716
rect 12575 30685 12587 30688
rect 12529 30679 12587 30685
rect 12618 30676 12624 30688
rect 12676 30716 12682 30728
rect 13740 30716 13768 30744
rect 12676 30688 13768 30716
rect 14360 30719 14418 30725
rect 12676 30676 12682 30688
rect 14360 30685 14372 30719
rect 14406 30716 14418 30719
rect 14642 30716 14648 30728
rect 14406 30688 14648 30716
rect 14406 30685 14418 30688
rect 14360 30679 14418 30685
rect 14642 30676 14648 30688
rect 14700 30676 14706 30728
rect 12796 30651 12854 30657
rect 12796 30617 12808 30651
rect 12842 30648 12854 30651
rect 13446 30648 13452 30660
rect 12842 30620 13452 30648
rect 12842 30617 12854 30620
rect 12796 30611 12854 30617
rect 13446 30608 13452 30620
rect 13504 30608 13510 30660
rect 14734 30608 14740 30660
rect 14792 30648 14798 30660
rect 15764 30648 15792 30756
rect 16040 30725 16068 30756
rect 16114 30744 16120 30796
rect 16172 30744 16178 30796
rect 16960 30793 16988 30824
rect 16945 30787 17003 30793
rect 16945 30753 16957 30787
rect 16991 30753 17003 30787
rect 16945 30747 17003 30753
rect 19610 30744 19616 30796
rect 19668 30744 19674 30796
rect 20625 30787 20683 30793
rect 20625 30753 20637 30787
rect 20671 30784 20683 30787
rect 21910 30784 21916 30796
rect 20671 30756 21916 30784
rect 20671 30753 20683 30756
rect 20625 30747 20683 30753
rect 21910 30744 21916 30756
rect 21968 30744 21974 30796
rect 23569 30787 23627 30793
rect 23569 30753 23581 30787
rect 23615 30784 23627 30787
rect 24688 30784 24716 30892
rect 26602 30880 26608 30892
rect 26660 30880 26666 30932
rect 27617 30923 27675 30929
rect 27617 30889 27629 30923
rect 27663 30920 27675 30923
rect 27982 30920 27988 30932
rect 27663 30892 27988 30920
rect 27663 30889 27675 30892
rect 27617 30883 27675 30889
rect 27982 30880 27988 30892
rect 28040 30920 28046 30932
rect 28626 30920 28632 30932
rect 28040 30892 28632 30920
rect 28040 30880 28046 30892
rect 28626 30880 28632 30892
rect 28684 30880 28690 30932
rect 28994 30880 29000 30932
rect 29052 30920 29058 30932
rect 29089 30923 29147 30929
rect 29089 30920 29101 30923
rect 29052 30892 29101 30920
rect 29052 30880 29058 30892
rect 29089 30889 29101 30892
rect 29135 30920 29147 30923
rect 29914 30920 29920 30932
rect 29135 30892 29920 30920
rect 29135 30889 29147 30892
rect 29089 30883 29147 30889
rect 29914 30880 29920 30892
rect 29972 30880 29978 30932
rect 33134 30920 33140 30932
rect 30576 30892 33140 30920
rect 23615 30756 24716 30784
rect 23615 30753 23627 30756
rect 23569 30747 23627 30753
rect 16025 30719 16083 30725
rect 16025 30685 16037 30719
rect 16071 30685 16083 30719
rect 16025 30679 16083 30685
rect 17218 30676 17224 30728
rect 17276 30716 17282 30728
rect 17681 30719 17739 30725
rect 17681 30716 17693 30719
rect 17276 30688 17693 30716
rect 17276 30676 17282 30688
rect 17681 30685 17693 30688
rect 17727 30716 17739 30719
rect 18230 30716 18236 30728
rect 17727 30688 18236 30716
rect 17727 30685 17739 30688
rect 17681 30679 17739 30685
rect 18230 30676 18236 30688
rect 18288 30676 18294 30728
rect 17954 30657 17960 30660
rect 14792 30620 15792 30648
rect 15933 30651 15991 30657
rect 14792 30608 14798 30620
rect 15933 30617 15945 30651
rect 15979 30648 15991 30651
rect 16393 30651 16451 30657
rect 16393 30648 16405 30651
rect 15979 30620 16405 30648
rect 15979 30617 15991 30620
rect 15933 30611 15991 30617
rect 16393 30617 16405 30620
rect 16439 30617 16451 30651
rect 16393 30611 16451 30617
rect 17948 30611 17960 30657
rect 17954 30608 17960 30611
rect 18012 30608 18018 30660
rect 19628 30648 19656 30744
rect 20369 30719 20427 30725
rect 20369 30685 20381 30719
rect 20415 30716 20427 30719
rect 20530 30716 20536 30728
rect 20415 30688 20536 30716
rect 20415 30685 20427 30688
rect 20369 30679 20427 30685
rect 20530 30676 20536 30688
rect 20588 30676 20594 30728
rect 21269 30719 21327 30725
rect 21269 30685 21281 30719
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 21821 30719 21879 30725
rect 21821 30685 21833 30719
rect 21867 30716 21879 30719
rect 22462 30716 22468 30728
rect 21867 30688 22468 30716
rect 21867 30685 21879 30688
rect 21821 30679 21879 30685
rect 21284 30648 21312 30679
rect 22462 30676 22468 30688
rect 22520 30716 22526 30728
rect 23584 30716 23612 30747
rect 29454 30744 29460 30796
rect 29512 30784 29518 30796
rect 30009 30787 30067 30793
rect 30009 30784 30021 30787
rect 29512 30756 30021 30784
rect 29512 30744 29518 30756
rect 30009 30753 30021 30756
rect 30055 30753 30067 30787
rect 30009 30747 30067 30753
rect 30101 30787 30159 30793
rect 30101 30753 30113 30787
rect 30147 30784 30159 30787
rect 30147 30756 30181 30784
rect 30147 30753 30159 30756
rect 30101 30747 30159 30753
rect 22520 30688 23612 30716
rect 23753 30719 23811 30725
rect 22520 30676 22526 30688
rect 23753 30685 23765 30719
rect 23799 30716 23811 30719
rect 24394 30716 24400 30728
rect 23799 30688 24400 30716
rect 23799 30685 23811 30688
rect 23753 30679 23811 30685
rect 24394 30676 24400 30688
rect 24452 30676 24458 30728
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 25777 30719 25835 30725
rect 25777 30716 25789 30719
rect 25004 30688 25789 30716
rect 25004 30676 25010 30688
rect 25777 30685 25789 30688
rect 25823 30716 25835 30719
rect 26142 30716 26148 30728
rect 25823 30688 26148 30716
rect 25823 30685 25835 30688
rect 25777 30679 25835 30685
rect 26142 30676 26148 30688
rect 26200 30716 26206 30728
rect 26237 30719 26295 30725
rect 26237 30716 26249 30719
rect 26200 30688 26249 30716
rect 26200 30676 26206 30688
rect 26237 30685 26249 30688
rect 26283 30716 26295 30719
rect 27709 30719 27767 30725
rect 27709 30716 27721 30719
rect 26283 30688 27721 30716
rect 26283 30685 26295 30688
rect 26237 30679 26295 30685
rect 27709 30685 27721 30688
rect 27755 30685 27767 30719
rect 27709 30679 27767 30685
rect 27976 30719 28034 30725
rect 27976 30685 27988 30719
rect 28022 30716 28034 30719
rect 28534 30716 28540 30728
rect 28022 30688 28540 30716
rect 28022 30685 28034 30688
rect 27976 30679 28034 30685
rect 28534 30676 28540 30688
rect 28592 30676 28598 30728
rect 30116 30716 30144 30747
rect 30576 30725 30604 30892
rect 33134 30880 33140 30892
rect 33192 30880 33198 30932
rect 36357 30923 36415 30929
rect 36357 30889 36369 30923
rect 36403 30920 36415 30923
rect 36446 30920 36452 30932
rect 36403 30892 36452 30920
rect 36403 30889 36415 30892
rect 36357 30883 36415 30889
rect 36446 30880 36452 30892
rect 36504 30880 36510 30932
rect 37918 30880 37924 30932
rect 37976 30880 37982 30932
rect 33781 30855 33839 30861
rect 33781 30821 33793 30855
rect 33827 30821 33839 30855
rect 33781 30815 33839 30821
rect 33796 30784 33824 30815
rect 33962 30784 33968 30796
rect 33796 30756 33968 30784
rect 33962 30744 33968 30756
rect 34020 30784 34026 30796
rect 34425 30787 34483 30793
rect 34425 30784 34437 30787
rect 34020 30756 34437 30784
rect 34020 30744 34026 30756
rect 34425 30753 34437 30756
rect 34471 30753 34483 30787
rect 34425 30747 34483 30753
rect 30561 30719 30619 30725
rect 30561 30716 30573 30719
rect 29380 30688 30573 30716
rect 18064 30620 19472 30648
rect 19628 30620 21312 30648
rect 22180 30651 22238 30657
rect 16114 30580 16120 30592
rect 12406 30552 16120 30580
rect 16114 30540 16120 30552
rect 16172 30540 16178 30592
rect 16574 30540 16580 30592
rect 16632 30580 16638 30592
rect 17589 30583 17647 30589
rect 17589 30580 17601 30583
rect 16632 30552 17601 30580
rect 16632 30540 16638 30552
rect 17589 30549 17601 30552
rect 17635 30580 17647 30583
rect 18064 30580 18092 30620
rect 19444 30592 19472 30620
rect 22180 30617 22192 30651
rect 22226 30648 22238 30651
rect 23566 30648 23572 30660
rect 22226 30620 23572 30648
rect 22226 30617 22238 30620
rect 22180 30611 22238 30617
rect 23566 30608 23572 30620
rect 23624 30608 23630 30660
rect 25406 30608 25412 30660
rect 25464 30648 25470 30660
rect 25510 30651 25568 30657
rect 25510 30648 25522 30651
rect 25464 30620 25522 30648
rect 25464 30608 25470 30620
rect 25510 30617 25522 30620
rect 25556 30617 25568 30651
rect 25510 30611 25568 30617
rect 26326 30608 26332 30660
rect 26384 30648 26390 30660
rect 26482 30651 26540 30657
rect 26482 30648 26494 30651
rect 26384 30620 26494 30648
rect 26384 30608 26390 30620
rect 26482 30617 26494 30620
rect 26528 30617 26540 30651
rect 26482 30611 26540 30617
rect 29380 30592 29408 30688
rect 30561 30685 30573 30688
rect 30607 30685 30619 30719
rect 30561 30679 30619 30685
rect 30929 30719 30987 30725
rect 30929 30685 30941 30719
rect 30975 30716 30987 30719
rect 31018 30716 31024 30728
rect 30975 30688 31024 30716
rect 30975 30685 30987 30688
rect 30929 30679 30987 30685
rect 31018 30676 31024 30688
rect 31076 30676 31082 30728
rect 32306 30676 32312 30728
rect 32364 30716 32370 30728
rect 32401 30719 32459 30725
rect 32401 30716 32413 30719
rect 32364 30688 32413 30716
rect 32364 30676 32370 30688
rect 32401 30685 32413 30688
rect 32447 30685 32459 30719
rect 32401 30679 32459 30685
rect 34977 30719 35035 30725
rect 34977 30685 34989 30719
rect 35023 30716 35035 30719
rect 35802 30716 35808 30728
rect 35023 30688 35808 30716
rect 35023 30685 35035 30688
rect 34977 30679 35035 30685
rect 35802 30676 35808 30688
rect 35860 30716 35866 30728
rect 37829 30719 37887 30725
rect 37829 30716 37841 30719
rect 35860 30688 37841 30716
rect 35860 30676 35866 30688
rect 37829 30685 37841 30688
rect 37875 30685 37887 30719
rect 37829 30679 37887 30685
rect 29917 30651 29975 30657
rect 29917 30617 29929 30651
rect 29963 30648 29975 30651
rect 30466 30648 30472 30660
rect 29963 30620 30472 30648
rect 29963 30617 29975 30620
rect 29917 30611 29975 30617
rect 30466 30608 30472 30620
rect 30524 30608 30530 30660
rect 31196 30651 31254 30657
rect 31196 30617 31208 30651
rect 31242 30648 31254 30651
rect 31294 30648 31300 30660
rect 31242 30620 31300 30648
rect 31242 30617 31254 30620
rect 31196 30611 31254 30617
rect 31294 30608 31300 30620
rect 31352 30608 31358 30660
rect 32668 30651 32726 30657
rect 32668 30617 32680 30651
rect 32714 30648 32726 30651
rect 33226 30648 33232 30660
rect 32714 30620 33232 30648
rect 32714 30617 32726 30620
rect 32668 30611 32726 30617
rect 33226 30608 33232 30620
rect 33284 30608 33290 30660
rect 35244 30651 35302 30657
rect 35244 30617 35256 30651
rect 35290 30648 35302 30651
rect 35342 30648 35348 30660
rect 35290 30620 35348 30648
rect 35290 30617 35302 30620
rect 35244 30611 35302 30617
rect 35342 30608 35348 30620
rect 35400 30608 35406 30660
rect 36906 30608 36912 30660
rect 36964 30608 36970 30660
rect 37584 30651 37642 30657
rect 37584 30617 37596 30651
rect 37630 30648 37642 30651
rect 37936 30648 37964 30880
rect 37630 30620 37964 30648
rect 37630 30617 37642 30620
rect 37584 30611 37642 30617
rect 17635 30552 18092 30580
rect 19061 30583 19119 30589
rect 17635 30549 17647 30552
rect 17589 30543 17647 30549
rect 19061 30549 19073 30583
rect 19107 30580 19119 30583
rect 19334 30580 19340 30592
rect 19107 30552 19340 30580
rect 19107 30549 19119 30552
rect 19061 30543 19119 30549
rect 19334 30540 19340 30552
rect 19392 30540 19398 30592
rect 19426 30540 19432 30592
rect 19484 30540 19490 30592
rect 20714 30540 20720 30592
rect 20772 30540 20778 30592
rect 23658 30540 23664 30592
rect 23716 30540 23722 30592
rect 24118 30540 24124 30592
rect 24176 30540 24182 30592
rect 29362 30540 29368 30592
rect 29420 30540 29426 30592
rect 29546 30540 29552 30592
rect 29604 30540 29610 30592
rect 32309 30583 32367 30589
rect 32309 30549 32321 30583
rect 32355 30580 32367 30583
rect 33042 30580 33048 30592
rect 32355 30552 33048 30580
rect 32355 30549 32367 30552
rect 32309 30543 32367 30549
rect 33042 30540 33048 30552
rect 33100 30540 33106 30592
rect 33870 30540 33876 30592
rect 33928 30540 33934 30592
rect 36449 30583 36507 30589
rect 36449 30549 36461 30583
rect 36495 30580 36507 30583
rect 36924 30580 36952 30608
rect 36495 30552 36952 30580
rect 36495 30549 36507 30552
rect 36449 30543 36507 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 11422 30376 11428 30388
rect 11164 30348 11428 30376
rect 8288 30311 8346 30317
rect 8288 30277 8300 30311
rect 8334 30308 8346 30311
rect 8754 30308 8760 30320
rect 8334 30280 8760 30308
rect 8334 30277 8346 30280
rect 8288 30271 8346 30277
rect 8754 30268 8760 30280
rect 8812 30268 8818 30320
rect 11164 30252 11192 30348
rect 11422 30336 11428 30348
rect 11480 30336 11486 30388
rect 11977 30379 12035 30385
rect 11977 30345 11989 30379
rect 12023 30376 12035 30379
rect 12158 30376 12164 30388
rect 12023 30348 12164 30376
rect 12023 30345 12035 30348
rect 11977 30339 12035 30345
rect 12158 30336 12164 30348
rect 12216 30336 12222 30388
rect 13906 30336 13912 30388
rect 13964 30376 13970 30388
rect 14001 30379 14059 30385
rect 14001 30376 14013 30379
rect 13964 30348 14013 30376
rect 13964 30336 13970 30348
rect 14001 30345 14013 30348
rect 14047 30376 14059 30379
rect 14918 30376 14924 30388
rect 14047 30348 14924 30376
rect 14047 30345 14059 30348
rect 14001 30339 14059 30345
rect 14918 30336 14924 30348
rect 14976 30336 14982 30388
rect 16114 30336 16120 30388
rect 16172 30376 16178 30388
rect 16209 30379 16267 30385
rect 16209 30376 16221 30379
rect 16172 30348 16221 30376
rect 16172 30336 16178 30348
rect 16209 30345 16221 30348
rect 16255 30345 16267 30379
rect 19242 30376 19248 30388
rect 16209 30339 16267 30345
rect 18800 30348 19248 30376
rect 12894 30317 12900 30320
rect 12888 30308 12900 30317
rect 12855 30280 12900 30308
rect 12888 30271 12900 30280
rect 12894 30268 12900 30271
rect 12952 30268 12958 30320
rect 10410 30200 10416 30252
rect 10468 30200 10474 30252
rect 11146 30200 11152 30252
rect 11204 30200 11210 30252
rect 11333 30243 11391 30249
rect 11333 30209 11345 30243
rect 11379 30240 11391 30243
rect 11514 30240 11520 30252
rect 11379 30212 11520 30240
rect 11379 30209 11391 30212
rect 11333 30203 11391 30209
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 11606 30200 11612 30252
rect 11664 30240 11670 30252
rect 11885 30243 11943 30249
rect 11885 30240 11897 30243
rect 11664 30212 11897 30240
rect 11664 30200 11670 30212
rect 11885 30209 11897 30212
rect 11931 30209 11943 30243
rect 11885 30203 11943 30209
rect 12618 30200 12624 30252
rect 12676 30200 12682 30252
rect 14918 30249 14924 30252
rect 14896 30243 14924 30249
rect 14896 30209 14908 30243
rect 14896 30203 14924 30209
rect 14918 30200 14924 30203
rect 14976 30200 14982 30252
rect 15010 30200 15016 30252
rect 15068 30200 15074 30252
rect 15746 30200 15752 30252
rect 15804 30200 15810 30252
rect 15838 30200 15844 30252
rect 15896 30240 15902 30252
rect 15933 30243 15991 30249
rect 15933 30240 15945 30243
rect 15896 30212 15945 30240
rect 15896 30200 15902 30212
rect 15933 30209 15945 30212
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 17129 30243 17187 30249
rect 17129 30209 17141 30243
rect 17175 30240 17187 30243
rect 17218 30240 17224 30252
rect 17175 30212 17224 30240
rect 17175 30209 17187 30212
rect 17129 30203 17187 30209
rect 17218 30200 17224 30212
rect 17276 30200 17282 30252
rect 17402 30249 17408 30252
rect 17396 30203 17408 30249
rect 17402 30200 17408 30203
rect 17460 30200 17466 30252
rect 18800 30249 18828 30348
rect 19242 30336 19248 30348
rect 19300 30336 19306 30388
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 22189 30379 22247 30385
rect 19392 30348 20392 30376
rect 19392 30336 19398 30348
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 19794 30200 19800 30252
rect 19852 30200 19858 30252
rect 20364 30240 20392 30348
rect 22189 30345 22201 30379
rect 22235 30376 22247 30379
rect 22278 30376 22284 30388
rect 22235 30348 22284 30376
rect 22235 30345 22247 30348
rect 22189 30339 22247 30345
rect 22278 30336 22284 30348
rect 22336 30336 22342 30388
rect 24578 30336 24584 30388
rect 24636 30336 24642 30388
rect 24946 30336 24952 30388
rect 25004 30336 25010 30388
rect 30466 30336 30472 30388
rect 30524 30336 30530 30388
rect 31018 30336 31024 30388
rect 31076 30376 31082 30388
rect 32306 30376 32312 30388
rect 31076 30348 32312 30376
rect 31076 30336 31082 30348
rect 32306 30336 32312 30348
rect 32364 30336 32370 30388
rect 33318 30336 33324 30388
rect 33376 30376 33382 30388
rect 33594 30376 33600 30388
rect 33376 30348 33600 30376
rect 33376 30336 33382 30348
rect 33594 30336 33600 30348
rect 33652 30376 33658 30388
rect 34422 30376 34428 30388
rect 33652 30348 34428 30376
rect 33652 30336 33658 30348
rect 34422 30336 34428 30348
rect 34480 30336 34486 30388
rect 36906 30336 36912 30388
rect 36964 30336 36970 30388
rect 23750 30249 23756 30252
rect 21085 30243 21143 30249
rect 21085 30240 21097 30243
rect 20364 30212 21097 30240
rect 21085 30209 21097 30212
rect 21131 30209 21143 30243
rect 21085 30203 21143 30209
rect 23728 30243 23756 30249
rect 23728 30209 23740 30243
rect 23728 30203 23756 30209
rect 23750 30200 23756 30203
rect 23808 30200 23814 30252
rect 23842 30200 23848 30252
rect 23900 30200 23906 30252
rect 24596 30240 24624 30336
rect 24964 30308 24992 30336
rect 25041 30311 25099 30317
rect 25041 30308 25053 30311
rect 24964 30280 25053 30308
rect 25041 30277 25053 30280
rect 25087 30277 25099 30311
rect 31036 30308 31064 30336
rect 25041 30271 25099 30277
rect 30576 30280 31064 30308
rect 24765 30243 24823 30249
rect 24765 30240 24777 30243
rect 24596 30212 24777 30240
rect 24765 30209 24777 30212
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 24854 30200 24860 30252
rect 24912 30200 24918 30252
rect 26418 30200 26424 30252
rect 26476 30240 26482 30252
rect 26789 30243 26847 30249
rect 26789 30240 26801 30243
rect 26476 30212 26801 30240
rect 26476 30200 26482 30212
rect 26789 30209 26801 30212
rect 26835 30209 26847 30243
rect 26789 30203 26847 30209
rect 27798 30200 27804 30252
rect 27856 30200 27862 30252
rect 27982 30249 27988 30252
rect 27960 30243 27988 30249
rect 27960 30209 27972 30243
rect 27960 30203 27988 30209
rect 27982 30200 27988 30203
rect 28040 30200 28046 30252
rect 28074 30200 28080 30252
rect 28132 30200 28138 30252
rect 28810 30200 28816 30252
rect 28868 30240 28874 30252
rect 28868 30212 29132 30240
rect 28868 30200 28874 30212
rect 7834 30132 7840 30184
rect 7892 30172 7898 30184
rect 8021 30175 8079 30181
rect 8021 30172 8033 30175
rect 7892 30144 8033 30172
rect 7892 30132 7898 30144
rect 8021 30141 8033 30144
rect 8067 30141 8079 30175
rect 8021 30135 8079 30141
rect 10134 30132 10140 30184
rect 10192 30132 10198 30184
rect 10296 30175 10354 30181
rect 10296 30141 10308 30175
rect 10342 30172 10354 30175
rect 10594 30172 10600 30184
rect 10342 30144 10600 30172
rect 10342 30141 10354 30144
rect 10296 30135 10354 30141
rect 10594 30132 10600 30144
rect 10652 30132 10658 30184
rect 11238 30132 11244 30184
rect 11296 30132 11302 30184
rect 12161 30175 12219 30181
rect 12161 30141 12173 30175
rect 12207 30172 12219 30175
rect 12207 30144 12664 30172
rect 12207 30141 12219 30144
rect 12161 30135 12219 30141
rect 9401 30107 9459 30113
rect 9401 30073 9413 30107
rect 9447 30104 9459 30107
rect 10689 30107 10747 30113
rect 9447 30076 9812 30104
rect 9447 30073 9459 30076
rect 9401 30067 9459 30073
rect 9490 29996 9496 30048
rect 9548 29996 9554 30048
rect 9784 30036 9812 30076
rect 10689 30073 10701 30107
rect 10735 30104 10747 30107
rect 10778 30104 10784 30116
rect 10735 30076 10784 30104
rect 10735 30073 10747 30076
rect 10689 30067 10747 30073
rect 10778 30064 10784 30076
rect 10836 30064 10842 30116
rect 11256 30104 11284 30132
rect 11517 30107 11575 30113
rect 11517 30104 11529 30107
rect 11256 30076 11529 30104
rect 11517 30073 11529 30076
rect 11563 30073 11575 30107
rect 11517 30067 11575 30073
rect 10410 30036 10416 30048
rect 9784 30008 10416 30036
rect 10410 29996 10416 30008
rect 10468 29996 10474 30048
rect 12636 30036 12664 30144
rect 14550 30132 14556 30184
rect 14608 30172 14614 30184
rect 14727 30175 14785 30181
rect 14727 30172 14739 30175
rect 14608 30144 14739 30172
rect 14608 30132 14614 30144
rect 14727 30141 14739 30144
rect 14773 30141 14785 30175
rect 14727 30135 14785 30141
rect 18601 30175 18659 30181
rect 18601 30141 18613 30175
rect 18647 30172 18659 30175
rect 19150 30172 19156 30184
rect 18647 30144 19156 30172
rect 18647 30141 18659 30144
rect 18601 30135 18659 30141
rect 19150 30132 19156 30144
rect 19208 30132 19214 30184
rect 19334 30132 19340 30184
rect 19392 30172 19398 30184
rect 19521 30175 19579 30181
rect 19521 30172 19533 30175
rect 19392 30144 19533 30172
rect 19392 30132 19398 30144
rect 19521 30141 19533 30144
rect 19567 30141 19579 30175
rect 19521 30135 19579 30141
rect 19610 30132 19616 30184
rect 19668 30181 19674 30184
rect 19668 30175 19696 30181
rect 19684 30141 19696 30175
rect 19668 30135 19696 30141
rect 19668 30132 19674 30135
rect 22738 30132 22744 30184
rect 22796 30132 22802 30184
rect 23569 30175 23627 30181
rect 23569 30141 23581 30175
rect 23615 30172 23627 30175
rect 24581 30175 24639 30181
rect 23615 30144 24072 30172
rect 23615 30141 23627 30144
rect 23569 30135 23627 30141
rect 15194 30064 15200 30116
rect 15252 30104 15258 30116
rect 15289 30107 15347 30113
rect 15289 30104 15301 30107
rect 15252 30076 15301 30104
rect 15252 30064 15258 30076
rect 15289 30073 15301 30076
rect 15335 30104 15347 30107
rect 16945 30107 17003 30113
rect 16945 30104 16957 30107
rect 15335 30076 16957 30104
rect 15335 30073 15347 30076
rect 15289 30067 15347 30073
rect 16945 30073 16957 30076
rect 16991 30073 17003 30107
rect 19245 30107 19303 30113
rect 19245 30104 19257 30107
rect 16945 30067 17003 30073
rect 18064 30076 19257 30104
rect 12894 30036 12900 30048
rect 12636 30008 12900 30036
rect 12894 29996 12900 30008
rect 12952 29996 12958 30048
rect 14093 30039 14151 30045
rect 14093 30005 14105 30039
rect 14139 30036 14151 30039
rect 16022 30036 16028 30048
rect 14139 30008 16028 30036
rect 14139 30005 14151 30008
rect 14093 29999 14151 30005
rect 16022 29996 16028 30008
rect 16080 29996 16086 30048
rect 16960 30036 16988 30067
rect 18064 30036 18092 30076
rect 19245 30073 19257 30076
rect 19291 30073 19303 30107
rect 19245 30067 19303 30073
rect 20441 30107 20499 30113
rect 20441 30073 20453 30107
rect 20487 30104 20499 30107
rect 21082 30104 21088 30116
rect 20487 30076 21088 30104
rect 20487 30073 20499 30076
rect 20441 30067 20499 30073
rect 21082 30064 21088 30076
rect 21140 30064 21146 30116
rect 16960 30008 18092 30036
rect 18509 30039 18567 30045
rect 18509 30005 18521 30039
rect 18555 30036 18567 30039
rect 19610 30036 19616 30048
rect 18555 30008 19616 30036
rect 18555 30005 18567 30008
rect 18509 29999 18567 30005
rect 19610 29996 19616 30008
rect 19668 29996 19674 30048
rect 19702 29996 19708 30048
rect 19760 30036 19766 30048
rect 20533 30039 20591 30045
rect 20533 30036 20545 30039
rect 19760 30008 20545 30036
rect 19760 29996 19766 30008
rect 20533 30005 20545 30008
rect 20579 30005 20591 30039
rect 20533 29999 20591 30005
rect 22925 30039 22983 30045
rect 22925 30005 22937 30039
rect 22971 30036 22983 30039
rect 23842 30036 23848 30048
rect 22971 30008 23848 30036
rect 22971 30005 22983 30008
rect 22925 29999 22983 30005
rect 23842 29996 23848 30008
rect 23900 29996 23906 30048
rect 24044 30036 24072 30144
rect 24581 30141 24593 30175
rect 24627 30172 24639 30175
rect 24872 30172 24900 30200
rect 28353 30175 28411 30181
rect 28353 30172 28365 30175
rect 24627 30144 24900 30172
rect 26252 30144 28365 30172
rect 24627 30141 24639 30144
rect 24581 30135 24639 30141
rect 26252 30116 26280 30144
rect 28353 30141 28365 30144
rect 28399 30141 28411 30175
rect 28353 30135 28411 30141
rect 28994 30132 29000 30184
rect 29052 30132 29058 30184
rect 29104 30172 29132 30212
rect 29546 30200 29552 30252
rect 29604 30240 29610 30252
rect 30576 30249 30604 30280
rect 34698 30268 34704 30320
rect 34756 30308 34762 30320
rect 34793 30311 34851 30317
rect 34793 30308 34805 30311
rect 34756 30280 34805 30308
rect 34756 30268 34762 30280
rect 34793 30277 34805 30280
rect 34839 30277 34851 30311
rect 34793 30271 34851 30277
rect 29641 30243 29699 30249
rect 29641 30240 29653 30243
rect 29604 30212 29653 30240
rect 29604 30200 29610 30212
rect 29641 30209 29653 30212
rect 29687 30209 29699 30243
rect 29641 30203 29699 30209
rect 30561 30243 30619 30249
rect 30561 30209 30573 30243
rect 30607 30209 30619 30243
rect 30561 30203 30619 30209
rect 30650 30200 30656 30252
rect 30708 30240 30714 30252
rect 32950 30249 32956 30252
rect 30817 30243 30875 30249
rect 30817 30240 30829 30243
rect 30708 30212 30829 30240
rect 30708 30200 30714 30212
rect 30817 30209 30829 30212
rect 30863 30209 30875 30243
rect 30817 30203 30875 30209
rect 32928 30243 32956 30249
rect 32928 30209 32940 30243
rect 32928 30203 32956 30209
rect 32950 30200 32956 30203
rect 33008 30200 33014 30252
rect 33042 30200 33048 30252
rect 33100 30200 33106 30252
rect 33778 30200 33784 30252
rect 33836 30200 33842 30252
rect 33962 30200 33968 30252
rect 34020 30200 34026 30252
rect 36170 30200 36176 30252
rect 36228 30200 36234 30252
rect 36924 30240 36952 30336
rect 37734 30268 37740 30320
rect 37792 30268 37798 30320
rect 37093 30243 37151 30249
rect 37093 30240 37105 30243
rect 36924 30212 37105 30240
rect 37093 30209 37105 30212
rect 37139 30209 37151 30243
rect 37093 30203 37151 30209
rect 37458 30200 37464 30252
rect 37516 30200 37522 30252
rect 37642 30200 37648 30252
rect 37700 30200 37706 30252
rect 29825 30175 29883 30181
rect 29825 30172 29837 30175
rect 29104 30144 29837 30172
rect 29825 30141 29837 30144
rect 29871 30141 29883 30175
rect 29825 30135 29883 30141
rect 32766 30132 32772 30184
rect 32824 30172 32830 30184
rect 34241 30175 34299 30181
rect 34241 30172 34253 30175
rect 32824 30144 34253 30172
rect 32824 30132 32830 30144
rect 34241 30141 34253 30144
rect 34287 30141 34299 30175
rect 34241 30135 34299 30141
rect 24121 30107 24179 30113
rect 24121 30073 24133 30107
rect 24167 30104 24179 30107
rect 26234 30104 26240 30116
rect 24167 30076 26240 30104
rect 24167 30073 24179 30076
rect 24121 30067 24179 30073
rect 26234 30064 26240 30076
rect 26292 30064 26298 30116
rect 33318 30064 33324 30116
rect 33376 30064 33382 30116
rect 34256 30104 34284 30135
rect 34606 30132 34612 30184
rect 34664 30132 34670 30184
rect 34698 30132 34704 30184
rect 34756 30132 34762 30184
rect 35897 30175 35955 30181
rect 35897 30172 35909 30175
rect 34808 30144 35909 30172
rect 34808 30116 34836 30144
rect 35897 30141 35909 30144
rect 35943 30141 35955 30175
rect 35897 30135 35955 30141
rect 36056 30175 36114 30181
rect 36056 30141 36068 30175
rect 36102 30172 36114 30175
rect 36354 30172 36360 30184
rect 36102 30144 36360 30172
rect 36102 30141 36114 30144
rect 36056 30135 36114 30141
rect 36354 30132 36360 30144
rect 36412 30132 36418 30184
rect 36909 30175 36967 30181
rect 36909 30141 36921 30175
rect 36955 30172 36967 30175
rect 37476 30172 37504 30200
rect 36955 30144 37504 30172
rect 36955 30141 36967 30144
rect 36909 30135 36967 30141
rect 37826 30132 37832 30184
rect 37884 30172 37890 30184
rect 38289 30175 38347 30181
rect 38289 30172 38301 30175
rect 37884 30144 38301 30172
rect 37884 30132 37890 30144
rect 38289 30141 38301 30144
rect 38335 30141 38347 30175
rect 38289 30135 38347 30141
rect 34790 30104 34796 30116
rect 34256 30076 34796 30104
rect 34790 30064 34796 30076
rect 34848 30064 34854 30116
rect 35161 30107 35219 30113
rect 35161 30073 35173 30107
rect 35207 30104 35219 30107
rect 35434 30104 35440 30116
rect 35207 30076 35440 30104
rect 35207 30073 35219 30076
rect 35161 30067 35219 30073
rect 35434 30064 35440 30076
rect 35492 30064 35498 30116
rect 36449 30107 36507 30113
rect 36449 30073 36461 30107
rect 36495 30073 36507 30107
rect 36449 30067 36507 30073
rect 37277 30107 37335 30113
rect 37277 30073 37289 30107
rect 37323 30104 37335 30107
rect 37366 30104 37372 30116
rect 37323 30076 37372 30104
rect 37323 30073 37335 30076
rect 37277 30067 37335 30073
rect 24578 30036 24584 30048
rect 24044 30008 24584 30036
rect 24578 29996 24584 30008
rect 24636 29996 24642 30048
rect 27157 30039 27215 30045
rect 27157 30005 27169 30039
rect 27203 30036 27215 30039
rect 27982 30036 27988 30048
rect 27203 30008 27988 30036
rect 27203 30005 27215 30008
rect 27157 29999 27215 30005
rect 27982 29996 27988 30008
rect 28040 29996 28046 30048
rect 29086 29996 29092 30048
rect 29144 29996 29150 30048
rect 31941 30039 31999 30045
rect 31941 30005 31953 30039
rect 31987 30036 31999 30039
rect 32030 30036 32036 30048
rect 31987 30008 32036 30036
rect 31987 30005 31999 30008
rect 31941 29999 31999 30005
rect 32030 29996 32036 30008
rect 32088 29996 32094 30048
rect 32125 30039 32183 30045
rect 32125 30005 32137 30039
rect 32171 30036 32183 30039
rect 33410 30036 33416 30048
rect 32171 30008 33416 30036
rect 32171 30005 32183 30008
rect 32125 29999 32183 30005
rect 33410 29996 33416 30008
rect 33468 29996 33474 30048
rect 35253 30039 35311 30045
rect 35253 30005 35265 30039
rect 35299 30036 35311 30039
rect 35710 30036 35716 30048
rect 35299 30008 35716 30036
rect 35299 30005 35311 30008
rect 35253 29999 35311 30005
rect 35710 29996 35716 30008
rect 35768 29996 35774 30048
rect 35894 29996 35900 30048
rect 35952 30036 35958 30048
rect 36464 30036 36492 30067
rect 37366 30064 37372 30076
rect 37424 30064 37430 30116
rect 35952 30008 36492 30036
rect 35952 29996 35958 30008
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 9490 29792 9496 29844
rect 9548 29832 9554 29844
rect 10965 29835 11023 29841
rect 9548 29804 10916 29832
rect 9548 29792 9554 29804
rect 10888 29764 10916 29804
rect 10965 29801 10977 29835
rect 11011 29832 11023 29835
rect 11146 29832 11152 29844
rect 11011 29804 11152 29832
rect 11011 29801 11023 29804
rect 10965 29795 11023 29801
rect 11146 29792 11152 29804
rect 11204 29792 11210 29844
rect 13541 29835 13599 29841
rect 13541 29801 13553 29835
rect 13587 29832 13599 29835
rect 14550 29832 14556 29844
rect 13587 29804 14556 29832
rect 13587 29801 13599 29804
rect 13541 29795 13599 29801
rect 14550 29792 14556 29804
rect 14608 29832 14614 29844
rect 16574 29832 16580 29844
rect 14608 29804 16580 29832
rect 14608 29792 14614 29804
rect 16574 29792 16580 29804
rect 16632 29792 16638 29844
rect 17402 29792 17408 29844
rect 17460 29832 17466 29844
rect 17589 29835 17647 29841
rect 17589 29832 17601 29835
rect 17460 29804 17601 29832
rect 17460 29792 17466 29804
rect 17589 29801 17601 29804
rect 17635 29801 17647 29835
rect 17589 29795 17647 29801
rect 19058 29792 19064 29844
rect 19116 29832 19122 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 19116 29804 19257 29832
rect 19116 29792 19122 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 19245 29795 19303 29801
rect 22738 29792 22744 29844
rect 22796 29792 22802 29844
rect 23566 29792 23572 29844
rect 23624 29792 23630 29844
rect 24857 29835 24915 29841
rect 24857 29801 24869 29835
rect 24903 29832 24915 29835
rect 25222 29832 25228 29844
rect 24903 29804 25228 29832
rect 24903 29801 24915 29804
rect 24857 29795 24915 29801
rect 25222 29792 25228 29804
rect 25280 29792 25286 29844
rect 28537 29835 28595 29841
rect 28537 29801 28549 29835
rect 28583 29832 28595 29835
rect 28810 29832 28816 29844
rect 28583 29804 28816 29832
rect 28583 29801 28595 29804
rect 28537 29795 28595 29801
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 29086 29792 29092 29844
rect 29144 29792 29150 29844
rect 30650 29792 30656 29844
rect 30708 29792 30714 29844
rect 32030 29792 32036 29844
rect 32088 29832 32094 29844
rect 32950 29832 32956 29844
rect 32088 29804 32956 29832
rect 32088 29792 32094 29804
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 33226 29792 33232 29844
rect 33284 29792 33290 29844
rect 33781 29835 33839 29841
rect 33781 29801 33793 29835
rect 33827 29832 33839 29835
rect 34146 29832 34152 29844
rect 33827 29804 34152 29832
rect 33827 29801 33839 29804
rect 33781 29795 33839 29801
rect 34146 29792 34152 29804
rect 34204 29792 34210 29844
rect 37277 29835 37335 29841
rect 37277 29832 37289 29835
rect 35176 29804 37289 29832
rect 11238 29764 11244 29776
rect 10888 29736 11244 29764
rect 11238 29724 11244 29736
rect 11296 29724 11302 29776
rect 27062 29764 27068 29776
rect 14568 29736 19012 29764
rect 11609 29699 11667 29705
rect 11609 29665 11621 29699
rect 11655 29696 11667 29699
rect 11655 29668 11689 29696
rect 11655 29665 11667 29668
rect 11609 29659 11667 29665
rect 5994 29588 6000 29640
rect 6052 29588 6058 29640
rect 6362 29588 6368 29640
rect 6420 29628 6426 29640
rect 6733 29631 6791 29637
rect 6733 29628 6745 29631
rect 6420 29600 6745 29628
rect 6420 29588 6426 29600
rect 6733 29597 6745 29600
rect 6779 29597 6791 29631
rect 6733 29591 6791 29597
rect 8754 29588 8760 29640
rect 8812 29628 8818 29640
rect 9306 29628 9312 29640
rect 8812 29600 9312 29628
rect 8812 29588 8818 29600
rect 9306 29588 9312 29600
rect 9364 29628 9370 29640
rect 9585 29631 9643 29637
rect 9585 29628 9597 29631
rect 9364 29600 9597 29628
rect 9364 29588 9370 29600
rect 9585 29597 9597 29600
rect 9631 29597 9643 29631
rect 9585 29591 9643 29597
rect 9852 29631 9910 29637
rect 9852 29597 9864 29631
rect 9898 29628 9910 29631
rect 10318 29628 10324 29640
rect 9898 29600 10324 29628
rect 9898 29597 9910 29600
rect 9852 29591 9910 29597
rect 10318 29588 10324 29600
rect 10376 29588 10382 29640
rect 11624 29628 11652 29659
rect 11790 29656 11796 29708
rect 11848 29696 11854 29708
rect 12437 29699 12495 29705
rect 12437 29696 12449 29699
rect 11848 29668 12449 29696
rect 11848 29656 11854 29668
rect 12437 29665 12449 29668
rect 12483 29665 12495 29699
rect 12437 29659 12495 29665
rect 12894 29656 12900 29708
rect 12952 29696 12958 29708
rect 13354 29696 13360 29708
rect 12952 29668 13360 29696
rect 12952 29656 12958 29668
rect 13354 29656 13360 29668
rect 13412 29696 13418 29708
rect 14568 29705 14596 29736
rect 13909 29699 13967 29705
rect 13909 29696 13921 29699
rect 13412 29668 13921 29696
rect 13412 29656 13418 29668
rect 13909 29665 13921 29668
rect 13955 29696 13967 29699
rect 14553 29699 14611 29705
rect 14553 29696 14565 29699
rect 13955 29668 14565 29696
rect 13955 29665 13967 29668
rect 13909 29659 13967 29665
rect 14553 29665 14565 29668
rect 14599 29665 14611 29699
rect 14553 29659 14611 29665
rect 14645 29699 14703 29705
rect 14645 29665 14657 29699
rect 14691 29696 14703 29699
rect 15286 29696 15292 29708
rect 14691 29668 15292 29696
rect 14691 29665 14703 29668
rect 14645 29659 14703 29665
rect 15286 29656 15292 29668
rect 15344 29656 15350 29708
rect 18785 29699 18843 29705
rect 18785 29665 18797 29699
rect 18831 29665 18843 29699
rect 18785 29659 18843 29665
rect 13722 29628 13728 29640
rect 11164 29600 13728 29628
rect 9493 29563 9551 29569
rect 9493 29529 9505 29563
rect 9539 29560 9551 29563
rect 11164 29560 11192 29600
rect 13722 29588 13728 29600
rect 13780 29588 13786 29640
rect 18138 29588 18144 29640
rect 18196 29588 18202 29640
rect 18800 29628 18828 29659
rect 18874 29656 18880 29708
rect 18932 29656 18938 29708
rect 18984 29696 19012 29736
rect 23952 29736 27068 29764
rect 23952 29708 23980 29736
rect 27062 29724 27068 29736
rect 27120 29724 27126 29776
rect 19889 29699 19947 29705
rect 19889 29696 19901 29699
rect 18984 29668 19901 29696
rect 19889 29665 19901 29668
rect 19935 29696 19947 29699
rect 20257 29699 20315 29705
rect 20257 29696 20269 29699
rect 19935 29668 20269 29696
rect 19935 29665 19947 29668
rect 19889 29659 19947 29665
rect 20257 29665 20269 29668
rect 20303 29665 20315 29699
rect 20257 29659 20315 29665
rect 20714 29656 20720 29708
rect 20772 29656 20778 29708
rect 23385 29699 23443 29705
rect 23385 29665 23397 29699
rect 23431 29696 23443 29699
rect 23934 29696 23940 29708
rect 23431 29668 23940 29696
rect 23431 29665 23443 29668
rect 23385 29659 23443 29665
rect 23934 29656 23940 29668
rect 23992 29656 23998 29708
rect 24118 29656 24124 29708
rect 24176 29656 24182 29708
rect 24670 29656 24676 29708
rect 24728 29656 24734 29708
rect 24762 29656 24768 29708
rect 24820 29696 24826 29708
rect 25409 29699 25467 29705
rect 25409 29696 25421 29699
rect 24820 29668 25421 29696
rect 24820 29656 24826 29668
rect 25409 29665 25421 29668
rect 25455 29665 25467 29699
rect 25409 29659 25467 29665
rect 26142 29656 26148 29708
rect 26200 29696 26206 29708
rect 26970 29696 26976 29708
rect 26200 29668 26976 29696
rect 26200 29656 26206 29668
rect 26970 29656 26976 29668
rect 27028 29696 27034 29708
rect 27157 29699 27215 29705
rect 27157 29696 27169 29699
rect 27028 29668 27169 29696
rect 27028 29656 27034 29668
rect 27157 29665 27169 29668
rect 27203 29665 27215 29699
rect 27157 29659 27215 29665
rect 19610 29628 19616 29640
rect 18800 29600 19616 29628
rect 19610 29588 19616 29600
rect 19668 29588 19674 29640
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29628 19763 29631
rect 20732 29628 20760 29656
rect 19751 29600 20760 29628
rect 23201 29631 23259 29637
rect 19751 29597 19763 29600
rect 19705 29591 19763 29597
rect 23201 29597 23213 29631
rect 23247 29628 23259 29631
rect 24688 29628 24716 29656
rect 23247 29600 24716 29628
rect 25225 29631 25283 29637
rect 23247 29597 23259 29600
rect 23201 29591 23259 29597
rect 25225 29597 25237 29631
rect 25271 29628 25283 29631
rect 25866 29628 25872 29640
rect 25271 29600 25872 29628
rect 25271 29597 25283 29600
rect 25225 29591 25283 29597
rect 25866 29588 25872 29600
rect 25924 29588 25930 29640
rect 27424 29631 27482 29637
rect 27424 29597 27436 29631
rect 27470 29628 27482 29631
rect 29104 29628 29132 29792
rect 31389 29767 31447 29773
rect 31389 29733 31401 29767
rect 31435 29733 31447 29767
rect 33244 29764 33272 29792
rect 33873 29767 33931 29773
rect 33873 29764 33885 29767
rect 33244 29736 33885 29764
rect 31389 29727 31447 29733
rect 33873 29733 33885 29736
rect 33919 29733 33931 29767
rect 33873 29727 33931 29733
rect 31297 29699 31355 29705
rect 31297 29665 31309 29699
rect 31343 29696 31355 29699
rect 31404 29696 31432 29727
rect 32033 29699 32091 29705
rect 32033 29696 32045 29699
rect 31343 29668 31432 29696
rect 31680 29668 32045 29696
rect 31343 29665 31355 29668
rect 31297 29659 31355 29665
rect 27470 29600 29132 29628
rect 27470 29597 27482 29600
rect 27424 29591 27482 29597
rect 9539 29532 11192 29560
rect 9539 29529 9551 29532
rect 9493 29523 9551 29529
rect 11164 29504 11192 29532
rect 11425 29563 11483 29569
rect 11425 29529 11437 29563
rect 11471 29560 11483 29563
rect 11885 29563 11943 29569
rect 11885 29560 11897 29563
rect 11471 29532 11897 29560
rect 11471 29529 11483 29532
rect 11425 29523 11483 29529
rect 11885 29529 11897 29532
rect 11931 29529 11943 29563
rect 11885 29523 11943 29529
rect 16850 29520 16856 29572
rect 16908 29560 16914 29572
rect 17497 29563 17555 29569
rect 17497 29560 17509 29563
rect 16908 29532 17509 29560
rect 16908 29520 16914 29532
rect 17497 29529 17509 29532
rect 17543 29560 17555 29563
rect 18874 29560 18880 29572
rect 17543 29532 18880 29560
rect 17543 29529 17555 29532
rect 17497 29523 17555 29529
rect 18874 29520 18880 29532
rect 18932 29520 18938 29572
rect 19794 29520 19800 29572
rect 19852 29560 19858 29572
rect 20070 29560 20076 29572
rect 19852 29532 20076 29560
rect 19852 29520 19858 29532
rect 20070 29520 20076 29532
rect 20128 29520 20134 29572
rect 23109 29563 23167 29569
rect 23109 29529 23121 29563
rect 23155 29560 23167 29563
rect 23658 29560 23664 29572
rect 23155 29532 23664 29560
rect 23155 29529 23167 29532
rect 23109 29523 23167 29529
rect 23658 29520 23664 29532
rect 23716 29560 23722 29572
rect 26789 29563 26847 29569
rect 26789 29560 26801 29563
rect 23716 29532 24992 29560
rect 23716 29520 23722 29532
rect 24964 29504 24992 29532
rect 26252 29532 26801 29560
rect 26252 29504 26280 29532
rect 26789 29529 26801 29532
rect 26835 29529 26847 29563
rect 26789 29523 26847 29529
rect 30561 29563 30619 29569
rect 30561 29529 30573 29563
rect 30607 29560 30619 29563
rect 31680 29560 31708 29668
rect 32033 29665 32045 29668
rect 32079 29665 32091 29699
rect 32033 29659 32091 29665
rect 31754 29588 31760 29640
rect 31812 29588 31818 29640
rect 32048 29628 32076 29659
rect 32766 29656 32772 29708
rect 32824 29656 32830 29708
rect 33134 29656 33140 29708
rect 33192 29656 33198 29708
rect 35176 29705 35204 29804
rect 37277 29801 37289 29804
rect 37323 29801 37335 29835
rect 37277 29795 37335 29801
rect 37458 29792 37464 29844
rect 37516 29792 37522 29844
rect 37185 29767 37243 29773
rect 37185 29733 37197 29767
rect 37231 29764 37243 29767
rect 37476 29764 37504 29792
rect 37231 29736 37504 29764
rect 37231 29733 37243 29736
rect 37185 29727 37243 29733
rect 35161 29699 35219 29705
rect 35161 29665 35173 29699
rect 35207 29665 35219 29699
rect 35161 29659 35219 29665
rect 37274 29656 37280 29708
rect 37332 29696 37338 29708
rect 37829 29699 37887 29705
rect 37829 29696 37841 29699
rect 37332 29668 37841 29696
rect 37332 29656 37338 29668
rect 37829 29665 37841 29668
rect 37875 29696 37887 29699
rect 38289 29699 38347 29705
rect 38289 29696 38301 29699
rect 37875 29668 38301 29696
rect 37875 29665 37887 29668
rect 37829 29659 37887 29665
rect 38289 29665 38301 29668
rect 38335 29665 38347 29699
rect 38289 29659 38347 29665
rect 33413 29631 33471 29637
rect 32048 29600 32803 29628
rect 30607 29532 31708 29560
rect 31849 29563 31907 29569
rect 30607 29529 30619 29532
rect 30561 29523 30619 29529
rect 31849 29529 31861 29563
rect 31895 29560 31907 29563
rect 32775 29560 32803 29600
rect 33413 29597 33425 29631
rect 33459 29628 33471 29631
rect 34330 29628 34336 29640
rect 33459 29600 34336 29628
rect 33459 29597 33471 29600
rect 33413 29591 33471 29597
rect 34330 29588 34336 29600
rect 34388 29588 34394 29640
rect 34422 29588 34428 29640
rect 34480 29588 34486 29640
rect 35802 29588 35808 29640
rect 35860 29628 35866 29640
rect 36630 29628 36636 29640
rect 35860 29600 36636 29628
rect 35860 29588 35866 29600
rect 36630 29588 36636 29600
rect 36688 29588 36694 29640
rect 37645 29631 37703 29637
rect 37645 29597 37657 29631
rect 37691 29628 37703 29631
rect 38102 29628 38108 29640
rect 37691 29600 38108 29628
rect 37691 29597 37703 29600
rect 37645 29591 37703 29597
rect 38102 29588 38108 29600
rect 38160 29588 38166 29640
rect 31895 29532 32628 29560
rect 32775 29532 32904 29560
rect 31895 29529 31907 29532
rect 31849 29523 31907 29529
rect 32600 29504 32628 29532
rect 5350 29452 5356 29504
rect 5408 29452 5414 29504
rect 6178 29452 6184 29504
rect 6236 29452 6242 29504
rect 8202 29452 8208 29504
rect 8260 29492 8266 29504
rect 8757 29495 8815 29501
rect 8757 29492 8769 29495
rect 8260 29464 8769 29492
rect 8260 29452 8266 29464
rect 8757 29461 8769 29464
rect 8803 29492 8815 29495
rect 9858 29492 9864 29504
rect 8803 29464 9864 29492
rect 8803 29461 8815 29464
rect 8757 29455 8815 29461
rect 9858 29452 9864 29464
rect 9916 29492 9922 29504
rect 10778 29492 10784 29504
rect 9916 29464 10784 29492
rect 9916 29452 9922 29464
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 11054 29452 11060 29504
rect 11112 29452 11118 29504
rect 11146 29452 11152 29504
rect 11204 29452 11210 29504
rect 11330 29452 11336 29504
rect 11388 29492 11394 29504
rect 11517 29495 11575 29501
rect 11517 29492 11529 29495
rect 11388 29464 11529 29492
rect 11388 29452 11394 29464
rect 11517 29461 11529 29464
rect 11563 29492 11575 29495
rect 11606 29492 11612 29504
rect 11563 29464 11612 29492
rect 11563 29461 11575 29464
rect 11517 29455 11575 29461
rect 11606 29452 11612 29464
rect 11664 29452 11670 29504
rect 14734 29452 14740 29504
rect 14792 29452 14798 29504
rect 15102 29452 15108 29504
rect 15160 29452 15166 29504
rect 18322 29452 18328 29504
rect 18380 29452 18386 29504
rect 18693 29495 18751 29501
rect 18693 29461 18705 29495
rect 18739 29492 18751 29495
rect 19334 29492 19340 29504
rect 18739 29464 19340 29492
rect 18739 29461 18751 29464
rect 18693 29455 18751 29461
rect 19334 29452 19340 29464
rect 19392 29492 19398 29504
rect 19613 29495 19671 29501
rect 19613 29492 19625 29495
rect 19392 29464 19625 29492
rect 19392 29452 19398 29464
rect 19613 29461 19625 29464
rect 19659 29492 19671 29495
rect 19978 29492 19984 29504
rect 19659 29464 19984 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 19978 29452 19984 29464
rect 20036 29452 20042 29504
rect 24118 29452 24124 29504
rect 24176 29492 24182 29504
rect 24673 29495 24731 29501
rect 24673 29492 24685 29495
rect 24176 29464 24685 29492
rect 24176 29452 24182 29464
rect 24673 29461 24685 29464
rect 24719 29492 24731 29495
rect 24762 29492 24768 29504
rect 24719 29464 24768 29492
rect 24719 29461 24731 29464
rect 24673 29455 24731 29461
rect 24762 29452 24768 29464
rect 24820 29452 24826 29504
rect 24946 29452 24952 29504
rect 25004 29492 25010 29504
rect 25317 29495 25375 29501
rect 25317 29492 25329 29495
rect 25004 29464 25329 29492
rect 25004 29452 25010 29464
rect 25317 29461 25329 29464
rect 25363 29461 25375 29495
rect 25317 29455 25375 29461
rect 25961 29495 26019 29501
rect 25961 29461 25973 29495
rect 26007 29492 26019 29495
rect 26234 29492 26240 29504
rect 26007 29464 26240 29492
rect 26007 29461 26019 29464
rect 25961 29455 26019 29461
rect 26234 29452 26240 29464
rect 26292 29452 26298 29504
rect 26418 29452 26424 29504
rect 26476 29452 26482 29504
rect 32214 29452 32220 29504
rect 32272 29452 32278 29504
rect 32582 29452 32588 29504
rect 32640 29452 32646 29504
rect 32674 29452 32680 29504
rect 32732 29452 32738 29504
rect 32876 29492 32904 29532
rect 32950 29520 32956 29572
rect 33008 29560 33014 29572
rect 33321 29563 33379 29569
rect 33321 29560 33333 29563
rect 33008 29532 33333 29560
rect 33008 29520 33014 29532
rect 33321 29529 33333 29532
rect 33367 29529 33379 29563
rect 33321 29523 33379 29529
rect 34698 29520 34704 29572
rect 34756 29560 34762 29572
rect 35713 29563 35771 29569
rect 34756 29532 35020 29560
rect 34756 29520 34762 29532
rect 34606 29492 34612 29504
rect 32876 29464 34612 29492
rect 34606 29452 34612 29464
rect 34664 29492 34670 29504
rect 34885 29495 34943 29501
rect 34885 29492 34897 29495
rect 34664 29464 34897 29492
rect 34664 29452 34670 29464
rect 34885 29461 34897 29464
rect 34931 29461 34943 29495
rect 34992 29492 35020 29532
rect 35713 29529 35725 29563
rect 35759 29560 35771 29563
rect 36050 29563 36108 29569
rect 36050 29560 36062 29563
rect 35759 29532 36062 29560
rect 35759 29529 35771 29532
rect 35713 29523 35771 29529
rect 36050 29529 36062 29532
rect 36096 29529 36108 29563
rect 36050 29523 36108 29529
rect 36446 29492 36452 29504
rect 34992 29464 36452 29492
rect 34885 29455 34943 29461
rect 36446 29452 36452 29464
rect 36504 29492 36510 29504
rect 37642 29492 37648 29504
rect 36504 29464 37648 29492
rect 36504 29452 36510 29464
rect 37642 29452 37648 29464
rect 37700 29492 37706 29504
rect 37737 29495 37795 29501
rect 37737 29492 37749 29495
rect 37700 29464 37749 29492
rect 37700 29452 37706 29464
rect 37737 29461 37749 29464
rect 37783 29461 37795 29495
rect 37737 29455 37795 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5905 29291 5963 29297
rect 5905 29257 5917 29291
rect 5951 29288 5963 29291
rect 6178 29288 6184 29300
rect 5951 29260 6184 29288
rect 5951 29257 5963 29260
rect 5905 29251 5963 29257
rect 6178 29248 6184 29260
rect 6236 29248 6242 29300
rect 10137 29291 10195 29297
rect 10137 29257 10149 29291
rect 10183 29288 10195 29291
rect 10594 29288 10600 29300
rect 10183 29260 10600 29288
rect 10183 29257 10195 29260
rect 10137 29251 10195 29257
rect 10594 29248 10600 29260
rect 10652 29288 10658 29300
rect 11790 29288 11796 29300
rect 10652 29260 11796 29288
rect 10652 29248 10658 29260
rect 11790 29248 11796 29260
rect 11848 29248 11854 29300
rect 12618 29288 12624 29300
rect 12406 29260 12624 29288
rect 5074 29180 5080 29232
rect 5132 29220 5138 29232
rect 6365 29223 6423 29229
rect 6365 29220 6377 29223
rect 5132 29192 6377 29220
rect 5132 29180 5138 29192
rect 6365 29189 6377 29192
rect 6411 29189 6423 29223
rect 11517 29223 11575 29229
rect 11517 29220 11529 29223
rect 6365 29183 6423 29189
rect 8772 29192 11529 29220
rect 5810 29112 5816 29164
rect 5868 29112 5874 29164
rect 8772 29096 8800 29192
rect 11517 29189 11529 29192
rect 11563 29220 11575 29223
rect 12406 29220 12434 29260
rect 12618 29248 12624 29260
rect 12676 29248 12682 29300
rect 14090 29248 14096 29300
rect 14148 29288 14154 29300
rect 14277 29291 14335 29297
rect 14277 29288 14289 29291
rect 14148 29260 14289 29288
rect 14148 29248 14154 29260
rect 14277 29257 14289 29260
rect 14323 29257 14335 29291
rect 14277 29251 14335 29257
rect 17497 29291 17555 29297
rect 17497 29257 17509 29291
rect 17543 29288 17555 29291
rect 17954 29288 17960 29300
rect 17543 29260 17960 29288
rect 17543 29257 17555 29260
rect 17497 29251 17555 29257
rect 17954 29248 17960 29260
rect 18012 29248 18018 29300
rect 18138 29248 18144 29300
rect 18196 29288 18202 29300
rect 18233 29291 18291 29297
rect 18233 29288 18245 29291
rect 18196 29260 18245 29288
rect 18196 29248 18202 29260
rect 18233 29257 18245 29260
rect 18279 29257 18291 29291
rect 18233 29251 18291 29257
rect 18322 29248 18328 29300
rect 18380 29248 18386 29300
rect 18693 29291 18751 29297
rect 18693 29257 18705 29291
rect 18739 29288 18751 29291
rect 19334 29288 19340 29300
rect 18739 29260 19340 29288
rect 18739 29257 18751 29260
rect 18693 29251 18751 29257
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 19426 29248 19432 29300
rect 19484 29248 19490 29300
rect 31294 29248 31300 29300
rect 31352 29248 31358 29300
rect 32214 29248 32220 29300
rect 32272 29248 32278 29300
rect 32674 29248 32680 29300
rect 32732 29288 32738 29300
rect 32953 29291 33011 29297
rect 32953 29288 32965 29291
rect 32732 29260 32965 29288
rect 32732 29248 32738 29260
rect 32953 29257 32965 29260
rect 32999 29257 33011 29291
rect 32953 29251 33011 29257
rect 33870 29248 33876 29300
rect 33928 29248 33934 29300
rect 34422 29248 34428 29300
rect 34480 29248 34486 29300
rect 34514 29248 34520 29300
rect 34572 29288 34578 29300
rect 34885 29291 34943 29297
rect 34885 29288 34897 29291
rect 34572 29260 34897 29288
rect 34572 29248 34578 29260
rect 34885 29257 34897 29260
rect 34931 29257 34943 29291
rect 34885 29251 34943 29257
rect 36357 29291 36415 29297
rect 36357 29257 36369 29291
rect 36403 29288 36415 29291
rect 36722 29288 36728 29300
rect 36403 29260 36728 29288
rect 36403 29257 36415 29260
rect 36357 29251 36415 29257
rect 11563 29192 12434 29220
rect 11563 29189 11575 29192
rect 11517 29183 11575 29189
rect 13722 29180 13728 29232
rect 13780 29220 13786 29232
rect 13780 29192 17448 29220
rect 13780 29180 13786 29192
rect 9024 29155 9082 29161
rect 9024 29121 9036 29155
rect 9070 29152 9082 29155
rect 10229 29155 10287 29161
rect 10229 29152 10241 29155
rect 9070 29124 10241 29152
rect 9070 29121 9082 29124
rect 9024 29115 9082 29121
rect 10229 29121 10241 29124
rect 10275 29121 10287 29155
rect 10229 29115 10287 29121
rect 10873 29155 10931 29161
rect 10873 29121 10885 29155
rect 10919 29152 10931 29155
rect 11054 29152 11060 29164
rect 10919 29124 11060 29152
rect 10919 29121 10931 29124
rect 10873 29115 10931 29121
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 11333 29155 11391 29161
rect 11333 29121 11345 29155
rect 11379 29152 11391 29155
rect 13265 29155 13323 29161
rect 13265 29152 13277 29155
rect 11379 29124 13277 29152
rect 11379 29121 11391 29124
rect 11333 29115 11391 29121
rect 13265 29121 13277 29124
rect 13311 29152 13323 29155
rect 15194 29152 15200 29164
rect 13311 29124 15200 29152
rect 13311 29121 13323 29124
rect 13265 29115 13323 29121
rect 15194 29112 15200 29124
rect 15252 29112 15258 29164
rect 5353 29087 5411 29093
rect 5353 29053 5365 29087
rect 5399 29053 5411 29087
rect 5353 29047 5411 29053
rect 6089 29087 6147 29093
rect 6089 29053 6101 29087
rect 6135 29053 6147 29087
rect 6089 29047 6147 29053
rect 5368 29016 5396 29047
rect 5445 29019 5503 29025
rect 5445 29016 5457 29019
rect 5368 28988 5457 29016
rect 5445 28985 5457 28988
rect 5491 28985 5503 29019
rect 6104 29016 6132 29047
rect 6454 29044 6460 29096
rect 6512 29084 6518 29096
rect 6917 29087 6975 29093
rect 6917 29084 6929 29087
rect 6512 29056 6929 29084
rect 6512 29044 6518 29056
rect 6917 29053 6929 29056
rect 6963 29053 6975 29087
rect 6917 29047 6975 29053
rect 8754 29044 8760 29096
rect 8812 29044 8818 29096
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29084 14979 29087
rect 15102 29084 15108 29096
rect 14967 29056 15108 29084
rect 14967 29053 14979 29056
rect 14921 29047 14979 29053
rect 15102 29044 15108 29056
rect 15160 29044 15166 29096
rect 17420 29093 17448 29192
rect 18141 29155 18199 29161
rect 18141 29121 18153 29155
rect 18187 29152 18199 29155
rect 18340 29152 18368 29248
rect 18187 29124 18368 29152
rect 18601 29155 18659 29161
rect 18187 29121 18199 29124
rect 18141 29115 18199 29121
rect 18601 29121 18613 29155
rect 18647 29152 18659 29155
rect 19061 29155 19119 29161
rect 19061 29152 19073 29155
rect 18647 29124 19073 29152
rect 18647 29121 18659 29124
rect 18601 29115 18659 29121
rect 19061 29121 19073 29124
rect 19107 29121 19119 29155
rect 19444 29152 19472 29248
rect 19613 29155 19671 29161
rect 19613 29152 19625 29155
rect 19444 29124 19625 29152
rect 19061 29115 19119 29121
rect 19613 29121 19625 29124
rect 19659 29121 19671 29155
rect 19613 29115 19671 29121
rect 31941 29155 31999 29161
rect 31941 29121 31953 29155
rect 31987 29152 31999 29155
rect 32232 29152 32260 29248
rect 32401 29223 32459 29229
rect 32401 29189 32413 29223
rect 32447 29220 32459 29223
rect 33888 29220 33916 29248
rect 32447 29192 33916 29220
rect 32447 29189 32459 29192
rect 32401 29183 32459 29189
rect 31987 29124 32260 29152
rect 32493 29155 32551 29161
rect 31987 29121 31999 29124
rect 31941 29115 31999 29121
rect 32493 29121 32505 29155
rect 32539 29152 32551 29155
rect 32582 29152 32588 29164
rect 32539 29124 32588 29152
rect 32539 29121 32551 29124
rect 32493 29115 32551 29121
rect 32582 29112 32588 29124
rect 32640 29152 32646 29164
rect 32950 29152 32956 29164
rect 32640 29124 32956 29152
rect 32640 29112 32646 29124
rect 32950 29112 32956 29124
rect 33008 29112 33014 29164
rect 33042 29112 33048 29164
rect 33100 29152 33106 29164
rect 33505 29155 33563 29161
rect 33505 29152 33517 29155
rect 33100 29124 33517 29152
rect 33100 29112 33106 29124
rect 33505 29121 33517 29124
rect 33551 29121 33563 29155
rect 33505 29115 33563 29121
rect 17405 29087 17463 29093
rect 17405 29053 17417 29087
rect 17451 29084 17463 29087
rect 18785 29087 18843 29093
rect 18785 29084 18797 29087
rect 17451 29056 18797 29084
rect 17451 29053 17463 29056
rect 17405 29047 17463 29053
rect 18785 29053 18797 29056
rect 18831 29053 18843 29087
rect 32214 29084 32220 29096
rect 18785 29047 18843 29053
rect 31128 29056 32220 29084
rect 7377 29019 7435 29025
rect 7377 29016 7389 29019
rect 6104 28988 7389 29016
rect 5445 28979 5503 28985
rect 7377 28985 7389 28988
rect 7423 29016 7435 29019
rect 7926 29016 7932 29028
rect 7423 28988 7932 29016
rect 7423 28985 7435 28988
rect 7377 28979 7435 28985
rect 7926 28976 7932 28988
rect 7984 28976 7990 29028
rect 4614 28908 4620 28960
rect 4672 28908 4678 28960
rect 4706 28908 4712 28960
rect 4764 28908 4770 28960
rect 8018 28908 8024 28960
rect 8076 28948 8082 28960
rect 8772 28948 8800 29044
rect 31128 29028 31156 29056
rect 32214 29044 32220 29056
rect 32272 29044 32278 29096
rect 33134 29044 33140 29096
rect 33192 29084 33198 29096
rect 33873 29087 33931 29093
rect 33873 29084 33885 29087
rect 33192 29056 33885 29084
rect 33192 29044 33198 29056
rect 33873 29053 33885 29056
rect 33919 29053 33931 29087
rect 33873 29047 33931 29053
rect 23661 29019 23719 29025
rect 23661 28985 23673 29019
rect 23707 29016 23719 29019
rect 23934 29016 23940 29028
rect 23707 28988 23940 29016
rect 23707 28985 23719 28988
rect 23661 28979 23719 28985
rect 23934 28976 23940 28988
rect 23992 28976 23998 29028
rect 24578 28976 24584 29028
rect 24636 29016 24642 29028
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 24636 28988 24869 29016
rect 24636 28976 24642 28988
rect 24857 28985 24869 28988
rect 24903 29016 24915 29019
rect 27157 29019 27215 29025
rect 27157 29016 27169 29019
rect 24903 28988 27169 29016
rect 24903 28985 24915 28988
rect 24857 28979 24915 28985
rect 27157 28985 27169 28988
rect 27203 29016 27215 29019
rect 27798 29016 27804 29028
rect 27203 28988 27804 29016
rect 27203 28985 27215 28988
rect 27157 28979 27215 28985
rect 27798 28976 27804 28988
rect 27856 29016 27862 29028
rect 28534 29016 28540 29028
rect 27856 28988 28540 29016
rect 27856 28976 27862 28988
rect 28534 28976 28540 28988
rect 28592 28976 28598 29028
rect 30742 28976 30748 29028
rect 30800 29016 30806 29028
rect 30800 28988 31064 29016
rect 30800 28976 30806 28988
rect 8076 28920 8800 28948
rect 13725 28951 13783 28957
rect 8076 28908 8082 28920
rect 13725 28917 13737 28951
rect 13771 28948 13783 28951
rect 13814 28948 13820 28960
rect 13771 28920 13820 28948
rect 13771 28917 13783 28920
rect 13725 28911 13783 28917
rect 13814 28908 13820 28920
rect 13872 28908 13878 28960
rect 31036 28948 31064 28988
rect 31110 28976 31116 29028
rect 31168 28976 31174 29028
rect 32766 29016 32772 29028
rect 31220 28988 32772 29016
rect 31220 28948 31248 28988
rect 32766 28976 32772 28988
rect 32824 28976 32830 29028
rect 32861 29019 32919 29025
rect 32861 28985 32873 29019
rect 32907 29016 32919 29019
rect 34440 29016 34468 29248
rect 34790 29180 34796 29232
rect 34848 29180 34854 29232
rect 34900 29220 34928 29251
rect 36722 29248 36728 29260
rect 36780 29248 36786 29300
rect 36814 29248 36820 29300
rect 36872 29248 36878 29300
rect 35894 29220 35900 29232
rect 34900 29192 35900 29220
rect 35894 29180 35900 29192
rect 35952 29180 35958 29232
rect 34808 29152 34836 29180
rect 35253 29155 35311 29161
rect 35253 29152 35265 29155
rect 34808 29124 35265 29152
rect 35253 29121 35265 29124
rect 35299 29121 35311 29155
rect 35253 29115 35311 29121
rect 36078 29112 36084 29164
rect 36136 29152 36142 29164
rect 36446 29152 36452 29164
rect 36136 29124 36452 29152
rect 36136 29112 36142 29124
rect 36446 29112 36452 29124
rect 36504 29112 36510 29164
rect 36173 29087 36231 29093
rect 36173 29053 36185 29087
rect 36219 29053 36231 29087
rect 36173 29047 36231 29053
rect 32907 28988 34468 29016
rect 32907 28985 32919 28988
rect 32861 28979 32919 28985
rect 35894 28976 35900 29028
rect 35952 29016 35958 29028
rect 36188 29016 36216 29047
rect 37642 29044 37648 29096
rect 37700 29084 37706 29096
rect 37829 29087 37887 29093
rect 37829 29084 37841 29087
rect 37700 29056 37841 29084
rect 37700 29044 37706 29056
rect 37829 29053 37841 29056
rect 37875 29053 37887 29087
rect 37829 29047 37887 29053
rect 35952 28988 36216 29016
rect 35952 28976 35958 28988
rect 36262 28976 36268 29028
rect 36320 29016 36326 29028
rect 37277 29019 37335 29025
rect 37277 29016 37289 29019
rect 36320 28988 37289 29016
rect 36320 28976 36326 28988
rect 37277 28985 37289 28988
rect 37323 28985 37335 29019
rect 37277 28979 37335 28985
rect 31036 28920 31248 28948
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 10778 28704 10784 28756
rect 10836 28744 10842 28756
rect 15010 28744 15016 28756
rect 10836 28716 15016 28744
rect 10836 28704 10842 28716
rect 15010 28704 15016 28716
rect 15068 28704 15074 28756
rect 3786 28500 3792 28552
rect 3844 28500 3850 28552
rect 4706 28500 4712 28552
rect 4764 28500 4770 28552
rect 4985 28543 5043 28549
rect 4985 28509 4997 28543
rect 5031 28540 5043 28543
rect 6178 28540 6184 28552
rect 5031 28512 6184 28540
rect 5031 28509 5043 28512
rect 4985 28503 5043 28509
rect 6178 28500 6184 28512
rect 6236 28500 6242 28552
rect 6457 28543 6515 28549
rect 6457 28509 6469 28543
rect 6503 28509 6515 28543
rect 6457 28503 6515 28509
rect 4724 28472 4752 28500
rect 5230 28475 5288 28481
rect 5230 28472 5242 28475
rect 4724 28444 5242 28472
rect 5230 28441 5242 28444
rect 5276 28441 5288 28475
rect 5230 28435 5288 28441
rect 5442 28432 5448 28484
rect 5500 28472 5506 28484
rect 6472 28472 6500 28503
rect 7190 28500 7196 28552
rect 7248 28500 7254 28552
rect 9766 28500 9772 28552
rect 9824 28500 9830 28552
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 11057 28543 11115 28549
rect 11057 28540 11069 28543
rect 10008 28512 11069 28540
rect 10008 28500 10014 28512
rect 11057 28509 11069 28512
rect 11103 28509 11115 28543
rect 11057 28503 11115 28509
rect 14458 28500 14464 28552
rect 14516 28500 14522 28552
rect 18046 28500 18052 28552
rect 18104 28500 18110 28552
rect 19426 28500 19432 28552
rect 19484 28540 19490 28552
rect 19889 28543 19947 28549
rect 19889 28540 19901 28543
rect 19484 28512 19901 28540
rect 19484 28500 19490 28512
rect 19889 28509 19901 28512
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28540 23535 28543
rect 23566 28540 23572 28552
rect 23523 28512 23572 28540
rect 23523 28509 23535 28512
rect 23477 28503 23535 28509
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 23658 28500 23664 28552
rect 23716 28540 23722 28552
rect 24397 28543 24455 28549
rect 24397 28540 24409 28543
rect 23716 28512 24409 28540
rect 23716 28500 23722 28512
rect 24397 28509 24409 28512
rect 24443 28509 24455 28543
rect 24397 28503 24455 28509
rect 25038 28500 25044 28552
rect 25096 28500 25102 28552
rect 27338 28500 27344 28552
rect 27396 28500 27402 28552
rect 27430 28500 27436 28552
rect 27488 28540 27494 28552
rect 28077 28543 28135 28549
rect 28077 28540 28089 28543
rect 27488 28512 28089 28540
rect 27488 28500 27494 28512
rect 28077 28509 28089 28512
rect 28123 28509 28135 28543
rect 28077 28503 28135 28509
rect 28350 28500 28356 28552
rect 28408 28540 28414 28552
rect 28813 28543 28871 28549
rect 28813 28540 28825 28543
rect 28408 28512 28825 28540
rect 28408 28500 28414 28512
rect 28813 28509 28825 28512
rect 28859 28509 28871 28543
rect 28813 28503 28871 28509
rect 33134 28500 33140 28552
rect 33192 28540 33198 28552
rect 33505 28543 33563 28549
rect 33505 28540 33517 28543
rect 33192 28512 33517 28540
rect 33192 28500 33198 28512
rect 33505 28509 33517 28512
rect 33551 28509 33563 28543
rect 33505 28503 33563 28509
rect 34238 28500 34244 28552
rect 34296 28500 34302 28552
rect 37918 28500 37924 28552
rect 37976 28500 37982 28552
rect 5500 28444 6500 28472
rect 13633 28475 13691 28481
rect 5500 28432 5506 28444
rect 13633 28441 13645 28475
rect 13679 28472 13691 28475
rect 13814 28472 13820 28484
rect 13679 28444 13820 28472
rect 13679 28441 13691 28444
rect 13633 28435 13691 28441
rect 13814 28432 13820 28444
rect 13872 28472 13878 28484
rect 14642 28472 14648 28484
rect 13872 28444 14648 28472
rect 13872 28432 13878 28444
rect 14642 28432 14648 28444
rect 14700 28432 14706 28484
rect 31113 28475 31171 28481
rect 31113 28472 31125 28475
rect 31036 28444 31125 28472
rect 31036 28416 31064 28444
rect 31113 28441 31125 28444
rect 31159 28472 31171 28475
rect 35345 28475 35403 28481
rect 35345 28472 35357 28475
rect 31159 28444 35357 28472
rect 31159 28441 31171 28444
rect 31113 28435 31171 28441
rect 35345 28441 35357 28444
rect 35391 28472 35403 28475
rect 35529 28475 35587 28481
rect 35529 28472 35541 28475
rect 35391 28444 35541 28472
rect 35391 28441 35403 28444
rect 35345 28435 35403 28441
rect 35529 28441 35541 28444
rect 35575 28441 35587 28475
rect 35529 28435 35587 28441
rect 4433 28407 4491 28413
rect 4433 28373 4445 28407
rect 4479 28404 4491 28407
rect 4614 28404 4620 28416
rect 4479 28376 4620 28404
rect 4479 28373 4491 28376
rect 4433 28367 4491 28373
rect 4614 28364 4620 28376
rect 4672 28364 4678 28416
rect 4706 28364 4712 28416
rect 4764 28364 4770 28416
rect 5534 28364 5540 28416
rect 5592 28404 5598 28416
rect 6362 28404 6368 28416
rect 5592 28376 6368 28404
rect 5592 28364 5598 28376
rect 6362 28364 6368 28376
rect 6420 28364 6426 28416
rect 7098 28364 7104 28416
rect 7156 28364 7162 28416
rect 7650 28364 7656 28416
rect 7708 28404 7714 28416
rect 7837 28407 7895 28413
rect 7837 28404 7849 28407
rect 7708 28376 7849 28404
rect 7708 28364 7714 28376
rect 7837 28373 7849 28376
rect 7883 28373 7895 28407
rect 7837 28367 7895 28373
rect 10321 28407 10379 28413
rect 10321 28373 10333 28407
rect 10367 28404 10379 28407
rect 10410 28404 10416 28416
rect 10367 28376 10416 28404
rect 10367 28373 10379 28376
rect 10321 28367 10379 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 10502 28364 10508 28416
rect 10560 28364 10566 28416
rect 14369 28407 14427 28413
rect 14369 28373 14381 28407
rect 14415 28404 14427 28407
rect 15010 28404 15016 28416
rect 14415 28376 15016 28404
rect 14415 28373 14427 28376
rect 14369 28367 14427 28373
rect 15010 28364 15016 28376
rect 15068 28364 15074 28416
rect 15105 28407 15163 28413
rect 15105 28373 15117 28407
rect 15151 28404 15163 28407
rect 15286 28404 15292 28416
rect 15151 28376 15292 28404
rect 15151 28373 15163 28376
rect 15105 28367 15163 28373
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 18506 28364 18512 28416
rect 18564 28404 18570 28416
rect 18601 28407 18659 28413
rect 18601 28404 18613 28407
rect 18564 28376 18613 28404
rect 18564 28364 18570 28376
rect 18601 28373 18613 28376
rect 18647 28373 18659 28407
rect 18601 28367 18659 28373
rect 18966 28364 18972 28416
rect 19024 28364 19030 28416
rect 19334 28364 19340 28416
rect 19392 28364 19398 28416
rect 22830 28364 22836 28416
rect 22888 28364 22894 28416
rect 23750 28364 23756 28416
rect 23808 28364 23814 28416
rect 26786 28364 26792 28416
rect 26844 28364 26850 28416
rect 27522 28364 27528 28416
rect 27580 28364 27586 28416
rect 28258 28364 28264 28416
rect 28316 28364 28322 28416
rect 28626 28364 28632 28416
rect 28684 28404 28690 28416
rect 29181 28407 29239 28413
rect 29181 28404 29193 28407
rect 28684 28376 29193 28404
rect 28684 28364 28690 28376
rect 29181 28373 29193 28376
rect 29227 28373 29239 28407
rect 29181 28367 29239 28373
rect 31018 28364 31024 28416
rect 31076 28364 31082 28416
rect 32398 28364 32404 28416
rect 32456 28364 32462 28416
rect 32950 28364 32956 28416
rect 33008 28364 33014 28416
rect 33686 28364 33692 28416
rect 33744 28364 33750 28416
rect 36630 28364 36636 28416
rect 36688 28404 36694 28416
rect 36817 28407 36875 28413
rect 36817 28404 36829 28407
rect 36688 28376 36829 28404
rect 36688 28364 36694 28376
rect 36817 28373 36829 28376
rect 36863 28373 36875 28407
rect 36817 28367 36875 28373
rect 36906 28364 36912 28416
rect 36964 28404 36970 28416
rect 37369 28407 37427 28413
rect 37369 28404 37381 28407
rect 36964 28376 37381 28404
rect 36964 28364 36970 28376
rect 37369 28373 37381 28376
rect 37415 28373 37427 28407
rect 37369 28367 37427 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 4249 28203 4307 28209
rect 4249 28169 4261 28203
rect 4295 28200 4307 28203
rect 5350 28200 5356 28212
rect 4295 28172 5356 28200
rect 4295 28169 4307 28172
rect 4249 28163 4307 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 5994 28160 6000 28212
rect 6052 28200 6058 28212
rect 6365 28203 6423 28209
rect 6365 28200 6377 28203
rect 6052 28172 6377 28200
rect 6052 28160 6058 28172
rect 6365 28169 6377 28172
rect 6411 28169 6423 28203
rect 6365 28163 6423 28169
rect 7190 28160 7196 28212
rect 7248 28160 7254 28212
rect 7650 28160 7656 28212
rect 7708 28160 7714 28212
rect 8113 28203 8171 28209
rect 8113 28169 8125 28203
rect 8159 28200 8171 28203
rect 8202 28200 8208 28212
rect 8159 28172 8208 28200
rect 8159 28169 8171 28172
rect 8113 28163 8171 28169
rect 8202 28160 8208 28172
rect 8260 28160 8266 28212
rect 9766 28160 9772 28212
rect 9824 28160 9830 28212
rect 10229 28203 10287 28209
rect 10229 28169 10241 28203
rect 10275 28200 10287 28203
rect 10502 28200 10508 28212
rect 10275 28172 10508 28200
rect 10275 28169 10287 28172
rect 10229 28163 10287 28169
rect 10502 28160 10508 28172
rect 10560 28160 10566 28212
rect 14458 28160 14464 28212
rect 14516 28160 14522 28212
rect 15194 28160 15200 28212
rect 15252 28200 15258 28212
rect 16853 28203 16911 28209
rect 16853 28200 16865 28203
rect 15252 28172 16865 28200
rect 15252 28160 15258 28172
rect 16853 28169 16865 28172
rect 16899 28200 16911 28203
rect 16899 28172 17080 28200
rect 16899 28169 16911 28172
rect 16853 28163 16911 28169
rect 5718 28132 5724 28144
rect 4540 28104 5724 28132
rect 3694 28024 3700 28076
rect 3752 28064 3758 28076
rect 4341 28067 4399 28073
rect 4341 28064 4353 28067
rect 3752 28036 4353 28064
rect 3752 28024 3758 28036
rect 4341 28033 4353 28036
rect 4387 28033 4399 28067
rect 4341 28027 4399 28033
rect 4540 28008 4568 28104
rect 5718 28092 5724 28104
rect 5776 28092 5782 28144
rect 7208 28132 7236 28160
rect 5828 28104 7236 28132
rect 7500 28135 7558 28141
rect 5828 28064 5856 28104
rect 7500 28101 7512 28135
rect 7546 28132 7558 28135
rect 7668 28132 7696 28160
rect 14734 28132 14740 28144
rect 7546 28104 7696 28132
rect 14016 28104 14740 28132
rect 7546 28101 7558 28104
rect 7500 28095 7558 28101
rect 5184 28036 5856 28064
rect 5925 28067 5983 28073
rect 2409 27999 2467 28005
rect 2409 27965 2421 27999
rect 2455 27996 2467 27999
rect 2774 27996 2780 28008
rect 2455 27968 2780 27996
rect 2455 27965 2467 27968
rect 2409 27959 2467 27965
rect 2774 27956 2780 27968
rect 2832 27956 2838 28008
rect 3602 27956 3608 28008
rect 3660 27956 3666 28008
rect 4157 27999 4215 28005
rect 4157 27965 4169 27999
rect 4203 27996 4215 27999
rect 4522 27996 4528 28008
rect 4203 27968 4528 27996
rect 4203 27965 4215 27968
rect 4157 27959 4215 27965
rect 4522 27956 4528 27968
rect 4580 27956 4586 28008
rect 4709 27931 4767 27937
rect 4709 27897 4721 27931
rect 4755 27928 4767 27931
rect 5184 27928 5212 28036
rect 5925 28033 5937 28067
rect 5971 28064 5983 28067
rect 6914 28064 6920 28076
rect 5971 28036 6920 28064
rect 5971 28033 5983 28036
rect 5925 28027 5983 28033
rect 6914 28024 6920 28036
rect 6972 28024 6978 28076
rect 10137 28067 10195 28073
rect 10137 28033 10149 28067
rect 10183 28064 10195 28067
rect 11330 28064 11336 28076
rect 10183 28036 11336 28064
rect 10183 28033 10195 28036
rect 10137 28027 10195 28033
rect 10704 28008 10732 28036
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 14016 28008 14044 28104
rect 14734 28092 14740 28104
rect 14792 28132 14798 28144
rect 17052 28141 17080 28172
rect 18230 28160 18236 28212
rect 18288 28200 18294 28212
rect 18325 28203 18383 28209
rect 18325 28200 18337 28203
rect 18288 28172 18337 28200
rect 18288 28160 18294 28172
rect 18325 28169 18337 28172
rect 18371 28169 18383 28203
rect 18325 28163 18383 28169
rect 19245 28203 19303 28209
rect 19245 28169 19257 28203
rect 19291 28200 19303 28203
rect 19334 28200 19340 28212
rect 19291 28172 19340 28200
rect 19291 28169 19303 28172
rect 19245 28163 19303 28169
rect 19334 28160 19340 28172
rect 19392 28160 19398 28212
rect 22465 28203 22523 28209
rect 22465 28169 22477 28203
rect 22511 28200 22523 28203
rect 22738 28200 22744 28212
rect 22511 28172 22744 28200
rect 22511 28169 22523 28172
rect 22465 28163 22523 28169
rect 22738 28160 22744 28172
rect 22796 28200 22802 28212
rect 22796 28172 24072 28200
rect 22796 28160 22802 28172
rect 14921 28135 14979 28141
rect 14921 28132 14933 28135
rect 14792 28104 14933 28132
rect 14792 28092 14798 28104
rect 14921 28101 14933 28104
rect 14967 28101 14979 28135
rect 14921 28095 14979 28101
rect 17037 28135 17095 28141
rect 17037 28101 17049 28135
rect 17083 28101 17095 28135
rect 23658 28132 23664 28144
rect 17037 28095 17095 28101
rect 23584 28104 23664 28132
rect 14829 28067 14887 28073
rect 14829 28033 14841 28067
rect 14875 28064 14887 28067
rect 15289 28067 15347 28073
rect 15289 28064 15301 28067
rect 14875 28036 15301 28064
rect 14875 28033 14887 28036
rect 14829 28027 14887 28033
rect 15289 28033 15301 28036
rect 15335 28033 15347 28067
rect 15289 28027 15347 28033
rect 19334 28024 19340 28076
rect 19392 28024 19398 28076
rect 23584 28073 23612 28104
rect 23658 28092 23664 28104
rect 23716 28092 23722 28144
rect 23578 28067 23636 28073
rect 23578 28033 23590 28067
rect 23624 28033 23636 28067
rect 24044 28064 24072 28172
rect 27522 28160 27528 28212
rect 27580 28160 27586 28212
rect 27982 28160 27988 28212
rect 28040 28200 28046 28212
rect 28813 28203 28871 28209
rect 28813 28200 28825 28203
rect 28040 28172 28825 28200
rect 28040 28160 28046 28172
rect 28813 28169 28825 28172
rect 28859 28169 28871 28203
rect 28813 28163 28871 28169
rect 32585 28203 32643 28209
rect 32585 28169 32597 28203
rect 32631 28200 32643 28203
rect 32950 28200 32956 28212
rect 32631 28172 32956 28200
rect 32631 28169 32643 28172
rect 32585 28163 32643 28169
rect 32950 28160 32956 28172
rect 33008 28160 33014 28212
rect 36262 28160 36268 28212
rect 36320 28160 36326 28212
rect 27240 28135 27298 28141
rect 27240 28101 27252 28135
rect 27286 28132 27298 28135
rect 27540 28132 27568 28160
rect 27286 28104 27568 28132
rect 35069 28135 35127 28141
rect 27286 28101 27298 28104
rect 27240 28095 27298 28101
rect 35069 28101 35081 28135
rect 35115 28132 35127 28135
rect 37734 28132 37740 28144
rect 35115 28104 37740 28132
rect 35115 28101 35127 28104
rect 35069 28095 35127 28101
rect 37734 28092 37740 28104
rect 37792 28092 37798 28144
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 24044 28036 24685 28064
rect 23578 28027 23636 28033
rect 24673 28033 24685 28036
rect 24719 28033 24731 28067
rect 24673 28027 24731 28033
rect 26970 28024 26976 28076
rect 27028 28024 27034 28076
rect 28074 28024 28080 28076
rect 28132 28064 28138 28076
rect 28905 28067 28963 28073
rect 28132 28036 28764 28064
rect 28132 28024 28138 28036
rect 6178 27956 6184 28008
rect 6236 27956 6242 28008
rect 7745 27999 7803 28005
rect 7745 27965 7757 27999
rect 7791 27996 7803 27999
rect 8018 27996 8024 28008
rect 7791 27968 8024 27996
rect 7791 27965 7803 27968
rect 7745 27959 7803 27965
rect 8018 27956 8024 27968
rect 8076 27956 8082 28008
rect 9674 27956 9680 28008
rect 9732 27956 9738 28008
rect 10413 27999 10471 28005
rect 10413 27965 10425 27999
rect 10459 27965 10471 27999
rect 10413 27959 10471 27965
rect 4755 27900 5212 27928
rect 8941 27931 8999 27937
rect 4755 27897 4767 27900
rect 4709 27891 4767 27897
rect 8941 27897 8953 27931
rect 8987 27928 8999 27931
rect 10428 27928 10456 27959
rect 10686 27956 10692 28008
rect 10744 27956 10750 28008
rect 11054 27956 11060 28008
rect 11112 27996 11118 28008
rect 11149 27999 11207 28005
rect 11149 27996 11161 27999
rect 11112 27968 11161 27996
rect 11112 27956 11118 27968
rect 11149 27965 11161 27968
rect 11195 27965 11207 27999
rect 11149 27959 11207 27965
rect 11514 27956 11520 28008
rect 11572 27956 11578 28008
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 13814 27996 13820 28008
rect 13679 27968 13820 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 13814 27956 13820 27968
rect 13872 27956 13878 28008
rect 13998 27956 14004 28008
rect 14056 27956 14062 28008
rect 14369 27999 14427 28005
rect 14369 27965 14381 27999
rect 14415 27965 14427 27999
rect 14369 27959 14427 27965
rect 8987 27900 14320 27928
rect 8987 27897 8999 27900
rect 8941 27891 8999 27897
rect 14292 27872 14320 27900
rect 2958 27820 2964 27872
rect 3016 27820 3022 27872
rect 3050 27820 3056 27872
rect 3108 27820 3114 27872
rect 4801 27863 4859 27869
rect 4801 27829 4813 27863
rect 4847 27860 4859 27863
rect 5442 27860 5448 27872
rect 4847 27832 5448 27860
rect 4847 27829 4859 27832
rect 4801 27823 4859 27829
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 9030 27820 9036 27872
rect 9088 27820 9094 27872
rect 10594 27820 10600 27872
rect 10652 27820 10658 27872
rect 12158 27820 12164 27872
rect 12216 27820 12222 27872
rect 12526 27820 12532 27872
rect 12584 27860 12590 27872
rect 12805 27863 12863 27869
rect 12805 27860 12817 27863
rect 12584 27832 12817 27860
rect 12584 27820 12590 27832
rect 12805 27829 12817 27832
rect 12851 27829 12863 27863
rect 12805 27823 12863 27829
rect 12986 27820 12992 27872
rect 13044 27820 13050 27872
rect 13538 27820 13544 27872
rect 13596 27860 13602 27872
rect 13725 27863 13783 27869
rect 13725 27860 13737 27863
rect 13596 27832 13737 27860
rect 13596 27820 13602 27832
rect 13725 27829 13737 27832
rect 13771 27829 13783 27863
rect 13725 27823 13783 27829
rect 14274 27820 14280 27872
rect 14332 27820 14338 27872
rect 14384 27860 14412 27959
rect 15010 27956 15016 28008
rect 15068 27956 15074 28008
rect 15562 27956 15568 28008
rect 15620 27996 15626 28008
rect 15841 27999 15899 28005
rect 15841 27996 15853 27999
rect 15620 27968 15853 27996
rect 15620 27956 15626 27968
rect 15841 27965 15853 27968
rect 15887 27965 15899 27999
rect 15841 27959 15899 27965
rect 18138 27956 18144 28008
rect 18196 27996 18202 28008
rect 18966 27996 18972 28008
rect 18196 27968 18972 27996
rect 18196 27956 18202 27968
rect 18966 27956 18972 27968
rect 19024 27996 19030 28008
rect 19061 27999 19119 28005
rect 19061 27996 19073 27999
rect 19024 27968 19073 27996
rect 19024 27956 19030 27968
rect 19061 27965 19073 27968
rect 19107 27965 19119 27999
rect 20073 27999 20131 28005
rect 20073 27996 20085 27999
rect 19061 27959 19119 27965
rect 19720 27968 20085 27996
rect 19720 27937 19748 27968
rect 20073 27965 20085 27968
rect 20119 27965 20131 27999
rect 20073 27959 20131 27965
rect 23845 27999 23903 28005
rect 23845 27965 23857 27999
rect 23891 27965 23903 27999
rect 23845 27959 23903 27965
rect 19705 27931 19763 27937
rect 19705 27897 19717 27931
rect 19751 27897 19763 27931
rect 19705 27891 19763 27897
rect 14918 27860 14924 27872
rect 14384 27832 14924 27860
rect 14918 27820 14924 27832
rect 14976 27820 14982 27872
rect 20714 27820 20720 27872
rect 20772 27820 20778 27872
rect 22370 27820 22376 27872
rect 22428 27820 22434 27872
rect 23474 27820 23480 27872
rect 23532 27860 23538 27872
rect 23860 27860 23888 27959
rect 24486 27956 24492 28008
rect 24544 27956 24550 28008
rect 26142 27956 26148 28008
rect 26200 27996 26206 28008
rect 26605 27999 26663 28005
rect 26605 27996 26617 27999
rect 26200 27968 26617 27996
rect 26200 27956 26206 27968
rect 26605 27965 26617 27968
rect 26651 27965 26663 27999
rect 26605 27959 26663 27965
rect 28626 27956 28632 28008
rect 28684 27956 28690 28008
rect 28736 27996 28764 28036
rect 28905 28033 28917 28067
rect 28951 28064 28963 28067
rect 28994 28064 29000 28076
rect 28951 28036 29000 28064
rect 28951 28033 28963 28036
rect 28905 28027 28963 28033
rect 28994 28024 29000 28036
rect 29052 28024 29058 28076
rect 29178 28024 29184 28076
rect 29236 28064 29242 28076
rect 31113 28067 31171 28073
rect 31113 28064 31125 28067
rect 29236 28036 31125 28064
rect 29236 28024 29242 28036
rect 31113 28033 31125 28036
rect 31159 28064 31171 28067
rect 32493 28067 32551 28073
rect 31159 28036 32076 28064
rect 31159 28033 31171 28036
rect 31113 28027 31171 28033
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 28736 27968 29929 27996
rect 29917 27965 29929 27968
rect 29963 27965 29975 27999
rect 29917 27959 29975 27965
rect 31941 27999 31999 28005
rect 31941 27965 31953 27999
rect 31987 27965 31999 27999
rect 32048 27996 32076 28036
rect 32493 28033 32505 28067
rect 32539 28064 32551 28067
rect 32582 28064 32588 28076
rect 32539 28036 32588 28064
rect 32539 28033 32551 28036
rect 32493 28027 32551 28033
rect 32582 28024 32588 28036
rect 32640 28024 32646 28076
rect 36078 28024 36084 28076
rect 36136 28064 36142 28076
rect 36357 28067 36415 28073
rect 36357 28064 36369 28067
rect 36136 28036 36369 28064
rect 36136 28024 36142 28036
rect 36357 28033 36369 28036
rect 36403 28033 36415 28067
rect 36357 28027 36415 28033
rect 32677 27999 32735 28005
rect 32677 27996 32689 27999
rect 32048 27968 32689 27996
rect 31941 27959 31999 27965
rect 32677 27965 32689 27968
rect 32723 27965 32735 27999
rect 32677 27959 32735 27965
rect 24670 27888 24676 27940
rect 24728 27928 24734 27940
rect 25593 27931 25651 27937
rect 25593 27928 25605 27931
rect 24728 27900 25605 27928
rect 24728 27888 24734 27900
rect 25593 27897 25605 27900
rect 25639 27897 25651 27931
rect 25593 27891 25651 27897
rect 28350 27888 28356 27940
rect 28408 27888 28414 27940
rect 28718 27888 28724 27940
rect 28776 27928 28782 27940
rect 29365 27931 29423 27937
rect 29365 27928 29377 27931
rect 28776 27900 29377 27928
rect 28776 27888 28782 27900
rect 29365 27897 29377 27900
rect 29411 27897 29423 27931
rect 31956 27928 31984 27959
rect 33226 27956 33232 28008
rect 33284 27996 33290 28008
rect 33505 27999 33563 28005
rect 33505 27996 33517 27999
rect 33284 27968 33517 27996
rect 33284 27956 33290 27968
rect 33505 27965 33517 27968
rect 33551 27965 33563 27999
rect 33505 27959 33563 27965
rect 33778 27956 33784 28008
rect 33836 27956 33842 28008
rect 34514 27956 34520 28008
rect 34572 27956 34578 28008
rect 35253 27999 35311 28005
rect 35253 27965 35265 27999
rect 35299 27996 35311 27999
rect 35342 27996 35348 28008
rect 35299 27968 35348 27996
rect 35299 27965 35311 27968
rect 35253 27959 35311 27965
rect 35342 27956 35348 27968
rect 35400 27956 35406 28008
rect 35894 27956 35900 28008
rect 35952 27996 35958 28008
rect 36173 27999 36231 28005
rect 36173 27996 36185 27999
rect 35952 27968 36185 27996
rect 35952 27956 35958 27968
rect 36173 27965 36185 27968
rect 36219 27996 36231 27999
rect 37001 27999 37059 28005
rect 37001 27996 37013 27999
rect 36219 27968 37013 27996
rect 36219 27965 36231 27968
rect 36173 27959 36231 27965
rect 37001 27965 37013 27968
rect 37047 27965 37059 27999
rect 37001 27959 37059 27965
rect 37829 27999 37887 28005
rect 37829 27965 37841 27999
rect 37875 27965 37887 27999
rect 37829 27959 37887 27965
rect 32125 27931 32183 27937
rect 32125 27928 32137 27931
rect 31956 27900 32137 27928
rect 29365 27891 29423 27897
rect 32125 27897 32137 27900
rect 32171 27897 32183 27931
rect 32125 27891 32183 27897
rect 36725 27931 36783 27937
rect 36725 27897 36737 27931
rect 36771 27928 36783 27931
rect 37844 27928 37872 27959
rect 36771 27900 37872 27928
rect 36771 27897 36783 27900
rect 36725 27891 36783 27897
rect 23532 27832 23888 27860
rect 23937 27863 23995 27869
rect 23532 27820 23538 27832
rect 23937 27829 23949 27863
rect 23983 27860 23995 27863
rect 24026 27860 24032 27872
rect 23983 27832 24032 27860
rect 23983 27829 23995 27832
rect 23937 27823 23995 27829
rect 24026 27820 24032 27832
rect 24084 27820 24090 27872
rect 25314 27820 25320 27872
rect 25372 27820 25378 27872
rect 26050 27820 26056 27872
rect 26108 27820 26114 27872
rect 27706 27820 27712 27872
rect 27764 27860 27770 27872
rect 28368 27860 28396 27888
rect 27764 27832 28396 27860
rect 27764 27820 27770 27832
rect 29270 27820 29276 27872
rect 29328 27820 29334 27872
rect 31297 27863 31355 27869
rect 31297 27829 31309 27863
rect 31343 27860 31355 27863
rect 31386 27860 31392 27872
rect 31343 27832 31392 27860
rect 31343 27829 31355 27832
rect 31297 27823 31355 27829
rect 31386 27820 31392 27832
rect 31444 27820 31450 27872
rect 32950 27820 32956 27872
rect 33008 27820 33014 27872
rect 34330 27820 34336 27872
rect 34388 27820 34394 27872
rect 35802 27820 35808 27872
rect 35860 27820 35866 27872
rect 37277 27863 37335 27869
rect 37277 27829 37289 27863
rect 37323 27860 37335 27863
rect 37366 27860 37372 27872
rect 37323 27832 37372 27860
rect 37323 27829 37335 27832
rect 37277 27823 37335 27829
rect 37366 27820 37372 27832
rect 37424 27820 37430 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2774 27616 2780 27668
rect 2832 27616 2838 27668
rect 5828 27628 6776 27656
rect 4982 27588 4988 27600
rect 3344 27560 4988 27588
rect 3344 27529 3372 27560
rect 4982 27548 4988 27560
rect 5040 27548 5046 27600
rect 5077 27591 5135 27597
rect 5077 27557 5089 27591
rect 5123 27588 5135 27591
rect 5828 27588 5856 27628
rect 5123 27560 5856 27588
rect 5123 27557 5135 27560
rect 5077 27551 5135 27557
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 3329 27523 3387 27529
rect 3329 27520 3341 27523
rect 1995 27492 3341 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 3329 27489 3341 27492
rect 3375 27489 3387 27523
rect 3329 27483 3387 27489
rect 4249 27523 4307 27529
rect 4249 27489 4261 27523
rect 4295 27520 4307 27523
rect 4433 27523 4491 27529
rect 4433 27520 4445 27523
rect 4295 27492 4445 27520
rect 4295 27489 4307 27492
rect 4249 27483 4307 27489
rect 4433 27489 4445 27492
rect 4479 27520 4491 27523
rect 5258 27520 5264 27532
rect 4479 27492 5264 27520
rect 4479 27489 4491 27492
rect 4433 27483 4491 27489
rect 5258 27480 5264 27492
rect 5316 27480 5322 27532
rect 5353 27523 5411 27529
rect 5353 27489 5365 27523
rect 5399 27520 5411 27523
rect 5442 27520 5448 27532
rect 5399 27492 5448 27520
rect 5399 27489 5411 27492
rect 5353 27483 5411 27489
rect 5442 27480 5448 27492
rect 5500 27480 5506 27532
rect 5813 27523 5871 27529
rect 5813 27489 5825 27523
rect 5859 27520 5871 27523
rect 5902 27520 5908 27532
rect 5859 27492 5908 27520
rect 5859 27489 5871 27492
rect 5813 27483 5871 27489
rect 5902 27480 5908 27492
rect 5960 27480 5966 27532
rect 6227 27523 6285 27529
rect 6227 27489 6239 27523
rect 6273 27520 6285 27523
rect 6546 27520 6552 27532
rect 6273 27492 6552 27520
rect 6273 27489 6285 27492
rect 6227 27483 6285 27489
rect 6546 27480 6552 27492
rect 6604 27480 6610 27532
rect 6748 27520 6776 27628
rect 6914 27616 6920 27668
rect 6972 27656 6978 27668
rect 9950 27656 9956 27668
rect 6972 27628 7880 27656
rect 6972 27616 6978 27628
rect 7852 27597 7880 27628
rect 9784 27628 9956 27656
rect 7837 27591 7895 27597
rect 7837 27557 7849 27591
rect 7883 27557 7895 27591
rect 7837 27551 7895 27557
rect 9309 27591 9367 27597
rect 9309 27557 9321 27591
rect 9355 27588 9367 27591
rect 9784 27588 9812 27628
rect 9950 27616 9956 27628
rect 10008 27616 10014 27668
rect 10870 27656 10876 27668
rect 10704 27628 10876 27656
rect 9355 27560 9812 27588
rect 9355 27557 9367 27560
rect 9309 27551 9367 27557
rect 10704 27529 10732 27628
rect 10870 27616 10876 27628
rect 10928 27656 10934 27668
rect 12618 27656 12624 27668
rect 10928 27628 12624 27656
rect 10928 27616 10934 27628
rect 12618 27616 12624 27628
rect 12676 27616 12682 27668
rect 14734 27616 14740 27668
rect 14792 27656 14798 27668
rect 14792 27628 15516 27656
rect 14792 27616 14798 27628
rect 15488 27588 15516 27628
rect 18046 27616 18052 27668
rect 18104 27656 18110 27668
rect 18325 27659 18383 27665
rect 18325 27656 18337 27659
rect 18104 27628 18337 27656
rect 18104 27616 18110 27628
rect 18325 27625 18337 27628
rect 18371 27625 18383 27659
rect 18325 27619 18383 27625
rect 19426 27616 19432 27668
rect 19484 27616 19490 27668
rect 23106 27616 23112 27668
rect 23164 27656 23170 27668
rect 24026 27656 24032 27668
rect 23164 27628 24032 27656
rect 23164 27616 23170 27628
rect 24026 27616 24032 27628
rect 24084 27616 24090 27668
rect 24213 27659 24271 27665
rect 24213 27625 24225 27659
rect 24259 27656 24271 27659
rect 24486 27656 24492 27668
rect 24259 27628 24492 27656
rect 24259 27625 24271 27628
rect 24213 27619 24271 27625
rect 24486 27616 24492 27628
rect 24544 27616 24550 27668
rect 27065 27659 27123 27665
rect 27065 27625 27077 27659
rect 27111 27656 27123 27659
rect 27338 27656 27344 27668
rect 27111 27628 27344 27656
rect 27111 27625 27123 27628
rect 27065 27619 27123 27625
rect 27338 27616 27344 27628
rect 27396 27616 27402 27668
rect 28994 27616 29000 27668
rect 29052 27616 29058 27668
rect 29365 27659 29423 27665
rect 29365 27656 29377 27659
rect 29288 27628 29377 27656
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 11164 27560 14504 27588
rect 15488 27560 17509 27588
rect 7101 27523 7159 27529
rect 7101 27520 7113 27523
rect 6748 27492 7113 27520
rect 7101 27489 7113 27492
rect 7147 27489 7159 27523
rect 7101 27483 7159 27489
rect 10689 27523 10747 27529
rect 10689 27489 10701 27523
rect 10735 27489 10747 27523
rect 10689 27483 10747 27489
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27421 2099 27455
rect 2041 27415 2099 27421
rect 4709 27455 4767 27461
rect 4709 27421 4721 27455
rect 4755 27452 4767 27455
rect 5074 27452 5080 27464
rect 4755 27424 5080 27452
rect 4755 27421 4767 27424
rect 4709 27415 4767 27421
rect 2056 27328 2084 27415
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 5169 27455 5227 27461
rect 5169 27421 5181 27455
rect 5215 27452 5227 27455
rect 5534 27452 5540 27464
rect 5215 27424 5540 27452
rect 5215 27421 5227 27424
rect 5169 27415 5227 27421
rect 5534 27412 5540 27424
rect 5592 27412 5598 27464
rect 6086 27412 6092 27464
rect 6144 27412 6150 27464
rect 6362 27412 6368 27464
rect 6420 27412 6426 27464
rect 8386 27412 8392 27464
rect 8444 27412 8450 27464
rect 10410 27412 10416 27464
rect 10468 27461 10474 27464
rect 10468 27452 10480 27461
rect 10468 27424 10513 27452
rect 10468 27415 10480 27424
rect 10468 27412 10474 27415
rect 2685 27387 2743 27393
rect 2685 27353 2697 27387
rect 2731 27384 2743 27387
rect 3145 27387 3203 27393
rect 3145 27384 3157 27387
rect 2731 27356 3157 27384
rect 2731 27353 2743 27356
rect 2685 27347 2743 27353
rect 3145 27353 3157 27356
rect 3191 27353 3203 27387
rect 3145 27347 3203 27353
rect 9214 27344 9220 27396
rect 9272 27384 9278 27396
rect 11164 27384 11192 27560
rect 11238 27480 11244 27532
rect 11296 27480 11302 27532
rect 11348 27529 11376 27560
rect 11333 27523 11391 27529
rect 11333 27489 11345 27523
rect 11379 27489 11391 27523
rect 13725 27523 13783 27529
rect 13725 27520 13737 27523
rect 11333 27483 11391 27489
rect 13004 27492 13737 27520
rect 12250 27412 12256 27464
rect 12308 27412 12314 27464
rect 12526 27412 12532 27464
rect 12584 27452 12590 27464
rect 13004 27452 13032 27492
rect 13725 27489 13737 27492
rect 13771 27489 13783 27523
rect 13725 27483 13783 27489
rect 12584 27424 13032 27452
rect 12584 27412 12590 27424
rect 13078 27412 13084 27464
rect 13136 27412 13142 27464
rect 13538 27412 13544 27464
rect 13596 27412 13602 27464
rect 14476 27452 14504 27560
rect 17497 27557 17509 27560
rect 17543 27588 17555 27591
rect 19245 27591 19303 27597
rect 17543 27560 18920 27588
rect 17543 27557 17555 27560
rect 17497 27551 17555 27557
rect 15387 27492 15976 27520
rect 15387 27452 15415 27492
rect 14476 27424 15415 27452
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27421 15531 27455
rect 15948 27452 15976 27492
rect 16022 27480 16028 27532
rect 16080 27480 16086 27532
rect 18892 27529 18920 27560
rect 19245 27557 19257 27591
rect 19291 27588 19303 27591
rect 19444 27588 19472 27616
rect 25682 27588 25688 27600
rect 19291 27560 19472 27588
rect 23768 27560 25688 27588
rect 19291 27557 19303 27560
rect 19245 27551 19303 27557
rect 23768 27532 23796 27560
rect 25682 27548 25688 27560
rect 25740 27548 25746 27600
rect 27356 27588 27384 27616
rect 27356 27560 27936 27588
rect 16117 27523 16175 27529
rect 16117 27489 16129 27523
rect 16163 27489 16175 27523
rect 18877 27523 18935 27529
rect 16117 27483 16175 27489
rect 16592 27492 18020 27520
rect 16132 27452 16160 27483
rect 16592 27461 16620 27492
rect 16577 27455 16635 27461
rect 16577 27452 16589 27455
rect 15948 27424 16589 27452
rect 15473 27415 15531 27421
rect 16577 27421 16589 27424
rect 16623 27421 16635 27455
rect 16577 27415 16635 27421
rect 17681 27455 17739 27461
rect 17681 27421 17693 27455
rect 17727 27421 17739 27455
rect 17992 27452 18020 27492
rect 18877 27489 18889 27523
rect 18923 27489 18935 27523
rect 18877 27483 18935 27489
rect 20625 27523 20683 27529
rect 20625 27489 20637 27523
rect 20671 27520 20683 27523
rect 22005 27523 22063 27529
rect 22005 27520 22017 27523
rect 20671 27492 22017 27520
rect 20671 27489 20683 27492
rect 20625 27483 20683 27489
rect 22005 27489 22017 27492
rect 22051 27489 22063 27523
rect 22005 27483 22063 27489
rect 23661 27523 23719 27529
rect 23661 27489 23673 27523
rect 23707 27520 23719 27523
rect 23750 27520 23756 27532
rect 23707 27492 23756 27520
rect 23707 27489 23719 27492
rect 23661 27483 23719 27489
rect 20369 27455 20427 27461
rect 17992 27424 19334 27452
rect 17681 27415 17739 27421
rect 9272 27356 11192 27384
rect 13633 27387 13691 27393
rect 9272 27344 9278 27356
rect 13633 27353 13645 27387
rect 13679 27384 13691 27387
rect 13998 27384 14004 27396
rect 13679 27356 14004 27384
rect 13679 27353 13691 27356
rect 13633 27347 13691 27353
rect 13998 27344 14004 27356
rect 14056 27344 14062 27396
rect 15228 27387 15286 27393
rect 15228 27353 15240 27387
rect 15274 27384 15286 27387
rect 15378 27384 15384 27396
rect 15274 27356 15384 27384
rect 15274 27353 15286 27356
rect 15228 27347 15286 27353
rect 15378 27344 15384 27356
rect 15436 27344 15442 27396
rect 15488 27328 15516 27415
rect 17696 27328 17724 27415
rect 18233 27387 18291 27393
rect 18233 27353 18245 27387
rect 18279 27384 18291 27387
rect 18785 27387 18843 27393
rect 18785 27384 18797 27387
rect 18279 27356 18797 27384
rect 18279 27353 18291 27356
rect 18233 27347 18291 27353
rect 18785 27353 18797 27356
rect 18831 27353 18843 27387
rect 19306 27384 19334 27424
rect 20369 27421 20381 27455
rect 20415 27452 20427 27455
rect 20714 27452 20720 27464
rect 20415 27424 20720 27452
rect 20415 27421 20427 27424
rect 20369 27415 20427 27421
rect 20714 27412 20720 27424
rect 20772 27412 20778 27464
rect 21358 27412 21364 27464
rect 21416 27412 21422 27464
rect 22020 27452 22048 27483
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 23842 27480 23848 27532
rect 23900 27520 23906 27532
rect 24857 27523 24915 27529
rect 24857 27520 24869 27523
rect 23900 27492 24869 27520
rect 23900 27480 23906 27492
rect 24857 27489 24869 27492
rect 24903 27489 24915 27523
rect 24857 27483 24915 27489
rect 25041 27523 25099 27529
rect 25041 27489 25053 27523
rect 25087 27520 25099 27523
rect 25501 27523 25559 27529
rect 25501 27520 25513 27523
rect 25087 27492 25513 27520
rect 25087 27489 25099 27492
rect 25041 27483 25099 27489
rect 25501 27489 25513 27492
rect 25547 27489 25559 27523
rect 25501 27483 25559 27489
rect 22094 27452 22100 27464
rect 22020 27424 22100 27452
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 22272 27455 22330 27461
rect 22272 27421 22284 27455
rect 22318 27452 22330 27455
rect 22830 27452 22836 27464
rect 22318 27424 22836 27452
rect 22318 27421 22330 27424
rect 22272 27415 22330 27421
rect 22830 27412 22836 27424
rect 22888 27412 22894 27464
rect 23290 27412 23296 27464
rect 23348 27452 23354 27464
rect 25406 27452 25412 27464
rect 23348 27424 25412 27452
rect 23348 27412 23354 27424
rect 25406 27412 25412 27424
rect 25464 27412 25470 27464
rect 20901 27387 20959 27393
rect 20901 27384 20913 27387
rect 19306 27356 20913 27384
rect 18785 27347 18843 27353
rect 20901 27353 20913 27356
rect 20947 27384 20959 27387
rect 21266 27384 21272 27396
rect 20947 27356 21272 27384
rect 20947 27353 20959 27356
rect 20901 27347 20959 27353
rect 21266 27344 21272 27356
rect 21324 27344 21330 27396
rect 23845 27387 23903 27393
rect 23845 27384 23857 27387
rect 23216 27356 23857 27384
rect 2038 27276 2044 27328
rect 2096 27276 2102 27328
rect 3237 27319 3295 27325
rect 3237 27285 3249 27319
rect 3283 27316 3295 27319
rect 3694 27316 3700 27328
rect 3283 27288 3700 27316
rect 3283 27285 3295 27288
rect 3237 27279 3295 27285
rect 3694 27276 3700 27288
rect 3752 27316 3758 27328
rect 4617 27319 4675 27325
rect 4617 27316 4629 27319
rect 3752 27288 4629 27316
rect 3752 27276 3758 27288
rect 4617 27285 4629 27288
rect 4663 27285 4675 27319
rect 4617 27279 4675 27285
rect 7006 27276 7012 27328
rect 7064 27276 7070 27328
rect 7650 27276 7656 27328
rect 7708 27316 7714 27328
rect 7745 27319 7803 27325
rect 7745 27316 7757 27319
rect 7708 27288 7757 27316
rect 7708 27276 7714 27288
rect 7745 27285 7757 27288
rect 7791 27285 7803 27319
rect 7745 27279 7803 27285
rect 9398 27276 9404 27328
rect 9456 27316 9462 27328
rect 10410 27316 10416 27328
rect 9456 27288 10416 27316
rect 9456 27276 9462 27288
rect 10410 27276 10416 27288
rect 10468 27276 10474 27328
rect 10778 27276 10784 27328
rect 10836 27276 10842 27328
rect 11146 27276 11152 27328
rect 11204 27276 11210 27328
rect 11606 27276 11612 27328
rect 11664 27276 11670 27328
rect 12437 27319 12495 27325
rect 12437 27285 12449 27319
rect 12483 27316 12495 27319
rect 12710 27316 12716 27328
rect 12483 27288 12716 27316
rect 12483 27285 12495 27288
rect 12437 27279 12495 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 12802 27276 12808 27328
rect 12860 27316 12866 27328
rect 13173 27319 13231 27325
rect 13173 27316 13185 27319
rect 12860 27288 13185 27316
rect 12860 27276 12866 27288
rect 13173 27285 13185 27288
rect 13219 27285 13231 27319
rect 13173 27279 13231 27285
rect 13906 27276 13912 27328
rect 13964 27316 13970 27328
rect 14093 27319 14151 27325
rect 14093 27316 14105 27319
rect 13964 27288 14105 27316
rect 13964 27276 13970 27288
rect 14093 27285 14105 27288
rect 14139 27285 14151 27319
rect 14093 27279 14151 27285
rect 15470 27276 15476 27328
rect 15528 27276 15534 27328
rect 15565 27319 15623 27325
rect 15565 27285 15577 27319
rect 15611 27316 15623 27319
rect 15838 27316 15844 27328
rect 15611 27288 15844 27316
rect 15611 27285 15623 27288
rect 15565 27279 15623 27285
rect 15838 27276 15844 27288
rect 15896 27276 15902 27328
rect 15930 27276 15936 27328
rect 15988 27276 15994 27328
rect 17678 27276 17684 27328
rect 17736 27276 17742 27328
rect 18693 27319 18751 27325
rect 18693 27285 18705 27319
rect 18739 27316 18751 27319
rect 18966 27316 18972 27328
rect 18739 27288 18972 27316
rect 18739 27285 18751 27288
rect 18693 27279 18751 27285
rect 18966 27276 18972 27288
rect 19024 27316 19030 27328
rect 19334 27316 19340 27328
rect 19024 27288 19340 27316
rect 19024 27276 19030 27288
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 21910 27276 21916 27328
rect 21968 27276 21974 27328
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 23216 27316 23244 27356
rect 23845 27353 23857 27356
rect 23891 27384 23903 27387
rect 23891 27356 24992 27384
rect 23891 27353 23903 27356
rect 23845 27347 23903 27353
rect 24964 27328 24992 27356
rect 22336 27288 23244 27316
rect 22336 27276 22342 27288
rect 23382 27276 23388 27328
rect 23440 27276 23446 27328
rect 23750 27276 23756 27328
rect 23808 27276 23814 27328
rect 24394 27276 24400 27328
rect 24452 27276 24458 27328
rect 24762 27276 24768 27328
rect 24820 27276 24826 27328
rect 24946 27276 24952 27328
rect 25004 27276 25010 27328
rect 25516 27316 25544 27483
rect 26970 27480 26976 27532
rect 27028 27480 27034 27532
rect 27157 27523 27215 27529
rect 27157 27489 27169 27523
rect 27203 27520 27215 27523
rect 27706 27520 27712 27532
rect 27203 27492 27712 27520
rect 27203 27489 27215 27492
rect 27157 27483 27215 27489
rect 27706 27480 27712 27492
rect 27764 27480 27770 27532
rect 27798 27480 27804 27532
rect 27856 27480 27862 27532
rect 27908 27520 27936 27560
rect 28902 27548 28908 27600
rect 28960 27588 28966 27600
rect 29178 27588 29184 27600
rect 28960 27560 29184 27588
rect 28960 27548 28966 27560
rect 29178 27548 29184 27560
rect 29236 27548 29242 27600
rect 28194 27523 28252 27529
rect 28194 27520 28206 27523
rect 27908 27492 28206 27520
rect 28194 27489 28206 27492
rect 28240 27489 28252 27523
rect 28194 27483 28252 27489
rect 28353 27523 28411 27529
rect 28353 27489 28365 27523
rect 28399 27520 28411 27523
rect 28534 27520 28540 27532
rect 28399 27492 28540 27520
rect 28399 27489 28411 27492
rect 28353 27483 28411 27489
rect 28534 27480 28540 27492
rect 28592 27520 28598 27532
rect 28994 27520 29000 27532
rect 28592 27492 29000 27520
rect 28592 27480 28598 27492
rect 28994 27480 29000 27492
rect 29052 27520 29058 27532
rect 29288 27520 29316 27628
rect 29365 27625 29377 27628
rect 29411 27656 29423 27659
rect 31570 27656 31576 27668
rect 29411 27628 31576 27656
rect 29411 27625 29423 27628
rect 29365 27619 29423 27625
rect 31570 27616 31576 27628
rect 31628 27616 31634 27668
rect 35894 27656 35900 27668
rect 32876 27628 34284 27656
rect 32677 27591 32735 27597
rect 32677 27557 32689 27591
rect 32723 27588 32735 27591
rect 32723 27560 32812 27588
rect 32723 27557 32735 27560
rect 32677 27551 32735 27557
rect 31297 27523 31355 27529
rect 31297 27520 31309 27523
rect 29052 27492 29316 27520
rect 30576 27492 31309 27520
rect 29052 27480 29058 27492
rect 25685 27455 25743 27461
rect 25685 27421 25697 27455
rect 25731 27452 25743 27455
rect 26988 27452 27016 27480
rect 30576 27464 30604 27492
rect 31297 27489 31309 27492
rect 31343 27489 31355 27523
rect 31297 27483 31355 27489
rect 25731 27424 27016 27452
rect 25731 27421 25743 27424
rect 25685 27415 25743 27421
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27341 27455 27399 27461
rect 27341 27452 27353 27455
rect 27120 27424 27353 27452
rect 27120 27412 27126 27424
rect 27341 27421 27353 27424
rect 27387 27421 27399 27455
rect 27341 27415 27399 27421
rect 28074 27412 28080 27464
rect 28132 27412 28138 27464
rect 29178 27412 29184 27464
rect 29236 27452 29242 27464
rect 30101 27455 30159 27461
rect 30101 27452 30113 27455
rect 29236 27424 30113 27452
rect 29236 27412 29242 27424
rect 30101 27421 30113 27424
rect 30147 27421 30159 27455
rect 30101 27415 30159 27421
rect 30558 27412 30564 27464
rect 30616 27412 30622 27464
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27421 31263 27455
rect 31312 27452 31340 27483
rect 32398 27452 32404 27464
rect 31312 27424 32404 27452
rect 31205 27415 31263 27421
rect 25952 27387 26010 27393
rect 25952 27353 25964 27387
rect 25998 27384 26010 27387
rect 26050 27384 26056 27396
rect 25998 27356 26056 27384
rect 25998 27353 26010 27356
rect 25952 27347 26010 27353
rect 26050 27344 26056 27356
rect 26108 27344 26114 27396
rect 28626 27316 28632 27328
rect 25516 27288 28632 27316
rect 28626 27276 28632 27288
rect 28684 27276 28690 27328
rect 29546 27276 29552 27328
rect 29604 27276 29610 27328
rect 30561 27319 30619 27325
rect 30561 27285 30573 27319
rect 30607 27316 30619 27319
rect 30650 27316 30656 27328
rect 30607 27288 30656 27316
rect 30607 27285 30619 27288
rect 30561 27279 30619 27285
rect 30650 27276 30656 27288
rect 30708 27276 30714 27328
rect 31220 27316 31248 27415
rect 32398 27412 32404 27424
rect 32456 27412 32462 27464
rect 32784 27452 32812 27560
rect 32876 27529 32904 27628
rect 33336 27600 33364 27628
rect 33318 27548 33324 27600
rect 33376 27548 33382 27600
rect 33505 27591 33563 27597
rect 33505 27557 33517 27591
rect 33551 27588 33563 27591
rect 34256 27588 34284 27628
rect 35728 27628 35900 27656
rect 34977 27591 35035 27597
rect 34977 27588 34989 27591
rect 33551 27560 34192 27588
rect 34256 27560 34989 27588
rect 33551 27557 33563 27560
rect 33505 27551 33563 27557
rect 32861 27523 32919 27529
rect 32861 27489 32873 27523
rect 32907 27489 32919 27523
rect 32861 27483 32919 27489
rect 33045 27523 33103 27529
rect 33045 27489 33057 27523
rect 33091 27520 33103 27523
rect 33686 27520 33692 27532
rect 33091 27492 33692 27520
rect 33091 27489 33103 27492
rect 33045 27483 33103 27489
rect 33686 27480 33692 27492
rect 33744 27480 33750 27532
rect 34164 27529 34192 27560
rect 34977 27557 34989 27560
rect 35023 27588 35035 27591
rect 35728 27588 35756 27628
rect 35894 27616 35900 27628
rect 35952 27616 35958 27668
rect 35023 27560 35756 27588
rect 35023 27557 35035 27560
rect 34977 27551 35035 27557
rect 34149 27523 34207 27529
rect 34149 27489 34161 27523
rect 34195 27489 34207 27523
rect 34149 27483 34207 27489
rect 34238 27480 34244 27532
rect 34296 27480 34302 27532
rect 34256 27452 34284 27480
rect 32784 27424 34284 27452
rect 34790 27412 34796 27464
rect 34848 27452 34854 27464
rect 36630 27452 36636 27464
rect 34848 27424 36636 27452
rect 34848 27412 34854 27424
rect 36630 27412 36636 27424
rect 36688 27452 36694 27464
rect 38105 27455 38163 27461
rect 38105 27452 38117 27455
rect 36688 27424 38117 27452
rect 36688 27412 36694 27424
rect 38105 27421 38117 27424
rect 38151 27421 38163 27455
rect 38105 27415 38163 27421
rect 31564 27387 31622 27393
rect 31564 27353 31576 27387
rect 31610 27384 31622 27387
rect 33597 27387 33655 27393
rect 33597 27384 33609 27387
rect 31610 27356 33609 27384
rect 31610 27353 31622 27356
rect 31564 27347 31622 27353
rect 33597 27353 33609 27356
rect 33643 27353 33655 27387
rect 33597 27347 33655 27353
rect 36388 27387 36446 27393
rect 36388 27353 36400 27387
rect 36434 27384 36446 27387
rect 36906 27384 36912 27396
rect 36434 27356 36912 27384
rect 36434 27353 36446 27356
rect 36388 27347 36446 27353
rect 36906 27344 36912 27356
rect 36964 27344 36970 27396
rect 37860 27387 37918 27393
rect 37860 27353 37872 27387
rect 37906 27384 37918 27387
rect 38010 27384 38016 27396
rect 37906 27356 38016 27384
rect 37906 27353 37918 27356
rect 37860 27347 37918 27353
rect 38010 27344 38016 27356
rect 38068 27344 38074 27396
rect 32122 27316 32128 27328
rect 31220 27288 32128 27316
rect 32122 27276 32128 27288
rect 32180 27276 32186 27328
rect 32582 27276 32588 27328
rect 32640 27316 32646 27328
rect 33137 27319 33195 27325
rect 33137 27316 33149 27319
rect 32640 27288 33149 27316
rect 32640 27276 32646 27288
rect 33137 27285 33149 27288
rect 33183 27316 33195 27319
rect 34146 27316 34152 27328
rect 33183 27288 34152 27316
rect 33183 27285 33195 27288
rect 33137 27279 33195 27285
rect 34146 27276 34152 27288
rect 34204 27276 34210 27328
rect 34514 27276 34520 27328
rect 34572 27316 34578 27328
rect 35253 27319 35311 27325
rect 35253 27316 35265 27319
rect 34572 27288 35265 27316
rect 34572 27276 34578 27288
rect 35253 27285 35265 27288
rect 35299 27316 35311 27319
rect 36630 27316 36636 27328
rect 35299 27288 36636 27316
rect 35299 27285 35311 27288
rect 35253 27279 35311 27285
rect 36630 27276 36636 27288
rect 36688 27276 36694 27328
rect 36725 27319 36783 27325
rect 36725 27285 36737 27319
rect 36771 27316 36783 27319
rect 37090 27316 37096 27328
rect 36771 27288 37096 27316
rect 36771 27285 36783 27288
rect 36725 27279 36783 27285
rect 37090 27276 37096 27288
rect 37148 27276 37154 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 3513 27115 3571 27121
rect 3513 27081 3525 27115
rect 3559 27112 3571 27115
rect 3602 27112 3608 27124
rect 3559 27084 3608 27112
rect 3559 27081 3571 27084
rect 3513 27075 3571 27081
rect 3602 27072 3608 27084
rect 3660 27072 3666 27124
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27112 4031 27115
rect 4614 27112 4620 27124
rect 4019 27084 4620 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 4614 27072 4620 27084
rect 4672 27072 4678 27124
rect 6365 27115 6423 27121
rect 6365 27081 6377 27115
rect 6411 27112 6423 27115
rect 6454 27112 6460 27124
rect 6411 27084 6460 27112
rect 6411 27081 6423 27084
rect 6365 27075 6423 27081
rect 6454 27072 6460 27084
rect 6512 27072 6518 27124
rect 9398 27072 9404 27124
rect 9456 27072 9462 27124
rect 9950 27112 9956 27124
rect 9508 27084 9956 27112
rect 2958 27004 2964 27056
rect 3016 27044 3022 27056
rect 3154 27047 3212 27053
rect 3154 27044 3166 27047
rect 3016 27016 3166 27044
rect 3016 27004 3022 27016
rect 3154 27013 3166 27016
rect 3200 27013 3212 27047
rect 5350 27044 5356 27056
rect 3154 27007 3212 27013
rect 3436 27016 5356 27044
rect 3436 26985 3464 27016
rect 5350 27004 5356 27016
rect 5408 27044 5414 27056
rect 6178 27044 6184 27056
rect 5408 27016 6184 27044
rect 5408 27004 5414 27016
rect 6178 27004 6184 27016
rect 6236 27044 6242 27056
rect 8288 27047 8346 27053
rect 6236 27016 7788 27044
rect 6236 27004 6242 27016
rect 3421 26979 3479 26985
rect 3421 26945 3433 26979
rect 3467 26945 3479 26979
rect 3421 26939 3479 26945
rect 2038 26732 2044 26784
rect 2096 26732 2102 26784
rect 2314 26732 2320 26784
rect 2372 26772 2378 26784
rect 3436 26772 3464 26939
rect 3694 26936 3700 26988
rect 3752 26976 3758 26988
rect 3881 26979 3939 26985
rect 3881 26976 3893 26979
rect 3752 26948 3893 26976
rect 3752 26936 3758 26948
rect 3881 26945 3893 26948
rect 3927 26945 3939 26979
rect 3881 26939 3939 26945
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26976 4491 26979
rect 6086 26976 6092 26988
rect 4479 26948 6092 26976
rect 4479 26945 4491 26948
rect 4433 26939 4491 26945
rect 6086 26936 6092 26948
rect 6144 26936 6150 26988
rect 7489 26979 7547 26985
rect 7489 26945 7501 26979
rect 7535 26976 7547 26979
rect 7650 26976 7656 26988
rect 7535 26948 7656 26976
rect 7535 26945 7547 26948
rect 7489 26939 7547 26945
rect 7650 26936 7656 26948
rect 7708 26936 7714 26988
rect 7760 26985 7788 27016
rect 8288 27013 8300 27047
rect 8334 27044 8346 27047
rect 9030 27044 9036 27056
rect 8334 27016 9036 27044
rect 8334 27013 8346 27016
rect 8288 27007 8346 27013
rect 9030 27004 9036 27016
rect 9088 27004 9094 27056
rect 7745 26979 7803 26985
rect 7745 26945 7757 26979
rect 7791 26976 7803 26979
rect 7834 26976 7840 26988
rect 7791 26948 7840 26976
rect 7791 26945 7803 26948
rect 7745 26939 7803 26945
rect 7834 26936 7840 26948
rect 7892 26936 7898 26988
rect 8018 26936 8024 26988
rect 8076 26936 8082 26988
rect 9508 26985 9536 27084
rect 9950 27072 9956 27084
rect 10008 27072 10014 27124
rect 10410 27072 10416 27124
rect 10468 27112 10474 27124
rect 10962 27112 10968 27124
rect 10468 27084 10968 27112
rect 10468 27072 10474 27084
rect 10962 27072 10968 27084
rect 11020 27072 11026 27124
rect 11146 27072 11152 27124
rect 11204 27112 11210 27124
rect 11333 27115 11391 27121
rect 11333 27112 11345 27115
rect 11204 27084 11345 27112
rect 11204 27072 11210 27084
rect 11333 27081 11345 27084
rect 11379 27081 11391 27115
rect 11333 27075 11391 27081
rect 11606 27072 11612 27124
rect 11664 27072 11670 27124
rect 11885 27115 11943 27121
rect 11885 27081 11897 27115
rect 11931 27112 11943 27115
rect 12158 27112 12164 27124
rect 11931 27084 12164 27112
rect 11931 27081 11943 27084
rect 11885 27075 11943 27081
rect 12158 27072 12164 27084
rect 12216 27072 12222 27124
rect 12250 27072 12256 27124
rect 12308 27072 12314 27124
rect 12618 27072 12624 27124
rect 12676 27072 12682 27124
rect 12710 27072 12716 27124
rect 12768 27072 12774 27124
rect 13814 27072 13820 27124
rect 13872 27112 13878 27124
rect 14826 27112 14832 27124
rect 13872 27084 14832 27112
rect 13872 27072 13878 27084
rect 14826 27072 14832 27084
rect 14884 27072 14890 27124
rect 15378 27072 15384 27124
rect 15436 27112 15442 27124
rect 15749 27115 15807 27121
rect 15436 27084 15608 27112
rect 15436 27072 15442 27084
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 10410 26936 10416 26988
rect 10468 26936 10474 26988
rect 10502 26936 10508 26988
rect 10560 26985 10566 26988
rect 10560 26979 10588 26985
rect 10576 26945 10588 26979
rect 10560 26939 10588 26945
rect 10560 26936 10566 26939
rect 3602 26868 3608 26920
rect 3660 26908 3666 26920
rect 4065 26911 4123 26917
rect 4065 26908 4077 26911
rect 3660 26880 4077 26908
rect 3660 26868 3666 26880
rect 4065 26877 4077 26880
rect 4111 26908 4123 26911
rect 4706 26908 4712 26920
rect 4111 26880 4712 26908
rect 4111 26877 4123 26880
rect 4065 26871 4123 26877
rect 4706 26868 4712 26880
rect 4764 26868 4770 26920
rect 9582 26868 9588 26920
rect 9640 26908 9646 26920
rect 9677 26911 9735 26917
rect 9677 26908 9689 26911
rect 9640 26880 9689 26908
rect 9640 26868 9646 26880
rect 9677 26877 9689 26880
rect 9723 26877 9735 26911
rect 9677 26871 9735 26877
rect 9858 26868 9864 26920
rect 9916 26868 9922 26920
rect 10689 26911 10747 26917
rect 10689 26908 10701 26911
rect 10244 26880 10701 26908
rect 9876 26840 9904 26868
rect 10244 26852 10272 26880
rect 10689 26877 10701 26880
rect 10735 26877 10747 26911
rect 10689 26871 10747 26877
rect 11238 26868 11244 26920
rect 11296 26908 11302 26920
rect 11624 26908 11652 27072
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26976 12495 26979
rect 12636 26976 12664 27072
rect 12719 26985 12747 27072
rect 15580 27044 15608 27084
rect 15749 27081 15761 27115
rect 15795 27112 15807 27115
rect 15930 27112 15936 27124
rect 15795 27084 15936 27112
rect 15795 27081 15807 27084
rect 15749 27075 15807 27081
rect 15930 27072 15936 27084
rect 15988 27072 15994 27124
rect 16574 27072 16580 27124
rect 16632 27112 16638 27124
rect 17037 27115 17095 27121
rect 17037 27112 17049 27115
rect 16632 27084 17049 27112
rect 16632 27072 16638 27084
rect 17037 27081 17049 27084
rect 17083 27112 17095 27115
rect 18046 27112 18052 27124
rect 17083 27084 18052 27112
rect 17083 27081 17095 27084
rect 17037 27075 17095 27081
rect 18046 27072 18052 27084
rect 18104 27072 18110 27124
rect 18230 27072 18236 27124
rect 18288 27072 18294 27124
rect 19426 27112 19432 27124
rect 18708 27084 19432 27112
rect 15841 27047 15899 27053
rect 15841 27044 15853 27047
rect 15580 27016 15853 27044
rect 15841 27013 15853 27016
rect 15887 27013 15899 27047
rect 15841 27007 15899 27013
rect 12483 26948 12664 26976
rect 12704 26979 12762 26985
rect 12483 26945 12495 26948
rect 12437 26939 12495 26945
rect 12704 26945 12716 26979
rect 12750 26945 12762 26979
rect 12704 26939 12762 26945
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 11296 26880 11652 26908
rect 11296 26868 11302 26880
rect 11698 26868 11704 26920
rect 11756 26868 11762 26920
rect 11793 26911 11851 26917
rect 11793 26877 11805 26911
rect 11839 26877 11851 26911
rect 11793 26871 11851 26877
rect 10137 26843 10195 26849
rect 10137 26840 10149 26843
rect 9876 26812 10149 26840
rect 10137 26809 10149 26812
rect 10183 26809 10195 26843
rect 10137 26803 10195 26809
rect 10226 26800 10232 26852
rect 10284 26800 10290 26852
rect 11808 26784 11836 26871
rect 13906 26868 13912 26920
rect 13964 26868 13970 26920
rect 2372 26744 3464 26772
rect 2372 26732 2378 26744
rect 10686 26732 10692 26784
rect 10744 26772 10750 26784
rect 11790 26772 11796 26784
rect 10744 26744 11796 26772
rect 10744 26732 10750 26744
rect 11790 26732 11796 26744
rect 11848 26732 11854 26784
rect 13924 26772 13952 26868
rect 14108 26852 14136 26939
rect 14826 26936 14832 26988
rect 14884 26936 14890 26988
rect 14918 26936 14924 26988
rect 14976 26985 14982 26988
rect 14976 26979 15004 26985
rect 14992 26945 15004 26979
rect 16592 26976 16620 27072
rect 18248 27044 18276 27072
rect 18248 27016 18644 27044
rect 14976 26939 15004 26945
rect 15672 26948 16620 26976
rect 18345 26979 18403 26985
rect 14976 26936 14982 26939
rect 14182 26868 14188 26920
rect 14240 26908 14246 26920
rect 15105 26911 15163 26917
rect 15105 26908 15117 26911
rect 14240 26880 15117 26908
rect 14240 26868 14246 26880
rect 15105 26877 15117 26880
rect 15151 26908 15163 26911
rect 15672 26908 15700 26948
rect 18345 26945 18357 26979
rect 18391 26976 18403 26979
rect 18506 26976 18512 26988
rect 18391 26948 18512 26976
rect 18391 26945 18403 26948
rect 18345 26939 18403 26945
rect 18506 26936 18512 26948
rect 18564 26936 18570 26988
rect 18616 26985 18644 27016
rect 18708 26985 18736 27084
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 21082 27072 21088 27124
rect 21140 27072 21146 27124
rect 21358 27072 21364 27124
rect 21416 27112 21422 27124
rect 21821 27115 21879 27121
rect 21821 27112 21833 27115
rect 21416 27084 21833 27112
rect 21416 27072 21422 27084
rect 21821 27081 21833 27084
rect 21867 27081 21879 27115
rect 21821 27075 21879 27081
rect 22278 27072 22284 27124
rect 22336 27072 22342 27124
rect 24489 27115 24547 27121
rect 22388 27084 24440 27112
rect 18601 26979 18659 26985
rect 18601 26945 18613 26979
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18693 26979 18751 26985
rect 18693 26945 18705 26979
rect 18739 26945 18751 26979
rect 18693 26939 18751 26945
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 20533 26979 20591 26985
rect 20533 26945 20545 26979
rect 20579 26976 20591 26979
rect 20993 26979 21051 26985
rect 20993 26976 21005 26979
rect 20579 26948 21005 26976
rect 20579 26945 20591 26948
rect 20533 26939 20591 26945
rect 20993 26945 21005 26948
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 22189 26979 22247 26985
rect 22189 26945 22201 26979
rect 22235 26945 22247 26979
rect 22189 26939 22247 26945
rect 15151 26880 15700 26908
rect 15151 26877 15163 26880
rect 15105 26871 15163 26877
rect 16390 26868 16396 26920
rect 16448 26868 16454 26920
rect 18892 26852 18920 26939
rect 19613 26911 19671 26917
rect 19613 26908 19625 26911
rect 18984 26880 19625 26908
rect 14090 26800 14096 26852
rect 14148 26800 14154 26852
rect 14553 26843 14611 26849
rect 14553 26809 14565 26843
rect 14599 26840 14611 26843
rect 14642 26840 14648 26852
rect 14599 26812 14648 26840
rect 14599 26809 14611 26812
rect 14553 26803 14611 26809
rect 14642 26800 14648 26812
rect 14700 26800 14706 26852
rect 18874 26800 18880 26852
rect 18932 26800 18938 26852
rect 16114 26772 16120 26784
rect 13924 26744 16120 26772
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 17221 26775 17279 26781
rect 17221 26741 17233 26775
rect 17267 26772 17279 26775
rect 17678 26772 17684 26784
rect 17267 26744 17684 26772
rect 17267 26741 17279 26744
rect 17221 26735 17279 26741
rect 17678 26732 17684 26744
rect 17736 26772 17742 26784
rect 18984 26772 19012 26880
rect 19613 26877 19625 26880
rect 19659 26877 19671 26911
rect 19613 26871 19671 26877
rect 19702 26868 19708 26920
rect 19760 26917 19766 26920
rect 19760 26911 19788 26917
rect 19776 26877 19788 26911
rect 19760 26871 19788 26877
rect 19889 26911 19947 26917
rect 19889 26877 19901 26911
rect 19935 26908 19947 26911
rect 20070 26908 20076 26920
rect 19935 26880 20076 26908
rect 19935 26877 19947 26880
rect 19889 26871 19947 26877
rect 19760 26868 19766 26871
rect 20070 26868 20076 26880
rect 20128 26868 20134 26920
rect 21266 26868 21272 26920
rect 21324 26868 21330 26920
rect 19334 26800 19340 26852
rect 19392 26800 19398 26852
rect 17736 26744 19012 26772
rect 17736 26732 17742 26744
rect 20622 26732 20628 26784
rect 20680 26732 20686 26784
rect 22204 26772 22232 26939
rect 22388 26920 22416 27084
rect 24412 27044 24440 27084
rect 24489 27081 24501 27115
rect 24535 27112 24547 27115
rect 24762 27112 24768 27124
rect 24535 27084 24768 27112
rect 24535 27081 24547 27084
rect 24489 27075 24547 27081
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 24949 27115 25007 27121
rect 24949 27081 24961 27115
rect 24995 27112 25007 27115
rect 25314 27112 25320 27124
rect 24995 27084 25320 27112
rect 24995 27081 25007 27084
rect 24949 27075 25007 27081
rect 25314 27072 25320 27084
rect 25372 27072 25378 27124
rect 26053 27115 26111 27121
rect 26053 27081 26065 27115
rect 26099 27112 26111 27115
rect 26142 27112 26148 27124
rect 26099 27084 26148 27112
rect 26099 27081 26111 27084
rect 26053 27075 26111 27081
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 26421 27115 26479 27121
rect 26421 27081 26433 27115
rect 26467 27112 26479 27115
rect 26786 27112 26792 27124
rect 26467 27084 26792 27112
rect 26467 27081 26479 27084
rect 26421 27075 26479 27081
rect 26786 27072 26792 27084
rect 26844 27072 26850 27124
rect 28074 27072 28080 27124
rect 28132 27112 28138 27124
rect 28353 27115 28411 27121
rect 28353 27112 28365 27115
rect 28132 27084 28365 27112
rect 28132 27072 28138 27084
rect 28353 27081 28365 27084
rect 28399 27081 28411 27115
rect 28353 27075 28411 27081
rect 28718 27072 28724 27124
rect 28776 27072 28782 27124
rect 29178 27072 29184 27124
rect 29236 27072 29242 27124
rect 29546 27072 29552 27124
rect 29604 27072 29610 27124
rect 30650 27072 30656 27124
rect 30708 27072 30714 27124
rect 31941 27115 31999 27121
rect 31941 27081 31953 27115
rect 31987 27112 31999 27115
rect 33226 27112 33232 27124
rect 31987 27084 33232 27112
rect 31987 27081 31999 27084
rect 31941 27075 31999 27081
rect 33226 27072 33232 27084
rect 33284 27072 33290 27124
rect 34330 27072 34336 27124
rect 34388 27112 34394 27124
rect 34425 27115 34483 27121
rect 34425 27112 34437 27115
rect 34388 27084 34437 27112
rect 34388 27072 34394 27084
rect 34425 27081 34437 27084
rect 34471 27081 34483 27115
rect 34425 27075 34483 27081
rect 37277 27115 37335 27121
rect 37277 27081 37289 27115
rect 37323 27112 37335 27115
rect 37918 27112 37924 27124
rect 37323 27084 37924 27112
rect 37323 27081 37335 27084
rect 37277 27075 37335 27081
rect 37918 27072 37924 27084
rect 37976 27072 37982 27124
rect 26513 27047 26571 27053
rect 24412 27016 26188 27044
rect 22738 26936 22744 26988
rect 22796 26976 22802 26988
rect 22833 26979 22891 26985
rect 22833 26976 22845 26979
rect 22796 26948 22845 26976
rect 22796 26936 22802 26948
rect 22833 26945 22845 26948
rect 22879 26945 22891 26979
rect 22833 26939 22891 26945
rect 24578 26936 24584 26988
rect 24636 26976 24642 26988
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 24636 26948 25605 26976
rect 24636 26936 24642 26948
rect 25593 26945 25605 26948
rect 25639 26976 25651 26979
rect 26050 26976 26056 26988
rect 25639 26948 26056 26976
rect 25639 26945 25651 26948
rect 25593 26939 25651 26945
rect 26050 26936 26056 26948
rect 26108 26936 26114 26988
rect 22370 26868 22376 26920
rect 22428 26868 22434 26920
rect 22646 26868 22652 26920
rect 22704 26868 22710 26920
rect 23290 26868 23296 26920
rect 23348 26868 23354 26920
rect 23569 26911 23627 26917
rect 23569 26908 23581 26911
rect 23400 26880 23581 26908
rect 23400 26852 23428 26880
rect 23569 26877 23581 26880
rect 23615 26877 23627 26911
rect 23569 26871 23627 26877
rect 23658 26868 23664 26920
rect 23716 26917 23722 26920
rect 23716 26911 23744 26917
rect 23732 26877 23744 26911
rect 23716 26871 23744 26877
rect 23845 26911 23903 26917
rect 23845 26877 23857 26911
rect 23891 26908 23903 26911
rect 24026 26908 24032 26920
rect 23891 26880 24032 26908
rect 23891 26877 23903 26880
rect 23845 26871 23903 26877
rect 23716 26868 23722 26871
rect 24026 26868 24032 26880
rect 24084 26908 24090 26920
rect 24596 26908 24624 26936
rect 24084 26880 24624 26908
rect 24084 26868 24090 26880
rect 24670 26868 24676 26920
rect 24728 26868 24734 26920
rect 24857 26911 24915 26917
rect 24857 26877 24869 26911
rect 24903 26908 24915 26911
rect 24946 26908 24952 26920
rect 24903 26880 24952 26908
rect 24903 26877 24915 26880
rect 24857 26871 24915 26877
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 26160 26908 26188 27016
rect 26513 27013 26525 27047
rect 26559 27044 26571 27047
rect 27240 27047 27298 27053
rect 26559 27016 27200 27044
rect 26559 27013 26571 27016
rect 26513 27007 26571 27013
rect 26970 26936 26976 26988
rect 27028 26936 27034 26988
rect 27172 26976 27200 27016
rect 27240 27013 27252 27047
rect 27286 27044 27298 27047
rect 29564 27044 29592 27072
rect 27286 27016 29592 27044
rect 30668 27044 30696 27072
rect 30806 27047 30864 27053
rect 30806 27044 30818 27047
rect 30668 27016 30818 27044
rect 27286 27013 27298 27016
rect 27240 27007 27298 27013
rect 30806 27013 30818 27016
rect 30852 27013 30864 27047
rect 30806 27007 30864 27013
rect 35336 27047 35394 27053
rect 35336 27013 35348 27047
rect 35382 27044 35394 27047
rect 35802 27044 35808 27056
rect 35382 27016 35808 27044
rect 35382 27013 35394 27016
rect 35336 27007 35394 27013
rect 35802 27004 35808 27016
rect 35860 27004 35866 27056
rect 37734 27004 37740 27056
rect 37792 27004 37798 27056
rect 28813 26979 28871 26985
rect 28813 26976 28825 26979
rect 27172 26948 28825 26976
rect 28813 26945 28825 26948
rect 28859 26976 28871 26979
rect 29086 26976 29092 26988
rect 28859 26948 29092 26976
rect 28859 26945 28871 26948
rect 28813 26939 28871 26945
rect 29086 26936 29092 26948
rect 29144 26976 29150 26988
rect 29454 26976 29460 26988
rect 29144 26948 29460 26976
rect 29144 26936 29150 26948
rect 29454 26936 29460 26948
rect 29512 26976 29518 26988
rect 29549 26979 29607 26985
rect 29549 26976 29561 26979
rect 29512 26948 29561 26976
rect 29512 26936 29518 26948
rect 29549 26945 29561 26948
rect 29595 26945 29607 26979
rect 29549 26939 29607 26945
rect 29638 26936 29644 26988
rect 29696 26936 29702 26988
rect 32766 26936 32772 26988
rect 32824 26936 32830 26988
rect 32928 26979 32986 26985
rect 32928 26945 32940 26979
rect 32974 26976 32986 26979
rect 32974 26945 32996 26976
rect 32928 26939 32996 26945
rect 26510 26908 26516 26920
rect 26160 26880 26516 26908
rect 26510 26868 26516 26880
rect 26568 26908 26574 26920
rect 26605 26911 26663 26917
rect 26605 26908 26617 26911
rect 26568 26880 26617 26908
rect 26568 26868 26574 26880
rect 26605 26877 26617 26880
rect 26651 26877 26663 26911
rect 26605 26871 26663 26877
rect 28629 26911 28687 26917
rect 28629 26877 28641 26911
rect 28675 26908 28687 26911
rect 28902 26908 28908 26920
rect 28675 26880 28908 26908
rect 28675 26877 28687 26880
rect 28629 26871 28687 26877
rect 28902 26868 28908 26880
rect 28960 26868 28966 26920
rect 29365 26911 29423 26917
rect 29365 26908 29377 26911
rect 29012 26880 29377 26908
rect 23382 26800 23388 26852
rect 23440 26800 23446 26852
rect 23842 26772 23848 26784
rect 22204 26744 23848 26772
rect 23842 26732 23848 26744
rect 23900 26732 23906 26784
rect 24688 26772 24716 26868
rect 25038 26800 25044 26852
rect 25096 26840 25102 26852
rect 25317 26843 25375 26849
rect 25317 26840 25329 26843
rect 25096 26812 25329 26840
rect 25096 26800 25102 26812
rect 25317 26809 25329 26812
rect 25363 26809 25375 26843
rect 25317 26803 25375 26809
rect 27706 26772 27712 26784
rect 24688 26744 27712 26772
rect 27706 26732 27712 26744
rect 27764 26772 27770 26784
rect 29012 26772 29040 26880
rect 29365 26877 29377 26880
rect 29411 26908 29423 26911
rect 30282 26908 30288 26920
rect 29411 26880 30288 26908
rect 29411 26877 29423 26880
rect 29365 26871 29423 26877
rect 30282 26868 30288 26880
rect 30340 26868 30346 26920
rect 30561 26911 30619 26917
rect 30561 26877 30573 26911
rect 30607 26877 30619 26911
rect 30561 26871 30619 26877
rect 30576 26784 30604 26871
rect 31570 26868 31576 26920
rect 31628 26908 31634 26920
rect 32784 26908 32812 26936
rect 31628 26880 32812 26908
rect 32968 26908 32996 26939
rect 33042 26936 33048 26988
rect 33100 26936 33106 26988
rect 33965 26979 34023 26985
rect 33965 26945 33977 26979
rect 34011 26976 34023 26979
rect 34238 26976 34244 26988
rect 34011 26948 34244 26976
rect 34011 26945 34023 26948
rect 33965 26939 34023 26945
rect 34238 26936 34244 26948
rect 34296 26936 34302 26988
rect 36078 26936 36084 26988
rect 36136 26976 36142 26988
rect 37645 26979 37703 26985
rect 37645 26976 37657 26979
rect 36136 26948 37657 26976
rect 36136 26936 36142 26948
rect 37645 26945 37657 26948
rect 37691 26976 37703 26979
rect 37918 26976 37924 26988
rect 37691 26948 37924 26976
rect 37691 26945 37703 26948
rect 37645 26939 37703 26945
rect 37918 26936 37924 26948
rect 37976 26936 37982 26988
rect 33226 26908 33232 26920
rect 32968 26880 33232 26908
rect 31628 26868 31634 26880
rect 33226 26868 33232 26880
rect 33284 26868 33290 26920
rect 33778 26868 33784 26920
rect 33836 26868 33842 26920
rect 34517 26911 34575 26917
rect 34517 26908 34529 26911
rect 34256 26880 34529 26908
rect 34256 26852 34284 26880
rect 34517 26877 34529 26880
rect 34563 26877 34575 26911
rect 34517 26871 34575 26877
rect 34698 26868 34704 26920
rect 34756 26868 34762 26920
rect 34790 26868 34796 26920
rect 34848 26908 34854 26920
rect 35069 26911 35127 26917
rect 35069 26908 35081 26911
rect 34848 26880 35081 26908
rect 34848 26868 34854 26880
rect 35069 26877 35081 26880
rect 35115 26877 35127 26911
rect 35069 26871 35127 26877
rect 36262 26868 36268 26920
rect 36320 26908 36326 26920
rect 37829 26911 37887 26917
rect 37829 26908 37841 26911
rect 36320 26880 37841 26908
rect 36320 26868 36326 26880
rect 37829 26877 37841 26880
rect 37875 26908 37887 26911
rect 38289 26911 38347 26917
rect 38289 26908 38301 26911
rect 37875 26880 38301 26908
rect 37875 26877 37887 26880
rect 37829 26871 37887 26877
rect 38289 26877 38301 26880
rect 38335 26877 38347 26911
rect 38289 26871 38347 26877
rect 33321 26843 33379 26849
rect 33321 26809 33333 26843
rect 33367 26840 33379 26843
rect 33594 26840 33600 26852
rect 33367 26812 33600 26840
rect 33367 26809 33379 26812
rect 33321 26803 33379 26809
rect 33594 26800 33600 26812
rect 33652 26800 33658 26852
rect 34238 26800 34244 26852
rect 34296 26800 34302 26852
rect 36449 26843 36507 26849
rect 36449 26809 36461 26843
rect 36495 26840 36507 26843
rect 36495 26812 37320 26840
rect 36495 26809 36507 26812
rect 36449 26803 36507 26809
rect 37292 26784 37320 26812
rect 27764 26744 29040 26772
rect 27764 26732 27770 26744
rect 30006 26732 30012 26784
rect 30064 26732 30070 26784
rect 30558 26732 30564 26784
rect 30616 26732 30622 26784
rect 32125 26775 32183 26781
rect 32125 26741 32137 26775
rect 32171 26772 32183 26775
rect 33226 26772 33232 26784
rect 32171 26744 33232 26772
rect 32171 26741 32183 26744
rect 32125 26735 32183 26741
rect 33226 26732 33232 26744
rect 33284 26732 33290 26784
rect 34057 26775 34115 26781
rect 34057 26741 34069 26775
rect 34103 26772 34115 26775
rect 34514 26772 34520 26784
rect 34103 26744 34520 26772
rect 34103 26741 34115 26744
rect 34057 26735 34115 26741
rect 34514 26732 34520 26744
rect 34572 26732 34578 26784
rect 36538 26732 36544 26784
rect 36596 26772 36602 26784
rect 36725 26775 36783 26781
rect 36725 26772 36737 26775
rect 36596 26744 36737 26772
rect 36596 26732 36602 26744
rect 36725 26741 36737 26744
rect 36771 26741 36783 26775
rect 36725 26735 36783 26741
rect 37274 26732 37280 26784
rect 37332 26732 37338 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 2038 26528 2044 26580
rect 2096 26568 2102 26580
rect 5902 26568 5908 26580
rect 2096 26540 3924 26568
rect 2096 26528 2102 26540
rect 3605 26503 3663 26509
rect 3605 26469 3617 26503
rect 3651 26500 3663 26503
rect 3651 26472 3832 26500
rect 3651 26469 3663 26472
rect 3605 26463 3663 26469
rect 3804 26444 3832 26472
rect 3786 26392 3792 26444
rect 3844 26392 3850 26444
rect 3896 26432 3924 26540
rect 4540 26540 5908 26568
rect 4433 26503 4491 26509
rect 4433 26469 4445 26503
rect 4479 26500 4491 26503
rect 4540 26500 4568 26540
rect 5902 26528 5908 26540
rect 5960 26568 5966 26580
rect 7101 26571 7159 26577
rect 5960 26540 6040 26568
rect 5960 26528 5966 26540
rect 6012 26509 6040 26540
rect 7101 26537 7113 26571
rect 7147 26568 7159 26571
rect 8386 26568 8392 26580
rect 7147 26540 8392 26568
rect 7147 26537 7159 26540
rect 7101 26531 7159 26537
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 9493 26571 9551 26577
rect 9493 26537 9505 26571
rect 9539 26568 9551 26571
rect 9582 26568 9588 26580
rect 9539 26540 9588 26568
rect 9539 26537 9551 26540
rect 9493 26531 9551 26537
rect 9582 26528 9588 26540
rect 9640 26568 9646 26580
rect 11514 26568 11520 26580
rect 9640 26540 11520 26568
rect 9640 26528 9646 26540
rect 11514 26528 11520 26540
rect 11572 26528 11578 26580
rect 12802 26528 12808 26580
rect 12860 26528 12866 26580
rect 13078 26528 13084 26580
rect 13136 26568 13142 26580
rect 13173 26571 13231 26577
rect 13173 26568 13185 26571
rect 13136 26540 13185 26568
rect 13136 26528 13142 26540
rect 13173 26537 13185 26540
rect 13219 26537 13231 26571
rect 13173 26531 13231 26537
rect 14090 26528 14096 26580
rect 14148 26568 14154 26580
rect 15562 26568 15568 26580
rect 14148 26540 15568 26568
rect 14148 26528 14154 26540
rect 15562 26528 15568 26540
rect 15620 26528 15626 26580
rect 17494 26528 17500 26580
rect 17552 26568 17558 26580
rect 17589 26571 17647 26577
rect 17589 26568 17601 26571
rect 17552 26540 17601 26568
rect 17552 26528 17558 26540
rect 17589 26537 17601 26540
rect 17635 26568 17647 26571
rect 19334 26568 19340 26580
rect 17635 26540 19340 26568
rect 17635 26537 17647 26540
rect 17589 26531 17647 26537
rect 19334 26528 19340 26540
rect 19392 26528 19398 26580
rect 22094 26568 22100 26580
rect 21836 26540 22100 26568
rect 4479 26472 4568 26500
rect 5997 26503 6055 26509
rect 4479 26469 4491 26472
rect 4433 26463 4491 26469
rect 5997 26469 6009 26503
rect 6043 26500 6055 26503
rect 8757 26503 8815 26509
rect 8757 26500 8769 26503
rect 6043 26472 8769 26500
rect 6043 26469 6055 26472
rect 5997 26463 6055 26469
rect 8757 26469 8769 26472
rect 8803 26500 8815 26503
rect 9858 26500 9864 26512
rect 8803 26472 9864 26500
rect 8803 26469 8815 26472
rect 8757 26463 8815 26469
rect 9858 26460 9864 26472
rect 9916 26460 9922 26512
rect 11330 26500 11336 26512
rect 10980 26472 11336 26500
rect 4826 26435 4884 26441
rect 4826 26432 4838 26435
rect 3896 26404 4838 26432
rect 4826 26401 4838 26404
rect 4872 26401 4884 26435
rect 4826 26395 4884 26401
rect 4985 26435 5043 26441
rect 4985 26401 4997 26435
rect 5031 26432 5043 26435
rect 5534 26432 5540 26444
rect 5031 26404 5540 26432
rect 5031 26401 5043 26404
rect 4985 26395 5043 26401
rect 5534 26392 5540 26404
rect 5592 26432 5598 26444
rect 6362 26432 6368 26444
rect 5592 26404 6368 26432
rect 5592 26392 5598 26404
rect 6362 26392 6368 26404
rect 6420 26392 6426 26444
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26432 6607 26435
rect 10980 26432 11008 26472
rect 11330 26460 11336 26472
rect 11388 26460 11394 26512
rect 12526 26500 12532 26512
rect 11532 26472 12532 26500
rect 6595 26404 7512 26432
rect 6595 26401 6607 26404
rect 6549 26395 6607 26401
rect 2225 26367 2283 26373
rect 2225 26333 2237 26367
rect 2271 26364 2283 26367
rect 2314 26364 2320 26376
rect 2271 26336 2320 26364
rect 2271 26333 2283 26336
rect 2225 26327 2283 26333
rect 2314 26324 2320 26336
rect 2372 26324 2378 26376
rect 2492 26367 2550 26373
rect 2492 26333 2504 26367
rect 2538 26364 2550 26367
rect 3050 26364 3056 26376
rect 2538 26336 3056 26364
rect 2538 26333 2550 26336
rect 2492 26327 2550 26333
rect 3050 26324 3056 26336
rect 3108 26324 3114 26376
rect 3970 26324 3976 26376
rect 4028 26324 4034 26376
rect 4706 26324 4712 26376
rect 4764 26324 4770 26376
rect 6733 26367 6791 26373
rect 6733 26333 6745 26367
rect 6779 26364 6791 26367
rect 7098 26364 7104 26376
rect 6779 26336 7104 26364
rect 6779 26333 6791 26336
rect 6733 26327 6791 26333
rect 7098 26324 7104 26336
rect 7156 26324 7162 26376
rect 7484 26373 7512 26404
rect 10796 26404 11008 26432
rect 7469 26367 7527 26373
rect 7469 26333 7481 26367
rect 7515 26364 7527 26367
rect 9490 26364 9496 26376
rect 7515 26336 9496 26364
rect 7515 26333 7527 26336
rect 7469 26327 7527 26333
rect 9490 26324 9496 26336
rect 9548 26364 9554 26376
rect 10796 26364 10824 26404
rect 11422 26392 11428 26444
rect 11480 26432 11486 26444
rect 11532 26441 11560 26472
rect 12526 26460 12532 26472
rect 12584 26460 12590 26512
rect 11517 26435 11575 26441
rect 11517 26432 11529 26435
rect 11480 26404 11529 26432
rect 11480 26392 11486 26404
rect 11517 26401 11529 26404
rect 11563 26401 11575 26435
rect 11517 26395 11575 26401
rect 9548 26336 10824 26364
rect 9548 26324 9554 26336
rect 10870 26324 10876 26376
rect 10928 26324 10934 26376
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26364 12587 26367
rect 12820 26364 12848 26528
rect 19061 26503 19119 26509
rect 19061 26469 19073 26503
rect 19107 26469 19119 26503
rect 19061 26463 19119 26469
rect 12986 26392 12992 26444
rect 13044 26432 13050 26444
rect 13633 26435 13691 26441
rect 13633 26432 13645 26435
rect 13044 26404 13645 26432
rect 13044 26392 13050 26404
rect 13633 26401 13645 26404
rect 13679 26401 13691 26435
rect 13633 26395 13691 26401
rect 13725 26435 13783 26441
rect 13725 26401 13737 26435
rect 13771 26401 13783 26435
rect 13725 26395 13783 26401
rect 12575 26336 12848 26364
rect 13740 26364 13768 26395
rect 15470 26392 15476 26444
rect 15528 26432 15534 26444
rect 19076 26432 19104 26463
rect 19426 26432 19432 26444
rect 15528 26404 17724 26432
rect 19076 26404 19432 26432
rect 15528 26392 15534 26404
rect 14734 26364 14740 26376
rect 13740 26336 14740 26364
rect 12575 26333 12587 26336
rect 12529 26327 12587 26333
rect 5810 26296 5816 26308
rect 5460 26268 5816 26296
rect 3694 26188 3700 26240
rect 3752 26228 3758 26240
rect 5460 26228 5488 26268
rect 5810 26256 5816 26268
rect 5868 26296 5874 26308
rect 6641 26299 6699 26305
rect 6641 26296 6653 26299
rect 5868 26268 6653 26296
rect 5868 26256 5874 26268
rect 6641 26265 6653 26268
rect 6687 26265 6699 26299
rect 6641 26259 6699 26265
rect 8754 26256 8760 26308
rect 8812 26296 8818 26308
rect 9309 26299 9367 26305
rect 9309 26296 9321 26299
rect 8812 26268 9321 26296
rect 8812 26256 8818 26268
rect 9309 26265 9321 26268
rect 9355 26296 9367 26299
rect 10226 26296 10232 26308
rect 9355 26268 10232 26296
rect 9355 26265 9367 26268
rect 9309 26259 9367 26265
rect 10226 26256 10232 26268
rect 10284 26256 10290 26308
rect 10628 26299 10686 26305
rect 10628 26265 10640 26299
rect 10674 26296 10686 26299
rect 11238 26296 11244 26308
rect 10674 26268 11244 26296
rect 10674 26265 10686 26268
rect 10628 26259 10686 26265
rect 11238 26256 11244 26268
rect 11296 26256 11302 26308
rect 11790 26296 11796 26308
rect 11532 26268 11796 26296
rect 3752 26200 5488 26228
rect 3752 26188 3758 26200
rect 5626 26188 5632 26240
rect 5684 26188 5690 26240
rect 7650 26188 7656 26240
rect 7708 26228 7714 26240
rect 7745 26231 7803 26237
rect 7745 26228 7757 26231
rect 7708 26200 7757 26228
rect 7708 26188 7714 26200
rect 7745 26197 7757 26200
rect 7791 26197 7803 26231
rect 7745 26191 7803 26197
rect 10962 26188 10968 26240
rect 11020 26188 11026 26240
rect 11146 26188 11152 26240
rect 11204 26228 11210 26240
rect 11333 26231 11391 26237
rect 11333 26228 11345 26231
rect 11204 26200 11345 26228
rect 11204 26188 11210 26200
rect 11333 26197 11345 26200
rect 11379 26197 11391 26231
rect 11333 26191 11391 26197
rect 11425 26231 11483 26237
rect 11425 26197 11437 26231
rect 11471 26228 11483 26231
rect 11532 26228 11560 26268
rect 11790 26256 11796 26268
rect 11848 26256 11854 26308
rect 12253 26299 12311 26305
rect 12253 26296 12265 26299
rect 12211 26268 12265 26296
rect 12253 26265 12265 26268
rect 12299 26296 12311 26299
rect 13740 26296 13768 26336
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 15206 26367 15264 26373
rect 15206 26333 15218 26367
rect 15252 26333 15264 26367
rect 15206 26327 15264 26333
rect 12299 26268 13768 26296
rect 12299 26265 12311 26268
rect 12253 26259 12311 26265
rect 11471 26200 11560 26228
rect 11471 26197 11483 26200
rect 11425 26191 11483 26197
rect 11606 26188 11612 26240
rect 11664 26228 11670 26240
rect 12268 26228 12296 26259
rect 14642 26256 14648 26308
rect 14700 26296 14706 26308
rect 15212 26296 15240 26327
rect 16114 26324 16120 26376
rect 16172 26324 16178 26376
rect 17494 26324 17500 26376
rect 17552 26324 17558 26376
rect 17696 26373 17724 26404
rect 19426 26392 19432 26404
rect 19484 26392 19490 26444
rect 21836 26441 21864 26540
rect 22094 26528 22100 26540
rect 22152 26568 22158 26580
rect 23198 26568 23204 26580
rect 22152 26540 23204 26568
rect 22152 26528 22158 26540
rect 23198 26528 23204 26540
rect 23256 26568 23262 26580
rect 23474 26568 23480 26580
rect 23256 26540 23480 26568
rect 23256 26528 23262 26540
rect 23474 26528 23480 26540
rect 23532 26528 23538 26580
rect 23566 26528 23572 26580
rect 23624 26528 23630 26580
rect 23842 26528 23848 26580
rect 23900 26568 23906 26580
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 23900 26540 24409 26568
rect 23900 26528 23906 26540
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 24397 26531 24455 26537
rect 26510 26528 26516 26580
rect 26568 26528 26574 26580
rect 29181 26571 29239 26577
rect 29181 26537 29193 26571
rect 29227 26568 29239 26571
rect 29638 26568 29644 26580
rect 29227 26540 29644 26568
rect 29227 26537 29239 26540
rect 29181 26531 29239 26537
rect 29638 26528 29644 26540
rect 29696 26528 29702 26580
rect 30282 26528 30288 26580
rect 30340 26568 30346 26580
rect 32585 26571 32643 26577
rect 30340 26540 32444 26568
rect 30340 26528 30346 26540
rect 23293 26503 23351 26509
rect 23293 26469 23305 26503
rect 23339 26500 23351 26503
rect 23584 26500 23612 26528
rect 23339 26472 23612 26500
rect 23676 26472 25728 26500
rect 23339 26469 23351 26472
rect 23293 26463 23351 26469
rect 20625 26435 20683 26441
rect 20625 26401 20637 26435
rect 20671 26432 20683 26435
rect 21821 26435 21879 26441
rect 21821 26432 21833 26435
rect 20671 26404 21833 26432
rect 20671 26401 20683 26404
rect 20625 26395 20683 26401
rect 21821 26401 21833 26404
rect 21867 26401 21879 26435
rect 21821 26395 21879 26401
rect 23382 26392 23388 26444
rect 23440 26432 23446 26444
rect 23676 26432 23704 26472
rect 23440 26404 23704 26432
rect 23937 26435 23995 26441
rect 23440 26392 23446 26404
rect 23937 26401 23949 26435
rect 23983 26432 23995 26435
rect 24210 26432 24216 26444
rect 23983 26404 24216 26432
rect 23983 26401 23995 26404
rect 23937 26395 23995 26401
rect 24210 26392 24216 26404
rect 24268 26392 24274 26444
rect 25700 26441 25728 26472
rect 27062 26460 27068 26512
rect 27120 26460 27126 26512
rect 25685 26435 25743 26441
rect 25685 26401 25697 26435
rect 25731 26401 25743 26435
rect 25685 26395 25743 26401
rect 17681 26367 17739 26373
rect 17681 26333 17693 26367
rect 17727 26364 17739 26367
rect 18230 26364 18236 26376
rect 17727 26336 18236 26364
rect 17727 26333 17739 26336
rect 17681 26327 17739 26333
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 21266 26324 21272 26376
rect 21324 26324 21330 26376
rect 21910 26324 21916 26376
rect 21968 26364 21974 26376
rect 22077 26367 22135 26373
rect 22077 26364 22089 26367
rect 21968 26336 22089 26364
rect 21968 26324 21974 26336
rect 22077 26333 22089 26336
rect 22123 26333 22135 26367
rect 23658 26364 23664 26376
rect 22077 26327 22135 26333
rect 23216 26336 23664 26364
rect 15286 26296 15292 26308
rect 14700 26268 15148 26296
rect 15212 26268 15292 26296
rect 14700 26256 14706 26268
rect 11664 26200 12296 26228
rect 11664 26188 11670 26200
rect 13078 26188 13084 26240
rect 13136 26188 13142 26240
rect 13541 26231 13599 26237
rect 13541 26197 13553 26231
rect 13587 26228 13599 26231
rect 13998 26228 14004 26240
rect 13587 26200 14004 26228
rect 13587 26197 13599 26200
rect 13541 26191 13599 26197
rect 13998 26188 14004 26200
rect 14056 26228 14062 26240
rect 14550 26228 14556 26240
rect 14056 26200 14556 26228
rect 14056 26188 14062 26200
rect 14550 26188 14556 26200
rect 14608 26188 14614 26240
rect 15120 26228 15148 26268
rect 15286 26256 15292 26268
rect 15344 26256 15350 26308
rect 17512 26296 17540 26324
rect 17954 26305 17960 26308
rect 15396 26268 17540 26296
rect 15396 26228 15424 26268
rect 17948 26259 17960 26305
rect 17954 26256 17960 26259
rect 18012 26256 18018 26308
rect 18874 26256 18880 26308
rect 18932 26296 18938 26308
rect 20380 26299 20438 26305
rect 18932 26268 19288 26296
rect 18932 26256 18938 26268
rect 15120 26200 15424 26228
rect 15562 26188 15568 26240
rect 15620 26188 15626 26240
rect 19260 26237 19288 26268
rect 20380 26265 20392 26299
rect 20426 26296 20438 26299
rect 20717 26299 20775 26305
rect 20717 26296 20729 26299
rect 20426 26268 20729 26296
rect 20426 26265 20438 26268
rect 20380 26259 20438 26265
rect 20717 26265 20729 26268
rect 20763 26265 20775 26299
rect 20717 26259 20775 26265
rect 19245 26231 19303 26237
rect 19245 26197 19257 26231
rect 19291 26228 19303 26231
rect 20254 26228 20260 26240
rect 19291 26200 20260 26228
rect 19291 26197 19303 26200
rect 19245 26191 19303 26197
rect 20254 26188 20260 26200
rect 20312 26188 20318 26240
rect 23216 26237 23244 26336
rect 23658 26324 23664 26336
rect 23716 26364 23722 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 23716 26336 24961 26364
rect 23716 26324 23722 26336
rect 24949 26333 24961 26336
rect 24995 26333 25007 26367
rect 27080 26364 27108 26460
rect 28445 26435 28503 26441
rect 28445 26401 28457 26435
rect 28491 26432 28503 26435
rect 30558 26432 30564 26444
rect 28491 26404 30564 26432
rect 28491 26401 28503 26404
rect 28445 26395 28503 26401
rect 30558 26392 30564 26404
rect 30616 26432 30622 26444
rect 31113 26435 31171 26441
rect 31113 26432 31125 26435
rect 30616 26404 31125 26432
rect 30616 26392 30622 26404
rect 31113 26401 31125 26404
rect 31159 26401 31171 26435
rect 31113 26395 31171 26401
rect 28537 26367 28595 26373
rect 28537 26364 28549 26367
rect 27080 26336 28549 26364
rect 24949 26327 25007 26333
rect 28537 26333 28549 26336
rect 28583 26333 28595 26367
rect 28537 26327 28595 26333
rect 28718 26324 28724 26376
rect 28776 26364 28782 26376
rect 28776 26336 29868 26364
rect 28776 26324 28782 26336
rect 23753 26299 23811 26305
rect 23753 26265 23765 26299
rect 23799 26296 23811 26299
rect 25133 26299 25191 26305
rect 25133 26296 25145 26299
rect 23799 26268 25145 26296
rect 23799 26265 23811 26268
rect 23753 26259 23811 26265
rect 25133 26265 25145 26268
rect 25179 26265 25191 26299
rect 25133 26259 25191 26265
rect 25406 26256 25412 26308
rect 25464 26296 25470 26308
rect 26053 26299 26111 26305
rect 26053 26296 26065 26299
rect 25464 26268 26065 26296
rect 25464 26256 25470 26268
rect 26053 26265 26065 26268
rect 26099 26296 26111 26299
rect 26234 26296 26240 26308
rect 26099 26268 26240 26296
rect 26099 26265 26111 26268
rect 26053 26259 26111 26265
rect 26234 26256 26240 26268
rect 26292 26296 26298 26308
rect 26789 26299 26847 26305
rect 26789 26296 26801 26299
rect 26292 26268 26801 26296
rect 26292 26256 26298 26268
rect 26789 26265 26801 26268
rect 26835 26296 26847 26299
rect 27798 26296 27804 26308
rect 26835 26268 27804 26296
rect 26835 26265 26847 26268
rect 26789 26259 26847 26265
rect 27798 26256 27804 26268
rect 27856 26256 27862 26308
rect 28200 26299 28258 26305
rect 28200 26265 28212 26299
rect 28246 26296 28258 26299
rect 29549 26299 29607 26305
rect 29549 26296 29561 26299
rect 28246 26268 29561 26296
rect 28246 26265 28258 26268
rect 28200 26259 28258 26265
rect 29549 26265 29561 26268
rect 29595 26265 29607 26299
rect 29840 26296 29868 26336
rect 30006 26324 30012 26376
rect 30064 26364 30070 26376
rect 31386 26373 31392 26376
rect 30101 26367 30159 26373
rect 30101 26364 30113 26367
rect 30064 26336 30113 26364
rect 30064 26324 30070 26336
rect 30101 26333 30113 26336
rect 30147 26333 30159 26367
rect 31380 26364 31392 26373
rect 31347 26336 31392 26364
rect 30101 26327 30159 26333
rect 31380 26327 31392 26336
rect 31386 26324 31392 26327
rect 31444 26324 31450 26376
rect 30929 26299 30987 26305
rect 30929 26296 30941 26299
rect 29840 26268 30941 26296
rect 29549 26259 29607 26265
rect 30929 26265 30941 26268
rect 30975 26296 30987 26299
rect 32416 26296 32444 26540
rect 32585 26537 32597 26571
rect 32631 26568 32643 26571
rect 33778 26568 33784 26580
rect 32631 26540 33784 26568
rect 32631 26537 32643 26540
rect 32585 26531 32643 26537
rect 33778 26528 33784 26540
rect 33836 26528 33842 26580
rect 34977 26571 35035 26577
rect 34977 26537 34989 26571
rect 35023 26568 35035 26571
rect 35342 26568 35348 26580
rect 35023 26540 35348 26568
rect 35023 26537 35035 26540
rect 34977 26531 35035 26537
rect 35342 26528 35348 26540
rect 35400 26528 35406 26580
rect 35452 26540 37964 26568
rect 32493 26503 32551 26509
rect 32493 26469 32505 26503
rect 32539 26469 32551 26503
rect 32493 26463 32551 26469
rect 32508 26364 32536 26463
rect 33965 26435 34023 26441
rect 33965 26401 33977 26435
rect 34011 26432 34023 26435
rect 34790 26432 34796 26444
rect 34011 26404 34796 26432
rect 34011 26401 34023 26404
rect 33965 26395 34023 26401
rect 34790 26392 34796 26404
rect 34848 26392 34854 26444
rect 33134 26364 33140 26376
rect 32508 26336 33140 26364
rect 33134 26324 33140 26336
rect 33192 26324 33198 26376
rect 34241 26367 34299 26373
rect 34241 26364 34253 26367
rect 33612 26336 34253 26364
rect 33612 26296 33640 26336
rect 34241 26333 34253 26336
rect 34287 26364 34299 26367
rect 34698 26364 34704 26376
rect 34287 26336 34704 26364
rect 34287 26333 34299 26336
rect 34241 26327 34299 26333
rect 34698 26324 34704 26336
rect 34756 26364 34762 26376
rect 35452 26364 35480 26540
rect 37274 26500 37280 26512
rect 36924 26472 37280 26500
rect 35526 26392 35532 26444
rect 35584 26392 35590 26444
rect 36078 26432 36084 26444
rect 35912 26404 36084 26432
rect 35912 26364 35940 26404
rect 36078 26392 36084 26404
rect 36136 26392 36142 26444
rect 36446 26392 36452 26444
rect 36504 26392 36510 26444
rect 36608 26435 36666 26441
rect 36608 26401 36620 26435
rect 36654 26432 36666 26435
rect 36924 26432 36952 26472
rect 37274 26460 37280 26472
rect 37332 26500 37338 26512
rect 37332 26472 37872 26500
rect 37332 26460 37338 26472
rect 36654 26404 36952 26432
rect 36654 26401 36666 26404
rect 36608 26395 36666 26401
rect 36998 26392 37004 26444
rect 37056 26392 37062 26444
rect 37090 26392 37096 26444
rect 37148 26432 37154 26444
rect 37461 26435 37519 26441
rect 37461 26432 37473 26435
rect 37148 26404 37473 26432
rect 37148 26392 37154 26404
rect 37461 26401 37473 26404
rect 37507 26401 37519 26435
rect 37461 26395 37519 26401
rect 37642 26392 37648 26444
rect 37700 26392 37706 26444
rect 37844 26376 37872 26472
rect 37936 26432 37964 26540
rect 38194 26432 38200 26444
rect 37936 26404 38200 26432
rect 38194 26392 38200 26404
rect 38252 26432 38258 26444
rect 38289 26435 38347 26441
rect 38289 26432 38301 26435
rect 38252 26404 38301 26432
rect 38252 26392 38258 26404
rect 38289 26401 38301 26404
rect 38335 26401 38347 26435
rect 38289 26395 38347 26401
rect 34756 26336 35480 26364
rect 35728 26336 35940 26364
rect 34756 26324 34762 26336
rect 30975 26268 32352 26296
rect 32416 26268 33640 26296
rect 33720 26299 33778 26305
rect 30975 26265 30987 26268
rect 30929 26259 30987 26265
rect 23201 26231 23259 26237
rect 23201 26197 23213 26231
rect 23247 26197 23259 26231
rect 23201 26191 23259 26197
rect 23661 26231 23719 26237
rect 23661 26197 23673 26231
rect 23707 26228 23719 26231
rect 24946 26228 24952 26240
rect 23707 26200 24952 26228
rect 23707 26197 23719 26200
rect 23661 26191 23719 26197
rect 24946 26188 24952 26200
rect 25004 26188 25010 26240
rect 32324 26228 32352 26268
rect 33720 26265 33732 26299
rect 33766 26296 33778 26299
rect 33962 26296 33968 26308
rect 33766 26268 33968 26296
rect 33766 26265 33778 26268
rect 33720 26259 33778 26265
rect 33962 26256 33968 26268
rect 34020 26256 34026 26308
rect 35342 26256 35348 26308
rect 35400 26256 35406 26308
rect 35728 26296 35756 26336
rect 36722 26324 36728 26376
rect 36780 26324 36786 26376
rect 37826 26324 37832 26376
rect 37884 26324 37890 26376
rect 37918 26324 37924 26376
rect 37976 26364 37982 26376
rect 37976 26336 38240 26364
rect 37976 26324 37982 26336
rect 35452 26268 35756 26296
rect 35805 26299 35863 26305
rect 33594 26228 33600 26240
rect 32324 26200 33600 26228
rect 33594 26188 33600 26200
rect 33652 26188 33658 26240
rect 35452 26237 35480 26268
rect 35805 26265 35817 26299
rect 35851 26296 35863 26299
rect 35894 26296 35900 26308
rect 35851 26268 35900 26296
rect 35851 26265 35863 26268
rect 35805 26259 35863 26265
rect 35894 26256 35900 26268
rect 35952 26256 35958 26308
rect 38212 26305 38240 26336
rect 38105 26299 38163 26305
rect 38105 26296 38117 26299
rect 37476 26268 38117 26296
rect 35437 26231 35495 26237
rect 35437 26197 35449 26231
rect 35483 26197 35495 26231
rect 35437 26191 35495 26197
rect 37182 26188 37188 26240
rect 37240 26228 37246 26240
rect 37476 26228 37504 26268
rect 38105 26265 38117 26268
rect 38151 26265 38163 26299
rect 38105 26259 38163 26265
rect 38197 26299 38255 26305
rect 38197 26265 38209 26299
rect 38243 26265 38255 26299
rect 38197 26259 38255 26265
rect 37240 26200 37504 26228
rect 37240 26188 37246 26200
rect 37734 26188 37740 26240
rect 37792 26188 37798 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 3421 26027 3479 26033
rect 3421 25993 3433 26027
rect 3467 26024 3479 26027
rect 3467 25996 4016 26024
rect 3467 25993 3479 25996
rect 3421 25987 3479 25993
rect 3988 25968 4016 25996
rect 5626 25984 5632 26036
rect 5684 26024 5690 26036
rect 6733 26027 6791 26033
rect 6733 26024 6745 26027
rect 5684 25996 6745 26024
rect 5684 25984 5690 25996
rect 6733 25993 6745 25996
rect 6779 25993 6791 26027
rect 6733 25987 6791 25993
rect 6825 26027 6883 26033
rect 6825 25993 6837 26027
rect 6871 26024 6883 26027
rect 7006 26024 7012 26036
rect 6871 25996 7012 26024
rect 6871 25993 6883 25996
rect 6825 25987 6883 25993
rect 7006 25984 7012 25996
rect 7064 25984 7070 26036
rect 7469 26027 7527 26033
rect 7469 25993 7481 26027
rect 7515 26024 7527 26027
rect 8110 26024 8116 26036
rect 7515 25996 8116 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 2314 25956 2320 25968
rect 1964 25928 2320 25956
rect 1964 25897 1992 25928
rect 2314 25916 2320 25928
rect 2372 25916 2378 25968
rect 3970 25916 3976 25968
rect 4028 25956 4034 25968
rect 4028 25928 5488 25956
rect 4028 25916 4034 25928
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25857 2007 25891
rect 1949 25851 2007 25857
rect 2038 25848 2044 25900
rect 2096 25888 2102 25900
rect 2205 25891 2263 25897
rect 2205 25888 2217 25891
rect 2096 25860 2217 25888
rect 2096 25848 2102 25860
rect 2205 25857 2217 25860
rect 2251 25857 2263 25891
rect 2205 25851 2263 25857
rect 4545 25891 4603 25897
rect 4545 25857 4557 25891
rect 4591 25888 4603 25891
rect 4706 25888 4712 25900
rect 4591 25860 4712 25888
rect 4591 25857 4603 25860
rect 4545 25851 4603 25857
rect 4706 25848 4712 25860
rect 4764 25848 4770 25900
rect 4801 25891 4859 25897
rect 4801 25857 4813 25891
rect 4847 25888 4859 25891
rect 5350 25888 5356 25900
rect 4847 25860 5356 25888
rect 4847 25857 4859 25860
rect 4801 25851 4859 25857
rect 5350 25848 5356 25860
rect 5408 25848 5414 25900
rect 5460 25897 5488 25928
rect 5445 25891 5503 25897
rect 5445 25857 5457 25891
rect 5491 25857 5503 25891
rect 5445 25851 5503 25857
rect 7009 25823 7067 25829
rect 7009 25789 7021 25823
rect 7055 25820 7067 25823
rect 7484 25820 7512 25987
rect 8110 25984 8116 25996
rect 8168 26024 8174 26036
rect 9214 26024 9220 26036
rect 8168 25996 9220 26024
rect 8168 25984 8174 25996
rect 9214 25984 9220 25996
rect 9272 25984 9278 26036
rect 9674 25984 9680 26036
rect 9732 26024 9738 26036
rect 10229 26027 10287 26033
rect 10229 26024 10241 26027
rect 9732 25996 10241 26024
rect 9732 25984 9738 25996
rect 10229 25993 10241 25996
rect 10275 25993 10287 26027
rect 10229 25987 10287 25993
rect 10594 25984 10600 26036
rect 10652 26024 10658 26036
rect 10689 26027 10747 26033
rect 10689 26024 10701 26027
rect 10652 25996 10701 26024
rect 10652 25984 10658 25996
rect 10689 25993 10701 25996
rect 10735 25993 10747 26027
rect 10689 25987 10747 25993
rect 11146 25984 11152 26036
rect 11204 26024 11210 26036
rect 11517 26027 11575 26033
rect 11517 26024 11529 26027
rect 11204 25996 11529 26024
rect 11204 25984 11210 25996
rect 11517 25993 11529 25996
rect 11563 25993 11575 26027
rect 11517 25987 11575 25993
rect 11698 25984 11704 26036
rect 11756 25984 11762 26036
rect 13078 25984 13084 26036
rect 13136 25984 13142 26036
rect 14829 26027 14887 26033
rect 14829 25993 14841 26027
rect 14875 26024 14887 26027
rect 15562 26024 15568 26036
rect 14875 25996 15568 26024
rect 14875 25993 14887 25996
rect 14829 25987 14887 25993
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 17589 26027 17647 26033
rect 17589 25993 17601 26027
rect 17635 26024 17647 26027
rect 17954 26024 17960 26036
rect 17635 25996 17960 26024
rect 17635 25993 17647 25996
rect 17589 25987 17647 25993
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 20073 26027 20131 26033
rect 20073 25993 20085 26027
rect 20119 26024 20131 26027
rect 21266 26024 21272 26036
rect 20119 25996 21272 26024
rect 20119 25993 20131 25996
rect 20073 25987 20131 25993
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 25682 25984 25688 26036
rect 25740 26024 25746 26036
rect 27157 26027 27215 26033
rect 27157 26024 27169 26027
rect 25740 25996 27169 26024
rect 25740 25984 25746 25996
rect 27157 25993 27169 25996
rect 27203 25993 27215 26027
rect 27157 25987 27215 25993
rect 27341 26027 27399 26033
rect 27341 25993 27353 26027
rect 27387 26024 27399 26027
rect 27430 26024 27436 26036
rect 27387 25996 27436 26024
rect 27387 25993 27399 25996
rect 27341 25987 27399 25993
rect 11238 25916 11244 25968
rect 11296 25956 11302 25968
rect 11716 25956 11744 25984
rect 11296 25928 11744 25956
rect 13096 25956 13124 25984
rect 13326 25959 13384 25965
rect 13326 25956 13338 25959
rect 13096 25928 13338 25956
rect 11296 25916 11302 25928
rect 13326 25925 13338 25928
rect 13372 25925 13384 25959
rect 13326 25919 13384 25925
rect 13538 25916 13544 25968
rect 13596 25916 13602 25968
rect 22956 25959 23014 25965
rect 22956 25925 22968 25959
rect 23002 25956 23014 25959
rect 23106 25956 23112 25968
rect 23002 25928 23112 25956
rect 23002 25925 23014 25928
rect 22956 25919 23014 25925
rect 23106 25916 23112 25928
rect 23164 25916 23170 25968
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 8757 25891 8815 25897
rect 8757 25888 8769 25891
rect 7892 25860 8769 25888
rect 7892 25848 7898 25860
rect 8757 25857 8769 25860
rect 8803 25857 8815 25891
rect 8757 25851 8815 25857
rect 9024 25891 9082 25897
rect 9024 25857 9036 25891
rect 9070 25888 9082 25891
rect 10042 25888 10048 25900
rect 9070 25860 10048 25888
rect 9070 25857 9082 25860
rect 9024 25851 9082 25857
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25888 10655 25891
rect 10686 25888 10692 25900
rect 10643 25860 10692 25888
rect 10643 25857 10655 25860
rect 10597 25851 10655 25857
rect 7055 25792 7512 25820
rect 7055 25789 7067 25792
rect 7009 25783 7067 25789
rect 9766 25780 9772 25832
rect 9824 25820 9830 25832
rect 10612 25820 10640 25851
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25888 13139 25891
rect 13556 25888 13584 25916
rect 13127 25860 13584 25888
rect 13127 25857 13139 25860
rect 13081 25851 13139 25857
rect 14550 25848 14556 25900
rect 14608 25888 14614 25900
rect 14921 25891 14979 25897
rect 14921 25888 14933 25891
rect 14608 25860 14933 25888
rect 14608 25848 14614 25860
rect 14921 25857 14933 25860
rect 14967 25888 14979 25891
rect 15286 25888 15292 25900
rect 14967 25860 15292 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 15672 25860 18184 25888
rect 9824 25792 10640 25820
rect 10873 25823 10931 25829
rect 9824 25780 9830 25792
rect 10873 25789 10885 25823
rect 10919 25820 10931 25823
rect 11146 25820 11152 25832
rect 10919 25792 11152 25820
rect 10919 25789 10931 25792
rect 10873 25783 10931 25789
rect 11146 25780 11152 25792
rect 11204 25820 11210 25832
rect 11606 25820 11612 25832
rect 11204 25792 11612 25820
rect 11204 25780 11210 25792
rect 11606 25780 11612 25792
rect 11664 25780 11670 25832
rect 12069 25823 12127 25829
rect 12069 25789 12081 25823
rect 12115 25789 12127 25823
rect 12069 25783 12127 25789
rect 4798 25712 4804 25764
rect 4856 25712 4862 25764
rect 10137 25755 10195 25761
rect 10137 25721 10149 25755
rect 10183 25752 10195 25755
rect 10502 25752 10508 25764
rect 10183 25724 10508 25752
rect 10183 25721 10195 25724
rect 10137 25715 10195 25721
rect 10502 25712 10508 25724
rect 10560 25752 10566 25764
rect 12084 25752 12112 25783
rect 14274 25780 14280 25832
rect 14332 25820 14338 25832
rect 14734 25820 14740 25832
rect 14332 25792 14740 25820
rect 14332 25780 14338 25792
rect 14734 25780 14740 25792
rect 14792 25820 14798 25832
rect 15672 25820 15700 25860
rect 18156 25832 18184 25860
rect 18690 25848 18696 25900
rect 18748 25848 18754 25900
rect 18785 25891 18843 25897
rect 18785 25857 18797 25891
rect 18831 25888 18843 25891
rect 18966 25888 18972 25900
rect 18831 25860 18972 25888
rect 18831 25857 18843 25860
rect 18785 25851 18843 25857
rect 18966 25848 18972 25860
rect 19024 25888 19030 25900
rect 19705 25891 19763 25897
rect 19024 25860 19656 25888
rect 19024 25848 19030 25860
rect 14792 25792 15700 25820
rect 14792 25780 14798 25792
rect 16390 25780 16396 25832
rect 16448 25780 16454 25832
rect 18138 25780 18144 25832
rect 18196 25780 18202 25832
rect 19628 25829 19656 25860
rect 19705 25857 19717 25891
rect 19751 25888 19763 25891
rect 20165 25891 20223 25897
rect 20165 25888 20177 25891
rect 19751 25860 20177 25888
rect 19751 25857 19763 25860
rect 19705 25851 19763 25857
rect 20165 25857 20177 25860
rect 20211 25857 20223 25891
rect 20165 25851 20223 25857
rect 20254 25848 20260 25900
rect 20312 25888 20318 25900
rect 20717 25891 20775 25897
rect 20717 25888 20729 25891
rect 20312 25860 20729 25888
rect 20312 25848 20318 25860
rect 20717 25857 20729 25860
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25888 23351 25891
rect 23339 25860 24900 25888
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 18233 25823 18291 25829
rect 18233 25789 18245 25823
rect 18279 25820 18291 25823
rect 18877 25823 18935 25829
rect 18279 25792 18368 25820
rect 18279 25789 18291 25792
rect 18233 25783 18291 25789
rect 10560 25724 12112 25752
rect 14461 25755 14519 25761
rect 10560 25712 10566 25724
rect 14461 25721 14473 25755
rect 14507 25752 14519 25755
rect 14918 25752 14924 25764
rect 14507 25724 14924 25752
rect 14507 25721 14519 25724
rect 14461 25715 14519 25721
rect 14918 25712 14924 25724
rect 14976 25712 14982 25764
rect 15289 25755 15347 25761
rect 15289 25721 15301 25755
rect 15335 25752 15347 25755
rect 16408 25752 16436 25780
rect 18340 25761 18368 25792
rect 18877 25789 18889 25823
rect 18923 25789 18935 25823
rect 19429 25823 19487 25829
rect 19429 25820 19441 25823
rect 18877 25783 18935 25789
rect 18984 25792 19441 25820
rect 15335 25724 16436 25752
rect 18325 25755 18383 25761
rect 15335 25721 15347 25724
rect 15289 25715 15347 25721
rect 18325 25721 18337 25755
rect 18371 25721 18383 25755
rect 18325 25715 18383 25721
rect 3329 25687 3387 25693
rect 3329 25653 3341 25687
rect 3375 25684 3387 25687
rect 4816 25684 4844 25712
rect 3375 25656 4844 25684
rect 3375 25653 3387 25656
rect 3329 25647 3387 25653
rect 4890 25644 4896 25696
rect 4948 25644 4954 25696
rect 6086 25644 6092 25696
rect 6144 25644 6150 25696
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6730 25684 6736 25696
rect 6411 25656 6736 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6730 25644 6736 25656
rect 6788 25644 6794 25696
rect 17126 25644 17132 25696
rect 17184 25684 17190 25696
rect 17405 25687 17463 25693
rect 17405 25684 17417 25687
rect 17184 25656 17417 25684
rect 17184 25644 17190 25656
rect 17405 25653 17417 25656
rect 17451 25684 17463 25687
rect 18892 25684 18920 25783
rect 18984 25764 19012 25792
rect 19429 25789 19441 25792
rect 19475 25789 19487 25823
rect 19429 25783 19487 25789
rect 19613 25823 19671 25829
rect 19613 25789 19625 25823
rect 19659 25820 19671 25823
rect 19659 25792 20300 25820
rect 19659 25789 19671 25792
rect 19613 25783 19671 25789
rect 20272 25764 20300 25792
rect 23198 25780 23204 25832
rect 23256 25820 23262 25832
rect 23256 25792 24808 25820
rect 23256 25780 23262 25792
rect 18966 25712 18972 25764
rect 19024 25712 19030 25764
rect 20254 25712 20260 25764
rect 20312 25712 20318 25764
rect 24780 25696 24808 25792
rect 24872 25696 24900 25860
rect 27172 25820 27200 25987
rect 27430 25984 27436 25996
rect 27488 25984 27494 26036
rect 27801 26027 27859 26033
rect 27801 25993 27813 26027
rect 27847 26024 27859 26027
rect 28258 26024 28264 26036
rect 27847 25996 28264 26024
rect 27847 25993 27859 25996
rect 27801 25987 27859 25993
rect 28258 25984 28264 25996
rect 28316 25984 28322 26036
rect 28442 25984 28448 26036
rect 28500 26024 28506 26036
rect 28902 26024 28908 26036
rect 28500 25996 28908 26024
rect 28500 25984 28506 25996
rect 28902 25984 28908 25996
rect 28960 25984 28966 26036
rect 31570 25984 31576 26036
rect 31628 25984 31634 26036
rect 32122 25984 32128 26036
rect 32180 25984 32186 26036
rect 32493 26027 32551 26033
rect 32493 25993 32505 26027
rect 32539 26024 32551 26027
rect 32950 26024 32956 26036
rect 32539 25996 32956 26024
rect 32539 25993 32551 25996
rect 32493 25987 32551 25993
rect 32950 25984 32956 25996
rect 33008 25984 33014 26036
rect 33226 25984 33232 26036
rect 33284 26024 33290 26036
rect 33321 26027 33379 26033
rect 33321 26024 33333 26027
rect 33284 25996 33333 26024
rect 33284 25984 33290 25996
rect 33321 25993 33333 25996
rect 33367 25993 33379 26027
rect 33321 25987 33379 25993
rect 33594 25984 33600 26036
rect 33652 25984 33658 26036
rect 33962 25984 33968 26036
rect 34020 25984 34026 26036
rect 35342 25984 35348 26036
rect 35400 26024 35406 26036
rect 37277 26027 37335 26033
rect 37277 26024 37289 26027
rect 35400 25996 37289 26024
rect 35400 25984 35406 25996
rect 37277 25993 37289 25996
rect 37323 25993 37335 26027
rect 37277 25987 37335 25993
rect 38194 25984 38200 26036
rect 38252 25984 38258 26036
rect 28626 25916 28632 25968
rect 28684 25956 28690 25968
rect 28684 25928 31524 25956
rect 28684 25916 28690 25928
rect 27709 25891 27767 25897
rect 27709 25857 27721 25891
rect 27755 25888 27767 25891
rect 29086 25888 29092 25900
rect 27755 25860 29092 25888
rect 27755 25857 27767 25860
rect 27709 25851 27767 25857
rect 29086 25848 29092 25860
rect 29144 25848 29150 25900
rect 31496 25888 31524 25928
rect 32582 25916 32588 25968
rect 32640 25916 32646 25968
rect 33612 25956 33640 25984
rect 35434 25956 35440 25968
rect 33612 25928 35440 25956
rect 35434 25916 35440 25928
rect 35492 25956 35498 25968
rect 35888 25959 35946 25965
rect 35492 25928 35848 25956
rect 35492 25916 35498 25928
rect 32858 25888 32864 25900
rect 31496 25860 32864 25888
rect 32858 25848 32864 25860
rect 32916 25888 32922 25900
rect 32916 25860 33088 25888
rect 32916 25848 32922 25860
rect 27614 25820 27620 25832
rect 27172 25792 27620 25820
rect 27614 25780 27620 25792
rect 27672 25820 27678 25832
rect 33060 25829 33088 25860
rect 34514 25848 34520 25900
rect 34572 25848 34578 25900
rect 34790 25848 34796 25900
rect 34848 25888 34854 25900
rect 35621 25891 35679 25897
rect 35621 25888 35633 25891
rect 34848 25860 35633 25888
rect 34848 25848 34854 25860
rect 35621 25857 35633 25860
rect 35667 25857 35679 25891
rect 35820 25888 35848 25928
rect 35888 25925 35900 25959
rect 35934 25956 35946 25959
rect 37366 25956 37372 25968
rect 35934 25928 37372 25956
rect 35934 25925 35946 25928
rect 35888 25919 35946 25925
rect 37366 25916 37372 25928
rect 37424 25916 37430 25968
rect 36814 25888 36820 25900
rect 35820 25860 36820 25888
rect 35621 25851 35679 25857
rect 36814 25848 36820 25860
rect 36872 25888 36878 25900
rect 36998 25888 37004 25900
rect 36872 25860 37004 25888
rect 36872 25848 36878 25860
rect 36998 25848 37004 25860
rect 37056 25848 37062 25900
rect 37826 25848 37832 25900
rect 37884 25848 37890 25900
rect 27893 25823 27951 25829
rect 27893 25820 27905 25823
rect 27672 25792 27905 25820
rect 27672 25780 27678 25792
rect 27893 25789 27905 25792
rect 27939 25789 27951 25823
rect 27893 25783 27951 25789
rect 32677 25823 32735 25829
rect 32677 25789 32689 25823
rect 32723 25789 32735 25823
rect 32677 25783 32735 25789
rect 33045 25823 33103 25829
rect 33045 25789 33057 25823
rect 33091 25789 33103 25823
rect 33045 25783 33103 25789
rect 33229 25823 33287 25829
rect 33229 25789 33241 25823
rect 33275 25820 33287 25823
rect 33410 25820 33416 25832
rect 33275 25792 33416 25820
rect 33275 25789 33287 25792
rect 33229 25783 33287 25789
rect 32692 25752 32720 25783
rect 33410 25780 33416 25792
rect 33468 25780 33474 25832
rect 37642 25780 37648 25832
rect 37700 25780 37706 25832
rect 34885 25755 34943 25761
rect 34885 25752 34897 25755
rect 31956 25724 34897 25752
rect 31956 25696 31984 25724
rect 34885 25721 34897 25724
rect 34931 25752 34943 25755
rect 35526 25752 35532 25764
rect 34931 25724 35532 25752
rect 34931 25721 34943 25724
rect 34885 25715 34943 25721
rect 35526 25712 35532 25724
rect 35584 25712 35590 25764
rect 37001 25755 37059 25761
rect 37001 25721 37013 25755
rect 37047 25752 37059 25755
rect 37660 25752 37688 25780
rect 37047 25724 37688 25752
rect 37047 25721 37059 25724
rect 37001 25715 37059 25721
rect 17451 25656 18920 25684
rect 21821 25687 21879 25693
rect 17451 25653 17463 25656
rect 17405 25647 17463 25653
rect 21821 25653 21833 25687
rect 21867 25684 21879 25687
rect 22554 25684 22560 25696
rect 21867 25656 22560 25684
rect 21867 25653 21879 25656
rect 21821 25647 21879 25653
rect 22554 25644 22560 25656
rect 22612 25644 22618 25696
rect 24762 25644 24768 25696
rect 24820 25644 24826 25696
rect 24854 25644 24860 25696
rect 24912 25684 24918 25696
rect 25317 25687 25375 25693
rect 25317 25684 25329 25687
rect 24912 25656 25329 25684
rect 24912 25644 24918 25656
rect 25317 25653 25329 25656
rect 25363 25684 25375 25687
rect 26418 25684 26424 25696
rect 25363 25656 26424 25684
rect 25363 25653 25375 25656
rect 25317 25647 25375 25653
rect 26418 25644 26424 25656
rect 26476 25644 26482 25696
rect 31938 25644 31944 25696
rect 31996 25644 32002 25696
rect 33686 25644 33692 25696
rect 33744 25644 33750 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2038 25440 2044 25492
rect 2096 25440 2102 25492
rect 4890 25480 4896 25492
rect 4356 25452 4896 25480
rect 2777 25415 2835 25421
rect 2777 25381 2789 25415
rect 2823 25381 2835 25415
rect 2777 25375 2835 25381
rect 2685 25347 2743 25353
rect 2685 25313 2697 25347
rect 2731 25344 2743 25347
rect 2792 25344 2820 25375
rect 3970 25372 3976 25424
rect 4028 25372 4034 25424
rect 2731 25316 2820 25344
rect 3421 25347 3479 25353
rect 2731 25313 2743 25316
rect 2685 25307 2743 25313
rect 3421 25313 3433 25347
rect 3467 25344 3479 25347
rect 3878 25344 3884 25356
rect 3467 25316 3884 25344
rect 3467 25313 3479 25316
rect 3421 25307 3479 25313
rect 3878 25304 3884 25316
rect 3936 25304 3942 25356
rect 4356 25285 4384 25452
rect 4890 25440 4896 25452
rect 4948 25440 4954 25492
rect 5534 25440 5540 25492
rect 5592 25480 5598 25492
rect 5813 25483 5871 25489
rect 5813 25480 5825 25483
rect 5592 25452 5825 25480
rect 5592 25440 5598 25452
rect 5813 25449 5825 25452
rect 5859 25480 5871 25483
rect 7650 25480 7656 25492
rect 5859 25452 7656 25480
rect 5859 25449 5871 25452
rect 5813 25443 5871 25449
rect 7650 25440 7656 25452
rect 7708 25440 7714 25492
rect 10042 25440 10048 25492
rect 10100 25440 10106 25492
rect 14182 25480 14188 25492
rect 13832 25452 14188 25480
rect 5074 25412 5080 25424
rect 4632 25384 5080 25412
rect 4632 25353 4660 25384
rect 5074 25372 5080 25384
rect 5132 25412 5138 25424
rect 13832 25421 13860 25452
rect 14182 25440 14188 25452
rect 14240 25440 14246 25492
rect 14458 25440 14464 25492
rect 14516 25480 14522 25492
rect 14734 25480 14740 25492
rect 14516 25452 14740 25480
rect 14516 25440 14522 25452
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 15010 25440 15016 25492
rect 15068 25480 15074 25492
rect 15068 25452 18000 25480
rect 15068 25440 15074 25452
rect 13817 25415 13875 25421
rect 5132 25384 11284 25412
rect 5132 25372 5138 25384
rect 11256 25356 11284 25384
rect 13817 25381 13829 25415
rect 13863 25381 13875 25415
rect 17972 25412 18000 25452
rect 18690 25440 18696 25492
rect 18748 25480 18754 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 18748 25452 19257 25480
rect 18748 25440 18754 25452
rect 19245 25449 19257 25452
rect 19291 25449 19303 25483
rect 19245 25443 19303 25449
rect 23569 25483 23627 25489
rect 23569 25449 23581 25483
rect 23615 25480 23627 25483
rect 23750 25480 23756 25492
rect 23615 25452 23756 25480
rect 23615 25449 23627 25452
rect 23569 25443 23627 25449
rect 23750 25440 23756 25452
rect 23808 25440 23814 25492
rect 24210 25440 24216 25492
rect 24268 25480 24274 25492
rect 24673 25483 24731 25489
rect 24673 25480 24685 25483
rect 24268 25452 24685 25480
rect 24268 25440 24274 25452
rect 24673 25449 24685 25452
rect 24719 25480 24731 25483
rect 25222 25480 25228 25492
rect 24719 25452 25228 25480
rect 24719 25449 24731 25452
rect 24673 25443 24731 25449
rect 25222 25440 25228 25452
rect 25280 25480 25286 25492
rect 28442 25480 28448 25492
rect 25280 25452 28448 25480
rect 25280 25440 25286 25452
rect 28442 25440 28448 25452
rect 28500 25440 28506 25492
rect 32858 25440 32864 25492
rect 32916 25480 32922 25492
rect 35069 25483 35127 25489
rect 35069 25480 35081 25483
rect 32916 25452 35081 25480
rect 32916 25440 32922 25452
rect 35069 25449 35081 25452
rect 35115 25449 35127 25483
rect 35069 25443 35127 25449
rect 18966 25412 18972 25424
rect 17972 25384 18972 25412
rect 13817 25375 13875 25381
rect 18966 25372 18972 25384
rect 19024 25372 19030 25424
rect 4617 25347 4675 25353
rect 4617 25313 4629 25347
rect 4663 25313 4675 25347
rect 4617 25307 4675 25313
rect 4798 25304 4804 25356
rect 4856 25344 4862 25356
rect 5353 25347 5411 25353
rect 5353 25344 5365 25347
rect 4856 25316 5365 25344
rect 4856 25304 4862 25316
rect 5353 25313 5365 25316
rect 5399 25313 5411 25347
rect 5353 25307 5411 25313
rect 10689 25347 10747 25353
rect 10689 25313 10701 25347
rect 10735 25344 10747 25347
rect 10962 25344 10968 25356
rect 10735 25316 10968 25344
rect 10735 25313 10747 25316
rect 10689 25307 10747 25313
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11238 25304 11244 25356
rect 11296 25304 11302 25356
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 19797 25347 19855 25353
rect 19797 25344 19809 25347
rect 19484 25316 19809 25344
rect 19484 25304 19490 25316
rect 19797 25313 19809 25316
rect 19843 25313 19855 25347
rect 19797 25307 19855 25313
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 22925 25347 22983 25353
rect 22925 25344 22937 25347
rect 22704 25316 22937 25344
rect 22704 25304 22710 25316
rect 22925 25313 22937 25316
rect 22971 25313 22983 25347
rect 22925 25307 22983 25313
rect 23934 25304 23940 25356
rect 23992 25344 23998 25356
rect 29365 25347 29423 25353
rect 29365 25344 29377 25347
rect 23992 25316 29377 25344
rect 23992 25304 23998 25316
rect 29365 25313 29377 25316
rect 29411 25344 29423 25347
rect 29638 25344 29644 25356
rect 29411 25316 29644 25344
rect 29411 25313 29423 25316
rect 29365 25307 29423 25313
rect 29638 25304 29644 25316
rect 29696 25344 29702 25356
rect 30742 25344 30748 25356
rect 29696 25316 30748 25344
rect 29696 25304 29702 25316
rect 30742 25304 30748 25316
rect 30800 25304 30806 25356
rect 4341 25279 4399 25285
rect 4341 25245 4353 25279
rect 4387 25245 4399 25279
rect 4341 25239 4399 25245
rect 7006 25236 7012 25288
rect 7064 25236 7070 25288
rect 8386 25236 8392 25288
rect 8444 25236 8450 25288
rect 13262 25236 13268 25288
rect 13320 25236 13326 25288
rect 16758 25236 16764 25288
rect 16816 25276 16822 25288
rect 16945 25279 17003 25285
rect 16945 25276 16957 25279
rect 16816 25248 16957 25276
rect 16816 25236 16822 25248
rect 16945 25245 16957 25248
rect 16991 25245 17003 25279
rect 16945 25239 17003 25245
rect 18046 25236 18052 25288
rect 18104 25236 18110 25288
rect 26418 25236 26424 25288
rect 26476 25236 26482 25288
rect 28997 25279 29055 25285
rect 28997 25245 29009 25279
rect 29043 25276 29055 25279
rect 29270 25276 29276 25288
rect 29043 25248 29276 25276
rect 29043 25245 29055 25248
rect 28997 25239 29055 25245
rect 29270 25236 29276 25248
rect 29328 25236 29334 25288
rect 30190 25236 30196 25288
rect 30248 25236 30254 25288
rect 35084 25276 35112 25443
rect 35434 25440 35440 25492
rect 35492 25440 35498 25492
rect 36265 25483 36323 25489
rect 36265 25449 36277 25483
rect 36311 25480 36323 25483
rect 37182 25480 37188 25492
rect 36311 25452 37188 25480
rect 36311 25449 36323 25452
rect 36265 25443 36323 25449
rect 37182 25440 37188 25452
rect 37240 25440 37246 25492
rect 38010 25440 38016 25492
rect 38068 25440 38074 25492
rect 37090 25412 37096 25424
rect 35728 25384 37096 25412
rect 35728 25353 35756 25384
rect 37090 25372 37096 25384
rect 37148 25372 37154 25424
rect 35713 25347 35771 25353
rect 35713 25313 35725 25347
rect 35759 25313 35771 25347
rect 36449 25347 36507 25353
rect 36449 25344 36461 25347
rect 35713 25307 35771 25313
rect 35811 25316 36461 25344
rect 35811 25276 35839 25316
rect 36449 25313 36461 25316
rect 36495 25313 36507 25347
rect 36449 25307 36507 25313
rect 37461 25347 37519 25353
rect 37461 25313 37473 25347
rect 37507 25344 37519 25347
rect 37734 25344 37740 25356
rect 37507 25316 37740 25344
rect 37507 25313 37519 25316
rect 37461 25307 37519 25313
rect 37734 25304 37740 25316
rect 37792 25304 37798 25356
rect 35084 25248 35839 25276
rect 35894 25236 35900 25288
rect 35952 25276 35958 25288
rect 36725 25279 36783 25285
rect 36725 25276 36737 25279
rect 35952 25248 36737 25276
rect 35952 25236 35958 25248
rect 36725 25245 36737 25248
rect 36771 25245 36783 25279
rect 36725 25239 36783 25245
rect 3237 25211 3295 25217
rect 3237 25177 3249 25211
rect 3283 25208 3295 25211
rect 4801 25211 4859 25217
rect 4801 25208 4813 25211
rect 3283 25180 4813 25208
rect 3283 25177 3295 25180
rect 3237 25171 3295 25177
rect 4801 25177 4813 25180
rect 4847 25177 4859 25211
rect 4801 25171 4859 25177
rect 9953 25211 10011 25217
rect 9953 25177 9965 25211
rect 9999 25208 10011 25211
rect 11146 25208 11152 25220
rect 9999 25180 11152 25208
rect 9999 25177 10011 25180
rect 9953 25171 10011 25177
rect 11146 25168 11152 25180
rect 11204 25168 11210 25220
rect 35710 25168 35716 25220
rect 35768 25208 35774 25220
rect 36633 25211 36691 25217
rect 36633 25208 36645 25211
rect 35768 25180 36645 25208
rect 35768 25168 35774 25180
rect 36633 25177 36645 25180
rect 36679 25177 36691 25211
rect 36633 25171 36691 25177
rect 3145 25143 3203 25149
rect 3145 25109 3157 25143
rect 3191 25140 3203 25143
rect 3694 25140 3700 25152
rect 3191 25112 3700 25140
rect 3191 25109 3203 25112
rect 3145 25103 3203 25109
rect 3694 25100 3700 25112
rect 3752 25140 3758 25152
rect 4433 25143 4491 25149
rect 4433 25140 4445 25143
rect 3752 25112 4445 25140
rect 3752 25100 3758 25112
rect 4433 25109 4445 25112
rect 4479 25140 4491 25143
rect 4890 25140 4896 25152
rect 4479 25112 4896 25140
rect 4479 25109 4491 25112
rect 4433 25103 4491 25109
rect 4890 25100 4896 25112
rect 4948 25100 4954 25152
rect 7558 25100 7564 25152
rect 7616 25100 7622 25152
rect 7742 25100 7748 25152
rect 7800 25100 7806 25152
rect 11057 25143 11115 25149
rect 11057 25109 11069 25143
rect 11103 25140 11115 25143
rect 11422 25140 11428 25152
rect 11103 25112 11428 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11422 25100 11428 25112
rect 11480 25100 11486 25152
rect 12710 25100 12716 25152
rect 12768 25100 12774 25152
rect 16390 25100 16396 25152
rect 16448 25100 16454 25152
rect 18601 25143 18659 25149
rect 18601 25109 18613 25143
rect 18647 25140 18659 25143
rect 18690 25140 18696 25152
rect 18647 25112 18696 25140
rect 18647 25109 18659 25112
rect 18601 25103 18659 25109
rect 18690 25100 18696 25112
rect 18748 25100 18754 25152
rect 25682 25100 25688 25152
rect 25740 25140 25746 25152
rect 25777 25143 25835 25149
rect 25777 25140 25789 25143
rect 25740 25112 25789 25140
rect 25740 25100 25746 25112
rect 25777 25109 25789 25112
rect 25823 25109 25835 25143
rect 25777 25103 25835 25109
rect 29546 25100 29552 25152
rect 29604 25100 29610 25152
rect 37093 25143 37151 25149
rect 37093 25109 37105 25143
rect 37139 25140 37151 25143
rect 38286 25140 38292 25152
rect 37139 25112 38292 25140
rect 37139 25109 37151 25112
rect 37093 25103 37151 25109
rect 38286 25100 38292 25112
rect 38344 25100 38350 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 4525 24939 4583 24945
rect 4525 24905 4537 24939
rect 4571 24936 4583 24939
rect 4706 24936 4712 24948
rect 4571 24908 4712 24936
rect 4571 24905 4583 24908
rect 4525 24899 4583 24905
rect 4706 24896 4712 24908
rect 4764 24896 4770 24948
rect 4893 24939 4951 24945
rect 4893 24905 4905 24939
rect 4939 24936 4951 24939
rect 5074 24936 5080 24948
rect 4939 24908 5080 24936
rect 4939 24905 4951 24908
rect 4893 24899 4951 24905
rect 5074 24896 5080 24908
rect 5132 24896 5138 24948
rect 5258 24896 5264 24948
rect 5316 24896 5322 24948
rect 7006 24896 7012 24948
rect 7064 24896 7070 24948
rect 12529 24939 12587 24945
rect 12529 24905 12541 24939
rect 12575 24936 12587 24939
rect 12710 24936 12716 24948
rect 12575 24908 12716 24936
rect 12575 24905 12587 24908
rect 12529 24899 12587 24905
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 29549 24939 29607 24945
rect 29549 24905 29561 24939
rect 29595 24936 29607 24939
rect 31110 24936 31116 24948
rect 29595 24908 31116 24936
rect 29595 24905 29607 24908
rect 29549 24899 29607 24905
rect 31110 24896 31116 24908
rect 31168 24896 31174 24948
rect 5276 24868 5304 24896
rect 8021 24871 8079 24877
rect 8021 24868 8033 24871
rect 5276 24840 8033 24868
rect 3970 24760 3976 24812
rect 4028 24760 4034 24812
rect 7374 24760 7380 24812
rect 7432 24760 7438 24812
rect 7006 24692 7012 24744
rect 7064 24732 7070 24744
rect 7576 24741 7604 24840
rect 8021 24837 8033 24840
rect 8067 24868 8079 24871
rect 24949 24871 25007 24877
rect 8067 24840 9674 24868
rect 8067 24837 8079 24840
rect 8021 24831 8079 24837
rect 7469 24735 7527 24741
rect 7469 24732 7481 24735
rect 7064 24704 7481 24732
rect 7064 24692 7070 24704
rect 7469 24701 7481 24704
rect 7515 24701 7527 24735
rect 7469 24695 7527 24701
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24701 7619 24735
rect 7561 24695 7619 24701
rect 8846 24692 8852 24744
rect 8904 24692 8910 24744
rect 8941 24735 8999 24741
rect 8941 24701 8953 24735
rect 8987 24701 8999 24735
rect 9646 24732 9674 24840
rect 24949 24837 24961 24871
rect 24995 24868 25007 24871
rect 26234 24868 26240 24880
rect 24995 24840 26240 24868
rect 24995 24837 25007 24840
rect 24949 24831 25007 24837
rect 26234 24828 26240 24840
rect 26292 24828 26298 24880
rect 28721 24871 28779 24877
rect 28721 24837 28733 24871
rect 28767 24868 28779 24871
rect 30009 24871 30067 24877
rect 30009 24868 30021 24871
rect 28767 24840 30021 24868
rect 28767 24837 28779 24840
rect 28721 24831 28779 24837
rect 30009 24837 30021 24840
rect 30055 24837 30067 24871
rect 30009 24831 30067 24837
rect 10134 24760 10140 24812
rect 10192 24800 10198 24812
rect 11885 24803 11943 24809
rect 11885 24800 11897 24803
rect 10192 24772 11897 24800
rect 10192 24760 10198 24772
rect 11885 24769 11897 24772
rect 11931 24769 11943 24803
rect 11885 24763 11943 24769
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24800 12495 24803
rect 13630 24800 13636 24812
rect 12483 24772 13636 24800
rect 12483 24769 12495 24772
rect 12437 24763 12495 24769
rect 11054 24732 11060 24744
rect 9646 24704 11060 24732
rect 8941 24695 8999 24701
rect 7190 24624 7196 24676
rect 7248 24664 7254 24676
rect 8956 24664 8984 24695
rect 7248 24636 8984 24664
rect 7248 24624 7254 24636
rect 10888 24608 10916 24704
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 11900 24732 11928 24763
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 17793 24803 17851 24809
rect 17793 24769 17805 24803
rect 17839 24800 17851 24803
rect 18049 24803 18107 24809
rect 17839 24772 18000 24800
rect 17839 24769 17851 24772
rect 17793 24763 17851 24769
rect 12713 24735 12771 24741
rect 12713 24732 12725 24735
rect 11900 24704 12725 24732
rect 12713 24701 12725 24704
rect 12759 24701 12771 24735
rect 12713 24695 12771 24701
rect 12728 24664 12756 24695
rect 12986 24692 12992 24744
rect 13044 24692 13050 24744
rect 13725 24735 13783 24741
rect 13725 24701 13737 24735
rect 13771 24732 13783 24735
rect 13906 24732 13912 24744
rect 13771 24704 13912 24732
rect 13771 24701 13783 24704
rect 13725 24695 13783 24701
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 16114 24692 16120 24744
rect 16172 24692 16178 24744
rect 16850 24692 16856 24744
rect 16908 24692 16914 24744
rect 17972 24732 18000 24772
rect 18049 24769 18061 24803
rect 18095 24800 18107 24803
rect 18230 24800 18236 24812
rect 18095 24772 18236 24800
rect 18095 24769 18107 24772
rect 18049 24763 18107 24769
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 25041 24803 25099 24809
rect 22520 24772 24716 24800
rect 22520 24760 22526 24772
rect 18325 24735 18383 24741
rect 18325 24732 18337 24735
rect 17972 24704 18337 24732
rect 18325 24701 18337 24704
rect 18371 24701 18383 24735
rect 18325 24695 18383 24701
rect 18874 24692 18880 24744
rect 18932 24692 18938 24744
rect 23750 24692 23756 24744
rect 23808 24692 23814 24744
rect 24489 24735 24547 24741
rect 24489 24701 24501 24735
rect 24535 24732 24547 24735
rect 24535 24704 24624 24732
rect 24535 24701 24547 24704
rect 24489 24695 24547 24701
rect 16868 24664 16896 24692
rect 12728 24636 16896 24664
rect 18046 24624 18052 24676
rect 18104 24624 18110 24676
rect 23768 24664 23796 24692
rect 24118 24664 24124 24676
rect 23768 24636 24124 24664
rect 24118 24624 24124 24636
rect 24176 24664 24182 24676
rect 24596 24673 24624 24704
rect 24581 24667 24639 24673
rect 24176 24636 24532 24664
rect 24176 24624 24182 24636
rect 3697 24599 3755 24605
rect 3697 24565 3709 24599
rect 3743 24596 3755 24599
rect 3878 24596 3884 24608
rect 3743 24568 3884 24596
rect 3743 24565 3755 24568
rect 3697 24559 3755 24565
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 8202 24556 8208 24608
rect 8260 24556 8266 24608
rect 9582 24556 9588 24608
rect 9640 24556 9646 24608
rect 10870 24556 10876 24608
rect 10928 24556 10934 24608
rect 12066 24556 12072 24608
rect 12124 24556 12130 24608
rect 13446 24556 13452 24608
rect 13504 24596 13510 24608
rect 13541 24599 13599 24605
rect 13541 24596 13553 24599
rect 13504 24568 13553 24596
rect 13504 24556 13510 24568
rect 13541 24565 13553 24568
rect 13587 24565 13599 24599
rect 13541 24559 13599 24565
rect 14274 24556 14280 24608
rect 14332 24556 14338 24608
rect 15378 24556 15384 24608
rect 15436 24596 15442 24608
rect 15565 24599 15623 24605
rect 15565 24596 15577 24599
rect 15436 24568 15577 24596
rect 15436 24556 15442 24568
rect 15565 24565 15577 24568
rect 15611 24565 15623 24599
rect 15565 24559 15623 24565
rect 16669 24599 16727 24605
rect 16669 24565 16681 24599
rect 16715 24596 16727 24599
rect 18064 24596 18092 24624
rect 16715 24568 18092 24596
rect 16715 24565 16727 24568
rect 16669 24559 16727 24565
rect 23842 24556 23848 24608
rect 23900 24556 23906 24608
rect 24504 24596 24532 24636
rect 24581 24633 24593 24667
rect 24627 24633 24639 24667
rect 24688 24664 24716 24772
rect 25041 24769 25053 24803
rect 25087 24800 25099 24803
rect 25409 24803 25467 24809
rect 25409 24800 25421 24803
rect 25087 24772 25421 24800
rect 25087 24769 25099 24772
rect 25041 24763 25099 24769
rect 25409 24769 25421 24772
rect 25455 24769 25467 24803
rect 26252 24800 26280 24828
rect 28813 24803 28871 24809
rect 28813 24800 28825 24803
rect 26252 24772 28825 24800
rect 25409 24763 25467 24769
rect 28813 24769 28825 24772
rect 28859 24800 28871 24803
rect 28859 24772 29040 24800
rect 28859 24769 28871 24772
rect 28813 24763 28871 24769
rect 25222 24692 25228 24744
rect 25280 24692 25286 24744
rect 25774 24692 25780 24744
rect 25832 24732 25838 24744
rect 25961 24735 26019 24741
rect 25961 24732 25973 24735
rect 25832 24704 25973 24732
rect 25832 24692 25838 24704
rect 25961 24701 25973 24704
rect 26007 24701 26019 24735
rect 25961 24695 26019 24701
rect 26142 24692 26148 24744
rect 26200 24692 26206 24744
rect 28905 24735 28963 24741
rect 28905 24732 28917 24735
rect 27816 24704 28917 24732
rect 27816 24673 27844 24704
rect 28905 24701 28917 24704
rect 28951 24701 28963 24735
rect 28905 24695 28963 24701
rect 27801 24667 27859 24673
rect 27801 24664 27813 24667
rect 24688 24636 27813 24664
rect 24581 24627 24639 24633
rect 27801 24633 27813 24636
rect 27847 24633 27859 24667
rect 27801 24627 27859 24633
rect 28261 24667 28319 24673
rect 28261 24633 28273 24667
rect 28307 24664 28319 24667
rect 29012 24664 29040 24772
rect 29362 24760 29368 24812
rect 29420 24800 29426 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 29420 24772 30573 24800
rect 29420 24760 29426 24772
rect 30561 24769 30573 24772
rect 30607 24769 30619 24803
rect 30561 24763 30619 24769
rect 29270 24692 29276 24744
rect 29328 24692 29334 24744
rect 29457 24735 29515 24741
rect 29457 24701 29469 24735
rect 29503 24701 29515 24735
rect 29457 24695 29515 24701
rect 29472 24664 29500 24695
rect 29822 24692 29828 24744
rect 29880 24732 29886 24744
rect 31297 24735 31355 24741
rect 31297 24732 31309 24735
rect 29880 24704 31309 24732
rect 29880 24692 29886 24704
rect 31297 24701 31309 24704
rect 31343 24701 31355 24735
rect 31297 24695 31355 24701
rect 34698 24692 34704 24744
rect 34756 24732 34762 24744
rect 35069 24735 35127 24741
rect 35069 24732 35081 24735
rect 34756 24704 35081 24732
rect 34756 24692 34762 24704
rect 35069 24701 35081 24704
rect 35115 24701 35127 24735
rect 35069 24695 35127 24701
rect 35894 24692 35900 24744
rect 35952 24692 35958 24744
rect 36998 24692 37004 24744
rect 37056 24692 37062 24744
rect 37090 24692 37096 24744
rect 37148 24732 37154 24744
rect 37829 24735 37887 24741
rect 37829 24732 37841 24735
rect 37148 24704 37841 24732
rect 37148 24692 37154 24704
rect 37829 24701 37841 24704
rect 37875 24701 37887 24735
rect 37829 24695 37887 24701
rect 29730 24664 29736 24676
rect 28307 24636 28764 24664
rect 29012 24636 29736 24664
rect 28307 24633 28319 24636
rect 28261 24627 28319 24633
rect 28736 24608 28764 24636
rect 29730 24624 29736 24636
rect 29788 24624 29794 24676
rect 26326 24596 26332 24608
rect 24504 24568 26332 24596
rect 26326 24556 26332 24568
rect 26384 24556 26390 24608
rect 26510 24556 26516 24608
rect 26568 24596 26574 24608
rect 26789 24599 26847 24605
rect 26789 24596 26801 24599
rect 26568 24568 26801 24596
rect 26568 24556 26574 24568
rect 26789 24565 26801 24568
rect 26835 24565 26847 24599
rect 26789 24559 26847 24565
rect 28350 24556 28356 24608
rect 28408 24556 28414 24608
rect 28718 24556 28724 24608
rect 28776 24556 28782 24608
rect 29914 24556 29920 24608
rect 29972 24556 29978 24608
rect 30742 24556 30748 24608
rect 30800 24556 30806 24608
rect 34330 24556 34336 24608
rect 34388 24596 34394 24608
rect 34517 24599 34575 24605
rect 34517 24596 34529 24599
rect 34388 24568 34529 24596
rect 34388 24556 34394 24568
rect 34517 24565 34529 24568
rect 34563 24565 34575 24599
rect 34517 24559 34575 24565
rect 35342 24556 35348 24608
rect 35400 24556 35406 24608
rect 36354 24556 36360 24608
rect 36412 24556 36418 24608
rect 36906 24556 36912 24608
rect 36964 24596 36970 24608
rect 37277 24599 37335 24605
rect 37277 24596 37289 24599
rect 36964 24568 37289 24596
rect 36964 24556 36970 24568
rect 37277 24565 37289 24568
rect 37323 24565 37335 24599
rect 37277 24559 37335 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 4801 24395 4859 24401
rect 4801 24361 4813 24395
rect 4847 24392 4859 24395
rect 5074 24392 5080 24404
rect 4847 24364 5080 24392
rect 4847 24361 4859 24364
rect 4801 24355 4859 24361
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 6917 24395 6975 24401
rect 6917 24361 6929 24395
rect 6963 24392 6975 24395
rect 7374 24392 7380 24404
rect 6963 24364 7380 24392
rect 6963 24361 6975 24364
rect 6917 24355 6975 24361
rect 7374 24352 7380 24364
rect 7432 24352 7438 24404
rect 11885 24395 11943 24401
rect 11885 24361 11897 24395
rect 11931 24392 11943 24395
rect 13906 24392 13912 24404
rect 11931 24364 13912 24392
rect 11931 24361 11943 24364
rect 11885 24355 11943 24361
rect 13906 24352 13912 24364
rect 13964 24352 13970 24404
rect 15749 24395 15807 24401
rect 15749 24361 15761 24395
rect 15795 24392 15807 24395
rect 16114 24392 16120 24404
rect 15795 24364 16120 24392
rect 15795 24361 15807 24364
rect 15749 24355 15807 24361
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 17310 24392 17316 24404
rect 16224 24364 17316 24392
rect 16224 24336 16252 24364
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 24026 24352 24032 24404
rect 24084 24392 24090 24404
rect 24121 24395 24179 24401
rect 24121 24392 24133 24395
rect 24084 24364 24133 24392
rect 24084 24352 24090 24364
rect 24121 24361 24133 24364
rect 24167 24361 24179 24395
rect 24121 24355 24179 24361
rect 24397 24395 24455 24401
rect 24397 24361 24409 24395
rect 24443 24392 24455 24395
rect 25038 24392 25044 24404
rect 24443 24364 25044 24392
rect 24443 24361 24455 24364
rect 24397 24355 24455 24361
rect 25038 24352 25044 24364
rect 25096 24392 25102 24404
rect 26142 24392 26148 24404
rect 25096 24364 26148 24392
rect 25096 24352 25102 24364
rect 26142 24352 26148 24364
rect 26200 24352 26206 24404
rect 26418 24352 26424 24404
rect 26476 24392 26482 24404
rect 26605 24395 26663 24401
rect 26605 24392 26617 24395
rect 26476 24364 26617 24392
rect 26476 24352 26482 24364
rect 26605 24361 26617 24364
rect 26651 24361 26663 24395
rect 26605 24355 26663 24361
rect 27614 24352 27620 24404
rect 27672 24392 27678 24404
rect 29365 24395 29423 24401
rect 27672 24364 28994 24392
rect 27672 24352 27678 24364
rect 12066 24324 12072 24336
rect 11256 24296 12072 24324
rect 11256 24265 11284 24296
rect 12066 24284 12072 24296
rect 12124 24284 12130 24336
rect 15657 24327 15715 24333
rect 15657 24293 15669 24327
rect 15703 24324 15715 24327
rect 16206 24324 16212 24336
rect 15703 24296 16212 24324
rect 15703 24293 15715 24296
rect 15657 24287 15715 24293
rect 16206 24284 16212 24296
rect 16264 24284 16270 24336
rect 27632 24324 27660 24352
rect 25976 24296 27660 24324
rect 28966 24324 28994 24364
rect 29365 24361 29377 24395
rect 29411 24392 29423 24395
rect 29822 24392 29828 24404
rect 29411 24364 29828 24392
rect 29411 24361 29423 24364
rect 29365 24355 29423 24361
rect 29822 24352 29828 24364
rect 29880 24352 29886 24404
rect 30190 24352 30196 24404
rect 30248 24392 30254 24404
rect 30285 24395 30343 24401
rect 30285 24392 30297 24395
rect 30248 24364 30297 24392
rect 30248 24352 30254 24364
rect 30285 24361 30297 24364
rect 30331 24361 30343 24395
rect 30285 24355 30343 24361
rect 31110 24352 31116 24404
rect 31168 24352 31174 24404
rect 34517 24395 34575 24401
rect 34517 24361 34529 24395
rect 34563 24392 34575 24395
rect 34606 24392 34612 24404
rect 34563 24364 34612 24392
rect 34563 24361 34575 24364
rect 34517 24355 34575 24361
rect 34606 24352 34612 24364
rect 34664 24352 34670 24404
rect 37734 24352 37740 24404
rect 37792 24392 37798 24404
rect 37792 24364 38424 24392
rect 37792 24352 37798 24364
rect 32582 24324 32588 24336
rect 28966 24296 32588 24324
rect 25976 24268 26004 24296
rect 32582 24284 32588 24296
rect 32640 24324 32646 24336
rect 33318 24324 33324 24336
rect 32640 24296 33324 24324
rect 32640 24284 32646 24296
rect 33318 24284 33324 24296
rect 33376 24284 33382 24336
rect 11241 24259 11299 24265
rect 11241 24225 11253 24259
rect 11287 24225 11299 24259
rect 15197 24259 15255 24265
rect 15197 24256 15209 24259
rect 11241 24219 11299 24225
rect 13188 24228 15209 24256
rect 3418 24148 3424 24200
rect 3476 24148 3482 24200
rect 4433 24191 4491 24197
rect 4433 24157 4445 24191
rect 4479 24188 4491 24191
rect 4614 24188 4620 24200
rect 4479 24160 4620 24188
rect 4479 24157 4491 24160
rect 4433 24151 4491 24157
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 6362 24148 6368 24200
rect 6420 24148 6426 24200
rect 7009 24191 7067 24197
rect 7009 24157 7021 24191
rect 7055 24188 7067 24191
rect 7098 24188 7104 24200
rect 7055 24160 7104 24188
rect 7055 24157 7067 24160
rect 7009 24151 7067 24157
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 9030 24148 9036 24200
rect 9088 24148 9094 24200
rect 10870 24148 10876 24200
rect 10928 24188 10934 24200
rect 13188 24188 13216 24228
rect 15197 24225 15209 24228
rect 15243 24256 15255 24259
rect 16301 24259 16359 24265
rect 16301 24256 16313 24259
rect 15243 24228 16313 24256
rect 15243 24225 15255 24228
rect 15197 24219 15255 24225
rect 16301 24225 16313 24228
rect 16347 24225 16359 24259
rect 18506 24256 18512 24268
rect 16301 24219 16359 24225
rect 17880 24228 18512 24256
rect 10928 24160 13216 24188
rect 13265 24191 13323 24197
rect 10928 24148 10934 24160
rect 13265 24157 13277 24191
rect 13311 24188 13323 24191
rect 13538 24188 13544 24200
rect 13311 24160 13544 24188
rect 13311 24157 13323 24160
rect 13265 24151 13323 24157
rect 13538 24148 13544 24160
rect 13596 24188 13602 24200
rect 14550 24188 14556 24200
rect 13596 24160 14556 24188
rect 13596 24148 13602 24160
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 14642 24148 14648 24200
rect 14700 24148 14706 24200
rect 16117 24191 16175 24197
rect 16117 24157 16129 24191
rect 16163 24188 16175 24191
rect 16390 24188 16396 24200
rect 16163 24160 16396 24188
rect 16163 24157 16175 24160
rect 16117 24151 16175 24157
rect 16390 24148 16396 24160
rect 16448 24148 16454 24200
rect 17880 24188 17908 24228
rect 18506 24216 18512 24228
rect 18564 24216 18570 24268
rect 25958 24216 25964 24268
rect 26016 24216 26022 24268
rect 27985 24259 28043 24265
rect 27985 24256 27997 24259
rect 26068 24228 27997 24256
rect 16684 24160 17908 24188
rect 6822 24080 6828 24132
rect 6880 24120 6886 24132
rect 7254 24123 7312 24129
rect 7254 24120 7266 24123
rect 6880 24092 7266 24120
rect 6880 24080 6886 24092
rect 7254 24089 7266 24092
rect 7300 24089 7312 24123
rect 13020 24123 13078 24129
rect 7254 24083 7312 24089
rect 11624 24092 12965 24120
rect 11624 24064 11652 24092
rect 2866 24012 2872 24064
rect 2924 24012 2930 24064
rect 3786 24012 3792 24064
rect 3844 24012 3850 24064
rect 5169 24055 5227 24061
rect 5169 24021 5181 24055
rect 5215 24052 5227 24055
rect 5258 24052 5264 24064
rect 5215 24024 5264 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 8662 24052 8668 24064
rect 8435 24024 8668 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 9306 24012 9312 24064
rect 9364 24052 9370 24064
rect 9677 24055 9735 24061
rect 9677 24052 9689 24055
rect 9364 24024 9689 24052
rect 9364 24012 9370 24024
rect 9677 24021 9689 24024
rect 9723 24021 9735 24055
rect 9677 24015 9735 24021
rect 11606 24012 11612 24064
rect 11664 24012 11670 24064
rect 11790 24012 11796 24064
rect 11848 24012 11854 24064
rect 12937 24052 12965 24092
rect 13020 24089 13032 24123
rect 13066 24120 13078 24123
rect 14093 24123 14151 24129
rect 14093 24120 14105 24123
rect 13066 24092 14105 24120
rect 13066 24089 13078 24092
rect 13020 24083 13078 24089
rect 14093 24089 14105 24092
rect 14139 24089 14151 24123
rect 14093 24083 14151 24089
rect 16209 24123 16267 24129
rect 16209 24089 16221 24123
rect 16255 24120 16267 24123
rect 16684 24120 16712 24160
rect 17954 24148 17960 24200
rect 18012 24148 18018 24200
rect 18598 24148 18604 24200
rect 18656 24148 18662 24200
rect 24762 24148 24768 24200
rect 24820 24188 24826 24200
rect 25777 24191 25835 24197
rect 25777 24188 25789 24191
rect 24820 24160 25789 24188
rect 24820 24148 24826 24160
rect 25777 24157 25789 24160
rect 25823 24188 25835 24191
rect 26068 24188 26096 24228
rect 27985 24225 27997 24228
rect 28031 24225 28043 24259
rect 27985 24219 28043 24225
rect 29638 24216 29644 24268
rect 29696 24216 29702 24268
rect 29730 24216 29736 24268
rect 29788 24216 29794 24268
rect 29914 24216 29920 24268
rect 29972 24256 29978 24268
rect 32401 24259 32459 24265
rect 32401 24256 32413 24259
rect 29972 24228 32413 24256
rect 29972 24216 29978 24228
rect 32401 24225 32413 24228
rect 32447 24225 32459 24259
rect 32401 24219 32459 24225
rect 35618 24216 35624 24268
rect 35676 24256 35682 24268
rect 38396 24265 38424 24364
rect 36357 24259 36415 24265
rect 36357 24256 36369 24259
rect 35676 24228 36369 24256
rect 35676 24216 35682 24228
rect 36357 24225 36369 24228
rect 36403 24225 36415 24259
rect 36357 24219 36415 24225
rect 38381 24259 38439 24265
rect 38381 24225 38393 24259
rect 38427 24225 38439 24259
rect 38381 24219 38439 24225
rect 25823 24160 26096 24188
rect 26145 24191 26203 24197
rect 25823 24157 25835 24160
rect 25777 24151 25835 24157
rect 26145 24157 26157 24191
rect 26191 24188 26203 24191
rect 26510 24188 26516 24200
rect 26191 24160 26516 24188
rect 26191 24157 26203 24160
rect 26145 24151 26203 24157
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 28252 24191 28310 24197
rect 28252 24157 28264 24191
rect 28298 24188 28310 24191
rect 29546 24188 29552 24200
rect 28298 24160 29552 24188
rect 28298 24157 28310 24160
rect 28252 24151 28310 24157
rect 16255 24092 16712 24120
rect 16255 24089 16267 24092
rect 16209 24083 16267 24089
rect 16758 24080 16764 24132
rect 16816 24120 16822 24132
rect 17712 24123 17770 24129
rect 16816 24092 17632 24120
rect 16816 24080 16822 24092
rect 13354 24052 13360 24064
rect 12937 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24052 13418 24064
rect 13633 24055 13691 24061
rect 13633 24052 13645 24055
rect 13412 24024 13645 24052
rect 13412 24012 13418 24024
rect 13633 24021 13645 24024
rect 13679 24052 13691 24055
rect 13722 24052 13728 24064
rect 13679 24024 13728 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 13722 24012 13728 24024
rect 13780 24052 13786 24064
rect 15562 24052 15568 24064
rect 13780 24024 15568 24052
rect 13780 24012 13786 24024
rect 15562 24012 15568 24024
rect 15620 24012 15626 24064
rect 16577 24055 16635 24061
rect 16577 24021 16589 24055
rect 16623 24052 16635 24055
rect 17034 24052 17040 24064
rect 16623 24024 17040 24052
rect 16623 24021 16635 24024
rect 16577 24015 16635 24021
rect 17034 24012 17040 24024
rect 17092 24012 17098 24064
rect 17604 24052 17632 24092
rect 17712 24089 17724 24123
rect 17758 24120 17770 24123
rect 18049 24123 18107 24129
rect 18049 24120 18061 24123
rect 17758 24092 18061 24120
rect 17758 24089 17770 24092
rect 17712 24083 17770 24089
rect 18049 24089 18061 24092
rect 18095 24089 18107 24123
rect 18049 24083 18107 24089
rect 25532 24123 25590 24129
rect 25532 24089 25544 24123
rect 25578 24120 25590 24123
rect 25682 24120 25688 24132
rect 25578 24092 25688 24120
rect 25578 24089 25590 24092
rect 25532 24083 25590 24089
rect 25682 24080 25688 24092
rect 25740 24080 25746 24132
rect 26712 24120 26740 24151
rect 29546 24148 29552 24160
rect 29604 24148 29610 24200
rect 29748 24120 29776 24216
rect 29825 24191 29883 24197
rect 29825 24157 29837 24191
rect 29871 24188 29883 24191
rect 30742 24188 30748 24200
rect 29871 24160 30748 24188
rect 29871 24157 29883 24160
rect 29825 24151 29883 24157
rect 30742 24148 30748 24160
rect 30800 24148 30806 24200
rect 30926 24148 30932 24200
rect 30984 24148 30990 24200
rect 31665 24191 31723 24197
rect 31665 24157 31677 24191
rect 31711 24157 31723 24191
rect 31665 24151 31723 24157
rect 29917 24123 29975 24129
rect 29917 24120 29929 24123
rect 25792 24092 26740 24120
rect 27264 24092 28396 24120
rect 29748 24092 29929 24120
rect 17862 24052 17868 24064
rect 17604 24024 17868 24052
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 25222 24012 25228 24064
rect 25280 24052 25286 24064
rect 25792 24052 25820 24092
rect 25280 24024 25820 24052
rect 25280 24012 25286 24024
rect 26234 24012 26240 24064
rect 26292 24012 26298 24064
rect 26326 24012 26332 24064
rect 26384 24052 26390 24064
rect 27264 24052 27292 24092
rect 26384 24024 27292 24052
rect 26384 24012 26390 24024
rect 27338 24012 27344 24064
rect 27396 24012 27402 24064
rect 28368 24052 28396 24092
rect 29917 24089 29929 24092
rect 29963 24089 29975 24123
rect 29917 24083 29975 24089
rect 30282 24080 30288 24132
rect 30340 24120 30346 24132
rect 31680 24120 31708 24151
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 33836 24160 34897 24188
rect 33836 24148 33842 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 35529 24191 35587 24197
rect 35529 24157 35541 24191
rect 35575 24188 35587 24191
rect 35710 24188 35716 24200
rect 35575 24160 35716 24188
rect 35575 24157 35587 24160
rect 35529 24151 35587 24157
rect 35710 24148 35716 24160
rect 35768 24148 35774 24200
rect 36170 24148 36176 24200
rect 36228 24148 36234 24200
rect 36624 24191 36682 24197
rect 36624 24157 36636 24191
rect 36670 24188 36682 24191
rect 36906 24188 36912 24200
rect 36670 24160 36912 24188
rect 36670 24157 36682 24160
rect 36624 24151 36682 24157
rect 36906 24148 36912 24160
rect 36964 24148 36970 24200
rect 30340 24092 31708 24120
rect 30340 24080 30346 24092
rect 29270 24052 29276 24064
rect 28368 24024 29276 24052
rect 29270 24012 29276 24024
rect 29328 24052 29334 24064
rect 30190 24052 30196 24064
rect 29328 24024 30196 24052
rect 29328 24012 29334 24024
rect 30190 24012 30196 24024
rect 30248 24012 30254 24064
rect 30374 24012 30380 24064
rect 30432 24012 30438 24064
rect 31846 24012 31852 24064
rect 31904 24012 31910 24064
rect 35621 24055 35679 24061
rect 35621 24021 35633 24055
rect 35667 24052 35679 24055
rect 35710 24052 35716 24064
rect 35667 24024 35716 24052
rect 35667 24021 35679 24024
rect 35621 24015 35679 24021
rect 35710 24012 35716 24024
rect 35768 24012 35774 24064
rect 36630 24012 36636 24064
rect 36688 24052 36694 24064
rect 37829 24055 37887 24061
rect 37829 24052 37841 24055
rect 36688 24024 37841 24052
rect 36688 24012 36694 24024
rect 37829 24021 37841 24024
rect 37875 24021 37887 24055
rect 37829 24015 37887 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 3237 23851 3295 23857
rect 3237 23817 3249 23851
rect 3283 23848 3295 23851
rect 3418 23848 3424 23860
rect 3283 23820 3424 23848
rect 3283 23817 3295 23820
rect 3237 23811 3295 23817
rect 3418 23808 3424 23820
rect 3476 23808 3482 23860
rect 4982 23808 4988 23860
rect 5040 23848 5046 23860
rect 5166 23848 5172 23860
rect 5040 23820 5172 23848
rect 5040 23808 5046 23820
rect 5166 23808 5172 23820
rect 5224 23848 5230 23860
rect 5224 23820 5488 23848
rect 5224 23808 5230 23820
rect 3605 23783 3663 23789
rect 3605 23749 3617 23783
rect 3651 23780 3663 23783
rect 5460 23780 5488 23820
rect 5718 23808 5724 23860
rect 5776 23848 5782 23860
rect 6089 23851 6147 23857
rect 6089 23848 6101 23851
rect 5776 23820 6101 23848
rect 5776 23808 5782 23820
rect 6089 23817 6101 23820
rect 6135 23817 6147 23851
rect 6089 23811 6147 23817
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 7742 23848 7748 23860
rect 6687 23820 7748 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 5813 23783 5871 23789
rect 5813 23780 5825 23783
rect 3651 23752 5396 23780
rect 5460 23752 5825 23780
rect 3651 23749 3663 23752
rect 3605 23743 3663 23749
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23712 3755 23715
rect 4706 23712 4712 23724
rect 3743 23684 4712 23712
rect 3743 23681 3755 23684
rect 3697 23675 3755 23681
rect 4706 23672 4712 23684
rect 4764 23672 4770 23724
rect 3050 23604 3056 23656
rect 3108 23604 3114 23656
rect 3878 23604 3884 23656
rect 3936 23604 3942 23656
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 4617 23647 4675 23653
rect 4617 23644 4629 23647
rect 4028 23616 4629 23644
rect 4028 23604 4034 23616
rect 4617 23613 4629 23616
rect 4663 23613 4675 23647
rect 4617 23607 4675 23613
rect 4798 23604 4804 23656
rect 4856 23604 4862 23656
rect 5258 23604 5264 23656
rect 5316 23604 5322 23656
rect 3896 23576 3924 23604
rect 5276 23576 5304 23604
rect 5368 23588 5396 23752
rect 5813 23749 5825 23752
rect 5859 23749 5871 23783
rect 5813 23743 5871 23749
rect 6104 23644 6132 23811
rect 7742 23808 7748 23820
rect 7800 23808 7806 23860
rect 8202 23808 8208 23860
rect 8260 23808 8266 23860
rect 8570 23808 8576 23860
rect 8628 23848 8634 23860
rect 9030 23848 9036 23860
rect 8628 23820 9036 23848
rect 8628 23808 8634 23820
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 9582 23808 9588 23860
rect 9640 23808 9646 23860
rect 13814 23848 13820 23860
rect 12728 23820 13820 23848
rect 7460 23783 7518 23789
rect 7460 23749 7472 23783
rect 7506 23780 7518 23783
rect 8220 23780 8248 23808
rect 7506 23752 8248 23780
rect 9600 23780 9628 23808
rect 9778 23783 9836 23789
rect 9778 23780 9790 23783
rect 9600 23752 9790 23780
rect 7506 23749 7518 23752
rect 7460 23743 7518 23749
rect 9778 23749 9790 23752
rect 9824 23749 9836 23783
rect 9778 23743 9836 23749
rect 10318 23740 10324 23792
rect 10376 23780 10382 23792
rect 11333 23783 11391 23789
rect 11333 23780 11345 23783
rect 10376 23752 11345 23780
rect 10376 23740 10382 23752
rect 11333 23749 11345 23752
rect 11379 23780 11391 23783
rect 12526 23780 12532 23792
rect 11379 23752 12532 23780
rect 11379 23749 11391 23752
rect 11333 23743 11391 23749
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 12728 23724 12756 23820
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 13909 23851 13967 23857
rect 13909 23817 13921 23851
rect 13955 23848 13967 23851
rect 14274 23848 14280 23860
rect 13955 23820 14280 23848
rect 13955 23817 13967 23820
rect 13909 23811 13967 23817
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 14369 23851 14427 23857
rect 14369 23817 14381 23851
rect 14415 23848 14427 23851
rect 14642 23848 14648 23860
rect 14415 23820 14648 23848
rect 14415 23817 14427 23820
rect 14369 23811 14427 23817
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 16485 23851 16543 23857
rect 16485 23817 16497 23851
rect 16531 23848 16543 23851
rect 16758 23848 16764 23860
rect 16531 23820 16764 23848
rect 16531 23817 16543 23820
rect 16485 23811 16543 23817
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 18046 23848 18052 23860
rect 16868 23820 18052 23848
rect 13296 23783 13354 23789
rect 13296 23749 13308 23783
rect 13342 23780 13354 23783
rect 13446 23780 13452 23792
rect 13342 23752 13452 23780
rect 13342 23749 13354 23752
rect 13296 23743 13354 23749
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 14550 23740 14556 23792
rect 14608 23780 14614 23792
rect 16298 23780 16304 23792
rect 14608 23752 16304 23780
rect 14608 23740 14614 23752
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23712 6791 23715
rect 7006 23712 7012 23724
rect 6779 23684 7012 23712
rect 6779 23681 6791 23684
rect 6733 23675 6791 23681
rect 6270 23644 6276 23656
rect 6104 23616 6276 23644
rect 6270 23604 6276 23616
rect 6328 23644 6334 23656
rect 6457 23647 6515 23653
rect 6457 23644 6469 23647
rect 6328 23616 6469 23644
rect 6328 23604 6334 23616
rect 6457 23613 6469 23616
rect 6503 23613 6515 23647
rect 6457 23607 6515 23613
rect 3896 23548 5304 23576
rect 5350 23536 5356 23588
rect 5408 23576 5414 23588
rect 6748 23576 6776 23675
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 11977 23715 12035 23721
rect 11977 23681 11989 23715
rect 12023 23712 12035 23715
rect 12710 23712 12716 23724
rect 12023 23684 12716 23712
rect 12023 23681 12035 23684
rect 11977 23675 12035 23681
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 14001 23715 14059 23721
rect 14001 23712 14013 23715
rect 13688 23684 14013 23712
rect 13688 23672 13694 23684
rect 14001 23681 14013 23684
rect 14047 23681 14059 23715
rect 14001 23675 14059 23681
rect 14182 23672 14188 23724
rect 14240 23712 14246 23724
rect 15120 23721 15148 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 15378 23721 15384 23724
rect 14921 23715 14979 23721
rect 14921 23712 14933 23715
rect 14240 23684 14933 23712
rect 14240 23672 14246 23684
rect 14921 23681 14933 23684
rect 14967 23681 14979 23715
rect 14921 23675 14979 23681
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 15372 23712 15384 23721
rect 15339 23684 15384 23712
rect 15105 23675 15163 23681
rect 15372 23675 15384 23684
rect 15378 23672 15384 23675
rect 15436 23672 15442 23724
rect 16868 23721 16896 23820
rect 18046 23808 18052 23820
rect 18104 23808 18110 23860
rect 18506 23808 18512 23860
rect 18564 23808 18570 23860
rect 18690 23808 18696 23860
rect 18748 23808 18754 23860
rect 18785 23851 18843 23857
rect 18785 23817 18797 23851
rect 18831 23848 18843 23851
rect 18874 23848 18880 23860
rect 18831 23820 18880 23848
rect 18831 23817 18843 23820
rect 18785 23811 18843 23817
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 22097 23851 22155 23857
rect 22097 23817 22109 23851
rect 22143 23848 22155 23851
rect 22186 23848 22192 23860
rect 22143 23820 22192 23848
rect 22143 23817 22155 23820
rect 22097 23811 22155 23817
rect 22186 23808 22192 23820
rect 22244 23848 22250 23860
rect 22462 23848 22468 23860
rect 22244 23820 22468 23848
rect 22244 23808 22250 23820
rect 22462 23808 22468 23820
rect 22520 23808 22526 23860
rect 23842 23808 23848 23860
rect 23900 23808 23906 23860
rect 25038 23808 25044 23860
rect 25096 23808 25102 23860
rect 26326 23808 26332 23860
rect 26384 23848 26390 23860
rect 26384 23820 27292 23848
rect 26384 23808 26390 23820
rect 18524 23780 18552 23808
rect 18708 23780 18736 23808
rect 19245 23783 19303 23789
rect 19245 23780 19257 23783
rect 18524 23752 18644 23780
rect 18708 23752 19257 23780
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17862 23672 17868 23724
rect 17920 23721 17926 23724
rect 17920 23715 17948 23721
rect 17936 23681 17948 23715
rect 17920 23675 17948 23681
rect 17920 23672 17926 23675
rect 18046 23672 18052 23724
rect 18104 23672 18110 23724
rect 18616 23712 18644 23752
rect 19245 23749 19257 23752
rect 19291 23749 19303 23783
rect 19245 23743 19303 23749
rect 23652 23783 23710 23789
rect 23652 23749 23664 23783
rect 23698 23780 23710 23783
rect 23860 23780 23888 23808
rect 23698 23752 23888 23780
rect 23698 23749 23710 23752
rect 23652 23743 23710 23749
rect 19153 23715 19211 23721
rect 19153 23712 19165 23715
rect 18616 23684 19165 23712
rect 19153 23681 19165 23684
rect 19199 23681 19211 23715
rect 19153 23675 19211 23681
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23712 24915 23715
rect 25056 23712 25084 23808
rect 27264 23780 27292 23820
rect 27338 23808 27344 23860
rect 27396 23808 27402 23860
rect 28350 23808 28356 23860
rect 28408 23808 28414 23860
rect 29730 23808 29736 23860
rect 29788 23848 29794 23860
rect 30469 23851 30527 23857
rect 29788 23820 30236 23848
rect 29788 23808 29794 23820
rect 27433 23783 27491 23789
rect 27433 23780 27445 23783
rect 27264 23752 27445 23780
rect 27433 23749 27445 23752
rect 27479 23780 27491 23783
rect 28166 23780 28172 23792
rect 27479 23752 28172 23780
rect 27479 23749 27491 23752
rect 27433 23743 27491 23749
rect 28166 23740 28172 23752
rect 28224 23740 28230 23792
rect 24903 23684 25084 23712
rect 24903 23681 24915 23684
rect 24857 23675 24915 23681
rect 25222 23672 25228 23724
rect 25280 23672 25286 23724
rect 25774 23672 25780 23724
rect 25832 23672 25838 23724
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 28368 23721 28396 23808
rect 30208 23780 30236 23820
rect 30469 23817 30481 23851
rect 30515 23848 30527 23851
rect 30926 23848 30932 23860
rect 30515 23820 30932 23848
rect 30515 23817 30527 23820
rect 30469 23811 30527 23817
rect 30926 23808 30932 23820
rect 30984 23808 30990 23860
rect 36909 23851 36967 23857
rect 36909 23817 36921 23851
rect 36955 23848 36967 23851
rect 36998 23848 37004 23860
rect 36955 23820 37004 23848
rect 36955 23817 36967 23820
rect 36909 23811 36967 23817
rect 36998 23808 37004 23820
rect 37056 23808 37062 23860
rect 30837 23783 30895 23789
rect 30837 23780 30849 23783
rect 30208 23752 30849 23780
rect 30837 23749 30849 23752
rect 30883 23749 30895 23783
rect 30837 23743 30895 23749
rect 34072 23752 35572 23780
rect 29362 23721 29368 23724
rect 28353 23715 28411 23721
rect 28353 23681 28365 23715
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 29340 23715 29368 23721
rect 29340 23681 29352 23715
rect 29340 23675 29368 23681
rect 29362 23672 29368 23675
rect 29420 23672 29426 23724
rect 30193 23715 30251 23721
rect 30193 23681 30205 23715
rect 30239 23712 30251 23715
rect 30282 23712 30288 23724
rect 30239 23684 30288 23712
rect 30239 23681 30251 23684
rect 30193 23675 30251 23681
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 34072 23721 34100 23752
rect 34330 23721 34336 23724
rect 30929 23715 30987 23721
rect 30929 23681 30941 23715
rect 30975 23712 30987 23715
rect 31297 23715 31355 23721
rect 31297 23712 31309 23715
rect 30975 23684 31309 23712
rect 30975 23681 30987 23684
rect 30929 23675 30987 23681
rect 31297 23681 31309 23684
rect 31343 23681 31355 23715
rect 31297 23675 31355 23681
rect 34057 23715 34115 23721
rect 34057 23681 34069 23715
rect 34103 23681 34115 23715
rect 34324 23712 34336 23721
rect 34291 23684 34336 23712
rect 34057 23675 34115 23681
rect 34324 23675 34336 23684
rect 34330 23672 34336 23675
rect 34388 23672 34394 23724
rect 35544 23721 35572 23752
rect 35529 23715 35587 23721
rect 35529 23681 35541 23715
rect 35575 23712 35587 23715
rect 35618 23712 35624 23724
rect 35575 23684 35624 23712
rect 35575 23681 35587 23684
rect 35529 23675 35587 23681
rect 35618 23672 35624 23684
rect 35676 23672 35682 23724
rect 35796 23715 35854 23721
rect 35796 23681 35808 23715
rect 35842 23712 35854 23715
rect 37277 23715 37335 23721
rect 37277 23712 37289 23715
rect 35842 23684 37289 23712
rect 35842 23681 35854 23684
rect 35796 23675 35854 23681
rect 37277 23681 37289 23684
rect 37323 23681 37335 23715
rect 37277 23675 37335 23681
rect 7098 23604 7104 23656
rect 7156 23644 7162 23656
rect 7193 23647 7251 23653
rect 7193 23644 7205 23647
rect 7156 23616 7205 23644
rect 7156 23604 7162 23616
rect 7193 23613 7205 23616
rect 7239 23613 7251 23647
rect 7193 23607 7251 23613
rect 5408 23548 6776 23576
rect 5408 23536 5414 23548
rect 2498 23468 2504 23520
rect 2556 23468 2562 23520
rect 4062 23468 4068 23520
rect 4120 23468 4126 23520
rect 5442 23468 5448 23520
rect 5500 23468 5506 23520
rect 7098 23468 7104 23520
rect 7156 23468 7162 23520
rect 7208 23508 7236 23607
rect 8386 23604 8392 23656
rect 8444 23604 8450 23656
rect 10045 23647 10103 23653
rect 10045 23613 10057 23647
rect 10091 23644 10103 23647
rect 10226 23644 10232 23656
rect 10091 23616 10232 23644
rect 10091 23613 10103 23616
rect 10045 23607 10103 23613
rect 10226 23604 10232 23616
rect 10284 23604 10290 23656
rect 13541 23647 13599 23653
rect 13541 23613 13553 23647
rect 13587 23613 13599 23647
rect 13541 23607 13599 23613
rect 8404 23576 8432 23604
rect 8665 23579 8723 23585
rect 8665 23576 8677 23579
rect 8404 23548 8677 23576
rect 8665 23545 8677 23548
rect 8711 23545 8723 23579
rect 13556 23576 13584 23607
rect 13722 23604 13728 23656
rect 13780 23604 13786 23656
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 14200 23644 14228 23672
rect 13872 23616 14228 23644
rect 13872 23604 13878 23616
rect 17034 23604 17040 23656
rect 17092 23644 17098 23656
rect 17773 23647 17831 23653
rect 17092 23616 17632 23644
rect 17092 23604 17098 23616
rect 14550 23576 14556 23588
rect 13556 23548 14556 23576
rect 8665 23539 8723 23545
rect 14550 23536 14556 23548
rect 14608 23536 14614 23588
rect 17494 23536 17500 23588
rect 17552 23536 17558 23588
rect 7834 23508 7840 23520
rect 7208 23480 7840 23508
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 12161 23511 12219 23517
rect 12161 23477 12173 23511
rect 12207 23508 12219 23511
rect 13722 23508 13728 23520
rect 12207 23480 13728 23508
rect 12207 23477 12219 23480
rect 12161 23471 12219 23477
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 16206 23508 16212 23520
rect 15436 23480 16212 23508
rect 15436 23468 15442 23480
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 17604 23508 17632 23616
rect 17773 23613 17785 23647
rect 17819 23644 17831 23647
rect 18230 23644 18236 23656
rect 17819 23616 18236 23644
rect 17819 23613 17831 23616
rect 17773 23607 17831 23613
rect 18230 23604 18236 23616
rect 18288 23604 18294 23656
rect 18690 23604 18696 23656
rect 18748 23644 18754 23656
rect 19337 23647 19395 23653
rect 19337 23644 19349 23647
rect 18748 23616 19349 23644
rect 18748 23604 18754 23616
rect 19337 23613 19349 23616
rect 19383 23613 19395 23647
rect 19337 23607 19395 23613
rect 20165 23647 20223 23653
rect 20165 23613 20177 23647
rect 20211 23613 20223 23647
rect 20165 23607 20223 23613
rect 20180 23576 20208 23607
rect 23382 23604 23388 23656
rect 23440 23604 23446 23656
rect 25041 23647 25099 23653
rect 25041 23613 25053 23647
rect 25087 23644 25099 23647
rect 25240 23644 25268 23672
rect 25792 23644 25820 23672
rect 25087 23616 25268 23644
rect 25424 23616 25820 23644
rect 25087 23613 25099 23616
rect 25041 23607 25099 23613
rect 18432 23548 20208 23576
rect 24765 23579 24823 23585
rect 18432 23508 18460 23548
rect 24765 23545 24777 23579
rect 24811 23576 24823 23579
rect 25424 23576 25452 23616
rect 25866 23604 25872 23656
rect 25924 23653 25930 23656
rect 25924 23647 25952 23653
rect 25940 23613 25952 23647
rect 25924 23607 25952 23613
rect 27525 23647 27583 23653
rect 27525 23613 27537 23647
rect 27571 23644 27583 23647
rect 27706 23644 27712 23656
rect 27571 23616 27712 23644
rect 27571 23613 27583 23616
rect 27525 23607 27583 23613
rect 25924 23604 25930 23607
rect 27706 23604 27712 23616
rect 27764 23604 27770 23656
rect 28994 23604 29000 23656
rect 29052 23644 29058 23656
rect 29181 23647 29239 23653
rect 29181 23644 29193 23647
rect 29052 23616 29193 23644
rect 29052 23604 29058 23616
rect 29181 23613 29193 23616
rect 29227 23613 29239 23647
rect 29181 23607 29239 23613
rect 29457 23647 29515 23653
rect 29457 23613 29469 23647
rect 29503 23644 29515 23647
rect 29822 23644 29828 23656
rect 29503 23616 29828 23644
rect 29503 23613 29515 23616
rect 29457 23607 29515 23613
rect 29822 23604 29828 23616
rect 29880 23604 29886 23656
rect 30098 23604 30104 23656
rect 30156 23644 30162 23656
rect 30377 23647 30435 23653
rect 30377 23644 30389 23647
rect 30156 23616 30389 23644
rect 30156 23604 30162 23616
rect 30377 23613 30389 23616
rect 30423 23613 30435 23647
rect 30377 23607 30435 23613
rect 24811 23548 25452 23576
rect 25501 23579 25559 23585
rect 24811 23545 24823 23548
rect 24765 23539 24823 23545
rect 25501 23545 25513 23579
rect 25547 23545 25559 23579
rect 25501 23539 25559 23545
rect 26697 23579 26755 23585
rect 26697 23545 26709 23579
rect 26743 23576 26755 23579
rect 27614 23576 27620 23588
rect 26743 23548 27620 23576
rect 26743 23545 26755 23548
rect 26697 23539 26755 23545
rect 17604 23480 18460 23508
rect 18693 23511 18751 23517
rect 18693 23477 18705 23511
rect 18739 23508 18751 23511
rect 19334 23508 19340 23520
rect 18739 23480 19340 23508
rect 18739 23477 18751 23480
rect 18693 23471 18751 23477
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 19610 23468 19616 23520
rect 19668 23468 19674 23520
rect 22462 23468 22468 23520
rect 22520 23508 22526 23520
rect 23750 23508 23756 23520
rect 22520 23480 23756 23508
rect 22520 23468 22526 23480
rect 23750 23468 23756 23480
rect 23808 23468 23814 23520
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25130 23508 25136 23520
rect 25004 23480 25136 23508
rect 25004 23468 25010 23480
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 25406 23468 25412 23520
rect 25464 23508 25470 23520
rect 25516 23508 25544 23539
rect 27614 23536 27620 23548
rect 27672 23536 27678 23588
rect 28718 23536 28724 23588
rect 28776 23536 28782 23588
rect 29733 23579 29791 23585
rect 29733 23545 29745 23579
rect 29779 23545 29791 23579
rect 30392 23576 30420 23607
rect 30466 23604 30472 23656
rect 30524 23644 30530 23656
rect 31021 23647 31079 23653
rect 31021 23644 31033 23647
rect 30524 23616 31033 23644
rect 30524 23604 30530 23616
rect 31021 23613 31033 23616
rect 31067 23644 31079 23647
rect 31110 23644 31116 23656
rect 31067 23616 31116 23644
rect 31067 23613 31079 23616
rect 31021 23607 31079 23613
rect 31110 23604 31116 23616
rect 31168 23604 31174 23656
rect 31849 23647 31907 23653
rect 31849 23644 31861 23647
rect 31726 23616 31861 23644
rect 31726 23576 31754 23616
rect 31849 23613 31861 23616
rect 31895 23613 31907 23647
rect 31849 23607 31907 23613
rect 33870 23604 33876 23656
rect 33928 23604 33934 23656
rect 36538 23604 36544 23656
rect 36596 23644 36602 23656
rect 37829 23647 37887 23653
rect 37829 23644 37841 23647
rect 36596 23616 37841 23644
rect 36596 23604 36602 23616
rect 37829 23613 37841 23616
rect 37875 23613 37887 23647
rect 37829 23607 37887 23613
rect 30392 23548 31754 23576
rect 29733 23539 29791 23545
rect 25464 23480 25544 23508
rect 25464 23468 25470 23480
rect 26970 23468 26976 23520
rect 27028 23468 27034 23520
rect 27801 23511 27859 23517
rect 27801 23477 27813 23511
rect 27847 23508 27859 23511
rect 27982 23508 27988 23520
rect 27847 23480 27988 23508
rect 27847 23477 27859 23480
rect 27801 23471 27859 23477
rect 27982 23468 27988 23480
rect 28040 23468 28046 23520
rect 28534 23468 28540 23520
rect 28592 23468 28598 23520
rect 28736 23508 28764 23536
rect 29748 23508 29776 23539
rect 28736 23480 29776 23508
rect 33318 23468 33324 23520
rect 33376 23468 33382 23520
rect 35437 23511 35495 23517
rect 35437 23477 35449 23511
rect 35483 23508 35495 23511
rect 35894 23508 35900 23520
rect 35483 23480 35900 23508
rect 35483 23477 35495 23480
rect 35437 23471 35495 23477
rect 35894 23468 35900 23480
rect 35952 23468 35958 23520
rect 36446 23468 36452 23520
rect 36504 23508 36510 23520
rect 38197 23511 38255 23517
rect 38197 23508 38209 23511
rect 36504 23480 38209 23508
rect 36504 23468 36510 23480
rect 38197 23477 38209 23480
rect 38243 23477 38255 23511
rect 38197 23471 38255 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 4614 23264 4620 23316
rect 4672 23264 4678 23316
rect 4706 23264 4712 23316
rect 4764 23304 4770 23316
rect 5445 23307 5503 23313
rect 5445 23304 5457 23307
rect 4764 23276 5457 23304
rect 4764 23264 4770 23276
rect 5445 23273 5457 23276
rect 5491 23273 5503 23307
rect 5445 23267 5503 23273
rect 6822 23264 6828 23316
rect 6880 23264 6886 23316
rect 7650 23304 7656 23316
rect 7208 23276 7656 23304
rect 4246 23236 4252 23248
rect 3988 23208 4252 23236
rect 3988 23177 4016 23208
rect 4246 23196 4252 23208
rect 4304 23196 4310 23248
rect 4338 23196 4344 23248
rect 4396 23236 4402 23248
rect 4396 23208 6040 23236
rect 4396 23196 4402 23208
rect 3973 23171 4031 23177
rect 3973 23137 3985 23171
rect 4019 23137 4031 23171
rect 3973 23131 4031 23137
rect 4065 23171 4123 23177
rect 4065 23137 4077 23171
rect 4111 23168 4123 23171
rect 4111 23140 4936 23168
rect 4111 23137 4123 23140
rect 4065 23131 4123 23137
rect 2038 23060 2044 23112
rect 2096 23100 2102 23112
rect 2225 23103 2283 23109
rect 2225 23100 2237 23103
rect 2096 23072 2237 23100
rect 2096 23060 2102 23072
rect 2225 23069 2237 23072
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2492 23103 2550 23109
rect 2492 23069 2504 23103
rect 2538 23100 2550 23103
rect 3786 23100 3792 23112
rect 2538 23072 3792 23100
rect 2538 23069 2550 23072
rect 2492 23063 2550 23069
rect 3786 23060 3792 23072
rect 3844 23060 3850 23112
rect 4154 23060 4160 23112
rect 4212 23060 4218 23112
rect 4430 23032 4436 23044
rect 3620 23004 4436 23032
rect 3620 22973 3648 23004
rect 4430 22992 4436 23004
rect 4488 23032 4494 23044
rect 4798 23032 4804 23044
rect 4488 23004 4804 23032
rect 4488 22992 4494 23004
rect 4798 22992 4804 23004
rect 4856 22992 4862 23044
rect 4908 23032 4936 23140
rect 5166 23128 5172 23180
rect 5224 23128 5230 23180
rect 6012 23177 6040 23208
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23137 6055 23171
rect 5997 23131 6055 23137
rect 6273 23171 6331 23177
rect 6273 23137 6285 23171
rect 6319 23168 6331 23171
rect 6914 23168 6920 23180
rect 6319 23140 6920 23168
rect 6319 23137 6331 23140
rect 6273 23131 6331 23137
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7208 23168 7236 23276
rect 7650 23264 7656 23276
rect 7708 23304 7714 23316
rect 7708 23276 8524 23304
rect 7708 23264 7714 23276
rect 8386 23236 8392 23248
rect 8036 23208 8392 23236
rect 7374 23168 7380 23180
rect 7208 23140 7380 23168
rect 7374 23128 7380 23140
rect 7432 23168 7438 23180
rect 7837 23171 7895 23177
rect 7432 23140 7604 23168
rect 7432 23128 7438 23140
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23100 5043 23103
rect 5442 23100 5448 23112
rect 5031 23072 5448 23100
rect 5031 23069 5043 23072
rect 4985 23063 5043 23069
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 7576 23109 7604 23140
rect 7837 23137 7849 23171
rect 7883 23168 7895 23171
rect 8036 23168 8064 23208
rect 8386 23196 8392 23208
rect 8444 23196 8450 23248
rect 8496 23236 8524 23276
rect 8846 23264 8852 23316
rect 8904 23304 8910 23316
rect 8941 23307 8999 23313
rect 8941 23304 8953 23307
rect 8904 23276 8953 23304
rect 8904 23264 8910 23276
rect 8941 23273 8953 23276
rect 8987 23273 8999 23307
rect 8941 23267 8999 23273
rect 9582 23264 9588 23316
rect 9640 23304 9646 23316
rect 9953 23307 10011 23313
rect 9953 23304 9965 23307
rect 9640 23276 9965 23304
rect 9640 23264 9646 23276
rect 9953 23273 9965 23276
rect 9999 23273 10011 23307
rect 9953 23267 10011 23273
rect 10413 23307 10471 23313
rect 10413 23273 10425 23307
rect 10459 23304 10471 23307
rect 12710 23304 12716 23316
rect 10459 23276 12716 23304
rect 10459 23273 10471 23276
rect 10413 23267 10471 23273
rect 10428 23236 10456 23267
rect 12710 23264 12716 23276
rect 12768 23264 12774 23316
rect 13262 23304 13268 23316
rect 13188 23276 13268 23304
rect 8496 23208 10456 23236
rect 11977 23239 12035 23245
rect 11977 23205 11989 23239
rect 12023 23205 12035 23239
rect 11977 23199 12035 23205
rect 7883 23140 8064 23168
rect 8113 23171 8171 23177
rect 7883 23137 7895 23140
rect 7837 23131 7895 23137
rect 8113 23137 8125 23171
rect 8159 23168 8171 23171
rect 8159 23140 8432 23168
rect 8159 23137 8171 23140
rect 8113 23131 8171 23137
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23069 7619 23103
rect 7561 23063 7619 23069
rect 7659 23060 7665 23112
rect 7717 23109 7723 23112
rect 7717 23103 7757 23109
rect 7745 23069 7757 23103
rect 8404 23100 8432 23140
rect 8570 23128 8576 23180
rect 8628 23128 8634 23180
rect 8662 23128 8668 23180
rect 8720 23168 8726 23180
rect 8757 23171 8815 23177
rect 8757 23168 8769 23171
rect 8720 23140 8769 23168
rect 8720 23128 8726 23140
rect 8757 23137 8769 23140
rect 8803 23137 8815 23171
rect 8757 23131 8815 23137
rect 9582 23128 9588 23180
rect 9640 23128 9646 23180
rect 11992 23168 12020 23199
rect 12989 23171 13047 23177
rect 11992 23140 12940 23168
rect 12912 23112 12940 23140
rect 12989 23137 13001 23171
rect 13035 23168 13047 23171
rect 13188 23168 13216 23276
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 15194 23264 15200 23316
rect 15252 23304 15258 23316
rect 15473 23307 15531 23313
rect 15473 23304 15485 23307
rect 15252 23276 15485 23304
rect 15252 23264 15258 23276
rect 15473 23273 15485 23276
rect 15519 23273 15531 23307
rect 15473 23267 15531 23273
rect 13354 23236 13360 23248
rect 13280 23208 13360 23236
rect 13280 23177 13308 23208
rect 13354 23196 13360 23208
rect 13412 23236 13418 23248
rect 15378 23236 15384 23248
rect 13412 23208 15384 23236
rect 13412 23196 13418 23208
rect 15378 23196 15384 23208
rect 15436 23196 15442 23248
rect 13035 23140 13216 23168
rect 13265 23171 13323 23177
rect 13035 23137 13047 23140
rect 12989 23131 13047 23137
rect 13265 23137 13277 23171
rect 13311 23137 13323 23171
rect 13265 23131 13323 23137
rect 13722 23128 13728 23180
rect 13780 23168 13786 23180
rect 14645 23171 14703 23177
rect 14645 23168 14657 23171
rect 13780 23140 14657 23168
rect 13780 23128 13786 23140
rect 14645 23137 14657 23140
rect 14691 23137 14703 23171
rect 14645 23131 14703 23137
rect 8404 23072 8616 23100
rect 7717 23063 7757 23069
rect 7717 23060 7723 23063
rect 5077 23035 5135 23041
rect 5077 23032 5089 23035
rect 4908 23004 5089 23032
rect 5077 23001 5089 23004
rect 5123 23032 5135 23035
rect 5350 23032 5356 23044
rect 5123 23004 5356 23032
rect 5123 23001 5135 23004
rect 5077 22995 5135 23001
rect 5350 22992 5356 23004
rect 5408 22992 5414 23044
rect 8588 23032 8616 23072
rect 9306 23060 9312 23112
rect 9364 23060 9370 23112
rect 10226 23060 10232 23112
rect 10284 23100 10290 23112
rect 10597 23103 10655 23109
rect 10597 23100 10609 23103
rect 10284 23072 10609 23100
rect 10284 23060 10290 23072
rect 10597 23069 10609 23072
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 12710 23060 12716 23112
rect 12768 23060 12774 23112
rect 12894 23109 12900 23112
rect 12872 23103 12900 23109
rect 12872 23069 12884 23103
rect 12872 23063 12900 23069
rect 12894 23060 12900 23063
rect 12952 23060 12958 23112
rect 13906 23060 13912 23112
rect 13964 23060 13970 23112
rect 15488 23100 15516 23267
rect 15562 23264 15568 23316
rect 15620 23264 15626 23316
rect 16298 23264 16304 23316
rect 16356 23304 16362 23316
rect 16945 23307 17003 23313
rect 16945 23304 16957 23307
rect 16356 23276 16957 23304
rect 16356 23264 16362 23276
rect 16945 23273 16957 23276
rect 16991 23304 17003 23307
rect 17954 23304 17960 23316
rect 16991 23276 17960 23304
rect 16991 23273 17003 23276
rect 16945 23267 17003 23273
rect 17954 23264 17960 23276
rect 18012 23264 18018 23316
rect 18417 23307 18475 23313
rect 18417 23273 18429 23307
rect 18463 23304 18475 23307
rect 18598 23304 18604 23316
rect 18463 23276 18604 23304
rect 18463 23273 18475 23276
rect 18417 23267 18475 23273
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 25406 23304 25412 23316
rect 24136 23276 25412 23304
rect 15580 23236 15608 23264
rect 18690 23236 18696 23248
rect 15580 23208 18696 23236
rect 18690 23196 18696 23208
rect 18748 23196 18754 23248
rect 17862 23128 17868 23180
rect 17920 23168 17926 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 17920 23140 19441 23168
rect 17920 23128 17926 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19429 23131 19487 23137
rect 21821 23171 21879 23177
rect 21821 23137 21833 23171
rect 21867 23168 21879 23171
rect 22462 23168 22468 23180
rect 21867 23140 22468 23168
rect 21867 23137 21879 23140
rect 21821 23131 21879 23137
rect 22462 23128 22468 23140
rect 22520 23128 22526 23180
rect 22738 23128 22744 23180
rect 22796 23168 22802 23180
rect 24136 23177 24164 23276
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 26602 23304 26608 23316
rect 25976 23276 26608 23304
rect 23753 23171 23811 23177
rect 23753 23168 23765 23171
rect 22796 23140 23765 23168
rect 22796 23128 22802 23140
rect 23753 23137 23765 23140
rect 23799 23168 23811 23171
rect 24121 23171 24179 23177
rect 24121 23168 24133 23171
rect 23799 23140 24133 23168
rect 23799 23137 23811 23140
rect 23753 23131 23811 23137
rect 24121 23137 24133 23140
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 25682 23128 25688 23180
rect 25740 23168 25746 23180
rect 25976 23177 26004 23276
rect 26602 23264 26608 23276
rect 26660 23264 26666 23316
rect 27706 23264 27712 23316
rect 27764 23264 27770 23316
rect 29273 23307 29331 23313
rect 29273 23273 29285 23307
rect 29319 23304 29331 23307
rect 29362 23304 29368 23316
rect 29319 23276 29368 23304
rect 29319 23273 29331 23276
rect 29273 23267 29331 23273
rect 29362 23264 29368 23276
rect 29420 23264 29426 23316
rect 29549 23307 29607 23313
rect 29549 23273 29561 23307
rect 29595 23304 29607 23307
rect 30282 23304 30288 23316
rect 29595 23276 30288 23304
rect 29595 23273 29607 23276
rect 29549 23267 29607 23273
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 32582 23264 32588 23316
rect 32640 23264 32646 23316
rect 34698 23264 34704 23316
rect 34756 23264 34762 23316
rect 34790 23264 34796 23316
rect 34848 23304 34854 23316
rect 36446 23304 36452 23316
rect 34848 23276 36452 23304
rect 34848 23264 34854 23276
rect 36446 23264 36452 23276
rect 36504 23264 36510 23316
rect 36998 23304 37004 23316
rect 36924 23276 37004 23304
rect 31110 23196 31116 23248
rect 31168 23236 31174 23248
rect 35986 23236 35992 23248
rect 31168 23208 35992 23236
rect 31168 23196 31174 23208
rect 35986 23196 35992 23208
rect 36044 23196 36050 23248
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 25740 23140 25973 23168
rect 25740 23128 25746 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 26145 23171 26203 23177
rect 26145 23137 26157 23171
rect 26191 23168 26203 23171
rect 26234 23168 26240 23180
rect 26191 23140 26240 23168
rect 26191 23137 26203 23140
rect 26145 23131 26203 23137
rect 26234 23128 26240 23140
rect 26292 23128 26298 23180
rect 26970 23128 26976 23180
rect 27028 23168 27034 23180
rect 27249 23171 27307 23177
rect 27249 23168 27261 23171
rect 27028 23140 27261 23168
rect 27028 23128 27034 23140
rect 27249 23137 27261 23140
rect 27295 23137 27307 23171
rect 27249 23131 27307 23137
rect 32582 23128 32588 23180
rect 32640 23168 32646 23180
rect 34057 23171 34115 23177
rect 34057 23168 34069 23171
rect 32640 23140 34069 23168
rect 32640 23128 32646 23140
rect 34057 23137 34069 23140
rect 34103 23137 34115 23171
rect 34057 23131 34115 23137
rect 34606 23128 34612 23180
rect 34664 23168 34670 23180
rect 35253 23171 35311 23177
rect 35253 23168 35265 23171
rect 34664 23140 35265 23168
rect 34664 23128 34670 23140
rect 35253 23137 35265 23140
rect 35299 23137 35311 23171
rect 35253 23131 35311 23137
rect 35894 23128 35900 23180
rect 35952 23168 35958 23180
rect 36587 23171 36645 23177
rect 36587 23168 36599 23171
rect 35952 23140 36599 23168
rect 35952 23128 35958 23140
rect 36587 23137 36599 23140
rect 36633 23137 36645 23171
rect 36587 23131 36645 23137
rect 36725 23171 36783 23177
rect 36725 23137 36737 23171
rect 36771 23168 36783 23171
rect 36924 23168 36952 23276
rect 36998 23264 37004 23276
rect 37056 23264 37062 23316
rect 36771 23140 36952 23168
rect 36771 23137 36783 23140
rect 36725 23131 36783 23137
rect 36998 23128 37004 23180
rect 37056 23128 37062 23180
rect 37645 23171 37703 23177
rect 37645 23137 37657 23171
rect 37691 23168 37703 23171
rect 37734 23168 37740 23180
rect 37691 23140 37740 23168
rect 37691 23137 37703 23140
rect 37645 23131 37703 23137
rect 37734 23128 37740 23140
rect 37792 23128 37798 23180
rect 15654 23100 15660 23112
rect 15488 23072 15660 23100
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 19610 23100 19616 23112
rect 18095 23072 19616 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 19610 23060 19616 23072
rect 19668 23060 19674 23112
rect 21266 23060 21272 23112
rect 21324 23060 21330 23112
rect 22094 23060 22100 23112
rect 22152 23100 22158 23112
rect 23017 23103 23075 23109
rect 23017 23100 23029 23103
rect 22152 23072 23029 23100
rect 22152 23060 22158 23072
rect 23017 23069 23029 23072
rect 23063 23069 23075 23103
rect 23017 23063 23075 23069
rect 23382 23060 23388 23112
rect 23440 23100 23446 23112
rect 24397 23103 24455 23109
rect 24397 23100 24409 23103
rect 23440 23072 24409 23100
rect 23440 23060 23446 23072
rect 24397 23069 24409 23072
rect 24443 23069 24455 23103
rect 24397 23063 24455 23069
rect 27890 23060 27896 23112
rect 27948 23060 27954 23112
rect 27982 23060 27988 23112
rect 28040 23100 28046 23112
rect 28149 23103 28207 23109
rect 28149 23100 28161 23103
rect 28040 23072 28161 23100
rect 28040 23060 28046 23072
rect 28149 23069 28161 23072
rect 28195 23069 28207 23103
rect 28149 23063 28207 23069
rect 30929 23103 30987 23109
rect 30929 23069 30941 23103
rect 30975 23100 30987 23103
rect 32306 23100 32312 23112
rect 30975 23072 32312 23100
rect 30975 23069 30987 23072
rect 30929 23063 30987 23069
rect 32306 23060 32312 23072
rect 32364 23060 32370 23112
rect 32766 23060 32772 23112
rect 32824 23100 32830 23112
rect 33229 23103 33287 23109
rect 33229 23100 33241 23103
rect 32824 23072 33241 23100
rect 32824 23060 32830 23072
rect 33229 23069 33241 23072
rect 33275 23069 33287 23103
rect 33229 23063 33287 23069
rect 35069 23103 35127 23109
rect 35069 23069 35081 23103
rect 35115 23100 35127 23103
rect 35342 23100 35348 23112
rect 35115 23072 35348 23100
rect 35115 23069 35127 23072
rect 35069 23063 35127 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 36446 23060 36452 23112
rect 36504 23060 36510 23112
rect 37458 23060 37464 23112
rect 37516 23060 37522 23112
rect 38381 23103 38439 23109
rect 38381 23069 38393 23103
rect 38427 23069 38439 23103
rect 38381 23063 38439 23069
rect 8588 23004 9904 23032
rect 9876 22976 9904 23004
rect 10686 22992 10692 23044
rect 10744 23032 10750 23044
rect 10842 23035 10900 23041
rect 10842 23032 10854 23035
rect 10744 23004 10854 23032
rect 10744 22992 10750 23004
rect 10842 23001 10854 23004
rect 10888 23001 10900 23035
rect 10842 22995 10900 23001
rect 22005 23035 22063 23041
rect 22005 23001 22017 23035
rect 22051 23032 22063 23035
rect 23290 23032 23296 23044
rect 22051 23004 23296 23032
rect 22051 23001 22063 23004
rect 22005 22995 22063 23001
rect 23290 22992 23296 23004
rect 23348 22992 23354 23044
rect 24664 23035 24722 23041
rect 24664 23001 24676 23035
rect 24710 23032 24722 23035
rect 26050 23032 26056 23044
rect 24710 23004 26056 23032
rect 24710 23001 24722 23004
rect 24664 22995 24722 23001
rect 26050 22992 26056 23004
rect 26108 22992 26114 23044
rect 26326 22992 26332 23044
rect 26384 23032 26390 23044
rect 26697 23035 26755 23041
rect 26697 23032 26709 23035
rect 26384 23004 26709 23032
rect 26384 22992 26390 23004
rect 26697 23001 26709 23004
rect 26743 23001 26755 23035
rect 26697 22995 26755 23001
rect 30684 23035 30742 23041
rect 30684 23001 30696 23035
rect 30730 23032 30742 23035
rect 31846 23032 31852 23044
rect 30730 23004 31852 23032
rect 30730 23001 30742 23004
rect 30684 22995 30742 23001
rect 31846 22992 31852 23004
rect 31904 22992 31910 23044
rect 33594 22992 33600 23044
rect 33652 23032 33658 23044
rect 33873 23035 33931 23041
rect 33873 23032 33885 23035
rect 33652 23004 33885 23032
rect 33652 22992 33658 23004
rect 33873 23001 33885 23004
rect 33919 23032 33931 23035
rect 33919 23004 35204 23032
rect 33919 23001 33931 23004
rect 33873 22995 33931 23001
rect 3605 22967 3663 22973
rect 3605 22933 3617 22967
rect 3651 22933 3663 22967
rect 3605 22927 3663 22933
rect 4522 22924 4528 22976
rect 4580 22924 4586 22976
rect 6914 22924 6920 22976
rect 6972 22924 6978 22976
rect 7006 22924 7012 22976
rect 7064 22964 7070 22976
rect 9401 22967 9459 22973
rect 9401 22964 9413 22967
rect 7064 22936 9413 22964
rect 7064 22924 7070 22936
rect 9401 22933 9413 22936
rect 9447 22933 9459 22967
rect 9401 22927 9459 22933
rect 9858 22924 9864 22976
rect 9916 22924 9922 22976
rect 12069 22967 12127 22973
rect 12069 22933 12081 22967
rect 12115 22964 12127 22967
rect 13170 22964 13176 22976
rect 12115 22936 13176 22964
rect 12115 22933 12127 22936
rect 12069 22927 12127 22933
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 14090 22924 14096 22976
rect 14148 22924 14154 22976
rect 17954 22924 17960 22976
rect 18012 22964 18018 22976
rect 18506 22964 18512 22976
rect 18012 22936 18512 22964
rect 18012 22924 18018 22936
rect 18506 22924 18512 22936
rect 18564 22924 18570 22976
rect 20714 22924 20720 22976
rect 20772 22924 20778 22976
rect 21910 22924 21916 22976
rect 21968 22924 21974 22976
rect 22370 22924 22376 22976
rect 22428 22924 22434 22976
rect 22462 22924 22468 22976
rect 22520 22924 22526 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23934 22964 23940 22976
rect 23532 22936 23940 22964
rect 23532 22924 23538 22936
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 25774 22924 25780 22976
rect 25832 22924 25838 22976
rect 26234 22924 26240 22976
rect 26292 22924 26298 22976
rect 26602 22924 26608 22976
rect 26660 22924 26666 22976
rect 32582 22924 32588 22976
rect 32640 22964 32646 22976
rect 32677 22967 32735 22973
rect 32677 22964 32689 22967
rect 32640 22936 32689 22964
rect 32640 22924 32646 22936
rect 32677 22933 32689 22936
rect 32723 22933 32735 22967
rect 32677 22927 32735 22933
rect 33042 22924 33048 22976
rect 33100 22964 33106 22976
rect 33505 22967 33563 22973
rect 33505 22964 33517 22967
rect 33100 22936 33517 22964
rect 33100 22924 33106 22936
rect 33505 22933 33517 22936
rect 33551 22933 33563 22967
rect 33505 22927 33563 22933
rect 33962 22924 33968 22976
rect 34020 22924 34026 22976
rect 35176 22973 35204 23004
rect 35161 22967 35219 22973
rect 35161 22933 35173 22967
rect 35207 22964 35219 22967
rect 35526 22964 35532 22976
rect 35207 22936 35532 22964
rect 35207 22933 35219 22936
rect 35161 22927 35219 22933
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 35805 22967 35863 22973
rect 35805 22933 35817 22967
rect 35851 22964 35863 22967
rect 36906 22964 36912 22976
rect 35851 22936 36912 22964
rect 35851 22933 35863 22936
rect 35805 22927 35863 22933
rect 36906 22924 36912 22936
rect 36964 22924 36970 22976
rect 37182 22924 37188 22976
rect 37240 22964 37246 22976
rect 37737 22967 37795 22973
rect 37737 22964 37749 22967
rect 37240 22936 37749 22964
rect 37240 22924 37246 22936
rect 37737 22933 37749 22936
rect 37783 22933 37795 22967
rect 38396 22964 38424 23063
rect 38396 22936 38884 22964
rect 37737 22927 37795 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 4522 22720 4528 22772
rect 4580 22760 4586 22772
rect 4580 22732 5948 22760
rect 4580 22720 4586 22732
rect 2216 22695 2274 22701
rect 2216 22661 2228 22695
rect 2262 22692 2274 22695
rect 2498 22692 2504 22704
rect 2262 22664 2504 22692
rect 2262 22661 2274 22664
rect 2216 22655 2274 22661
rect 2498 22652 2504 22664
rect 2556 22652 2562 22704
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22624 2007 22627
rect 2038 22624 2044 22636
rect 1995 22596 2044 22624
rect 1995 22593 2007 22596
rect 1949 22587 2007 22593
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 4338 22584 4344 22636
rect 4396 22584 4402 22636
rect 4430 22584 4436 22636
rect 4488 22633 4494 22636
rect 5920 22633 5948 22732
rect 6362 22720 6368 22772
rect 6420 22760 6426 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6420 22732 6561 22760
rect 6420 22720 6426 22732
rect 6549 22729 6561 22732
rect 6595 22729 6607 22763
rect 6549 22723 6607 22729
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 6972 22732 8493 22760
rect 6972 22720 6978 22732
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 8481 22723 8539 22729
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10318 22760 10324 22772
rect 9916 22732 10324 22760
rect 9916 22720 9922 22732
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 10686 22720 10692 22772
rect 10744 22720 10750 22772
rect 12986 22720 12992 22772
rect 13044 22720 13050 22772
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 14090 22760 14096 22772
rect 13403 22732 14096 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 17862 22720 17868 22772
rect 17920 22720 17926 22772
rect 18049 22763 18107 22769
rect 18049 22729 18061 22763
rect 18095 22760 18107 22763
rect 18230 22760 18236 22772
rect 18095 22732 18236 22760
rect 18095 22729 18107 22732
rect 18049 22723 18107 22729
rect 18230 22720 18236 22732
rect 18288 22720 18294 22772
rect 20901 22763 20959 22769
rect 20901 22729 20913 22763
rect 20947 22760 20959 22763
rect 21266 22760 21272 22772
rect 20947 22732 21272 22760
rect 20947 22729 20959 22732
rect 20901 22723 20959 22729
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 21358 22720 21364 22772
rect 21416 22760 21422 22772
rect 21910 22760 21916 22772
rect 21416 22732 21916 22760
rect 21416 22720 21422 22732
rect 21910 22720 21916 22732
rect 21968 22760 21974 22772
rect 22189 22763 22247 22769
rect 22189 22760 22201 22763
rect 21968 22732 22201 22760
rect 21968 22720 21974 22732
rect 22189 22729 22201 22732
rect 22235 22729 22247 22763
rect 22189 22723 22247 22729
rect 22281 22763 22339 22769
rect 22281 22729 22293 22763
rect 22327 22760 22339 22763
rect 22462 22760 22468 22772
rect 22327 22732 22468 22760
rect 22327 22729 22339 22732
rect 22281 22723 22339 22729
rect 22462 22720 22468 22732
rect 22520 22720 22526 22772
rect 25222 22720 25228 22772
rect 25280 22760 25286 22772
rect 25961 22763 26019 22769
rect 25961 22760 25973 22763
rect 25280 22732 25973 22760
rect 25280 22720 25286 22732
rect 25961 22729 25973 22732
rect 26007 22729 26019 22763
rect 25961 22723 26019 22729
rect 26050 22720 26056 22772
rect 26108 22720 26114 22772
rect 26326 22720 26332 22772
rect 26384 22720 26390 22772
rect 26602 22720 26608 22772
rect 26660 22720 26666 22772
rect 27614 22720 27620 22772
rect 27672 22720 27678 22772
rect 28077 22763 28135 22769
rect 28077 22729 28089 22763
rect 28123 22760 28135 22763
rect 28534 22760 28540 22772
rect 28123 22732 28540 22760
rect 28123 22729 28135 22732
rect 28077 22723 28135 22729
rect 28534 22720 28540 22732
rect 28592 22720 28598 22772
rect 28629 22763 28687 22769
rect 28629 22729 28641 22763
rect 28675 22760 28687 22763
rect 30098 22760 30104 22772
rect 28675 22732 30104 22760
rect 28675 22729 28687 22732
rect 28629 22723 28687 22729
rect 30098 22720 30104 22732
rect 30156 22720 30162 22772
rect 33778 22720 33784 22772
rect 33836 22720 33842 22772
rect 35342 22760 35348 22772
rect 35176 22732 35348 22760
rect 7558 22652 7564 22704
rect 7616 22692 7622 22704
rect 7662 22695 7720 22701
rect 7662 22692 7674 22695
rect 7616 22664 7674 22692
rect 7616 22652 7622 22664
rect 7662 22661 7674 22664
rect 7708 22661 7720 22695
rect 8389 22695 8447 22701
rect 8389 22692 8401 22695
rect 7662 22655 7720 22661
rect 7760 22664 8401 22692
rect 4488 22627 4516 22633
rect 4504 22593 4516 22627
rect 4488 22587 4516 22593
rect 5905 22627 5963 22633
rect 5905 22593 5917 22627
rect 5951 22593 5963 22627
rect 7760 22624 7788 22664
rect 8389 22661 8401 22664
rect 8435 22661 8447 22695
rect 8389 22655 8447 22661
rect 8570 22652 8576 22704
rect 8628 22692 8634 22704
rect 11606 22692 11612 22704
rect 8628 22664 11612 22692
rect 8628 22652 8634 22664
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 11790 22701 11796 22704
rect 11784 22692 11796 22701
rect 11751 22664 11796 22692
rect 11784 22655 11796 22664
rect 11790 22652 11796 22655
rect 11848 22652 11854 22704
rect 12434 22652 12440 22704
rect 12492 22692 12498 22704
rect 13449 22695 13507 22701
rect 13449 22692 13461 22695
rect 12492 22664 13461 22692
rect 12492 22652 12498 22664
rect 13449 22661 13461 22664
rect 13495 22692 13507 22695
rect 13630 22692 13636 22704
rect 13495 22664 13636 22692
rect 13495 22661 13507 22664
rect 13449 22655 13507 22661
rect 13630 22652 13636 22664
rect 13688 22652 13694 22704
rect 14001 22695 14059 22701
rect 14001 22661 14013 22695
rect 14047 22692 14059 22695
rect 17880 22692 17908 22720
rect 14047 22664 17908 22692
rect 14047 22661 14059 22664
rect 14001 22655 14059 22661
rect 5905 22587 5963 22593
rect 6840 22596 7788 22624
rect 4488 22584 4494 22587
rect 3421 22559 3479 22565
rect 3421 22525 3433 22559
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22556 3663 22559
rect 3970 22556 3976 22568
rect 3651 22528 3976 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 3329 22423 3387 22429
rect 3329 22389 3341 22423
rect 3375 22420 3387 22423
rect 3436 22420 3464 22519
rect 3970 22516 3976 22528
rect 4028 22516 4034 22568
rect 4617 22559 4675 22565
rect 4617 22525 4629 22559
rect 4663 22556 4675 22559
rect 5261 22559 5319 22565
rect 4663 22528 5212 22556
rect 4663 22525 4675 22528
rect 4617 22519 4675 22525
rect 3878 22448 3884 22500
rect 3936 22488 3942 22500
rect 4065 22491 4123 22497
rect 4065 22488 4077 22491
rect 3936 22460 4077 22488
rect 3936 22448 3942 22460
rect 4065 22457 4077 22460
rect 4111 22457 4123 22491
rect 5184 22488 5212 22528
rect 5261 22525 5273 22559
rect 5307 22556 5319 22559
rect 6840 22556 6868 22596
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 7892 22596 7941 22624
rect 7892 22584 7898 22596
rect 7929 22593 7941 22596
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 8662 22584 8668 22636
rect 8720 22624 8726 22636
rect 9401 22627 9459 22633
rect 9401 22624 9413 22627
rect 8720 22596 9413 22624
rect 8720 22584 8726 22596
rect 9401 22593 9413 22596
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 10226 22584 10232 22636
rect 10284 22624 10290 22636
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10284 22596 11529 22624
rect 10284 22584 10290 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 13354 22624 13360 22636
rect 12584 22596 13360 22624
rect 12584 22584 12590 22596
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 5307 22528 6868 22556
rect 5307 22525 5319 22528
rect 5261 22519 5319 22525
rect 8110 22516 8116 22568
rect 8168 22556 8174 22568
rect 8570 22556 8576 22568
rect 8168 22528 8576 22556
rect 8168 22516 8174 22528
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 11330 22516 11336 22568
rect 11388 22516 11394 22568
rect 13262 22516 13268 22568
rect 13320 22516 13326 22568
rect 13633 22559 13691 22565
rect 13633 22525 13645 22559
rect 13679 22556 13691 22559
rect 14016 22556 14044 22655
rect 16298 22584 16304 22636
rect 16356 22624 16362 22636
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16356 22596 16681 22624
rect 16356 22584 16362 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16936 22627 16994 22633
rect 16936 22593 16948 22627
rect 16982 22624 16994 22627
rect 17678 22624 17684 22636
rect 16982 22596 17684 22624
rect 16982 22593 16994 22596
rect 16936 22587 16994 22593
rect 17678 22584 17684 22596
rect 17736 22584 17742 22636
rect 18248 22624 18276 22720
rect 22370 22652 22376 22704
rect 22428 22692 22434 22704
rect 24848 22695 24906 22701
rect 22428 22664 23244 22692
rect 22428 22652 22434 22664
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 18248 22596 18705 22624
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22624 21327 22627
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 21315 22596 22661 22624
rect 21315 22593 21327 22596
rect 21269 22587 21327 22593
rect 22649 22593 22661 22596
rect 22695 22593 22707 22627
rect 23216 22624 23244 22664
rect 24848 22661 24860 22695
rect 24894 22692 24906 22695
rect 26344 22692 26372 22720
rect 24894 22664 26372 22692
rect 24894 22661 24906 22664
rect 24848 22655 24906 22661
rect 23216 22596 23336 22624
rect 22649 22587 22707 22593
rect 13679 22528 14044 22556
rect 20809 22559 20867 22565
rect 13679 22525 13691 22528
rect 13633 22519 13691 22525
rect 20809 22525 20821 22559
rect 20855 22525 20867 22559
rect 20809 22519 20867 22525
rect 6178 22488 6184 22500
rect 5184 22460 6184 22488
rect 4065 22451 4123 22457
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 8754 22488 8760 22500
rect 7944 22460 8760 22488
rect 4614 22420 4620 22432
rect 3375 22392 4620 22420
rect 3375 22389 3387 22392
rect 3329 22383 3387 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 5350 22380 5356 22432
rect 5408 22380 5414 22432
rect 6196 22420 6224 22448
rect 7944 22420 7972 22460
rect 8754 22448 8760 22460
rect 8812 22448 8818 22500
rect 12897 22491 12955 22497
rect 12897 22457 12909 22491
rect 12943 22488 12955 22491
rect 13280 22488 13308 22516
rect 12943 22460 13308 22488
rect 12943 22457 12955 22460
rect 12897 22451 12955 22457
rect 6196 22392 7972 22420
rect 8018 22380 8024 22432
rect 8076 22380 8082 22432
rect 8294 22380 8300 22432
rect 8352 22420 8358 22432
rect 8849 22423 8907 22429
rect 8849 22420 8861 22423
rect 8352 22392 8861 22420
rect 8352 22380 8358 22392
rect 8849 22389 8861 22392
rect 8895 22389 8907 22423
rect 8849 22383 8907 22389
rect 9582 22380 9588 22432
rect 9640 22420 9646 22432
rect 13648 22420 13676 22519
rect 20824 22488 20852 22519
rect 21358 22516 21364 22568
rect 21416 22516 21422 22568
rect 21545 22559 21603 22565
rect 21545 22525 21557 22559
rect 21591 22556 21603 22559
rect 22465 22559 22523 22565
rect 21591 22528 21956 22556
rect 21591 22525 21603 22528
rect 21545 22519 21603 22525
rect 21821 22491 21879 22497
rect 21821 22488 21833 22491
rect 20824 22460 21833 22488
rect 21821 22457 21833 22460
rect 21867 22457 21879 22491
rect 21821 22451 21879 22457
rect 9640 22392 13676 22420
rect 9640 22380 9646 22392
rect 18138 22380 18144 22432
rect 18196 22380 18202 22432
rect 20162 22380 20168 22432
rect 20220 22380 20226 22432
rect 21928 22420 21956 22528
rect 22465 22525 22477 22559
rect 22511 22525 22523 22559
rect 22465 22519 22523 22525
rect 22480 22488 22508 22519
rect 22554 22516 22560 22568
rect 22612 22556 22618 22568
rect 23201 22559 23259 22565
rect 23201 22556 23213 22559
rect 22612 22528 23213 22556
rect 22612 22516 22618 22528
rect 23201 22525 23213 22528
rect 23247 22525 23259 22559
rect 23308 22556 23336 22596
rect 23382 22584 23388 22636
rect 23440 22624 23446 22636
rect 26620 22633 26648 22720
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 23440 22596 24593 22624
rect 23440 22584 23446 22596
rect 24581 22593 24593 22596
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 26605 22627 26663 22633
rect 26605 22593 26617 22627
rect 26651 22593 26663 22627
rect 27632 22624 27660 22720
rect 27890 22652 27896 22704
rect 27948 22692 27954 22704
rect 28902 22692 28908 22704
rect 27948 22664 28908 22692
rect 27948 22652 27954 22664
rect 28902 22652 28908 22664
rect 28960 22692 28966 22704
rect 28960 22664 30052 22692
rect 28960 22652 28966 22664
rect 28169 22627 28227 22633
rect 28169 22624 28181 22627
rect 27632 22596 28181 22624
rect 26605 22587 26663 22593
rect 28169 22593 28181 22596
rect 28215 22593 28227 22627
rect 28169 22587 28227 22593
rect 28626 22584 28632 22636
rect 28684 22584 28690 22636
rect 30024 22633 30052 22664
rect 30374 22652 30380 22704
rect 30432 22652 30438 22704
rect 35176 22692 35204 22732
rect 35342 22720 35348 22732
rect 35400 22760 35406 22772
rect 35618 22760 35624 22772
rect 35400 22732 35624 22760
rect 35400 22720 35406 22732
rect 35618 22720 35624 22732
rect 35676 22720 35682 22772
rect 36081 22763 36139 22769
rect 36081 22729 36093 22763
rect 36127 22760 36139 22763
rect 36538 22760 36544 22772
rect 36127 22732 36544 22760
rect 36127 22729 36139 22732
rect 36081 22723 36139 22729
rect 36538 22720 36544 22732
rect 36596 22720 36602 22772
rect 36630 22720 36636 22772
rect 36688 22720 36694 22772
rect 37090 22720 37096 22772
rect 37148 22720 37154 22772
rect 38013 22763 38071 22769
rect 38013 22729 38025 22763
rect 38059 22760 38071 22763
rect 38856 22760 38884 22936
rect 38059 22732 38884 22760
rect 38059 22729 38071 22732
rect 38013 22723 38071 22729
rect 32324 22664 35204 22692
rect 29753 22627 29811 22633
rect 29753 22593 29765 22627
rect 29799 22624 29811 22627
rect 30009 22627 30067 22633
rect 29799 22596 29960 22624
rect 29799 22593 29811 22596
rect 29753 22587 29811 22593
rect 23937 22559 23995 22565
rect 23937 22556 23949 22559
rect 23308 22528 23949 22556
rect 23201 22519 23259 22525
rect 23937 22525 23949 22528
rect 23983 22525 23995 22559
rect 23937 22519 23995 22525
rect 27709 22559 27767 22565
rect 27709 22525 27721 22559
rect 27755 22556 27767 22559
rect 27985 22559 28043 22565
rect 27985 22556 27997 22559
rect 27755 22528 27997 22556
rect 27755 22525 27767 22528
rect 27709 22519 27767 22525
rect 27985 22525 27997 22528
rect 28031 22556 28043 22559
rect 28644 22556 28672 22584
rect 28994 22556 29000 22568
rect 28031 22528 29000 22556
rect 28031 22525 28043 22528
rect 27985 22519 28043 22525
rect 28994 22516 29000 22528
rect 29052 22516 29058 22568
rect 29932 22556 29960 22596
rect 30009 22593 30021 22627
rect 30055 22593 30067 22627
rect 30009 22587 30067 22593
rect 30392 22556 30420 22652
rect 32324 22636 32352 22664
rect 32306 22584 32312 22636
rect 32364 22584 32370 22636
rect 32582 22633 32588 22636
rect 32576 22624 32588 22633
rect 32543 22596 32588 22624
rect 32576 22587 32588 22596
rect 32582 22584 32588 22587
rect 32640 22584 32646 22636
rect 35176 22633 35204 22664
rect 35526 22652 35532 22704
rect 35584 22692 35590 22704
rect 35713 22695 35771 22701
rect 35713 22692 35725 22695
rect 35584 22664 35725 22692
rect 35584 22652 35590 22664
rect 35713 22661 35725 22664
rect 35759 22692 35771 22695
rect 36446 22692 36452 22704
rect 35759 22664 36452 22692
rect 35759 22661 35771 22664
rect 35713 22655 35771 22661
rect 36446 22652 36452 22664
rect 36504 22692 36510 22704
rect 36725 22695 36783 22701
rect 36725 22692 36737 22695
rect 36504 22664 36737 22692
rect 36504 22652 36510 22664
rect 36725 22661 36737 22664
rect 36771 22661 36783 22695
rect 36725 22655 36783 22661
rect 34905 22627 34963 22633
rect 34905 22593 34917 22627
rect 34951 22624 34963 22627
rect 35161 22627 35219 22633
rect 34951 22596 35112 22624
rect 34951 22593 34963 22596
rect 34905 22587 34963 22593
rect 29932 22528 30420 22556
rect 35084 22556 35112 22596
rect 35161 22593 35173 22627
rect 35207 22593 35219 22627
rect 35161 22587 35219 22593
rect 35986 22584 35992 22636
rect 36044 22624 36050 22636
rect 36740 22624 36768 22655
rect 36906 22652 36912 22704
rect 36964 22692 36970 22704
rect 37550 22692 37556 22704
rect 36964 22664 37556 22692
rect 36964 22652 36970 22664
rect 37550 22652 37556 22664
rect 37608 22652 37614 22704
rect 36044 22596 36492 22624
rect 36740 22596 37596 22624
rect 36044 22584 36050 22596
rect 35084 22528 35204 22556
rect 23474 22488 23480 22500
rect 22480 22460 23480 22488
rect 23474 22448 23480 22460
rect 23532 22488 23538 22500
rect 24210 22488 24216 22500
rect 23532 22460 24216 22488
rect 23532 22448 23538 22460
rect 24210 22448 24216 22460
rect 24268 22448 24274 22500
rect 35176 22488 35204 22528
rect 35434 22516 35440 22568
rect 35492 22516 35498 22568
rect 35621 22559 35679 22565
rect 35621 22525 35633 22559
rect 35667 22556 35679 22559
rect 36354 22556 36360 22568
rect 35667 22528 36360 22556
rect 35667 22525 35679 22528
rect 35621 22519 35679 22525
rect 36354 22516 36360 22528
rect 36412 22516 36418 22568
rect 36464 22565 36492 22596
rect 36449 22559 36507 22565
rect 36449 22525 36461 22559
rect 36495 22556 36507 22559
rect 36722 22556 36728 22568
rect 36495 22528 36728 22556
rect 36495 22525 36507 22528
rect 36449 22519 36507 22525
rect 36722 22516 36728 22528
rect 36780 22516 36786 22568
rect 37274 22516 37280 22568
rect 37332 22556 37338 22568
rect 37568 22565 37596 22596
rect 37642 22584 37648 22636
rect 37700 22584 37706 22636
rect 37369 22559 37427 22565
rect 37369 22556 37381 22559
rect 37332 22528 37381 22556
rect 37332 22516 37338 22528
rect 37369 22525 37381 22528
rect 37415 22525 37427 22559
rect 37369 22519 37427 22525
rect 37553 22559 37611 22565
rect 37553 22525 37565 22559
rect 37599 22556 37611 22559
rect 37734 22556 37740 22568
rect 37599 22528 37740 22556
rect 37599 22525 37611 22528
rect 37553 22519 37611 22525
rect 37734 22516 37740 22528
rect 37792 22516 37798 22568
rect 35710 22488 35716 22500
rect 35176 22460 35716 22488
rect 35710 22448 35716 22460
rect 35768 22448 35774 22500
rect 22186 22420 22192 22432
rect 21928 22392 22192 22420
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 22830 22380 22836 22432
rect 22888 22420 22894 22432
rect 23385 22423 23443 22429
rect 23385 22420 23397 22423
rect 22888 22392 23397 22420
rect 22888 22380 22894 22392
rect 23385 22389 23397 22392
rect 23431 22389 23443 22423
rect 23385 22383 23443 22389
rect 28534 22380 28540 22432
rect 28592 22380 28598 22432
rect 30374 22380 30380 22432
rect 30432 22380 30438 22432
rect 33689 22423 33747 22429
rect 33689 22389 33701 22423
rect 33735 22420 33747 22423
rect 33870 22420 33876 22432
rect 33735 22392 33876 22420
rect 33735 22389 33747 22392
rect 33689 22383 33747 22389
rect 33870 22380 33876 22392
rect 33928 22420 33934 22432
rect 34514 22420 34520 22432
rect 33928 22392 34520 22420
rect 33928 22380 33934 22392
rect 34514 22380 34520 22392
rect 34572 22380 34578 22432
rect 35434 22380 35440 22432
rect 35492 22420 35498 22432
rect 35618 22420 35624 22432
rect 35492 22392 35624 22420
rect 35492 22380 35498 22392
rect 35618 22380 35624 22392
rect 35676 22420 35682 22432
rect 38289 22423 38347 22429
rect 38289 22420 38301 22423
rect 35676 22392 38301 22420
rect 35676 22380 35682 22392
rect 38289 22389 38301 22392
rect 38335 22389 38347 22423
rect 38289 22383 38347 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3789 22219 3847 22225
rect 3789 22185 3801 22219
rect 3835 22216 3847 22219
rect 3970 22216 3976 22228
rect 3835 22188 3976 22216
rect 3835 22185 3847 22188
rect 3789 22179 3847 22185
rect 3970 22176 3976 22188
rect 4028 22176 4034 22228
rect 5626 22216 5632 22228
rect 4172 22188 5632 22216
rect 3878 22108 3884 22160
rect 3936 22148 3942 22160
rect 4172 22148 4200 22188
rect 5626 22176 5632 22188
rect 5684 22216 5690 22228
rect 5902 22216 5908 22228
rect 5684 22188 5908 22216
rect 5684 22176 5690 22188
rect 5902 22176 5908 22188
rect 5960 22176 5966 22228
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7377 22219 7435 22225
rect 7377 22216 7389 22219
rect 6972 22188 7389 22216
rect 6972 22176 6978 22188
rect 7377 22185 7389 22188
rect 7423 22185 7435 22219
rect 7377 22179 7435 22185
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 11793 22219 11851 22225
rect 11793 22216 11805 22219
rect 11388 22188 11805 22216
rect 11388 22176 11394 22188
rect 11793 22185 11805 22188
rect 11839 22185 11851 22219
rect 11793 22179 11851 22185
rect 16761 22219 16819 22225
rect 16761 22185 16773 22219
rect 16807 22216 16819 22219
rect 16850 22216 16856 22228
rect 16807 22188 16856 22216
rect 16807 22185 16819 22188
rect 16761 22179 16819 22185
rect 16850 22176 16856 22188
rect 16908 22176 16914 22228
rect 17678 22176 17684 22228
rect 17736 22176 17742 22228
rect 18046 22176 18052 22228
rect 18104 22216 18110 22228
rect 18104 22188 19334 22216
rect 18104 22176 18110 22188
rect 3936 22120 4200 22148
rect 10888 22120 12388 22148
rect 3936 22108 3942 22120
rect 10888 22092 10916 22120
rect 5166 22040 5172 22092
rect 5224 22080 5230 22092
rect 7834 22080 7840 22092
rect 5224 22052 7840 22080
rect 5224 22040 5230 22052
rect 7834 22040 7840 22052
rect 7892 22040 7898 22092
rect 7926 22040 7932 22092
rect 7984 22080 7990 22092
rect 8021 22083 8079 22089
rect 8021 22080 8033 22083
rect 7984 22052 8033 22080
rect 7984 22040 7990 22052
rect 8021 22049 8033 22052
rect 8067 22080 8079 22083
rect 8478 22080 8484 22092
rect 8067 22052 8484 22080
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 8478 22040 8484 22052
rect 8536 22040 8542 22092
rect 10870 22040 10876 22092
rect 10928 22040 10934 22092
rect 12360 22089 12388 22120
rect 12345 22083 12403 22089
rect 12345 22049 12357 22083
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12894 22040 12900 22092
rect 12952 22080 12958 22092
rect 13173 22083 13231 22089
rect 13173 22080 13185 22083
rect 12952 22052 13185 22080
rect 12952 22040 12958 22052
rect 13173 22049 13185 22052
rect 13219 22049 13231 22083
rect 16868 22080 16896 22176
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16868 22052 16957 22080
rect 13173 22043 13231 22049
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 18138 22080 18144 22092
rect 17175 22052 18144 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 19306 22080 19334 22188
rect 21818 22176 21824 22228
rect 21876 22216 21882 22228
rect 21876 22188 24072 22216
rect 21876 22176 21882 22188
rect 24044 22160 24072 22188
rect 25682 22176 25688 22228
rect 25740 22176 25746 22228
rect 26234 22176 26240 22228
rect 26292 22216 26298 22228
rect 26697 22219 26755 22225
rect 26697 22216 26709 22219
rect 26292 22188 26709 22216
rect 26292 22176 26298 22188
rect 26697 22185 26709 22188
rect 26743 22185 26755 22219
rect 28810 22216 28816 22228
rect 26697 22179 26755 22185
rect 28368 22188 28816 22216
rect 22554 22148 22560 22160
rect 22287 22120 22560 22148
rect 19705 22083 19763 22089
rect 19705 22080 19717 22083
rect 19306 22052 19717 22080
rect 19705 22049 19717 22052
rect 19751 22049 19763 22083
rect 22287 22080 22315 22120
rect 22554 22108 22560 22120
rect 22612 22108 22618 22160
rect 23014 22108 23020 22160
rect 23072 22148 23078 22160
rect 23072 22120 23796 22148
rect 23072 22108 23078 22120
rect 19705 22043 19763 22049
rect 22020 22052 22315 22080
rect 22393 22083 22451 22089
rect 2038 21972 2044 22024
rect 2096 22012 2102 22024
rect 2225 22015 2283 22021
rect 2225 22012 2237 22015
rect 2096 21984 2237 22012
rect 2096 21972 2102 21984
rect 2225 21981 2237 21984
rect 2271 22012 2283 22015
rect 5184 22012 5212 22040
rect 2271 21984 5212 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7745 22015 7803 22021
rect 7745 22012 7757 22015
rect 7156 21984 7757 22012
rect 7156 21972 7162 21984
rect 7745 21981 7757 21984
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 2492 21947 2550 21953
rect 2492 21913 2504 21947
rect 2538 21944 2550 21947
rect 2866 21944 2872 21956
rect 2538 21916 2872 21944
rect 2538 21913 2550 21916
rect 2492 21907 2550 21913
rect 2866 21904 2872 21916
rect 2924 21904 2930 21956
rect 4062 21904 4068 21956
rect 4120 21904 4126 21956
rect 4924 21947 4982 21953
rect 4924 21913 4936 21947
rect 4970 21944 4982 21947
rect 5350 21944 5356 21956
rect 4970 21916 5356 21944
rect 4970 21913 4982 21916
rect 4924 21907 4982 21913
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 5442 21904 5448 21956
rect 5500 21944 5506 21956
rect 5902 21944 5908 21956
rect 5500 21916 5908 21944
rect 5500 21904 5506 21916
rect 5902 21904 5908 21916
rect 5960 21904 5966 21956
rect 6270 21904 6276 21956
rect 6328 21944 6334 21956
rect 9950 21944 9956 21956
rect 6328 21916 9956 21944
rect 6328 21904 6334 21916
rect 9950 21904 9956 21916
rect 10008 21904 10014 21956
rect 3605 21879 3663 21885
rect 3605 21845 3617 21879
rect 3651 21876 3663 21879
rect 4080 21876 4108 21904
rect 3651 21848 4108 21876
rect 5997 21879 6055 21885
rect 3651 21845 3663 21848
rect 3605 21839 3663 21845
rect 5997 21845 6009 21879
rect 6043 21876 6055 21879
rect 6178 21876 6184 21888
rect 6043 21848 6184 21876
rect 6043 21845 6055 21848
rect 5997 21839 6055 21845
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 7837 21879 7895 21885
rect 7837 21845 7849 21879
rect 7883 21876 7895 21879
rect 8294 21876 8300 21888
rect 7883 21848 8300 21876
rect 7883 21845 7895 21848
rect 7837 21839 7895 21845
rect 8294 21836 8300 21848
rect 8352 21836 8358 21888
rect 10318 21836 10324 21888
rect 10376 21876 10382 21888
rect 10888 21885 10916 22040
rect 11606 21972 11612 22024
rect 11664 21972 11670 22024
rect 19978 22021 19984 22024
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 19972 21975 19984 22021
rect 12161 21947 12219 21953
rect 12161 21913 12173 21947
rect 12207 21944 12219 21947
rect 12621 21947 12679 21953
rect 12621 21944 12633 21947
rect 12207 21916 12633 21944
rect 12207 21913 12219 21916
rect 12161 21907 12219 21913
rect 12621 21913 12633 21916
rect 12667 21913 12679 21947
rect 12621 21907 12679 21913
rect 10873 21879 10931 21885
rect 10873 21876 10885 21879
rect 10376 21848 10885 21876
rect 10376 21836 10382 21848
rect 10873 21845 10885 21848
rect 10919 21845 10931 21879
rect 10873 21839 10931 21845
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 12253 21879 12311 21885
rect 12253 21845 12265 21879
rect 12299 21876 12311 21879
rect 12434 21876 12440 21888
rect 12299 21848 12440 21876
rect 12299 21845 12311 21848
rect 12253 21839 12311 21845
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 17218 21836 17224 21888
rect 17276 21836 17282 21888
rect 17589 21879 17647 21885
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 18248 21876 18276 21975
rect 19978 21972 19984 21975
rect 20036 21972 20042 22024
rect 21818 21972 21824 22024
rect 21876 21972 21882 22024
rect 22020 22021 22048 22052
rect 22393 22049 22405 22083
rect 22439 22080 22451 22083
rect 22738 22080 22744 22092
rect 22439 22052 22744 22080
rect 22439 22049 22451 22052
rect 22393 22043 22451 22049
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 22833 22083 22891 22089
rect 22833 22049 22845 22083
rect 22879 22080 22891 22083
rect 22879 22052 23152 22080
rect 22879 22049 22891 22052
rect 22833 22043 22891 22049
rect 21980 22015 22048 22021
rect 21980 21981 21992 22015
rect 22026 21984 22048 22015
rect 22026 21981 22038 21984
rect 21980 21975 22038 21981
rect 22094 21972 22100 22024
rect 22152 21972 22158 22024
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 21100 21916 21312 21944
rect 17635 21848 18276 21876
rect 18693 21879 18751 21885
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 18693 21845 18705 21879
rect 18739 21876 18751 21879
rect 18782 21876 18788 21888
rect 18739 21848 18788 21876
rect 18739 21845 18751 21848
rect 18693 21839 18751 21845
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 21100 21885 21128 21916
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21845 21143 21879
rect 21085 21839 21143 21845
rect 21174 21836 21180 21888
rect 21232 21836 21238 21888
rect 21284 21876 21312 21916
rect 23032 21888 23060 21975
rect 23124 21944 23152 22052
rect 23290 22040 23296 22092
rect 23348 22040 23354 22092
rect 23768 22089 23796 22120
rect 24026 22108 24032 22160
rect 24084 22108 24090 22160
rect 23753 22083 23811 22089
rect 23753 22049 23765 22083
rect 23799 22080 23811 22083
rect 24118 22080 24124 22092
rect 23799 22052 24124 22080
rect 23799 22049 23811 22052
rect 23753 22043 23811 22049
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 25774 22040 25780 22092
rect 25832 22080 25838 22092
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 25832 22052 26065 22080
rect 25832 22040 25838 22052
rect 26053 22049 26065 22052
rect 26099 22049 26111 22083
rect 26053 22043 26111 22049
rect 26142 22040 26148 22092
rect 26200 22080 26206 22092
rect 28368 22089 28396 22188
rect 28810 22176 28816 22188
rect 28868 22176 28874 22228
rect 29362 22176 29368 22228
rect 29420 22216 29426 22228
rect 34241 22219 34299 22225
rect 34241 22216 34253 22219
rect 29420 22188 34253 22216
rect 29420 22176 29426 22188
rect 34241 22185 34253 22188
rect 34287 22216 34299 22219
rect 34790 22216 34796 22228
rect 34287 22188 34796 22216
rect 34287 22185 34299 22188
rect 34241 22179 34299 22185
rect 34790 22176 34796 22188
rect 34848 22176 34854 22228
rect 35434 22176 35440 22228
rect 35492 22176 35498 22228
rect 37458 22176 37464 22228
rect 37516 22176 37522 22228
rect 37642 22176 37648 22228
rect 37700 22216 37706 22228
rect 37829 22219 37887 22225
rect 37829 22216 37841 22219
rect 37700 22188 37841 22216
rect 37700 22176 37706 22188
rect 37829 22185 37841 22188
rect 37875 22185 37887 22219
rect 37829 22179 37887 22185
rect 28442 22108 28448 22160
rect 28500 22148 28506 22160
rect 30374 22148 30380 22160
rect 28500 22120 30380 22148
rect 28500 22108 28506 22120
rect 30374 22108 30380 22120
rect 30432 22108 30438 22160
rect 33870 22108 33876 22160
rect 33928 22108 33934 22160
rect 36262 22148 36268 22160
rect 34808 22120 36268 22148
rect 28353 22083 28411 22089
rect 28353 22080 28365 22083
rect 26200 22052 28365 22080
rect 26200 22040 26206 22052
rect 28353 22049 28365 22052
rect 28399 22049 28411 22083
rect 28353 22043 28411 22049
rect 28828 22052 28994 22080
rect 23308 22012 23336 22040
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23308 21984 24409 22012
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 28828 22012 28856 22052
rect 24949 21975 25007 21981
rect 25700 21984 28856 22012
rect 23198 21944 23204 21956
rect 23124 21916 23204 21944
rect 23198 21904 23204 21916
rect 23256 21944 23262 21956
rect 24964 21944 24992 21975
rect 25700 21956 25728 21984
rect 23256 21916 24992 21944
rect 23256 21904 23262 21916
rect 25682 21904 25688 21956
rect 25740 21904 25746 21956
rect 28442 21904 28448 21956
rect 28500 21904 28506 21956
rect 28966 21944 28994 22052
rect 32214 22040 32220 22092
rect 32272 22080 32278 22092
rect 32493 22083 32551 22089
rect 32493 22080 32505 22083
rect 32272 22052 32505 22080
rect 32272 22040 32278 22052
rect 32493 22049 32505 22052
rect 32539 22049 32551 22083
rect 32493 22043 32551 22049
rect 34422 22040 34428 22092
rect 34480 22080 34486 22092
rect 34808 22089 34836 22120
rect 36262 22108 36268 22120
rect 36320 22108 36326 22160
rect 37476 22148 37504 22176
rect 37737 22151 37795 22157
rect 37737 22148 37749 22151
rect 37476 22120 37749 22148
rect 37737 22117 37749 22120
rect 37783 22117 37795 22151
rect 37737 22111 37795 22117
rect 34793 22083 34851 22089
rect 34793 22080 34805 22083
rect 34480 22052 34805 22080
rect 34480 22040 34486 22052
rect 34793 22049 34805 22052
rect 34839 22049 34851 22083
rect 34793 22043 34851 22049
rect 35713 22083 35771 22089
rect 35713 22049 35725 22083
rect 35759 22080 35771 22083
rect 35986 22080 35992 22092
rect 35759 22052 35992 22080
rect 35759 22049 35771 22052
rect 35713 22043 35771 22049
rect 35986 22040 35992 22052
rect 36044 22040 36050 22092
rect 37752 22080 37780 22111
rect 38381 22083 38439 22089
rect 38381 22080 38393 22083
rect 37752 22052 38393 22080
rect 38381 22049 38393 22052
rect 38427 22049 38439 22083
rect 38381 22043 38439 22049
rect 31849 22015 31907 22021
rect 31849 21981 31861 22015
rect 31895 22012 31907 22015
rect 33042 22012 33048 22024
rect 31895 21984 33048 22012
rect 31895 21981 31907 21984
rect 31849 21975 31907 21981
rect 33042 21972 33048 21984
rect 33100 21972 33106 22024
rect 35250 22012 35256 22024
rect 34164 21984 35256 22012
rect 31938 21944 31944 21956
rect 28966 21916 31944 21944
rect 31938 21904 31944 21916
rect 31996 21904 32002 21956
rect 32760 21947 32818 21953
rect 32760 21913 32772 21947
rect 32806 21944 32818 21947
rect 34164 21944 34192 21984
rect 35250 21972 35256 21984
rect 35308 21972 35314 22024
rect 35342 21972 35348 22024
rect 35400 22012 35406 22024
rect 36354 22012 36360 22024
rect 35400 21984 36360 22012
rect 35400 21972 35406 21984
rect 36354 21972 36360 21984
rect 36412 21972 36418 22024
rect 36624 22015 36682 22021
rect 36624 21981 36636 22015
rect 36670 22012 36682 22015
rect 37182 22012 37188 22024
rect 36670 21984 37188 22012
rect 36670 21981 36682 21984
rect 36624 21975 36682 21981
rect 37182 21972 37188 21984
rect 37240 21972 37246 22024
rect 32806 21916 34192 21944
rect 35069 21947 35127 21953
rect 32806 21913 32818 21916
rect 32760 21907 32818 21913
rect 35069 21913 35081 21947
rect 35115 21944 35127 21947
rect 35115 21916 35480 21944
rect 35115 21913 35127 21916
rect 35069 21907 35127 21913
rect 22094 21876 22100 21888
rect 21284 21848 22100 21876
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 23014 21836 23020 21888
rect 23072 21836 23078 21888
rect 23106 21836 23112 21888
rect 23164 21836 23170 21888
rect 23474 21836 23480 21888
rect 23532 21836 23538 21888
rect 23566 21836 23572 21888
rect 23624 21836 23630 21888
rect 24118 21836 24124 21888
rect 24176 21876 24182 21888
rect 24213 21879 24271 21885
rect 24213 21876 24225 21879
rect 24176 21848 24225 21876
rect 24176 21836 24182 21848
rect 24213 21845 24225 21848
rect 24259 21876 24271 21879
rect 28460 21876 28488 21904
rect 24259 21848 28488 21876
rect 24259 21845 24271 21848
rect 24213 21839 24271 21845
rect 28810 21836 28816 21888
rect 28868 21876 28874 21888
rect 29362 21876 29368 21888
rect 28868 21848 29368 21876
rect 28868 21836 28874 21848
rect 29362 21836 29368 21848
rect 29420 21836 29426 21888
rect 32398 21836 32404 21888
rect 32456 21836 32462 21888
rect 34974 21836 34980 21888
rect 35032 21836 35038 21888
rect 35452 21876 35480 21916
rect 35894 21904 35900 21956
rect 35952 21904 35958 21956
rect 36446 21944 36452 21956
rect 36004 21916 36452 21944
rect 35805 21879 35863 21885
rect 35805 21876 35817 21879
rect 35452 21848 35817 21876
rect 35805 21845 35817 21848
rect 35851 21876 35863 21879
rect 36004 21876 36032 21916
rect 36446 21904 36452 21916
rect 36504 21904 36510 21956
rect 35851 21848 36032 21876
rect 35851 21845 35863 21848
rect 35805 21839 35863 21845
rect 36170 21836 36176 21888
rect 36228 21876 36234 21888
rect 36265 21879 36323 21885
rect 36265 21876 36277 21879
rect 36228 21848 36277 21876
rect 36228 21836 36234 21848
rect 36265 21845 36277 21848
rect 36311 21845 36323 21879
rect 36265 21839 36323 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2961 21675 3019 21681
rect 2961 21641 2973 21675
rect 3007 21672 3019 21675
rect 3050 21672 3056 21684
rect 3007 21644 3056 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 3050 21632 3056 21644
rect 3108 21632 3114 21684
rect 4249 21675 4307 21681
rect 4249 21641 4261 21675
rect 4295 21672 4307 21675
rect 5166 21672 5172 21684
rect 4295 21644 5172 21672
rect 4295 21641 4307 21644
rect 4249 21635 4307 21641
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 7926 21632 7932 21684
rect 7984 21672 7990 21684
rect 8570 21672 8576 21684
rect 7984 21644 8576 21672
rect 7984 21632 7990 21644
rect 8570 21632 8576 21644
rect 8628 21672 8634 21684
rect 13722 21672 13728 21684
rect 8628 21644 13728 21672
rect 8628 21632 8634 21644
rect 13722 21632 13728 21644
rect 13780 21672 13786 21684
rect 13817 21675 13875 21681
rect 13817 21672 13829 21675
rect 13780 21644 13829 21672
rect 13780 21632 13786 21644
rect 13817 21641 13829 21644
rect 13863 21641 13875 21675
rect 13817 21635 13875 21641
rect 21174 21632 21180 21684
rect 21232 21632 21238 21684
rect 21637 21675 21695 21681
rect 21637 21641 21649 21675
rect 21683 21672 21695 21675
rect 22370 21672 22376 21684
rect 21683 21644 22376 21672
rect 21683 21641 21695 21644
rect 21637 21635 21695 21641
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 22554 21632 22560 21684
rect 22612 21672 22618 21684
rect 23382 21672 23388 21684
rect 22612 21644 23388 21672
rect 22612 21632 22618 21644
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 24026 21632 24032 21684
rect 24084 21672 24090 21684
rect 24121 21675 24179 21681
rect 24121 21672 24133 21675
rect 24084 21644 24133 21672
rect 24084 21632 24090 21644
rect 24121 21641 24133 21644
rect 24167 21672 24179 21675
rect 24302 21672 24308 21684
rect 24167 21644 24308 21672
rect 24167 21641 24179 21644
rect 24121 21635 24179 21641
rect 24302 21632 24308 21644
rect 24360 21632 24366 21684
rect 32766 21632 32772 21684
rect 32824 21632 32830 21684
rect 33137 21675 33195 21681
rect 33137 21641 33149 21675
rect 33183 21672 33195 21675
rect 33318 21672 33324 21684
rect 33183 21644 33324 21672
rect 33183 21641 33195 21644
rect 33137 21635 33195 21641
rect 33318 21632 33324 21644
rect 33376 21632 33382 21684
rect 33594 21632 33600 21684
rect 33652 21632 33658 21684
rect 35437 21675 35495 21681
rect 35437 21641 35449 21675
rect 35483 21641 35495 21675
rect 35437 21635 35495 21641
rect 3329 21607 3387 21613
rect 3329 21573 3341 21607
rect 3375 21604 3387 21607
rect 5902 21604 5908 21616
rect 3375 21576 5908 21604
rect 3375 21573 3387 21576
rect 3329 21567 3387 21573
rect 5902 21564 5908 21576
rect 5960 21564 5966 21616
rect 11698 21564 11704 21616
rect 11756 21604 11762 21616
rect 20524 21607 20582 21613
rect 11756 21576 13492 21604
rect 11756 21564 11762 21576
rect 5537 21539 5595 21545
rect 5537 21505 5549 21539
rect 5583 21536 5595 21539
rect 12161 21539 12219 21545
rect 5583 21508 5856 21536
rect 5583 21505 5595 21508
rect 5537 21499 5595 21505
rect 3418 21428 3424 21480
rect 3476 21428 3482 21480
rect 3602 21428 3608 21480
rect 3660 21428 3666 21480
rect 5828 21341 5856 21508
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 12434 21536 12440 21548
rect 12207 21508 12440 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 12434 21496 12440 21508
rect 12492 21536 12498 21548
rect 12618 21536 12624 21548
rect 12492 21508 12624 21536
rect 12492 21496 12498 21508
rect 12618 21496 12624 21508
rect 12676 21496 12682 21548
rect 13464 21545 13492 21576
rect 20524 21573 20536 21607
rect 20570 21604 20582 21607
rect 20714 21604 20720 21616
rect 20570 21576 20720 21604
rect 20570 21573 20582 21576
rect 20524 21567 20582 21573
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 21192 21604 21220 21632
rect 22462 21604 22468 21616
rect 21192 21576 22468 21604
rect 22462 21564 22468 21576
rect 22520 21564 22526 21616
rect 33229 21607 33287 21613
rect 33229 21573 33241 21607
rect 33275 21604 33287 21607
rect 33612 21604 33640 21632
rect 33275 21576 33640 21604
rect 35452 21604 35480 21635
rect 37550 21632 37556 21684
rect 37608 21632 37614 21684
rect 37645 21607 37703 21613
rect 37645 21604 37657 21607
rect 35452 21576 37657 21604
rect 33275 21573 33287 21576
rect 33229 21567 33287 21573
rect 37645 21573 37657 21576
rect 37691 21573 37703 21607
rect 37645 21567 37703 21573
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 16485 21539 16543 21545
rect 16485 21505 16497 21539
rect 16531 21536 16543 21539
rect 17129 21539 17187 21545
rect 17129 21536 17141 21539
rect 16531 21508 17141 21536
rect 16531 21505 16543 21508
rect 16485 21499 16543 21505
rect 17129 21505 17141 21508
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 17954 21536 17960 21548
rect 17276 21508 17960 21536
rect 17276 21496 17282 21508
rect 17954 21496 17960 21508
rect 18012 21536 18018 21548
rect 18509 21539 18567 21545
rect 18012 21508 18276 21536
rect 18012 21496 18018 21508
rect 18248 21480 18276 21508
rect 18509 21505 18521 21539
rect 18555 21536 18567 21539
rect 19978 21536 19984 21548
rect 18555 21508 19984 21536
rect 18555 21505 18567 21508
rect 18509 21499 18567 21505
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 29917 21539 29975 21545
rect 23891 21508 24624 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 10594 21428 10600 21480
rect 10652 21428 10658 21480
rect 11333 21471 11391 21477
rect 11333 21437 11345 21471
rect 11379 21468 11391 21471
rect 12253 21471 12311 21477
rect 11379 21440 11836 21468
rect 11379 21437 11391 21440
rect 11333 21431 11391 21437
rect 11808 21409 11836 21440
rect 12253 21437 12265 21471
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 11793 21403 11851 21409
rect 11793 21369 11805 21403
rect 11839 21369 11851 21403
rect 12268 21400 12296 21431
rect 12342 21428 12348 21480
rect 12400 21428 12406 21480
rect 15838 21428 15844 21480
rect 15896 21428 15902 21480
rect 17313 21471 17371 21477
rect 17313 21437 17325 21471
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 12434 21400 12440 21412
rect 12268 21372 12440 21400
rect 11793 21363 11851 21369
rect 12434 21360 12440 21372
rect 12492 21360 12498 21412
rect 15749 21403 15807 21409
rect 15749 21400 15761 21403
rect 12636 21372 15761 21400
rect 5813 21335 5871 21341
rect 5813 21301 5825 21335
rect 5859 21332 5871 21335
rect 6086 21332 6092 21344
rect 5859 21304 6092 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 6086 21292 6092 21304
rect 6144 21332 6150 21344
rect 8294 21332 8300 21344
rect 6144 21304 8300 21332
rect 6144 21292 6150 21304
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 9950 21292 9956 21344
rect 10008 21292 10014 21344
rect 10686 21292 10692 21344
rect 10744 21292 10750 21344
rect 11422 21292 11428 21344
rect 11480 21332 11486 21344
rect 12636 21332 12664 21372
rect 15749 21369 15761 21372
rect 15795 21400 15807 21403
rect 17218 21400 17224 21412
rect 15795 21372 17224 21400
rect 15795 21369 15807 21372
rect 15749 21363 15807 21369
rect 17218 21360 17224 21372
rect 17276 21400 17282 21412
rect 17328 21400 17356 21431
rect 17862 21428 17868 21480
rect 17920 21428 17926 21480
rect 18230 21428 18236 21480
rect 18288 21428 18294 21480
rect 19150 21428 19156 21480
rect 19208 21428 19214 21480
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 17276 21372 17356 21400
rect 17276 21360 17282 21372
rect 18322 21360 18328 21412
rect 18380 21400 18386 21412
rect 18601 21403 18659 21409
rect 18601 21400 18613 21403
rect 18380 21372 18613 21400
rect 18380 21360 18386 21372
rect 18601 21369 18613 21372
rect 18647 21369 18659 21403
rect 18601 21363 18659 21369
rect 11480 21304 12664 21332
rect 11480 21292 11486 21304
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 12897 21335 12955 21341
rect 12897 21332 12909 21335
rect 12768 21304 12909 21332
rect 12768 21292 12774 21304
rect 12897 21301 12909 21304
rect 12943 21301 12955 21335
rect 12897 21295 12955 21301
rect 16758 21292 16764 21344
rect 16816 21292 16822 21344
rect 19613 21335 19671 21341
rect 19613 21301 19625 21335
rect 19659 21332 19671 21335
rect 19886 21332 19892 21344
rect 19659 21304 19892 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 19886 21292 19892 21304
rect 19944 21292 19950 21344
rect 20272 21332 20300 21431
rect 20898 21332 20904 21344
rect 20272 21304 20904 21332
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 24596 21341 24624 21508
rect 29917 21505 29929 21539
rect 29963 21536 29975 21539
rect 30190 21536 30196 21548
rect 29963 21508 30196 21536
rect 29963 21505 29975 21508
rect 29917 21499 29975 21505
rect 30190 21496 30196 21508
rect 30248 21496 30254 21548
rect 31938 21496 31944 21548
rect 31996 21536 32002 21548
rect 32677 21539 32735 21545
rect 32677 21536 32689 21539
rect 31996 21508 32689 21536
rect 31996 21496 32002 21508
rect 32677 21505 32689 21508
rect 32723 21536 32735 21539
rect 32723 21508 33364 21536
rect 32723 21505 32735 21508
rect 32677 21499 32735 21505
rect 29641 21471 29699 21477
rect 29641 21468 29653 21471
rect 29380 21440 29653 21468
rect 24581 21335 24639 21341
rect 24581 21301 24593 21335
rect 24627 21332 24639 21335
rect 24854 21332 24860 21344
rect 24627 21304 24860 21332
rect 24627 21301 24639 21304
rect 24581 21295 24639 21301
rect 24854 21292 24860 21304
rect 24912 21332 24918 21344
rect 27982 21332 27988 21344
rect 24912 21304 27988 21332
rect 24912 21292 24918 21304
rect 27982 21292 27988 21304
rect 28040 21292 28046 21344
rect 29270 21292 29276 21344
rect 29328 21332 29334 21344
rect 29380 21341 29408 21440
rect 29641 21437 29653 21440
rect 29687 21437 29699 21471
rect 29641 21431 29699 21437
rect 29825 21471 29883 21477
rect 29825 21437 29837 21471
rect 29871 21468 29883 21471
rect 30377 21471 30435 21477
rect 30377 21468 30389 21471
rect 29871 21440 30389 21468
rect 29871 21437 29883 21440
rect 29825 21431 29883 21437
rect 30377 21437 30389 21440
rect 30423 21437 30435 21471
rect 30377 21431 30435 21437
rect 30466 21428 30472 21480
rect 30524 21468 30530 21480
rect 33336 21477 33364 21508
rect 33778 21496 33784 21548
rect 33836 21496 33842 21548
rect 34790 21496 34796 21548
rect 34848 21496 34854 21548
rect 35434 21496 35440 21548
rect 35492 21536 35498 21548
rect 36081 21539 36139 21545
rect 36081 21536 36093 21539
rect 35492 21508 36093 21536
rect 35492 21496 35498 21508
rect 36081 21505 36093 21508
rect 36127 21505 36139 21539
rect 36081 21499 36139 21505
rect 30929 21471 30987 21477
rect 30929 21468 30941 21471
rect 30524 21440 30941 21468
rect 30524 21428 30530 21440
rect 30929 21437 30941 21440
rect 30975 21437 30987 21471
rect 30929 21431 30987 21437
rect 31757 21471 31815 21477
rect 31757 21437 31769 21471
rect 31803 21437 31815 21471
rect 31757 21431 31815 21437
rect 33321 21471 33379 21477
rect 33321 21437 33333 21471
rect 33367 21437 33379 21471
rect 33321 21431 33379 21437
rect 33597 21471 33655 21477
rect 33597 21437 33609 21471
rect 33643 21468 33655 21471
rect 34146 21468 34152 21480
rect 33643 21440 34152 21468
rect 33643 21437 33655 21440
rect 33597 21431 33655 21437
rect 30285 21403 30343 21409
rect 30285 21369 30297 21403
rect 30331 21400 30343 21403
rect 31772 21400 31800 21431
rect 34146 21428 34152 21440
rect 34204 21428 34210 21480
rect 34517 21471 34575 21477
rect 34517 21468 34529 21471
rect 34348 21440 34529 21468
rect 30331 21372 31800 21400
rect 30331 21369 30343 21372
rect 30285 21363 30343 21369
rect 33410 21360 33416 21412
rect 33468 21400 33474 21412
rect 34241 21403 34299 21409
rect 34241 21400 34253 21403
rect 33468 21372 34253 21400
rect 33468 21360 33474 21372
rect 34241 21369 34253 21372
rect 34287 21369 34299 21403
rect 34241 21363 34299 21369
rect 29365 21335 29423 21341
rect 29365 21332 29377 21335
rect 29328 21304 29377 21332
rect 29328 21292 29334 21304
rect 29365 21301 29377 21304
rect 29411 21301 29423 21335
rect 29365 21295 29423 21301
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 31113 21335 31171 21341
rect 31113 21332 31125 21335
rect 30984 21304 31125 21332
rect 30984 21292 30990 21304
rect 31113 21301 31125 21304
rect 31159 21301 31171 21335
rect 31113 21295 31171 21301
rect 33870 21292 33876 21344
rect 33928 21332 33934 21344
rect 34348 21332 34376 21440
rect 34517 21437 34529 21440
rect 34563 21437 34575 21471
rect 34517 21431 34575 21437
rect 34606 21428 34612 21480
rect 34664 21477 34670 21480
rect 34664 21471 34692 21477
rect 34680 21437 34692 21471
rect 34664 21431 34692 21437
rect 34664 21428 34670 21431
rect 34974 21428 34980 21480
rect 35032 21468 35038 21480
rect 36265 21471 36323 21477
rect 36265 21468 36277 21471
rect 35032 21440 36277 21468
rect 35032 21428 35038 21440
rect 36265 21437 36277 21440
rect 36311 21437 36323 21471
rect 36265 21431 36323 21437
rect 36817 21471 36875 21477
rect 36817 21437 36829 21471
rect 36863 21437 36875 21471
rect 36817 21431 36875 21437
rect 35250 21360 35256 21412
rect 35308 21400 35314 21412
rect 35529 21403 35587 21409
rect 35529 21400 35541 21403
rect 35308 21372 35541 21400
rect 35308 21360 35314 21372
rect 35529 21369 35541 21372
rect 35575 21369 35587 21403
rect 35529 21363 35587 21369
rect 36832 21332 36860 21431
rect 37458 21428 37464 21480
rect 37516 21428 37522 21480
rect 33928 21304 36860 21332
rect 33928 21292 33934 21304
rect 38010 21292 38016 21344
rect 38068 21292 38074 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 3418 21088 3424 21140
rect 3476 21128 3482 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 3476 21100 3801 21128
rect 3476 21088 3482 21100
rect 3789 21097 3801 21100
rect 3835 21097 3847 21131
rect 3789 21091 3847 21097
rect 10594 21088 10600 21140
rect 10652 21128 10658 21140
rect 10873 21131 10931 21137
rect 10873 21128 10885 21131
rect 10652 21100 10885 21128
rect 10652 21088 10658 21100
rect 10873 21097 10885 21100
rect 10919 21097 10931 21131
rect 10873 21091 10931 21097
rect 11054 21088 11060 21140
rect 11112 21088 11118 21140
rect 11698 21088 11704 21140
rect 11756 21088 11762 21140
rect 16758 21088 16764 21140
rect 16816 21088 16822 21140
rect 16853 21131 16911 21137
rect 16853 21097 16865 21131
rect 16899 21128 16911 21131
rect 17126 21128 17132 21140
rect 16899 21100 17132 21128
rect 16899 21097 16911 21100
rect 16853 21091 16911 21097
rect 17126 21088 17132 21100
rect 17184 21128 17190 21140
rect 17862 21128 17868 21140
rect 17184 21100 17868 21128
rect 17184 21088 17190 21100
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18322 21088 18328 21140
rect 18380 21088 18386 21140
rect 21729 21131 21787 21137
rect 21729 21097 21741 21131
rect 21775 21128 21787 21131
rect 23014 21128 23020 21140
rect 21775 21100 23020 21128
rect 21775 21097 21787 21100
rect 21729 21091 21787 21097
rect 23014 21088 23020 21100
rect 23072 21128 23078 21140
rect 23072 21100 23336 21128
rect 23072 21088 23078 21100
rect 3602 21020 3608 21072
rect 3660 21060 3666 21072
rect 4890 21060 4896 21072
rect 3660 21032 4896 21060
rect 3660 21020 3666 21032
rect 4890 21020 4896 21032
rect 4948 21020 4954 21072
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20992 4491 20995
rect 4614 20992 4620 21004
rect 4479 20964 4620 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 5258 20992 5264 21004
rect 4816 20964 5264 20992
rect 4522 20748 4528 20800
rect 4580 20788 4586 20800
rect 4816 20797 4844 20964
rect 5258 20952 5264 20964
rect 5316 20992 5322 21004
rect 5316 20964 11008 20992
rect 5316 20952 5322 20964
rect 6638 20884 6644 20936
rect 6696 20884 6702 20936
rect 7742 20884 7748 20936
rect 7800 20924 7806 20936
rect 7837 20927 7895 20933
rect 7837 20924 7849 20927
rect 7800 20896 7849 20924
rect 7800 20884 7806 20896
rect 7837 20893 7849 20896
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 8297 20927 8355 20933
rect 8297 20893 8309 20927
rect 8343 20924 8355 20927
rect 8343 20896 8432 20924
rect 8343 20893 8355 20896
rect 8297 20887 8355 20893
rect 8404 20868 8432 20896
rect 6454 20816 6460 20868
rect 6512 20856 6518 20868
rect 7285 20859 7343 20865
rect 7285 20856 7297 20859
rect 6512 20828 7297 20856
rect 6512 20816 6518 20828
rect 7285 20825 7297 20828
rect 7331 20825 7343 20859
rect 7285 20819 7343 20825
rect 8386 20816 8392 20868
rect 8444 20816 8450 20868
rect 8941 20859 8999 20865
rect 8941 20825 8953 20859
rect 8987 20825 8999 20859
rect 10980 20856 11008 20964
rect 11072 20924 11100 21088
rect 11422 20952 11428 21004
rect 11480 20952 11486 21004
rect 13170 20952 13176 21004
rect 13228 20992 13234 21004
rect 13633 20995 13691 21001
rect 13633 20992 13645 20995
rect 13228 20964 13645 20992
rect 13228 20952 13234 20964
rect 13633 20961 13645 20964
rect 13679 20961 13691 20995
rect 13633 20955 13691 20961
rect 13722 20952 13728 21004
rect 13780 20952 13786 21004
rect 16776 21001 16804 21088
rect 16761 20995 16819 21001
rect 16761 20961 16773 20995
rect 16807 20961 16819 20995
rect 18340 20992 18368 21088
rect 19061 21063 19119 21069
rect 18524 21032 18828 21060
rect 18524 21001 18552 21032
rect 18800 21004 18828 21032
rect 19061 21029 19073 21063
rect 19107 21060 19119 21063
rect 19426 21060 19432 21072
rect 19107 21032 19432 21060
rect 19107 21029 19119 21032
rect 19061 21023 19119 21029
rect 19426 21020 19432 21032
rect 19484 21020 19490 21072
rect 23198 21020 23204 21072
rect 23256 21020 23262 21072
rect 16761 20955 16819 20961
rect 18156 20964 18368 20992
rect 18509 20995 18567 21001
rect 11241 20927 11299 20933
rect 11241 20924 11253 20927
rect 11072 20896 11253 20924
rect 11241 20893 11253 20896
rect 11287 20893 11299 20927
rect 11241 20887 11299 20893
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 13081 20927 13139 20933
rect 12492 20896 13032 20924
rect 12492 20884 12498 20896
rect 11054 20856 11060 20868
rect 10980 20828 11060 20856
rect 8941 20819 8999 20825
rect 4801 20791 4859 20797
rect 4801 20788 4813 20791
rect 4580 20760 4813 20788
rect 4580 20748 4586 20760
rect 4801 20757 4813 20760
rect 4847 20757 4859 20791
rect 4801 20751 4859 20757
rect 7190 20748 7196 20800
rect 7248 20748 7254 20800
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 8665 20791 8723 20797
rect 8665 20788 8677 20791
rect 8352 20760 8677 20788
rect 8352 20748 8358 20760
rect 8665 20757 8677 20760
rect 8711 20788 8723 20791
rect 8956 20788 8984 20819
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 11333 20859 11391 20865
rect 11333 20825 11345 20859
rect 11379 20856 11391 20859
rect 12618 20856 12624 20868
rect 11379 20828 12624 20856
rect 11379 20825 11391 20828
rect 11333 20819 11391 20825
rect 12618 20816 12624 20828
rect 12676 20816 12682 20868
rect 12802 20816 12808 20868
rect 12860 20865 12866 20868
rect 12860 20819 12872 20865
rect 13004 20856 13032 20896
rect 13081 20893 13093 20927
rect 13127 20924 13139 20927
rect 13446 20924 13452 20936
rect 13127 20896 13452 20924
rect 13127 20893 13139 20896
rect 13081 20887 13139 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 14645 20927 14703 20933
rect 14645 20924 14657 20927
rect 13872 20896 14657 20924
rect 13872 20884 13878 20896
rect 14645 20893 14657 20896
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 17977 20927 18035 20933
rect 17977 20893 17989 20927
rect 18023 20924 18035 20927
rect 18156 20924 18184 20964
rect 18509 20961 18521 20995
rect 18555 20961 18567 20995
rect 18509 20955 18567 20961
rect 18782 20952 18788 21004
rect 18840 20952 18846 21004
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 19392 20964 19717 20992
rect 19392 20952 19398 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 19886 20952 19892 21004
rect 19944 20992 19950 21004
rect 20254 20992 20260 21004
rect 19944 20964 20260 20992
rect 19944 20952 19950 20964
rect 20254 20952 20260 20964
rect 20312 20952 20318 21004
rect 23308 21001 23336 21100
rect 23566 21088 23572 21140
rect 23624 21128 23630 21140
rect 23937 21131 23995 21137
rect 23937 21128 23949 21131
rect 23624 21100 23949 21128
rect 23624 21088 23630 21100
rect 23937 21097 23949 21100
rect 23983 21097 23995 21131
rect 23937 21091 23995 21097
rect 29362 21088 29368 21140
rect 29420 21088 29426 21140
rect 30101 21131 30159 21137
rect 30101 21097 30113 21131
rect 30147 21128 30159 21131
rect 31294 21128 31300 21140
rect 30147 21100 31300 21128
rect 30147 21097 30159 21100
rect 30101 21091 30159 21097
rect 31294 21088 31300 21100
rect 31352 21088 31358 21140
rect 32398 21088 32404 21140
rect 32456 21088 32462 21140
rect 34146 21088 34152 21140
rect 34204 21128 34210 21140
rect 34606 21128 34612 21140
rect 34204 21100 34612 21128
rect 34204 21088 34210 21100
rect 34606 21088 34612 21100
rect 34664 21088 34670 21140
rect 35802 21088 35808 21140
rect 35860 21128 35866 21140
rect 36173 21131 36231 21137
rect 36173 21128 36185 21131
rect 35860 21100 36185 21128
rect 35860 21088 35866 21100
rect 36173 21097 36185 21100
rect 36219 21128 36231 21131
rect 36354 21128 36360 21140
rect 36219 21100 36360 21128
rect 36219 21097 36231 21100
rect 36173 21091 36231 21097
rect 36354 21088 36360 21100
rect 36412 21088 36418 21140
rect 36722 21088 36728 21140
rect 36780 21088 36786 21140
rect 37185 21131 37243 21137
rect 37185 21097 37197 21131
rect 37231 21128 37243 21131
rect 37274 21128 37280 21140
rect 37231 21100 37280 21128
rect 37231 21097 37243 21100
rect 37185 21091 37243 21097
rect 37274 21088 37280 21100
rect 37332 21088 37338 21140
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 27157 20995 27215 21001
rect 27157 20961 27169 20995
rect 27203 20992 27215 20995
rect 32416 20992 32444 21088
rect 37458 21020 37464 21072
rect 37516 21020 37522 21072
rect 27203 20964 27384 20992
rect 32416 20964 32904 20992
rect 27203 20961 27215 20964
rect 27157 20955 27215 20961
rect 27356 20936 27384 20964
rect 18023 20896 18184 20924
rect 18233 20927 18291 20933
rect 18023 20893 18035 20896
rect 17977 20887 18035 20893
rect 18233 20893 18245 20927
rect 18279 20924 18291 20927
rect 18598 20924 18604 20936
rect 18279 20896 18604 20924
rect 18279 20893 18291 20896
rect 18233 20887 18291 20893
rect 14093 20859 14151 20865
rect 14093 20856 14105 20859
rect 13004 20828 14105 20856
rect 14093 20825 14105 20828
rect 14139 20825 14151 20859
rect 14093 20819 14151 20825
rect 16025 20859 16083 20865
rect 16025 20825 16037 20859
rect 16071 20856 16083 20859
rect 16206 20856 16212 20868
rect 16071 20828 16212 20856
rect 16071 20825 16083 20828
rect 16025 20819 16083 20825
rect 12860 20816 12866 20819
rect 16206 20816 16212 20828
rect 16264 20856 16270 20868
rect 18248 20856 18276 20887
rect 18598 20884 18604 20896
rect 18656 20884 18662 20936
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 20898 20924 20904 20936
rect 20395 20896 20904 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 20898 20884 20904 20896
rect 20956 20924 20962 20936
rect 21542 20924 21548 20936
rect 20956 20896 21548 20924
rect 20956 20884 20962 20896
rect 21542 20884 21548 20896
rect 21600 20924 21606 20936
rect 21821 20927 21879 20933
rect 21821 20924 21833 20927
rect 21600 20896 21833 20924
rect 21600 20884 21606 20896
rect 21821 20893 21833 20896
rect 21867 20924 21879 20927
rect 22554 20924 22560 20936
rect 21867 20896 22560 20924
rect 21867 20893 21879 20896
rect 21821 20887 21879 20893
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 27246 20884 27252 20936
rect 27304 20884 27310 20936
rect 27338 20884 27344 20936
rect 27396 20884 27402 20936
rect 27430 20884 27436 20936
rect 27488 20924 27494 20936
rect 27488 20896 31340 20924
rect 27488 20884 27494 20896
rect 16264 20828 16528 20856
rect 16264 20816 16270 20828
rect 16500 20800 16528 20828
rect 18064 20828 18276 20856
rect 20616 20859 20674 20865
rect 18064 20800 18092 20828
rect 20616 20825 20628 20859
rect 20662 20856 20674 20859
rect 21910 20856 21916 20868
rect 20662 20828 21916 20856
rect 20662 20825 20674 20828
rect 20616 20819 20674 20825
rect 21910 20816 21916 20828
rect 21968 20816 21974 20868
rect 22088 20859 22146 20865
rect 22088 20825 22100 20859
rect 22134 20856 22146 20859
rect 22830 20856 22836 20868
rect 22134 20828 22836 20856
rect 22134 20825 22146 20828
rect 22088 20819 22146 20825
rect 22830 20816 22836 20828
rect 22888 20816 22894 20868
rect 24946 20816 24952 20868
rect 25004 20856 25010 20868
rect 25777 20859 25835 20865
rect 25777 20856 25789 20859
rect 25004 20828 25789 20856
rect 25004 20816 25010 20828
rect 25777 20825 25789 20828
rect 25823 20856 25835 20859
rect 27448 20856 27476 20884
rect 25823 20828 27476 20856
rect 25823 20825 25835 20828
rect 25777 20819 25835 20825
rect 31202 20816 31208 20868
rect 31260 20865 31266 20868
rect 31260 20819 31272 20865
rect 31312 20856 31340 20896
rect 31386 20884 31392 20936
rect 31444 20924 31450 20936
rect 31481 20927 31539 20933
rect 31481 20924 31493 20927
rect 31444 20896 31493 20924
rect 31444 20884 31450 20896
rect 31481 20893 31493 20896
rect 31527 20924 31539 20927
rect 32769 20927 32827 20933
rect 32769 20924 32781 20927
rect 31527 20896 32781 20924
rect 31527 20893 31539 20896
rect 31481 20887 31539 20893
rect 32769 20893 32781 20896
rect 32815 20893 32827 20927
rect 32876 20924 32904 20964
rect 33025 20927 33083 20933
rect 33025 20924 33037 20927
rect 32876 20896 33037 20924
rect 32769 20887 32827 20893
rect 33025 20893 33037 20896
rect 33071 20893 33083 20927
rect 34422 20924 34428 20936
rect 33025 20887 33083 20893
rect 33980 20896 34428 20924
rect 33980 20856 34008 20896
rect 34422 20884 34428 20896
rect 34480 20884 34486 20936
rect 34698 20856 34704 20868
rect 31312 20828 34008 20856
rect 34072 20828 34704 20856
rect 31260 20816 31266 20819
rect 8711 20760 8984 20788
rect 8711 20757 8723 20760
rect 8665 20751 8723 20757
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 10226 20788 10232 20800
rect 9732 20760 10232 20788
rect 9732 20748 9738 20760
rect 10226 20748 10232 20760
rect 10284 20748 10290 20800
rect 13170 20748 13176 20800
rect 13228 20748 13234 20800
rect 13538 20748 13544 20800
rect 13596 20748 13602 20800
rect 16114 20748 16120 20800
rect 16172 20748 16178 20800
rect 16482 20748 16488 20800
rect 16540 20748 16546 20800
rect 18046 20748 18052 20800
rect 18104 20748 18110 20800
rect 18230 20748 18236 20800
rect 18288 20788 18294 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18288 20760 18613 20788
rect 18288 20748 18294 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 18601 20751 18659 20757
rect 18690 20748 18696 20800
rect 18748 20748 18754 20800
rect 19242 20748 19248 20800
rect 19300 20748 19306 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19392 20760 19625 20788
rect 19392 20748 19398 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 19613 20751 19671 20757
rect 26510 20748 26516 20800
rect 26568 20748 26574 20800
rect 27890 20748 27896 20800
rect 27948 20748 27954 20800
rect 27982 20748 27988 20800
rect 28040 20788 28046 20800
rect 29917 20791 29975 20797
rect 29917 20788 29929 20791
rect 28040 20760 29929 20788
rect 28040 20748 28046 20760
rect 29917 20757 29929 20760
rect 29963 20788 29975 20791
rect 31018 20788 31024 20800
rect 29963 20760 31024 20788
rect 29963 20757 29975 20760
rect 29917 20751 29975 20757
rect 31018 20748 31024 20760
rect 31076 20788 31082 20800
rect 34072 20788 34100 20828
rect 34698 20816 34704 20828
rect 34756 20816 34762 20868
rect 31076 20760 34100 20788
rect 31076 20748 31082 20760
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 9769 20587 9827 20593
rect 9769 20584 9781 20587
rect 5276 20556 9781 20584
rect 5276 20528 5304 20556
rect 9769 20553 9781 20556
rect 9815 20584 9827 20587
rect 10410 20584 10416 20596
rect 9815 20556 10416 20584
rect 9815 20553 9827 20556
rect 9769 20547 9827 20553
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11054 20544 11060 20596
rect 11112 20544 11118 20596
rect 11333 20587 11391 20593
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 11606 20584 11612 20596
rect 11379 20556 11612 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 11606 20544 11612 20556
rect 11664 20584 11670 20596
rect 12894 20584 12900 20596
rect 11664 20556 12900 20584
rect 11664 20544 11670 20556
rect 12894 20544 12900 20556
rect 12952 20544 12958 20596
rect 13538 20544 13544 20596
rect 13596 20584 13602 20596
rect 13725 20587 13783 20593
rect 13725 20584 13737 20587
rect 13596 20556 13737 20584
rect 13596 20544 13602 20556
rect 13725 20553 13737 20556
rect 13771 20553 13783 20587
rect 13725 20547 13783 20553
rect 15105 20587 15163 20593
rect 15105 20553 15117 20587
rect 15151 20584 15163 20587
rect 15838 20584 15844 20596
rect 15151 20556 15844 20584
rect 15151 20553 15163 20556
rect 15105 20547 15163 20553
rect 15838 20544 15844 20556
rect 15896 20584 15902 20596
rect 18138 20584 18144 20596
rect 15896 20556 18144 20584
rect 15896 20544 15902 20556
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 19061 20587 19119 20593
rect 18288 20556 18828 20584
rect 18288 20544 18294 20556
rect 3513 20519 3571 20525
rect 3513 20485 3525 20519
rect 3559 20516 3571 20519
rect 3559 20488 5120 20516
rect 3559 20485 3571 20488
rect 3513 20479 3571 20485
rect 5092 20460 5120 20488
rect 5258 20476 5264 20528
rect 5316 20476 5322 20528
rect 6908 20519 6966 20525
rect 6908 20485 6920 20519
rect 6954 20516 6966 20519
rect 7190 20516 7196 20528
rect 6954 20488 7196 20516
rect 6954 20485 6966 20488
rect 6908 20479 6966 20485
rect 7190 20476 7196 20488
rect 7248 20476 7254 20528
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 10198 20519 10256 20525
rect 10198 20516 10210 20519
rect 10008 20488 10210 20516
rect 10008 20476 10014 20488
rect 10198 20485 10210 20488
rect 10244 20485 10256 20519
rect 10198 20479 10256 20485
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 3973 20451 4031 20457
rect 3973 20448 3985 20451
rect 3651 20420 3985 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 3973 20417 3985 20420
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 5074 20408 5080 20460
rect 5132 20408 5138 20460
rect 7466 20408 7472 20460
rect 7524 20448 7530 20460
rect 8113 20451 8171 20457
rect 8113 20448 8125 20451
rect 7524 20420 8125 20448
rect 7524 20408 7530 20420
rect 8113 20417 8125 20420
rect 8159 20448 8171 20451
rect 8386 20448 8392 20460
rect 8159 20420 8392 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 10428 20448 10456 20544
rect 11072 20516 11100 20544
rect 11793 20519 11851 20525
rect 11793 20516 11805 20519
rect 11072 20488 11805 20516
rect 11793 20485 11805 20488
rect 11839 20516 11851 20519
rect 11839 20488 12112 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 11422 20448 11428 20460
rect 10428 20420 11428 20448
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11756 20420 11897 20448
rect 11756 20408 11762 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 12084 20448 12112 20488
rect 16114 20476 16120 20528
rect 16172 20516 16178 20528
rect 16218 20519 16276 20525
rect 16218 20516 16230 20519
rect 16172 20488 16230 20516
rect 16172 20476 16178 20488
rect 16218 20485 16230 20488
rect 16264 20485 16276 20519
rect 16218 20479 16276 20485
rect 16482 20476 16488 20528
rect 16540 20516 16546 20528
rect 18800 20516 18828 20556
rect 19061 20553 19073 20587
rect 19107 20584 19119 20587
rect 19150 20584 19156 20596
rect 19107 20556 19156 20584
rect 19107 20553 19119 20556
rect 19061 20547 19119 20553
rect 19150 20544 19156 20556
rect 19208 20544 19214 20596
rect 19334 20544 19340 20596
rect 19392 20544 19398 20596
rect 19521 20587 19579 20593
rect 19521 20553 19533 20587
rect 19567 20584 19579 20587
rect 19978 20584 19984 20596
rect 19567 20556 19984 20584
rect 19567 20553 19579 20556
rect 19521 20547 19579 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 21910 20544 21916 20596
rect 21968 20544 21974 20596
rect 26329 20587 26387 20593
rect 26329 20553 26341 20587
rect 26375 20584 26387 20587
rect 26510 20584 26516 20596
rect 26375 20556 26516 20584
rect 26375 20553 26387 20556
rect 26329 20547 26387 20553
rect 26510 20544 26516 20556
rect 26568 20544 26574 20596
rect 29825 20587 29883 20593
rect 29825 20553 29837 20587
rect 29871 20584 29883 20587
rect 30466 20584 30472 20596
rect 29871 20556 30472 20584
rect 29871 20553 29883 20556
rect 29825 20547 29883 20553
rect 30466 20544 30472 20556
rect 30524 20544 30530 20596
rect 30576 20556 31156 20584
rect 18969 20519 19027 20525
rect 16540 20488 17264 20516
rect 18800 20488 18920 20516
rect 16540 20476 16546 20488
rect 12250 20448 12256 20460
rect 12084 20420 12256 20448
rect 11885 20411 11943 20417
rect 12250 20408 12256 20420
rect 12308 20408 12314 20460
rect 12894 20408 12900 20460
rect 12952 20457 12958 20460
rect 12952 20451 12980 20457
rect 12968 20417 12980 20451
rect 12952 20411 12980 20417
rect 12952 20408 12958 20411
rect 13078 20408 13084 20460
rect 13136 20408 13142 20460
rect 14182 20408 14188 20460
rect 14240 20408 14246 20460
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 17236 20448 17264 20488
rect 17236 20420 17448 20448
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20380 3111 20383
rect 3789 20383 3847 20389
rect 3099 20352 3188 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3160 20321 3188 20352
rect 3789 20349 3801 20383
rect 3835 20380 3847 20383
rect 3878 20380 3884 20392
rect 3835 20352 3884 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 3878 20340 3884 20352
rect 3936 20380 3942 20392
rect 4522 20380 4528 20392
rect 3936 20352 4528 20380
rect 3936 20340 3942 20352
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 4614 20340 4620 20392
rect 4672 20340 4678 20392
rect 6362 20340 6368 20392
rect 6420 20380 6426 20392
rect 6641 20383 6699 20389
rect 6641 20380 6653 20383
rect 6420 20352 6653 20380
rect 6420 20340 6426 20352
rect 6641 20349 6653 20352
rect 6687 20349 6699 20383
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 6641 20343 6699 20349
rect 7659 20352 8493 20380
rect 3145 20315 3203 20321
rect 3145 20281 3157 20315
rect 3191 20281 3203 20315
rect 3145 20275 3203 20281
rect 2409 20247 2467 20253
rect 2409 20213 2421 20247
rect 2455 20244 2467 20247
rect 2498 20244 2504 20256
rect 2455 20216 2504 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 4890 20204 4896 20256
rect 4948 20204 4954 20256
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 7659 20244 7687 20352
rect 8481 20349 8493 20352
rect 8527 20349 8539 20383
rect 8481 20343 8539 20349
rect 8496 20312 8524 20343
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 9732 20352 9965 20380
rect 9732 20340 9738 20352
rect 9953 20349 9965 20352
rect 9999 20349 10011 20383
rect 9953 20343 10011 20349
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20380 12127 20383
rect 12434 20380 12440 20392
rect 12115 20352 12440 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 12526 20340 12532 20392
rect 12584 20340 12590 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 12636 20352 12817 20380
rect 9858 20312 9864 20324
rect 8496 20284 9864 20312
rect 9858 20272 9864 20284
rect 9916 20272 9922 20324
rect 5592 20216 7687 20244
rect 5592 20204 5598 20216
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 8021 20247 8079 20253
rect 8021 20244 8033 20247
rect 7800 20216 8033 20244
rect 7800 20204 7806 20216
rect 8021 20213 8033 20216
rect 8067 20213 8079 20247
rect 8021 20207 8079 20213
rect 11974 20204 11980 20256
rect 12032 20244 12038 20256
rect 12636 20244 12664 20352
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13998 20340 14004 20392
rect 14056 20340 14062 20392
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 14274 20380 14280 20392
rect 14139 20352 14280 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20349 16543 20383
rect 17313 20383 17371 20389
rect 17313 20380 17325 20383
rect 16485 20343 16543 20349
rect 16960 20352 17325 20380
rect 13814 20244 13820 20256
rect 12032 20216 13820 20244
rect 12032 20204 12038 20216
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 14550 20204 14556 20256
rect 14608 20204 14614 20256
rect 15838 20204 15844 20256
rect 15896 20244 15902 20256
rect 16500 20244 16528 20343
rect 15896 20216 16528 20244
rect 16960 20244 16988 20352
rect 17313 20349 17325 20352
rect 17359 20349 17371 20383
rect 17420 20380 17448 20420
rect 18046 20408 18052 20460
rect 18104 20408 18110 20460
rect 18138 20408 18144 20460
rect 18196 20457 18202 20460
rect 18196 20451 18224 20457
rect 18212 20417 18224 20451
rect 18196 20411 18224 20417
rect 18196 20408 18202 20411
rect 18322 20408 18328 20460
rect 18380 20408 18386 20460
rect 18892 20448 18920 20488
rect 18969 20485 18981 20519
rect 19015 20516 19027 20519
rect 19352 20516 19380 20544
rect 19015 20488 19380 20516
rect 19015 20485 19027 20488
rect 18969 20479 19027 20485
rect 27706 20476 27712 20528
rect 27764 20516 27770 20528
rect 30576 20516 30604 20556
rect 27764 20488 30604 20516
rect 27764 20476 27770 20488
rect 30926 20476 30932 20528
rect 30984 20525 30990 20528
rect 30984 20519 31018 20525
rect 31006 20485 31018 20519
rect 31128 20516 31156 20556
rect 31202 20544 31208 20596
rect 31260 20584 31266 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 31260 20556 31309 20584
rect 31260 20544 31266 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 31297 20547 31355 20553
rect 33321 20587 33379 20593
rect 33321 20553 33333 20587
rect 33367 20584 33379 20587
rect 33410 20584 33416 20596
rect 33367 20556 33416 20584
rect 33367 20553 33379 20556
rect 33321 20547 33379 20553
rect 33410 20544 33416 20556
rect 33468 20544 33474 20596
rect 33962 20544 33968 20596
rect 34020 20584 34026 20596
rect 34057 20587 34115 20593
rect 34057 20584 34069 20587
rect 34020 20556 34069 20584
rect 34020 20544 34026 20556
rect 34057 20553 34069 20556
rect 34103 20553 34115 20587
rect 34057 20547 34115 20553
rect 34698 20544 34704 20596
rect 34756 20584 34762 20596
rect 34977 20587 35035 20593
rect 34977 20584 34989 20587
rect 34756 20556 34989 20584
rect 34756 20544 34762 20556
rect 34977 20553 34989 20556
rect 35023 20553 35035 20587
rect 34977 20547 35035 20553
rect 35345 20519 35403 20525
rect 35345 20516 35357 20519
rect 31128 20488 35357 20516
rect 30984 20479 31018 20485
rect 35345 20485 35357 20488
rect 35391 20516 35403 20519
rect 35986 20516 35992 20528
rect 35391 20488 35992 20516
rect 35391 20485 35403 20488
rect 35345 20479 35403 20485
rect 30984 20476 30990 20479
rect 35986 20476 35992 20488
rect 36044 20476 36050 20528
rect 19429 20451 19487 20457
rect 19429 20448 19441 20451
rect 18892 20420 19441 20448
rect 19429 20417 19441 20420
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 22557 20451 22615 20457
rect 22557 20417 22569 20451
rect 22603 20448 22615 20451
rect 23106 20448 23112 20460
rect 22603 20420 23112 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 27522 20448 27528 20460
rect 26283 20420 27528 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 27522 20408 27528 20420
rect 27580 20408 27586 20460
rect 27982 20408 27988 20460
rect 28040 20408 28046 20460
rect 31110 20408 31116 20460
rect 31168 20448 31174 20460
rect 33410 20448 33416 20460
rect 31168 20420 33416 20448
rect 31168 20408 31174 20420
rect 33410 20408 33416 20420
rect 33468 20408 33474 20460
rect 34606 20408 34612 20460
rect 34664 20408 34670 20460
rect 17773 20383 17831 20389
rect 17773 20380 17785 20383
rect 17420 20352 17785 20380
rect 17313 20343 17371 20349
rect 17773 20349 17785 20352
rect 17819 20349 17831 20383
rect 18340 20380 18368 20408
rect 17773 20343 17831 20349
rect 17880 20352 18368 20380
rect 17037 20315 17095 20321
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 17880 20312 17908 20352
rect 18966 20340 18972 20392
rect 19024 20380 19030 20392
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 19024 20352 19625 20380
rect 19024 20340 19030 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 23290 20340 23296 20392
rect 23348 20340 23354 20392
rect 23934 20340 23940 20392
rect 23992 20340 23998 20392
rect 25774 20340 25780 20392
rect 25832 20340 25838 20392
rect 26513 20383 26571 20389
rect 26513 20349 26525 20383
rect 26559 20380 26571 20383
rect 27430 20380 27436 20392
rect 26559 20352 27436 20380
rect 26559 20349 26571 20352
rect 26513 20343 26571 20349
rect 27430 20340 27436 20352
rect 27488 20340 27494 20392
rect 27614 20340 27620 20392
rect 27672 20340 27678 20392
rect 31205 20383 31263 20389
rect 31205 20349 31217 20383
rect 31251 20380 31263 20383
rect 31386 20380 31392 20392
rect 31251 20352 31392 20380
rect 31251 20349 31263 20352
rect 31205 20343 31263 20349
rect 17083 20284 17908 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 22922 20272 22928 20324
rect 22980 20312 22986 20324
rect 24397 20315 24455 20321
rect 24397 20312 24409 20315
rect 22980 20284 24409 20312
rect 22980 20272 22986 20284
rect 24397 20281 24409 20284
rect 24443 20312 24455 20315
rect 24443 20284 25728 20312
rect 24443 20281 24455 20284
rect 24397 20275 24455 20281
rect 25700 20256 25728 20284
rect 29288 20284 30328 20312
rect 18046 20244 18052 20256
rect 16960 20216 18052 20244
rect 15896 20204 15902 20216
rect 18046 20204 18052 20216
rect 18104 20204 18110 20256
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 18322 20244 18328 20256
rect 18196 20216 18328 20244
rect 18196 20204 18202 20216
rect 18322 20204 18328 20216
rect 18380 20204 18386 20256
rect 22646 20204 22652 20256
rect 22704 20204 22710 20256
rect 23382 20204 23388 20256
rect 23440 20204 23446 20256
rect 25133 20247 25191 20253
rect 25133 20213 25145 20247
rect 25179 20244 25191 20247
rect 25222 20244 25228 20256
rect 25179 20216 25228 20244
rect 25179 20213 25191 20216
rect 25133 20207 25191 20213
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 25682 20204 25688 20256
rect 25740 20204 25746 20256
rect 25866 20204 25872 20256
rect 25924 20204 25930 20256
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 28902 20204 28908 20256
rect 28960 20244 28966 20256
rect 29288 20253 29316 20284
rect 29273 20247 29331 20253
rect 29273 20244 29285 20247
rect 28960 20216 29285 20244
rect 28960 20204 28966 20216
rect 29273 20213 29285 20216
rect 29319 20213 29331 20247
rect 30300 20244 30328 20284
rect 31220 20244 31248 20343
rect 31386 20340 31392 20352
rect 31444 20340 31450 20392
rect 31754 20340 31760 20392
rect 31812 20380 31818 20392
rect 31849 20383 31907 20389
rect 31849 20380 31861 20383
rect 31812 20352 31861 20380
rect 31812 20340 31818 20352
rect 31849 20349 31861 20352
rect 31895 20349 31907 20383
rect 31849 20343 31907 20349
rect 30300 20216 31248 20244
rect 29273 20207 29331 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 3605 20043 3663 20049
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 4246 20040 4252 20052
rect 3651 20012 4252 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 4246 20000 4252 20012
rect 4304 20040 4310 20052
rect 4614 20040 4620 20052
rect 4304 20012 4620 20040
rect 4304 20000 4310 20012
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6696 20012 6837 20040
rect 6696 20000 6702 20012
rect 6825 20009 6837 20012
rect 6871 20009 6883 20043
rect 8846 20040 8852 20052
rect 6825 20003 6883 20009
rect 7392 20012 8852 20040
rect 7392 19972 7420 20012
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9858 20000 9864 20052
rect 9916 20000 9922 20052
rect 11974 20000 11980 20052
rect 12032 20000 12038 20052
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17954 20040 17960 20052
rect 17175 20012 17960 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 18966 20000 18972 20052
rect 19024 20000 19030 20052
rect 23198 20040 23204 20052
rect 22112 20012 23204 20040
rect 5920 19944 7420 19972
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 2225 19907 2283 19913
rect 2225 19904 2237 19907
rect 2096 19876 2237 19904
rect 2096 19864 2102 19876
rect 2225 19873 2237 19876
rect 2271 19873 2283 19907
rect 2225 19867 2283 19873
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 4890 19904 4896 19916
rect 4479 19876 4896 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 2498 19845 2504 19848
rect 2492 19836 2504 19845
rect 2459 19808 2504 19836
rect 2492 19799 2504 19808
rect 2498 19796 2504 19799
rect 2556 19796 2562 19848
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19836 4307 19839
rect 4614 19836 4620 19848
rect 4295 19808 4620 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 5166 19796 5172 19848
rect 5224 19796 5230 19848
rect 4157 19771 4215 19777
rect 4157 19737 4169 19771
rect 4203 19768 4215 19771
rect 4203 19740 5488 19768
rect 4203 19737 4215 19740
rect 4157 19731 4215 19737
rect 5092 19712 5120 19740
rect 3786 19660 3792 19712
rect 3844 19660 3850 19712
rect 4617 19703 4675 19709
rect 4617 19669 4629 19703
rect 4663 19700 4675 19703
rect 4706 19700 4712 19712
rect 4663 19672 4712 19700
rect 4663 19669 4675 19672
rect 4617 19663 4675 19669
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 5074 19660 5080 19712
rect 5132 19660 5138 19712
rect 5350 19660 5356 19712
rect 5408 19660 5414 19712
rect 5460 19700 5488 19740
rect 5920 19700 5948 19944
rect 6086 19864 6092 19916
rect 6144 19904 6150 19916
rect 6181 19907 6239 19913
rect 6181 19904 6193 19907
rect 6144 19876 6193 19904
rect 6144 19864 6150 19876
rect 6181 19873 6193 19876
rect 6227 19873 6239 19907
rect 6181 19867 6239 19873
rect 6362 19864 6368 19916
rect 6420 19864 6426 19916
rect 9674 19904 9680 19916
rect 8312 19876 9680 19904
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19805 6055 19839
rect 6380 19836 6408 19864
rect 8312 19845 8340 19876
rect 9674 19864 9680 19876
rect 9732 19904 9738 19916
rect 10597 19907 10655 19913
rect 10597 19904 10609 19907
rect 9732 19876 10609 19904
rect 9732 19864 9738 19876
rect 10597 19873 10609 19876
rect 10643 19873 10655 19907
rect 10597 19867 10655 19873
rect 13446 19864 13452 19916
rect 13504 19904 13510 19916
rect 13504 19876 15792 19904
rect 13504 19864 13510 19876
rect 8297 19839 8355 19845
rect 8297 19836 8309 19839
rect 6380 19808 8309 19836
rect 5997 19799 6055 19805
rect 8297 19805 8309 19808
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 6012 19768 6040 19799
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 10686 19796 10692 19848
rect 10744 19836 10750 19848
rect 10853 19839 10911 19845
rect 10853 19836 10865 19839
rect 10744 19808 10865 19836
rect 10744 19796 10750 19808
rect 10853 19805 10865 19808
rect 10899 19805 10911 19839
rect 10853 19799 10911 19805
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 14274 19836 14280 19848
rect 12676 19808 14280 19836
rect 12676 19796 12682 19808
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 15764 19845 15792 19876
rect 18598 19864 18604 19916
rect 18656 19864 18662 19916
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 22112 19913 22140 20012
rect 23198 20000 23204 20012
rect 23256 20000 23262 20052
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 23477 20043 23535 20049
rect 23477 20040 23489 20043
rect 23348 20012 23489 20040
rect 23348 20000 23354 20012
rect 23477 20009 23489 20012
rect 23523 20009 23535 20043
rect 23477 20003 23535 20009
rect 23934 20000 23940 20052
rect 23992 20000 23998 20052
rect 25866 20040 25872 20052
rect 24872 20012 25872 20040
rect 22649 19975 22707 19981
rect 22649 19941 22661 19975
rect 22695 19972 22707 19975
rect 23952 19972 23980 20000
rect 22695 19944 23980 19972
rect 22695 19941 22707 19944
rect 22649 19935 22707 19941
rect 22922 19913 22928 19916
rect 19797 19907 19855 19913
rect 19797 19904 19809 19907
rect 19484 19876 19809 19904
rect 19484 19864 19490 19876
rect 19797 19873 19809 19876
rect 19843 19873 19855 19907
rect 19797 19867 19855 19873
rect 22097 19907 22155 19913
rect 22097 19873 22109 19907
rect 22143 19873 22155 19907
rect 22097 19867 22155 19873
rect 22879 19907 22928 19913
rect 22879 19873 22891 19907
rect 22925 19873 22928 19907
rect 22879 19867 22928 19873
rect 22922 19864 22928 19867
rect 22980 19864 22986 19916
rect 23017 19907 23075 19913
rect 23017 19873 23029 19907
rect 23063 19904 23075 19907
rect 23106 19904 23112 19916
rect 23063 19876 23112 19904
rect 23063 19873 23075 19876
rect 23017 19867 23075 19873
rect 23106 19864 23112 19876
rect 23164 19904 23170 19916
rect 23474 19904 23480 19916
rect 23164 19876 23480 19904
rect 23164 19864 23170 19876
rect 23474 19864 23480 19876
rect 23532 19864 23538 19916
rect 24872 19913 24900 20012
rect 25866 20000 25872 20012
rect 25924 20000 25930 20052
rect 26881 20043 26939 20049
rect 26881 20009 26893 20043
rect 26927 20040 26939 20043
rect 27062 20040 27068 20052
rect 26927 20012 27068 20040
rect 26927 20009 26939 20012
rect 26881 20003 26939 20009
rect 27062 20000 27068 20012
rect 27120 20040 27126 20052
rect 27246 20040 27252 20052
rect 27120 20012 27252 20040
rect 27120 20000 27126 20012
rect 27246 20000 27252 20012
rect 27304 20000 27310 20052
rect 27614 20000 27620 20052
rect 27672 20040 27678 20052
rect 27709 20043 27767 20049
rect 27709 20040 27721 20043
rect 27672 20012 27721 20040
rect 27672 20000 27678 20012
rect 27709 20009 27721 20012
rect 27755 20009 27767 20043
rect 27709 20003 27767 20009
rect 29365 20043 29423 20049
rect 29365 20009 29377 20043
rect 29411 20040 29423 20043
rect 30374 20040 30380 20052
rect 29411 20012 30380 20040
rect 29411 20009 29423 20012
rect 29365 20003 29423 20009
rect 30374 20000 30380 20012
rect 30432 20040 30438 20052
rect 31846 20040 31852 20052
rect 30432 20012 31852 20040
rect 30432 20000 30438 20012
rect 31846 20000 31852 20012
rect 31904 20000 31910 20052
rect 30650 19932 30656 19984
rect 30708 19972 30714 19984
rect 30745 19975 30803 19981
rect 30745 19972 30757 19975
rect 30708 19944 30757 19972
rect 30708 19932 30714 19944
rect 30745 19941 30757 19944
rect 30791 19972 30803 19975
rect 31110 19972 31116 19984
rect 30791 19944 31116 19972
rect 30791 19941 30803 19944
rect 30745 19935 30803 19941
rect 31110 19932 31116 19944
rect 31168 19932 31174 19984
rect 31294 19932 31300 19984
rect 31352 19972 31358 19984
rect 31352 19944 31754 19972
rect 31352 19932 31358 19944
rect 24857 19907 24915 19913
rect 24857 19873 24869 19907
rect 24903 19873 24915 19907
rect 24857 19867 24915 19873
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 27065 19907 27123 19913
rect 27065 19904 27077 19907
rect 26752 19876 27077 19904
rect 26752 19864 26758 19876
rect 27065 19873 27077 19876
rect 27111 19873 27123 19907
rect 27065 19867 27123 19873
rect 27249 19907 27307 19913
rect 27249 19873 27261 19907
rect 27295 19904 27307 19907
rect 27890 19904 27896 19916
rect 27295 19876 27896 19904
rect 27295 19873 27307 19876
rect 27249 19867 27307 19873
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 29362 19864 29368 19916
rect 29420 19904 29426 19916
rect 30193 19907 30251 19913
rect 30193 19904 30205 19907
rect 29420 19876 30205 19904
rect 29420 19864 29426 19876
rect 30193 19873 30205 19876
rect 30239 19873 30251 19907
rect 30193 19867 30251 19873
rect 30466 19864 30472 19916
rect 30524 19864 30530 19916
rect 31389 19907 31447 19913
rect 31389 19904 31401 19907
rect 31036 19876 31401 19904
rect 31036 19848 31064 19876
rect 31389 19873 31401 19876
rect 31435 19873 31447 19907
rect 31726 19904 31754 19944
rect 33505 19907 33563 19913
rect 33505 19904 33517 19907
rect 31726 19876 33517 19904
rect 31389 19867 31447 19873
rect 33505 19873 33517 19876
rect 33551 19873 33563 19907
rect 33505 19867 33563 19873
rect 14645 19839 14703 19845
rect 14645 19836 14657 19839
rect 14608 19808 14657 19836
rect 14608 19796 14614 19808
rect 14645 19805 14657 19808
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19836 15807 19839
rect 15838 19836 15844 19848
rect 15795 19808 15844 19836
rect 15795 19805 15807 19808
rect 15749 19799 15807 19805
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 18782 19836 18788 19848
rect 17144 19808 18788 19836
rect 6270 19768 6276 19780
rect 6012 19740 6276 19768
rect 6270 19728 6276 19740
rect 6328 19728 6334 19780
rect 8052 19771 8110 19777
rect 8052 19737 8064 19771
rect 8098 19768 8110 19771
rect 8941 19771 8999 19777
rect 8941 19768 8953 19771
rect 8098 19740 8953 19768
rect 8098 19737 8110 19740
rect 8052 19731 8110 19737
rect 8941 19737 8953 19740
rect 8987 19737 8999 19771
rect 8941 19731 8999 19737
rect 13204 19771 13262 19777
rect 13204 19737 13216 19771
rect 13250 19768 13262 19771
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13250 19740 14105 19768
rect 13250 19737 13262 19740
rect 13204 19731 13262 19737
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14093 19731 14151 19737
rect 16016 19771 16074 19777
rect 16016 19737 16028 19771
rect 16062 19768 16074 19771
rect 16482 19768 16488 19780
rect 16062 19740 16488 19768
rect 16062 19737 16074 19740
rect 16016 19731 16074 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 6365 19703 6423 19709
rect 6365 19700 6377 19703
rect 5460 19672 6377 19700
rect 6365 19669 6377 19672
rect 6411 19669 6423 19703
rect 6365 19663 6423 19669
rect 6454 19660 6460 19712
rect 6512 19660 6518 19712
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 8570 19700 8576 19712
rect 6972 19672 8576 19700
rect 6972 19660 6978 19672
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 8665 19703 8723 19709
rect 8665 19669 8677 19703
rect 8711 19700 8723 19703
rect 10226 19700 10232 19712
rect 8711 19672 10232 19700
rect 8711 19669 8723 19672
rect 8665 19663 8723 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 12069 19703 12127 19709
rect 12069 19669 12081 19703
rect 12115 19700 12127 19703
rect 12434 19700 12440 19712
rect 12115 19672 12440 19700
rect 12115 19669 12127 19672
rect 12069 19663 12127 19669
rect 12434 19660 12440 19672
rect 12492 19700 12498 19712
rect 12894 19700 12900 19712
rect 12492 19672 12900 19700
rect 12492 19660 12498 19672
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13817 19703 13875 19709
rect 13817 19669 13829 19703
rect 13863 19700 13875 19703
rect 13998 19700 14004 19712
rect 13863 19672 14004 19700
rect 13863 19669 13875 19672
rect 13817 19663 13875 19669
rect 13998 19660 14004 19672
rect 14056 19700 14062 19712
rect 17144 19700 17172 19808
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 21266 19796 21272 19848
rect 21324 19796 21330 19848
rect 22281 19839 22339 19845
rect 22281 19836 22293 19839
rect 21376 19808 22293 19836
rect 18356 19771 18414 19777
rect 18356 19737 18368 19771
rect 18402 19768 18414 19771
rect 19245 19771 19303 19777
rect 19245 19768 19257 19771
rect 18402 19740 19257 19768
rect 18402 19737 18414 19740
rect 18356 19731 18414 19737
rect 19245 19737 19257 19740
rect 19291 19737 19303 19771
rect 19245 19731 19303 19737
rect 21376 19712 21404 19808
rect 22281 19805 22293 19808
rect 22327 19836 22339 19839
rect 22554 19836 22560 19848
rect 22327 19808 22560 19836
rect 22327 19805 22339 19808
rect 22281 19799 22339 19805
rect 22554 19796 22560 19808
rect 22612 19796 22618 19848
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 24121 19839 24179 19845
rect 24121 19836 24133 19839
rect 23348 19808 24133 19836
rect 23348 19796 23354 19808
rect 24121 19805 24133 19808
rect 24167 19805 24179 19839
rect 24121 19799 24179 19805
rect 25130 19796 25136 19848
rect 25188 19836 25194 19848
rect 25501 19839 25559 19845
rect 25501 19836 25513 19839
rect 25188 19808 25513 19836
rect 25188 19796 25194 19808
rect 25501 19805 25513 19808
rect 25547 19836 25559 19839
rect 27985 19839 28043 19845
rect 27985 19836 27997 19839
rect 25547 19808 27997 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 27985 19805 27997 19808
rect 28031 19836 28043 19839
rect 28074 19836 28080 19848
rect 28031 19808 28080 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 30374 19845 30380 19848
rect 30352 19839 30380 19845
rect 30352 19805 30364 19839
rect 30352 19799 30380 19805
rect 30374 19796 30380 19799
rect 30432 19796 30438 19848
rect 31018 19796 31024 19848
rect 31076 19796 31082 19848
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19836 31263 19839
rect 31294 19836 31300 19848
rect 31251 19808 31300 19836
rect 31251 19805 31263 19808
rect 31205 19799 31263 19805
rect 31294 19796 31300 19808
rect 31352 19796 31358 19848
rect 23109 19771 23167 19777
rect 23109 19737 23121 19771
rect 23155 19768 23167 19771
rect 23569 19771 23627 19777
rect 23569 19768 23581 19771
rect 23155 19740 23581 19768
rect 23155 19737 23167 19740
rect 23109 19731 23167 19737
rect 23569 19737 23581 19740
rect 23615 19737 23627 19771
rect 23569 19731 23627 19737
rect 24673 19771 24731 19777
rect 24673 19737 24685 19771
rect 24719 19768 24731 19771
rect 25768 19771 25826 19777
rect 24719 19740 25728 19768
rect 24719 19737 24731 19740
rect 24673 19731 24731 19737
rect 14056 19672 17172 19700
rect 17221 19703 17279 19709
rect 14056 19660 14062 19672
rect 17221 19669 17233 19703
rect 17267 19700 17279 19703
rect 18046 19700 18052 19712
rect 17267 19672 18052 19700
rect 17267 19669 17279 19672
rect 17221 19663 17279 19669
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 20717 19703 20775 19709
rect 20717 19669 20729 19703
rect 20763 19700 20775 19703
rect 20806 19700 20812 19712
rect 20763 19672 20812 19700
rect 20763 19669 20775 19672
rect 20717 19663 20775 19669
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 21358 19660 21364 19712
rect 21416 19660 21422 19712
rect 21726 19660 21732 19712
rect 21784 19660 21790 19712
rect 22186 19660 22192 19712
rect 22244 19660 22250 19712
rect 23198 19660 23204 19712
rect 23256 19700 23262 19712
rect 24688 19700 24716 19731
rect 23256 19672 24716 19700
rect 25409 19703 25467 19709
rect 23256 19660 23262 19672
rect 25409 19669 25421 19703
rect 25455 19700 25467 19703
rect 25498 19700 25504 19712
rect 25455 19672 25504 19700
rect 25455 19669 25467 19672
rect 25409 19663 25467 19669
rect 25498 19660 25504 19672
rect 25556 19660 25562 19712
rect 25700 19700 25728 19740
rect 25768 19737 25780 19771
rect 25814 19768 25826 19771
rect 26970 19768 26976 19780
rect 25814 19740 26976 19768
rect 25814 19737 25826 19740
rect 25768 19731 25826 19737
rect 26970 19728 26976 19740
rect 27028 19728 27034 19780
rect 28252 19771 28310 19777
rect 28252 19737 28264 19771
rect 28298 19768 28310 19771
rect 28534 19768 28540 19780
rect 28298 19740 28540 19768
rect 28298 19737 28310 19740
rect 28252 19731 28310 19737
rect 28534 19728 28540 19740
rect 28592 19728 28598 19780
rect 31404 19768 31432 19867
rect 32030 19796 32036 19848
rect 32088 19796 32094 19848
rect 32769 19839 32827 19845
rect 32769 19805 32781 19839
rect 32815 19805 32827 19839
rect 32769 19799 32827 19805
rect 34517 19839 34575 19845
rect 34517 19805 34529 19839
rect 34563 19836 34575 19839
rect 34882 19836 34888 19848
rect 34563 19808 34888 19836
rect 34563 19805 34575 19808
rect 34517 19799 34575 19805
rect 32784 19768 32812 19799
rect 34882 19796 34888 19808
rect 34940 19796 34946 19848
rect 35342 19796 35348 19848
rect 35400 19796 35406 19848
rect 36081 19839 36139 19845
rect 36081 19805 36093 19839
rect 36127 19836 36139 19839
rect 36446 19836 36452 19848
rect 36127 19808 36452 19836
rect 36127 19805 36139 19808
rect 36081 19799 36139 19805
rect 36446 19796 36452 19808
rect 36504 19796 36510 19848
rect 36814 19796 36820 19848
rect 36872 19796 36878 19848
rect 38470 19796 38476 19848
rect 38528 19796 38534 19848
rect 31404 19740 32812 19768
rect 25958 19700 25964 19712
rect 25700 19672 25964 19700
rect 25958 19660 25964 19672
rect 26016 19660 26022 19712
rect 27341 19703 27399 19709
rect 27341 19669 27353 19703
rect 27387 19700 27399 19703
rect 27522 19700 27528 19712
rect 27387 19672 27528 19700
rect 27387 19669 27399 19672
rect 27341 19663 27399 19669
rect 27522 19660 27528 19672
rect 27580 19660 27586 19712
rect 29549 19703 29607 19709
rect 29549 19669 29561 19703
rect 29595 19700 29607 19703
rect 29914 19700 29920 19712
rect 29595 19672 29920 19700
rect 29595 19669 29607 19672
rect 29549 19663 29607 19669
rect 29914 19660 29920 19672
rect 29972 19660 29978 19712
rect 30374 19660 30380 19712
rect 30432 19700 30438 19712
rect 31481 19703 31539 19709
rect 31481 19700 31493 19703
rect 30432 19672 31493 19700
rect 30432 19660 30438 19672
rect 31481 19669 31493 19672
rect 31527 19669 31539 19703
rect 31481 19663 31539 19669
rect 32214 19660 32220 19712
rect 32272 19660 32278 19712
rect 32950 19660 32956 19712
rect 33008 19660 33014 19712
rect 33778 19660 33784 19712
rect 33836 19700 33842 19712
rect 33873 19703 33931 19709
rect 33873 19700 33885 19703
rect 33836 19672 33885 19700
rect 33836 19660 33842 19672
rect 33873 19669 33885 19672
rect 33919 19669 33931 19703
rect 33873 19663 33931 19669
rect 34698 19660 34704 19712
rect 34756 19660 34762 19712
rect 35434 19660 35440 19712
rect 35492 19660 35498 19712
rect 36170 19660 36176 19712
rect 36228 19660 36234 19712
rect 37826 19660 37832 19712
rect 37884 19660 37890 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 2038 19456 2044 19508
rect 2096 19456 2102 19508
rect 3237 19499 3295 19505
rect 3237 19465 3249 19499
rect 3283 19496 3295 19499
rect 5166 19496 5172 19508
rect 3283 19468 5172 19496
rect 3283 19465 3295 19468
rect 3237 19459 3295 19465
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19360 1915 19363
rect 2056 19360 2084 19456
rect 1903 19332 2084 19360
rect 2124 19363 2182 19369
rect 1903 19329 1915 19332
rect 1857 19323 1915 19329
rect 2124 19329 2136 19363
rect 2170 19360 2182 19363
rect 2958 19360 2964 19372
rect 2170 19332 2964 19360
rect 2170 19329 2182 19332
rect 2124 19323 2182 19329
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3375 19332 3464 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3436 19304 3464 19332
rect 3418 19252 3424 19304
rect 3476 19252 3482 19304
rect 3528 19301 3556 19468
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 5721 19499 5779 19505
rect 5721 19496 5733 19499
rect 5408 19468 5733 19496
rect 5408 19456 5414 19468
rect 5721 19465 5733 19468
rect 5767 19465 5779 19499
rect 5721 19459 5779 19465
rect 6181 19499 6239 19505
rect 6181 19465 6193 19499
rect 6227 19496 6239 19499
rect 9490 19496 9496 19508
rect 6227 19468 9496 19496
rect 6227 19465 6239 19468
rect 6181 19459 6239 19465
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 12161 19499 12219 19505
rect 12161 19465 12173 19499
rect 12207 19496 12219 19499
rect 12250 19496 12256 19508
rect 12207 19468 12256 19496
rect 12207 19465 12219 19468
rect 12161 19459 12219 19465
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 12406 19468 12664 19496
rect 5074 19388 5080 19440
rect 5132 19428 5138 19440
rect 5813 19431 5871 19437
rect 5813 19428 5825 19431
rect 5132 19400 5825 19428
rect 5132 19388 5138 19400
rect 5813 19397 5825 19400
rect 5859 19397 5871 19431
rect 5813 19391 5871 19397
rect 6270 19388 6276 19440
rect 6328 19428 6334 19440
rect 6914 19428 6920 19440
rect 6328 19400 6920 19428
rect 6328 19388 6334 19400
rect 6914 19388 6920 19400
rect 6972 19388 6978 19440
rect 8588 19400 9812 19428
rect 8588 19372 8616 19400
rect 4246 19320 4252 19372
rect 4304 19320 4310 19372
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 7742 19369 7748 19372
rect 7720 19363 7748 19369
rect 5684 19332 7052 19360
rect 5684 19320 5690 19332
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19261 3571 19295
rect 4366 19295 4424 19301
rect 4366 19292 4378 19295
rect 3513 19255 3571 19261
rect 4080 19264 4378 19292
rect 4080 19236 4108 19264
rect 4366 19261 4378 19264
rect 4412 19261 4424 19295
rect 4366 19255 4424 19261
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 5537 19295 5595 19301
rect 4571 19264 5488 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 3973 19227 4031 19233
rect 3973 19193 3985 19227
rect 4019 19193 4031 19227
rect 3973 19187 4031 19193
rect 3988 19156 4016 19187
rect 4062 19184 4068 19236
rect 4120 19184 4126 19236
rect 5460 19224 5488 19264
rect 5537 19261 5549 19295
rect 5583 19292 5595 19295
rect 5583 19264 6500 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 5092 19196 5396 19224
rect 5460 19196 5672 19224
rect 5092 19156 5120 19196
rect 3988 19128 5120 19156
rect 5166 19116 5172 19168
rect 5224 19116 5230 19168
rect 5368 19156 5396 19196
rect 5644 19168 5672 19196
rect 5534 19156 5540 19168
rect 5368 19128 5540 19156
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 5626 19116 5632 19168
rect 5684 19116 5690 19168
rect 6472 19156 6500 19264
rect 6914 19252 6920 19304
rect 6972 19252 6978 19304
rect 7024 19292 7052 19332
rect 7720 19329 7732 19363
rect 7720 19323 7748 19329
rect 7742 19320 7748 19323
rect 7800 19320 7806 19372
rect 8570 19320 8576 19372
rect 8628 19320 8634 19372
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8720 19332 8769 19360
rect 8720 19320 8726 19332
rect 8757 19329 8769 19332
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 8846 19320 8852 19372
rect 8904 19360 8910 19372
rect 9217 19363 9275 19369
rect 8904 19332 9168 19360
rect 8904 19320 8910 19332
rect 7024 19264 7236 19292
rect 6641 19159 6699 19165
rect 6641 19156 6653 19159
rect 6472 19128 6653 19156
rect 6641 19125 6653 19128
rect 6687 19156 6699 19159
rect 7098 19156 7104 19168
rect 6687 19128 7104 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7208 19156 7236 19264
rect 7558 19252 7564 19304
rect 7616 19252 7622 19304
rect 7834 19252 7840 19304
rect 7892 19252 7898 19304
rect 9140 19292 9168 19332
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9677 19363 9735 19369
rect 9677 19360 9689 19363
rect 9263 19332 9689 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9677 19329 9689 19332
rect 9723 19329 9735 19363
rect 9677 19323 9735 19329
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9140 19264 9321 19292
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 9309 19255 9367 19261
rect 9490 19252 9496 19304
rect 9548 19252 9554 19304
rect 9784 19292 9812 19400
rect 12406 19360 12434 19468
rect 12636 19428 12664 19468
rect 12710 19456 12716 19508
rect 12768 19456 12774 19508
rect 13078 19456 13084 19508
rect 13136 19456 13142 19508
rect 13817 19499 13875 19505
rect 13817 19465 13829 19499
rect 13863 19496 13875 19499
rect 14182 19496 14188 19508
rect 13863 19468 14188 19496
rect 13863 19465 13875 19468
rect 13817 19459 13875 19465
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 18690 19456 18696 19508
rect 18748 19456 18754 19508
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 21266 19496 21272 19508
rect 20947 19468 21272 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22244 19468 24072 19496
rect 22244 19456 22250 19468
rect 13096 19428 13124 19456
rect 12636 19400 13124 19428
rect 14366 19388 14372 19440
rect 14424 19428 14430 19440
rect 14461 19431 14519 19437
rect 14461 19428 14473 19431
rect 14424 19400 14473 19428
rect 14424 19388 14430 19400
rect 14461 19397 14473 19400
rect 14507 19428 14519 19431
rect 15654 19428 15660 19440
rect 14507 19400 15660 19428
rect 14507 19397 14519 19400
rect 14461 19391 14519 19397
rect 15654 19388 15660 19400
rect 15712 19388 15718 19440
rect 17313 19431 17371 19437
rect 17313 19397 17325 19431
rect 17359 19428 17371 19431
rect 22088 19431 22146 19437
rect 17359 19400 18276 19428
rect 17359 19397 17371 19400
rect 17313 19391 17371 19397
rect 18248 19372 18276 19400
rect 21284 19400 22048 19428
rect 12084 19332 12434 19360
rect 10229 19295 10287 19301
rect 10229 19292 10241 19295
rect 9784 19264 10241 19292
rect 10229 19261 10241 19264
rect 10275 19261 10287 19295
rect 10229 19255 10287 19261
rect 11333 19295 11391 19301
rect 11333 19261 11345 19295
rect 11379 19292 11391 19295
rect 11882 19292 11888 19304
rect 11379 19264 11888 19292
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 11882 19252 11888 19264
rect 11940 19252 11946 19304
rect 8113 19227 8171 19233
rect 8113 19193 8125 19227
rect 8159 19193 8171 19227
rect 8113 19187 8171 19193
rect 8128 19156 8156 19187
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 11514 19224 11520 19236
rect 8352 19196 11520 19224
rect 8352 19184 8358 19196
rect 11514 19184 11520 19196
rect 11572 19184 11578 19236
rect 7208 19128 8156 19156
rect 8846 19116 8852 19168
rect 8904 19116 8910 19168
rect 10689 19159 10747 19165
rect 10689 19125 10701 19159
rect 10735 19156 10747 19159
rect 11701 19159 11759 19165
rect 11701 19156 11713 19159
rect 10735 19128 11713 19156
rect 10735 19125 10747 19128
rect 10689 19119 10747 19125
rect 11701 19125 11713 19128
rect 11747 19156 11759 19159
rect 12084 19156 12112 19332
rect 12618 19320 12624 19372
rect 12676 19320 12682 19372
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 13173 19363 13231 19369
rect 13173 19360 13185 19363
rect 12952 19332 13185 19360
rect 12952 19320 12958 19332
rect 13173 19329 13185 19332
rect 13219 19329 13231 19363
rect 13173 19323 13231 19329
rect 15856 19332 18000 19360
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12308 19264 12817 19292
rect 12308 19252 12314 19264
rect 12805 19261 12817 19264
rect 12851 19292 12863 19295
rect 13814 19292 13820 19304
rect 12851 19264 13820 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 13814 19252 13820 19264
rect 13872 19292 13878 19304
rect 14458 19292 14464 19304
rect 13872 19264 14464 19292
rect 13872 19252 13878 19264
rect 14458 19252 14464 19264
rect 14516 19292 14522 19304
rect 15856 19292 15884 19332
rect 14516 19264 15884 19292
rect 14516 19252 14522 19264
rect 17402 19252 17408 19304
rect 17460 19252 17466 19304
rect 17586 19252 17592 19304
rect 17644 19252 17650 19304
rect 17972 19292 18000 19332
rect 18046 19320 18052 19372
rect 18104 19320 18110 19372
rect 18230 19320 18236 19372
rect 18288 19320 18294 19372
rect 18874 19360 18880 19372
rect 18340 19332 18880 19360
rect 18340 19292 18368 19332
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 21284 19369 21312 19400
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19329 21327 19363
rect 21269 19323 21327 19329
rect 21358 19320 21364 19372
rect 21416 19320 21422 19372
rect 21542 19320 21548 19372
rect 21600 19360 21606 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21600 19332 21833 19360
rect 21600 19320 21606 19332
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 22020 19360 22048 19400
rect 22088 19397 22100 19431
rect 22134 19428 22146 19431
rect 22646 19428 22652 19440
rect 22134 19400 22652 19428
rect 22134 19397 22146 19400
rect 22088 19391 22146 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 24044 19437 24072 19468
rect 25222 19456 25228 19508
rect 25280 19456 25286 19508
rect 25958 19456 25964 19508
rect 26016 19496 26022 19508
rect 26418 19496 26424 19508
rect 26016 19468 26424 19496
rect 26016 19456 26022 19468
rect 26418 19456 26424 19468
rect 26476 19496 26482 19508
rect 26694 19496 26700 19508
rect 26476 19468 26700 19496
rect 26476 19456 26482 19468
rect 26694 19456 26700 19468
rect 26752 19456 26758 19508
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28902 19496 28908 19508
rect 28132 19468 28908 19496
rect 28132 19456 28138 19468
rect 28902 19456 28908 19468
rect 28960 19496 28966 19508
rect 29362 19496 29368 19508
rect 28960 19468 29040 19496
rect 28960 19456 28966 19468
rect 23293 19431 23351 19437
rect 23293 19397 23305 19431
rect 23339 19397 23351 19431
rect 23293 19391 23351 19397
rect 24029 19431 24087 19437
rect 24029 19397 24041 19431
rect 24075 19397 24087 19431
rect 24029 19391 24087 19397
rect 23308 19360 23336 19391
rect 22020 19332 23336 19360
rect 25041 19363 25099 19369
rect 21821 19323 21879 19329
rect 25041 19329 25053 19363
rect 25087 19360 25099 19363
rect 25130 19360 25136 19372
rect 25087 19332 25136 19360
rect 25087 19329 25099 19332
rect 25041 19323 25099 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25240 19360 25268 19456
rect 25297 19363 25355 19369
rect 25297 19360 25309 19363
rect 25240 19332 25309 19360
rect 25297 19329 25309 19332
rect 25343 19329 25355 19363
rect 25297 19323 25355 19329
rect 26973 19363 27031 19369
rect 26973 19329 26985 19363
rect 27019 19360 27031 19363
rect 27062 19360 27068 19372
rect 27019 19332 27068 19360
rect 27019 19329 27031 19332
rect 26973 19323 27031 19329
rect 27062 19320 27068 19332
rect 27120 19320 27126 19372
rect 27154 19320 27160 19372
rect 27212 19320 27218 19372
rect 27890 19320 27896 19372
rect 27948 19320 27954 19372
rect 29012 19369 29040 19468
rect 29104 19468 29368 19496
rect 28997 19363 29055 19369
rect 28997 19329 29009 19363
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 17972 19264 18368 19292
rect 21453 19295 21511 19301
rect 21453 19261 21465 19295
rect 21499 19292 21511 19295
rect 21726 19292 21732 19304
rect 21499 19264 21732 19292
rect 21499 19261 21511 19264
rect 21453 19255 21511 19261
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 23290 19252 23296 19304
rect 23348 19252 23354 19304
rect 23845 19295 23903 19301
rect 23845 19261 23857 19295
rect 23891 19261 23903 19295
rect 23845 19255 23903 19261
rect 11747 19128 12112 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 12250 19116 12256 19168
rect 12308 19116 12314 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15896 19128 15945 19156
rect 15896 19116 15902 19128
rect 15933 19125 15945 19128
rect 15979 19156 15991 19159
rect 16022 19156 16028 19168
rect 15979 19128 16028 19156
rect 15979 19125 15991 19128
rect 15933 19119 15991 19125
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16942 19116 16948 19168
rect 17000 19116 17006 19168
rect 21744 19156 21772 19252
rect 23201 19227 23259 19233
rect 23201 19193 23213 19227
rect 23247 19224 23259 19227
rect 23308 19224 23336 19252
rect 23247 19196 23336 19224
rect 23247 19193 23259 19196
rect 23201 19187 23259 19193
rect 22554 19156 22560 19168
rect 21744 19128 22560 19156
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 22830 19116 22836 19168
rect 22888 19156 22894 19168
rect 23860 19156 23888 19255
rect 24578 19252 24584 19304
rect 24636 19252 24642 19304
rect 26878 19292 26884 19304
rect 26436 19264 26884 19292
rect 26436 19233 26464 19264
rect 26878 19252 26884 19264
rect 26936 19292 26942 19304
rect 28010 19295 28068 19301
rect 28010 19292 28022 19295
rect 26936 19264 28022 19292
rect 26936 19252 26942 19264
rect 28010 19261 28022 19264
rect 28056 19261 28068 19295
rect 28010 19255 28068 19261
rect 28166 19252 28172 19304
rect 28224 19292 28230 19304
rect 29104 19292 29132 19468
rect 29362 19456 29368 19468
rect 29420 19456 29426 19508
rect 30374 19456 30380 19508
rect 30432 19456 30438 19508
rect 30745 19499 30803 19505
rect 30745 19465 30757 19499
rect 30791 19496 30803 19499
rect 32214 19496 32220 19508
rect 30791 19468 32220 19496
rect 30791 19465 30803 19468
rect 30745 19459 30803 19465
rect 32214 19456 32220 19468
rect 32272 19456 32278 19508
rect 34425 19499 34483 19505
rect 34425 19465 34437 19499
rect 34471 19496 34483 19499
rect 34698 19496 34704 19508
rect 34471 19468 34704 19496
rect 34471 19465 34483 19468
rect 34425 19459 34483 19465
rect 34698 19456 34704 19468
rect 34756 19456 34762 19508
rect 34882 19456 34888 19508
rect 34940 19456 34946 19508
rect 35345 19499 35403 19505
rect 35345 19465 35357 19499
rect 35391 19496 35403 19499
rect 35434 19496 35440 19508
rect 35391 19468 35440 19496
rect 35391 19465 35403 19468
rect 35345 19459 35403 19465
rect 35434 19456 35440 19468
rect 35492 19456 35498 19508
rect 35989 19499 36047 19505
rect 35989 19465 36001 19499
rect 36035 19496 36047 19499
rect 36170 19496 36176 19508
rect 36035 19468 36176 19496
rect 36035 19465 36047 19468
rect 35989 19459 36047 19465
rect 36170 19456 36176 19468
rect 36228 19456 36234 19508
rect 36449 19499 36507 19505
rect 36449 19465 36461 19499
rect 36495 19465 36507 19499
rect 36449 19459 36507 19465
rect 29264 19431 29322 19437
rect 29264 19397 29276 19431
rect 29310 19428 29322 19431
rect 30392 19428 30420 19456
rect 31018 19428 31024 19440
rect 29310 19400 30420 19428
rect 30760 19400 31024 19428
rect 29310 19397 29322 19400
rect 29264 19391 29322 19397
rect 30760 19360 30788 19400
rect 31018 19388 31024 19400
rect 31076 19388 31082 19440
rect 32030 19428 32036 19440
rect 31220 19400 32036 19428
rect 28224 19264 29132 19292
rect 30392 19332 30788 19360
rect 30837 19363 30895 19369
rect 28224 19252 28230 19264
rect 26421 19227 26479 19233
rect 26421 19193 26433 19227
rect 26467 19193 26479 19227
rect 26421 19187 26479 19193
rect 27617 19227 27675 19233
rect 27617 19193 27629 19227
rect 27663 19193 27675 19227
rect 28902 19224 28908 19236
rect 27617 19187 27675 19193
rect 28552 19196 28908 19224
rect 22888 19128 23888 19156
rect 22888 19116 22894 19128
rect 25406 19116 25412 19168
rect 25464 19156 25470 19168
rect 27632 19156 27660 19187
rect 28552 19156 28580 19196
rect 28902 19184 28908 19196
rect 28960 19184 28966 19236
rect 30392 19233 30420 19332
rect 30837 19329 30849 19363
rect 30883 19360 30895 19363
rect 30926 19360 30932 19372
rect 30883 19332 30932 19360
rect 30883 19329 30895 19332
rect 30837 19323 30895 19329
rect 30926 19320 30932 19332
rect 30984 19320 30990 19372
rect 30653 19295 30711 19301
rect 30653 19261 30665 19295
rect 30699 19292 30711 19295
rect 30742 19292 30748 19304
rect 30699 19264 30748 19292
rect 30699 19261 30711 19264
rect 30653 19255 30711 19261
rect 30742 19252 30748 19264
rect 30800 19252 30806 19304
rect 31220 19233 31248 19400
rect 32030 19388 32036 19400
rect 32088 19388 32094 19440
rect 31846 19320 31852 19372
rect 31904 19320 31910 19372
rect 34517 19363 34575 19369
rect 34517 19329 34529 19363
rect 34563 19360 34575 19363
rect 34698 19360 34704 19372
rect 34563 19332 34704 19360
rect 34563 19329 34575 19332
rect 34517 19323 34575 19329
rect 34698 19320 34704 19332
rect 34756 19360 34762 19372
rect 35253 19363 35311 19369
rect 35253 19360 35265 19363
rect 34756 19332 35265 19360
rect 34756 19320 34762 19332
rect 35253 19329 35265 19332
rect 35299 19360 35311 19363
rect 36081 19363 36139 19369
rect 36081 19360 36093 19363
rect 35299 19332 36093 19360
rect 35299 19329 35311 19332
rect 35253 19323 35311 19329
rect 36081 19329 36093 19332
rect 36127 19329 36139 19363
rect 36464 19360 36492 19459
rect 36538 19388 36544 19440
rect 36596 19428 36602 19440
rect 37277 19431 37335 19437
rect 37277 19428 37289 19431
rect 36596 19400 37289 19428
rect 36596 19388 36602 19400
rect 37277 19397 37289 19400
rect 37323 19397 37335 19431
rect 37277 19391 37335 19397
rect 36464 19332 37872 19360
rect 36081 19323 36139 19329
rect 33965 19295 34023 19301
rect 33965 19261 33977 19295
rect 34011 19292 34023 19295
rect 34609 19295 34667 19301
rect 34011 19264 34100 19292
rect 34011 19261 34023 19264
rect 33965 19255 34023 19261
rect 34072 19233 34100 19264
rect 34609 19261 34621 19295
rect 34655 19261 34667 19295
rect 35437 19295 35495 19301
rect 35437 19292 35449 19295
rect 34609 19255 34667 19261
rect 34716 19264 35449 19292
rect 30377 19227 30435 19233
rect 30377 19193 30389 19227
rect 30423 19193 30435 19227
rect 30377 19187 30435 19193
rect 31205 19227 31263 19233
rect 31205 19193 31217 19227
rect 31251 19193 31263 19227
rect 31205 19187 31263 19193
rect 33229 19227 33287 19233
rect 33229 19193 33241 19227
rect 33275 19224 33287 19227
rect 34057 19227 34115 19233
rect 33275 19196 33456 19224
rect 33275 19193 33287 19196
rect 33229 19187 33287 19193
rect 33428 19168 33456 19196
rect 34057 19193 34069 19227
rect 34103 19193 34115 19227
rect 34624 19224 34652 19255
rect 34057 19187 34115 19193
rect 34440 19196 34652 19224
rect 25464 19128 28580 19156
rect 28813 19159 28871 19165
rect 25464 19116 25470 19128
rect 28813 19125 28825 19159
rect 28859 19156 28871 19159
rect 30006 19156 30012 19168
rect 28859 19128 30012 19156
rect 28859 19125 28871 19128
rect 28813 19119 28871 19125
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 31294 19116 31300 19168
rect 31352 19116 31358 19168
rect 33318 19116 33324 19168
rect 33376 19116 33382 19168
rect 33410 19116 33416 19168
rect 33468 19156 33474 19168
rect 34440 19156 34468 19196
rect 33468 19128 34468 19156
rect 33468 19116 33474 19128
rect 34606 19116 34612 19168
rect 34664 19156 34670 19168
rect 34716 19156 34744 19264
rect 35437 19261 35449 19264
rect 35483 19261 35495 19295
rect 35437 19255 35495 19261
rect 35897 19295 35955 19301
rect 35897 19261 35909 19295
rect 35943 19292 35955 19295
rect 35986 19292 35992 19304
rect 35943 19264 35992 19292
rect 35943 19261 35955 19264
rect 35897 19255 35955 19261
rect 35986 19252 35992 19264
rect 36044 19292 36050 19304
rect 37844 19301 37872 19332
rect 36725 19295 36783 19301
rect 36725 19292 36737 19295
rect 36044 19264 36737 19292
rect 36044 19252 36050 19264
rect 36725 19261 36737 19264
rect 36771 19261 36783 19295
rect 36725 19255 36783 19261
rect 37829 19295 37887 19301
rect 37829 19261 37841 19295
rect 37875 19261 37887 19295
rect 37829 19255 37887 19261
rect 34664 19128 34744 19156
rect 34664 19116 34670 19128
rect 35342 19116 35348 19168
rect 35400 19156 35406 19168
rect 35894 19156 35900 19168
rect 35400 19128 35900 19156
rect 35400 19116 35406 19128
rect 35894 19116 35900 19128
rect 35952 19116 35958 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 4614 18912 4620 18964
rect 4672 18912 4678 18964
rect 5166 18912 5172 18964
rect 5224 18912 5230 18964
rect 6914 18952 6920 18964
rect 5828 18924 6920 18952
rect 3418 18844 3424 18896
rect 3476 18884 3482 18896
rect 3605 18887 3663 18893
rect 3605 18884 3617 18887
rect 3476 18856 3617 18884
rect 3476 18844 3482 18856
rect 3605 18853 3617 18856
rect 3651 18884 3663 18887
rect 3651 18856 4844 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 2038 18776 2044 18828
rect 2096 18816 2102 18828
rect 2225 18819 2283 18825
rect 2225 18816 2237 18819
rect 2096 18788 2237 18816
rect 2096 18776 2102 18788
rect 2225 18785 2237 18788
rect 2271 18785 2283 18819
rect 2225 18779 2283 18785
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4614 18816 4620 18828
rect 4479 18788 4620 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 3786 18748 3792 18760
rect 1627 18720 3792 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 4706 18748 4712 18760
rect 4203 18720 4712 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 4816 18748 4844 18856
rect 5184 18816 5212 18912
rect 5828 18825 5856 18924
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 7926 18952 7932 18964
rect 7024 18924 7932 18952
rect 7024 18884 7052 18924
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 8389 18955 8447 18961
rect 8389 18921 8401 18955
rect 8435 18952 8447 18955
rect 8570 18952 8576 18964
rect 8435 18924 8576 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 8757 18955 8815 18961
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 10042 18952 10048 18964
rect 8803 18924 10048 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 6104 18856 7052 18884
rect 6104 18828 6132 18856
rect 5813 18819 5871 18825
rect 5184 18788 5764 18816
rect 5736 18757 5764 18788
rect 5813 18785 5825 18819
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18816 6055 18819
rect 6086 18816 6092 18828
rect 6043 18788 6092 18816
rect 6043 18785 6055 18788
rect 5997 18779 6055 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6825 18819 6883 18825
rect 6825 18785 6837 18819
rect 6871 18816 6883 18819
rect 6871 18788 7144 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 5169 18751 5227 18757
rect 5169 18748 5181 18751
rect 4816 18720 5181 18748
rect 5169 18717 5181 18720
rect 5215 18717 5227 18751
rect 5169 18711 5227 18717
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 6362 18708 6368 18760
rect 6420 18748 6426 18760
rect 7009 18751 7067 18757
rect 7009 18748 7021 18751
rect 6420 18720 7021 18748
rect 6420 18708 6426 18720
rect 7009 18717 7021 18720
rect 7055 18717 7067 18751
rect 7116 18748 7144 18788
rect 8570 18748 8576 18760
rect 7116 18720 8576 18748
rect 7009 18711 7067 18717
rect 8570 18708 8576 18720
rect 8628 18748 8634 18760
rect 8772 18748 8800 18915
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 12710 18952 12716 18964
rect 12406 18924 12716 18952
rect 12406 18884 12434 18924
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 12802 18912 12808 18964
rect 12860 18912 12866 18964
rect 16482 18912 16488 18964
rect 16540 18912 16546 18964
rect 17313 18955 17371 18961
rect 17313 18921 17325 18955
rect 17359 18952 17371 18955
rect 17402 18952 17408 18964
rect 17359 18924 17408 18952
rect 17359 18921 17371 18924
rect 17313 18915 17371 18921
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 21361 18955 21419 18961
rect 21361 18921 21373 18955
rect 21407 18952 21419 18955
rect 22370 18952 22376 18964
rect 21407 18924 22376 18952
rect 21407 18921 21419 18924
rect 21361 18915 21419 18921
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 23290 18912 23296 18964
rect 23348 18912 23354 18964
rect 23658 18912 23664 18964
rect 23716 18952 23722 18964
rect 24302 18952 24308 18964
rect 23716 18924 24308 18952
rect 23716 18912 23722 18924
rect 24302 18912 24308 18924
rect 24360 18912 24366 18964
rect 24578 18912 24584 18964
rect 24636 18912 24642 18964
rect 25133 18955 25191 18961
rect 25133 18952 25145 18955
rect 24688 18924 25145 18952
rect 22830 18884 22836 18896
rect 9876 18856 12434 18884
rect 22572 18856 22836 18884
rect 8846 18776 8852 18828
rect 8904 18816 8910 18828
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 8904 18788 9505 18816
rect 8904 18776 8910 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 8628 18720 8800 18748
rect 8628 18708 8634 18720
rect 2133 18683 2191 18689
rect 2133 18649 2145 18683
rect 2179 18680 2191 18683
rect 2470 18683 2528 18689
rect 2470 18680 2482 18683
rect 2179 18652 2482 18680
rect 2179 18649 2191 18652
rect 2133 18643 2191 18649
rect 2470 18649 2482 18652
rect 2516 18649 2528 18683
rect 6549 18683 6607 18689
rect 6549 18680 6561 18683
rect 2470 18643 2528 18649
rect 5092 18652 6561 18680
rect 5092 18624 5120 18652
rect 6549 18649 6561 18652
rect 6595 18649 6607 18683
rect 6549 18643 6607 18649
rect 7276 18683 7334 18689
rect 7276 18649 7288 18683
rect 7322 18680 7334 18683
rect 8941 18683 8999 18689
rect 8941 18680 8953 18683
rect 7322 18652 8953 18680
rect 7322 18649 7334 18652
rect 7276 18643 7334 18649
rect 8941 18649 8953 18652
rect 8987 18649 8999 18683
rect 8941 18643 8999 18649
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 5074 18612 5080 18624
rect 4304 18584 5080 18612
rect 4304 18572 4310 18584
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 5353 18615 5411 18621
rect 5353 18581 5365 18615
rect 5399 18612 5411 18615
rect 5718 18612 5724 18624
rect 5399 18584 5724 18612
rect 5399 18581 5411 18584
rect 5353 18575 5411 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 6178 18572 6184 18624
rect 6236 18572 6242 18624
rect 6641 18615 6699 18621
rect 6641 18581 6653 18615
rect 6687 18612 6699 18615
rect 6822 18612 6828 18624
rect 6687 18584 6828 18612
rect 6687 18581 6699 18584
rect 6641 18575 6699 18581
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9490 18612 9496 18624
rect 9272 18584 9496 18612
rect 9272 18572 9278 18584
rect 9490 18572 9496 18584
rect 9548 18612 9554 18624
rect 9876 18621 9904 18856
rect 12250 18776 12256 18828
rect 12308 18776 12314 18828
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 17037 18819 17095 18825
rect 17037 18816 17049 18819
rect 17000 18788 17049 18816
rect 17000 18776 17006 18788
rect 17037 18785 17049 18788
rect 17083 18785 17095 18819
rect 17037 18779 17095 18785
rect 17954 18776 17960 18828
rect 18012 18776 18018 18828
rect 21542 18776 21548 18828
rect 21600 18776 21606 18828
rect 22256 18819 22314 18825
rect 22256 18785 22268 18819
rect 22302 18816 22314 18819
rect 22572 18816 22600 18856
rect 22830 18844 22836 18856
rect 22888 18844 22894 18896
rect 22302 18788 22600 18816
rect 22649 18819 22707 18825
rect 22302 18785 22314 18788
rect 22256 18779 22314 18785
rect 22649 18785 22661 18819
rect 22695 18816 22707 18819
rect 23109 18819 23167 18825
rect 22695 18788 22968 18816
rect 22695 18785 22707 18788
rect 22649 18779 22707 18785
rect 11514 18708 11520 18760
rect 11572 18708 11578 18760
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 21560 18748 21588 18776
rect 22940 18760 22968 18788
rect 23109 18785 23121 18819
rect 23155 18816 23167 18819
rect 23308 18816 23336 18912
rect 23155 18788 23336 18816
rect 23155 18785 23167 18788
rect 23109 18779 23167 18785
rect 20027 18720 21588 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20088 18624 20116 18720
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 22922 18708 22928 18760
rect 22980 18748 22986 18760
rect 22980 18720 23152 18748
rect 22980 18708 22986 18720
rect 20248 18683 20306 18689
rect 20248 18649 20260 18683
rect 20294 18680 20306 18683
rect 20714 18680 20720 18692
rect 20294 18652 20720 18680
rect 20294 18649 20306 18652
rect 20248 18643 20306 18649
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 23124 18680 23152 18720
rect 23290 18708 23296 18760
rect 23348 18748 23354 18760
rect 24596 18748 24624 18912
rect 23348 18720 24624 18748
rect 23348 18708 23354 18720
rect 24026 18680 24032 18692
rect 23124 18652 24032 18680
rect 24026 18640 24032 18652
rect 24084 18680 24090 18692
rect 24688 18680 24716 18924
rect 25133 18921 25145 18924
rect 25179 18952 25191 18955
rect 25406 18952 25412 18964
rect 25179 18924 25412 18952
rect 25179 18921 25191 18924
rect 25133 18915 25191 18921
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 26605 18955 26663 18961
rect 26605 18921 26617 18955
rect 26651 18952 26663 18955
rect 27338 18952 27344 18964
rect 26651 18924 27344 18952
rect 26651 18921 26663 18924
rect 26605 18915 26663 18921
rect 27338 18912 27344 18924
rect 27396 18952 27402 18964
rect 27890 18952 27896 18964
rect 27396 18924 27896 18952
rect 27396 18912 27402 18924
rect 27890 18912 27896 18924
rect 27948 18912 27954 18964
rect 28810 18912 28816 18964
rect 28868 18952 28874 18964
rect 29273 18955 29331 18961
rect 29273 18952 29285 18955
rect 28868 18924 29285 18952
rect 28868 18912 28874 18924
rect 29273 18921 29285 18924
rect 29319 18952 29331 18955
rect 30650 18952 30656 18964
rect 29319 18924 30656 18952
rect 29319 18921 29331 18924
rect 29273 18915 29331 18921
rect 30650 18912 30656 18924
rect 30708 18912 30714 18964
rect 31113 18955 31171 18961
rect 31113 18921 31125 18955
rect 31159 18952 31171 18955
rect 31754 18952 31760 18964
rect 31159 18924 31760 18952
rect 31159 18921 31171 18924
rect 31113 18915 31171 18921
rect 31754 18912 31760 18924
rect 31812 18912 31818 18964
rect 34517 18955 34575 18961
rect 34517 18921 34529 18955
rect 34563 18952 34575 18955
rect 35342 18952 35348 18964
rect 34563 18924 35348 18952
rect 34563 18921 34575 18924
rect 34517 18915 34575 18921
rect 35342 18912 35348 18924
rect 35400 18912 35406 18964
rect 35434 18912 35440 18964
rect 35492 18952 35498 18964
rect 35802 18952 35808 18964
rect 35492 18924 35808 18952
rect 35492 18912 35498 18924
rect 35802 18912 35808 18924
rect 35860 18952 35866 18964
rect 35860 18924 37136 18952
rect 35860 18912 35866 18924
rect 28718 18844 28724 18896
rect 28776 18884 28782 18896
rect 28776 18856 31754 18884
rect 28776 18844 28782 18856
rect 31726 18828 31754 18856
rect 36814 18844 36820 18896
rect 36872 18844 36878 18896
rect 25130 18776 25136 18828
rect 25188 18816 25194 18828
rect 25225 18819 25283 18825
rect 25225 18816 25237 18819
rect 25188 18788 25237 18816
rect 25188 18776 25194 18788
rect 25225 18785 25237 18788
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 28074 18776 28080 18828
rect 28132 18776 28138 18828
rect 28810 18776 28816 18828
rect 28868 18816 28874 18828
rect 30101 18819 30159 18825
rect 30101 18816 30113 18819
rect 28868 18788 30113 18816
rect 28868 18776 28874 18788
rect 30101 18785 30113 18788
rect 30147 18785 30159 18819
rect 30101 18779 30159 18785
rect 30561 18819 30619 18825
rect 30561 18785 30573 18819
rect 30607 18816 30619 18819
rect 30834 18816 30840 18828
rect 30607 18788 30840 18816
rect 30607 18785 30619 18788
rect 30561 18779 30619 18785
rect 30834 18776 30840 18788
rect 30892 18816 30898 18828
rect 31389 18819 31447 18825
rect 31389 18816 31401 18819
rect 30892 18788 31401 18816
rect 30892 18776 30898 18788
rect 31389 18785 31401 18788
rect 31435 18785 31447 18819
rect 31726 18788 31760 18828
rect 31389 18779 31447 18785
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 35618 18816 35624 18828
rect 34164 18788 35624 18816
rect 25498 18757 25504 18760
rect 25492 18748 25504 18757
rect 25459 18720 25504 18748
rect 25492 18711 25504 18720
rect 25498 18708 25504 18711
rect 25556 18708 25562 18760
rect 28258 18708 28264 18760
rect 28316 18748 28322 18760
rect 28721 18751 28779 18757
rect 28721 18748 28733 18751
rect 28316 18720 28733 18748
rect 28316 18708 28322 18720
rect 28721 18717 28733 18720
rect 28767 18717 28779 18751
rect 28721 18711 28779 18717
rect 30745 18751 30803 18757
rect 30745 18717 30757 18751
rect 30791 18748 30803 18751
rect 32950 18748 32956 18760
rect 30791 18720 32956 18748
rect 30791 18717 30803 18720
rect 30745 18711 30803 18717
rect 32950 18708 32956 18720
rect 33008 18708 33014 18760
rect 33137 18751 33195 18757
rect 33137 18717 33149 18751
rect 33183 18748 33195 18751
rect 33226 18748 33232 18760
rect 33183 18720 33232 18748
rect 33183 18717 33195 18720
rect 33137 18711 33195 18717
rect 33226 18708 33232 18720
rect 33284 18708 33290 18760
rect 33404 18751 33462 18757
rect 33404 18717 33416 18751
rect 33450 18717 33462 18751
rect 34164 18748 34192 18788
rect 35618 18776 35624 18788
rect 35676 18816 35682 18828
rect 35805 18819 35863 18825
rect 35805 18816 35817 18819
rect 35676 18788 35817 18816
rect 35676 18776 35682 18788
rect 35805 18785 35817 18788
rect 35851 18785 35863 18819
rect 35805 18779 35863 18785
rect 35894 18776 35900 18828
rect 35952 18825 35958 18828
rect 35952 18819 36001 18825
rect 35952 18785 35955 18819
rect 35989 18785 36001 18819
rect 35952 18779 36001 18785
rect 36357 18819 36415 18825
rect 36357 18785 36369 18819
rect 36403 18816 36415 18819
rect 36722 18816 36728 18828
rect 36403 18788 36728 18816
rect 36403 18785 36415 18788
rect 36357 18779 36415 18785
rect 35952 18776 35958 18779
rect 36722 18776 36728 18788
rect 36780 18776 36786 18828
rect 36832 18816 36860 18844
rect 37108 18825 37136 18924
rect 38470 18912 38476 18964
rect 38528 18912 38534 18964
rect 37001 18819 37059 18825
rect 37001 18816 37013 18819
rect 36832 18788 37013 18816
rect 37001 18785 37013 18788
rect 37047 18785 37059 18819
rect 37001 18779 37059 18785
rect 37093 18819 37151 18825
rect 37093 18785 37105 18819
rect 37139 18785 37151 18819
rect 37093 18779 37151 18785
rect 33404 18711 33462 18717
rect 33520 18720 34192 18748
rect 24084 18652 24716 18680
rect 27832 18683 27890 18689
rect 24084 18640 24090 18652
rect 27832 18649 27844 18683
rect 27878 18680 27890 18683
rect 28169 18683 28227 18689
rect 28169 18680 28181 18683
rect 27878 18652 28181 18680
rect 27878 18649 27890 18652
rect 27832 18643 27890 18649
rect 28169 18649 28181 18652
rect 28215 18649 28227 18683
rect 29917 18683 29975 18689
rect 28169 18643 28227 18649
rect 28276 18652 29684 18680
rect 9861 18615 9919 18621
rect 9861 18612 9873 18615
rect 9548 18584 9873 18612
rect 9548 18572 9554 18584
rect 9861 18581 9873 18584
rect 9907 18581 9919 18615
rect 9861 18575 9919 18581
rect 10502 18572 10508 18624
rect 10560 18612 10566 18624
rect 10873 18615 10931 18621
rect 10873 18612 10885 18615
rect 10560 18584 10885 18612
rect 10560 18572 10566 18584
rect 10873 18581 10885 18584
rect 10919 18581 10931 18615
rect 10873 18575 10931 18581
rect 16393 18615 16451 18621
rect 16393 18581 16405 18615
rect 16439 18612 16451 18615
rect 17586 18612 17592 18624
rect 16439 18584 17592 18612
rect 16439 18581 16451 18584
rect 16393 18575 16451 18581
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 20070 18572 20076 18624
rect 20128 18572 20134 18624
rect 21453 18615 21511 18621
rect 21453 18581 21465 18615
rect 21499 18612 21511 18615
rect 22646 18612 22652 18624
rect 21499 18584 22652 18612
rect 21499 18581 21511 18584
rect 21453 18575 21511 18581
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 25590 18612 25596 18624
rect 22796 18584 25596 18612
rect 22796 18572 22802 18584
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 26697 18615 26755 18621
rect 26697 18581 26709 18615
rect 26743 18612 26755 18615
rect 27154 18612 27160 18624
rect 26743 18584 27160 18612
rect 26743 18581 26755 18584
rect 26697 18575 26755 18581
rect 27154 18572 27160 18584
rect 27212 18612 27218 18624
rect 27430 18612 27436 18624
rect 27212 18584 27436 18612
rect 27212 18572 27218 18584
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 27522 18572 27528 18624
rect 27580 18612 27586 18624
rect 28276 18612 28304 18652
rect 27580 18584 28304 18612
rect 27580 18572 27586 18584
rect 29546 18572 29552 18624
rect 29604 18572 29610 18624
rect 29656 18612 29684 18652
rect 29917 18649 29929 18683
rect 29963 18680 29975 18683
rect 31294 18680 31300 18692
rect 29963 18652 31300 18680
rect 29963 18649 29975 18652
rect 29917 18643 29975 18649
rect 31294 18640 31300 18652
rect 31352 18640 31358 18692
rect 33318 18640 33324 18692
rect 33376 18680 33382 18692
rect 33428 18680 33456 18711
rect 33376 18652 33456 18680
rect 33376 18640 33382 18652
rect 30009 18615 30067 18621
rect 30009 18612 30021 18615
rect 29656 18584 30021 18612
rect 30009 18581 30021 18584
rect 30055 18612 30067 18615
rect 30190 18612 30196 18624
rect 30055 18584 30196 18612
rect 30055 18581 30067 18584
rect 30009 18575 30067 18581
rect 30190 18572 30196 18584
rect 30248 18612 30254 18624
rect 30653 18615 30711 18621
rect 30653 18612 30665 18615
rect 30248 18584 30665 18612
rect 30248 18572 30254 18584
rect 30653 18581 30665 18584
rect 30699 18612 30711 18615
rect 30926 18612 30932 18624
rect 30699 18584 30932 18612
rect 30699 18581 30711 18584
rect 30653 18575 30711 18581
rect 30926 18572 30932 18584
rect 30984 18572 30990 18624
rect 33042 18572 33048 18624
rect 33100 18612 33106 18624
rect 33520 18612 33548 18720
rect 36078 18708 36084 18760
rect 36136 18708 36142 18760
rect 36817 18751 36875 18757
rect 36817 18717 36829 18751
rect 36863 18748 36875 18751
rect 38488 18748 38516 18912
rect 36863 18720 38516 18748
rect 36863 18717 36875 18720
rect 36817 18711 36875 18717
rect 37366 18689 37372 18692
rect 37360 18643 37372 18689
rect 37366 18640 37372 18643
rect 37424 18640 37430 18692
rect 33100 18584 33548 18612
rect 33100 18572 33106 18584
rect 34606 18572 34612 18624
rect 34664 18612 34670 18624
rect 34885 18615 34943 18621
rect 34885 18612 34897 18615
rect 34664 18584 34897 18612
rect 34664 18572 34670 18584
rect 34885 18581 34897 18584
rect 34931 18581 34943 18615
rect 34885 18575 34943 18581
rect 35161 18615 35219 18621
rect 35161 18581 35173 18615
rect 35207 18612 35219 18615
rect 37642 18612 37648 18624
rect 35207 18584 37648 18612
rect 35207 18581 35219 18584
rect 35161 18575 35219 18581
rect 37642 18572 37648 18584
rect 37700 18572 37706 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 4154 18408 4160 18420
rect 3896 18380 4160 18408
rect 2038 18232 2044 18284
rect 2096 18272 2102 18284
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 2096 18244 2329 18272
rect 2096 18232 2102 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 2584 18275 2642 18281
rect 2584 18241 2596 18275
rect 2630 18272 2642 18275
rect 3326 18272 3332 18284
rect 2630 18244 3332 18272
rect 2630 18241 2642 18244
rect 2584 18235 2642 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 3896 18213 3924 18380
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 7558 18408 7564 18420
rect 5684 18380 7564 18408
rect 5684 18368 5690 18380
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 7745 18411 7803 18417
rect 7745 18377 7757 18411
rect 7791 18408 7803 18411
rect 7834 18408 7840 18420
rect 7791 18380 7840 18408
rect 7791 18377 7803 18380
rect 7745 18371 7803 18377
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 10042 18368 10048 18420
rect 10100 18408 10106 18420
rect 10137 18411 10195 18417
rect 10137 18408 10149 18411
rect 10100 18380 10149 18408
rect 10100 18368 10106 18380
rect 10137 18377 10149 18380
rect 10183 18377 10195 18411
rect 10137 18371 10195 18377
rect 11514 18368 11520 18420
rect 11572 18368 11578 18420
rect 11977 18411 12035 18417
rect 11977 18377 11989 18411
rect 12023 18408 12035 18411
rect 12342 18408 12348 18420
rect 12023 18380 12348 18408
rect 12023 18377 12035 18380
rect 11977 18371 12035 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 21637 18411 21695 18417
rect 21637 18377 21649 18411
rect 21683 18377 21695 18411
rect 23658 18408 23664 18420
rect 21637 18371 21695 18377
rect 22296 18380 23664 18408
rect 4062 18340 4068 18352
rect 3988 18312 4068 18340
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 3697 18139 3755 18145
rect 3697 18105 3709 18139
rect 3743 18136 3755 18139
rect 3988 18136 4016 18312
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 9585 18343 9643 18349
rect 9585 18309 9597 18343
rect 9631 18340 9643 18343
rect 20898 18340 20904 18352
rect 9631 18312 20904 18340
rect 9631 18309 9643 18312
rect 9585 18303 9643 18309
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 4617 18275 4675 18281
rect 4617 18272 4629 18275
rect 4203 18244 4629 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4617 18241 4629 18244
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 6362 18232 6368 18284
rect 6420 18232 6426 18284
rect 6638 18281 6644 18284
rect 6632 18235 6644 18281
rect 6638 18232 6644 18235
rect 6696 18232 6702 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 11931 18244 13093 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 20070 18232 20076 18284
rect 20128 18272 20134 18284
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 20128 18244 20269 18272
rect 20128 18232 20134 18244
rect 20257 18241 20269 18244
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20524 18275 20582 18281
rect 20524 18241 20536 18275
rect 20570 18272 20582 18275
rect 20806 18272 20812 18284
rect 20570 18244 20812 18272
rect 20570 18241 20582 18244
rect 20524 18235 20582 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21652 18272 21680 18371
rect 22094 18300 22100 18352
rect 22152 18340 22158 18352
rect 22296 18340 22324 18380
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 25774 18368 25780 18420
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27249 18411 27307 18417
rect 27249 18408 27261 18411
rect 26283 18380 27261 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27249 18377 27261 18380
rect 27295 18408 27307 18411
rect 27522 18408 27528 18420
rect 27295 18380 27528 18408
rect 27295 18377 27307 18380
rect 27249 18371 27307 18377
rect 27522 18368 27528 18380
rect 27580 18368 27586 18420
rect 27709 18411 27767 18417
rect 27709 18377 27721 18411
rect 27755 18408 27767 18411
rect 28258 18408 28264 18420
rect 27755 18380 28264 18408
rect 27755 18377 27767 18380
rect 27709 18371 27767 18377
rect 28258 18368 28264 18380
rect 28316 18368 28322 18420
rect 28534 18368 28540 18420
rect 28592 18408 28598 18420
rect 28905 18411 28963 18417
rect 28905 18408 28917 18411
rect 28592 18380 28917 18408
rect 28592 18368 28598 18380
rect 28905 18377 28917 18380
rect 28951 18377 28963 18411
rect 28905 18371 28963 18377
rect 29546 18368 29552 18420
rect 29604 18368 29610 18420
rect 29914 18368 29920 18420
rect 29972 18368 29978 18420
rect 30006 18368 30012 18420
rect 30064 18368 30070 18420
rect 35434 18368 35440 18420
rect 35492 18368 35498 18420
rect 36449 18411 36507 18417
rect 36449 18377 36461 18411
rect 36495 18408 36507 18411
rect 36814 18408 36820 18420
rect 36495 18380 36820 18408
rect 36495 18377 36507 18380
rect 36449 18371 36507 18377
rect 36814 18368 36820 18380
rect 36872 18368 36878 18420
rect 37645 18411 37703 18417
rect 37645 18377 37657 18411
rect 37691 18408 37703 18411
rect 37826 18408 37832 18420
rect 37691 18380 37832 18408
rect 37691 18377 37703 18380
rect 37645 18371 37703 18377
rect 37826 18368 37832 18380
rect 37884 18368 37890 18420
rect 22152 18312 22324 18340
rect 22152 18300 22158 18312
rect 22830 18300 22836 18352
rect 22888 18300 22894 18352
rect 22956 18343 23014 18349
rect 22956 18309 22968 18343
rect 23002 18340 23014 18343
rect 23382 18340 23388 18352
rect 23002 18312 23388 18340
rect 23002 18309 23014 18312
rect 22956 18303 23014 18309
rect 23382 18300 23388 18312
rect 23440 18300 23446 18352
rect 24026 18300 24032 18352
rect 24084 18300 24090 18352
rect 26145 18343 26203 18349
rect 26145 18309 26157 18343
rect 26191 18340 26203 18343
rect 26326 18340 26332 18352
rect 26191 18312 26332 18340
rect 26191 18309 26203 18312
rect 26145 18303 26203 18309
rect 26326 18300 26332 18312
rect 26384 18300 26390 18352
rect 22848 18272 22876 18300
rect 21652 18244 22876 18272
rect 23290 18232 23296 18284
rect 23348 18232 23354 18284
rect 4065 18207 4123 18213
rect 4065 18173 4077 18207
rect 4111 18204 4123 18207
rect 4246 18204 4252 18216
rect 4111 18176 4252 18204
rect 4111 18173 4123 18176
rect 4065 18167 4123 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 4448 18176 5181 18204
rect 4448 18136 4476 18176
rect 5169 18173 5181 18176
rect 5215 18173 5227 18207
rect 5169 18167 5227 18173
rect 11330 18164 11336 18216
rect 11388 18164 11394 18216
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 3743 18108 4476 18136
rect 4525 18139 4583 18145
rect 3743 18105 3755 18108
rect 3697 18099 3755 18105
rect 4525 18105 4537 18139
rect 4571 18136 4583 18139
rect 4706 18136 4712 18148
rect 4571 18108 4712 18136
rect 4571 18105 4583 18108
rect 4525 18099 4583 18105
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 12084 18136 12112 18167
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12308 18176 12909 18204
rect 12308 18164 12314 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 13630 18164 13636 18216
rect 13688 18164 13694 18216
rect 15654 18164 15660 18216
rect 15712 18164 15718 18216
rect 16482 18164 16488 18216
rect 16540 18164 16546 18216
rect 17770 18164 17776 18216
rect 17828 18164 17834 18216
rect 23198 18164 23204 18216
rect 23256 18164 23262 18216
rect 14734 18136 14740 18148
rect 10520 18108 14740 18136
rect 6086 18028 6092 18080
rect 6144 18028 6150 18080
rect 8294 18028 8300 18080
rect 8352 18028 8358 18080
rect 10226 18028 10232 18080
rect 10284 18068 10290 18080
rect 10520 18077 10548 18108
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 16945 18139 17003 18145
rect 16945 18105 16957 18139
rect 16991 18136 17003 18139
rect 16991 18108 17908 18136
rect 16991 18105 17003 18108
rect 16945 18099 17003 18105
rect 17880 18080 17908 18108
rect 10505 18071 10563 18077
rect 10505 18068 10517 18071
rect 10284 18040 10517 18068
rect 10284 18028 10290 18040
rect 10505 18037 10517 18040
rect 10551 18037 10563 18071
rect 10505 18031 10563 18037
rect 10686 18028 10692 18080
rect 10744 18028 10750 18080
rect 12342 18028 12348 18080
rect 12400 18028 12406 18080
rect 15010 18028 15016 18080
rect 15068 18068 15074 18080
rect 15105 18071 15163 18077
rect 15105 18068 15117 18071
rect 15068 18040 15117 18068
rect 15068 18028 15074 18040
rect 15105 18037 15117 18040
rect 15151 18037 15163 18071
rect 15105 18031 15163 18037
rect 15838 18028 15844 18080
rect 15896 18028 15902 18080
rect 17218 18028 17224 18080
rect 17276 18028 17282 18080
rect 17862 18028 17868 18080
rect 17920 18028 17926 18080
rect 21821 18071 21879 18077
rect 21821 18037 21833 18071
rect 21867 18068 21879 18071
rect 23308 18068 23336 18232
rect 23937 18207 23995 18213
rect 23937 18173 23949 18207
rect 23983 18204 23995 18207
rect 24044 18204 24072 18300
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18272 24363 18275
rect 24578 18272 24584 18284
rect 24351 18244 24584 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 24578 18232 24584 18244
rect 24636 18232 24642 18284
rect 29564 18281 29592 18368
rect 33226 18300 33232 18352
rect 33284 18340 33290 18352
rect 35452 18340 35480 18368
rect 33284 18312 35480 18340
rect 33284 18300 33290 18312
rect 33520 18281 33548 18312
rect 33778 18281 33784 18284
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27801 18275 27859 18281
rect 27801 18272 27813 18275
rect 27387 18244 27813 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27801 18241 27813 18244
rect 27847 18241 27859 18275
rect 27801 18235 27859 18241
rect 29549 18275 29607 18281
rect 29549 18241 29561 18275
rect 29595 18241 29607 18275
rect 29549 18235 29607 18241
rect 33505 18275 33563 18281
rect 33505 18241 33517 18275
rect 33551 18241 33563 18275
rect 33772 18272 33784 18281
rect 33739 18244 33784 18272
rect 33505 18235 33563 18241
rect 33772 18235 33784 18244
rect 33778 18232 33784 18235
rect 33836 18232 33842 18284
rect 35084 18281 35112 18312
rect 35618 18300 35624 18352
rect 35676 18340 35682 18352
rect 36170 18340 36176 18352
rect 35676 18312 36176 18340
rect 35676 18300 35682 18312
rect 36170 18300 36176 18312
rect 36228 18300 36234 18352
rect 36538 18300 36544 18352
rect 36596 18300 36602 18352
rect 35069 18275 35127 18281
rect 35069 18241 35081 18275
rect 35115 18241 35127 18275
rect 35069 18235 35127 18241
rect 35336 18275 35394 18281
rect 35336 18241 35348 18275
rect 35382 18272 35394 18275
rect 36556 18272 36584 18300
rect 35382 18244 36584 18272
rect 35382 18241 35394 18244
rect 35336 18235 35394 18241
rect 23983 18176 24072 18204
rect 23983 18173 23995 18176
rect 23937 18167 23995 18173
rect 25590 18164 25596 18216
rect 25648 18204 25654 18216
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 25648 18176 25697 18204
rect 25648 18164 25654 18176
rect 25685 18173 25697 18176
rect 25731 18204 25743 18207
rect 26421 18207 26479 18213
rect 26421 18204 26433 18207
rect 25731 18176 26433 18204
rect 25731 18173 25743 18176
rect 25685 18167 25743 18173
rect 26421 18173 26433 18176
rect 26467 18204 26479 18207
rect 26510 18204 26516 18216
rect 26467 18176 26516 18204
rect 26467 18173 26479 18176
rect 26421 18167 26479 18173
rect 26510 18164 26516 18176
rect 26568 18164 26574 18216
rect 27157 18207 27215 18213
rect 27157 18173 27169 18207
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 27172 18136 27200 18167
rect 27430 18164 27436 18216
rect 27488 18204 27494 18216
rect 28353 18207 28411 18213
rect 28353 18204 28365 18207
rect 27488 18176 28365 18204
rect 27488 18164 27494 18176
rect 28353 18173 28365 18176
rect 28399 18173 28411 18207
rect 28353 18167 28411 18173
rect 28994 18164 29000 18216
rect 29052 18204 29058 18216
rect 29730 18204 29736 18216
rect 29052 18176 29736 18204
rect 29052 18164 29058 18176
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 37550 18164 37556 18216
rect 37608 18204 37614 18216
rect 37737 18207 37795 18213
rect 37737 18204 37749 18207
rect 37608 18176 37749 18204
rect 37608 18164 37614 18176
rect 37737 18173 37749 18176
rect 37783 18173 37795 18207
rect 37737 18167 37795 18173
rect 37826 18164 37832 18216
rect 37884 18204 37890 18216
rect 38289 18207 38347 18213
rect 38289 18204 38301 18207
rect 37884 18176 38301 18204
rect 37884 18164 37890 18176
rect 38289 18173 38301 18176
rect 38335 18173 38347 18207
rect 38289 18167 38347 18173
rect 27706 18136 27712 18148
rect 27172 18108 27712 18136
rect 27706 18096 27712 18108
rect 27764 18096 27770 18148
rect 21867 18040 23336 18068
rect 21867 18037 21879 18040
rect 21821 18031 21879 18037
rect 28718 18028 28724 18080
rect 28776 18028 28782 18080
rect 30374 18028 30380 18080
rect 30432 18028 30438 18080
rect 30742 18028 30748 18080
rect 30800 18028 30806 18080
rect 34885 18071 34943 18077
rect 34885 18037 34897 18071
rect 34931 18068 34943 18071
rect 36078 18068 36084 18080
rect 34931 18040 36084 18068
rect 34931 18037 34943 18040
rect 34885 18031 34943 18037
rect 36078 18028 36084 18040
rect 36136 18068 36142 18080
rect 36446 18068 36452 18080
rect 36136 18040 36452 18068
rect 36136 18028 36142 18040
rect 36446 18028 36452 18040
rect 36504 18028 36510 18080
rect 36722 18028 36728 18080
rect 36780 18028 36786 18080
rect 37274 18028 37280 18080
rect 37332 18028 37338 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 2958 17824 2964 17876
rect 3016 17824 3022 17876
rect 3326 17824 3332 17876
rect 3384 17864 3390 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3384 17836 3801 17864
rect 3384 17824 3390 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 3789 17827 3847 17833
rect 6638 17824 6644 17876
rect 6696 17864 6702 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 6696 17836 7113 17864
rect 6696 17824 6702 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 7101 17827 7159 17833
rect 15105 17867 15163 17873
rect 15105 17833 15117 17867
rect 15151 17864 15163 17867
rect 15654 17864 15660 17876
rect 15151 17836 15660 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 17405 17867 17463 17873
rect 17405 17833 17417 17867
rect 17451 17864 17463 17867
rect 17770 17864 17776 17876
rect 17451 17836 17776 17864
rect 17451 17833 17463 17836
rect 17405 17827 17463 17833
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 20898 17824 20904 17876
rect 20956 17824 20962 17876
rect 24673 17867 24731 17873
rect 24673 17864 24685 17867
rect 22296 17836 24685 17864
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 7193 17799 7251 17805
rect 7193 17796 7205 17799
rect 6880 17768 7205 17796
rect 6880 17756 6886 17768
rect 7193 17765 7205 17768
rect 7239 17765 7251 17799
rect 7193 17759 7251 17765
rect 10229 17799 10287 17805
rect 10229 17765 10241 17799
rect 10275 17765 10287 17799
rect 17313 17799 17371 17805
rect 10229 17759 10287 17765
rect 12452 17768 15976 17796
rect 3605 17731 3663 17737
rect 3605 17697 3617 17731
rect 3651 17728 3663 17731
rect 3786 17728 3792 17740
rect 3651 17700 3792 17728
rect 3651 17697 3663 17700
rect 3605 17691 3663 17697
rect 3786 17688 3792 17700
rect 3844 17688 3850 17740
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4706 17728 4712 17740
rect 4479 17700 4712 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 6178 17688 6184 17740
rect 6236 17728 6242 17740
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 6236 17700 6469 17728
rect 6236 17688 6242 17700
rect 6457 17697 6469 17700
rect 6503 17697 6515 17731
rect 6457 17691 6515 17697
rect 7834 17688 7840 17740
rect 7892 17688 7898 17740
rect 9585 17731 9643 17737
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 10244 17728 10272 17759
rect 9631 17700 10272 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 10686 17688 10692 17740
rect 10744 17688 10750 17740
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17697 10839 17731
rect 10781 17691 10839 17697
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 10796 17660 10824 17691
rect 10100 17632 10824 17660
rect 12181 17663 12239 17669
rect 10100 17620 10106 17632
rect 12181 17629 12193 17663
rect 12227 17660 12239 17663
rect 12342 17660 12348 17672
rect 12227 17632 12348 17660
rect 12227 17629 12239 17632
rect 12181 17623 12239 17629
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 12452 17669 12480 17768
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 14792 17700 15669 17728
rect 14792 17688 14798 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 4614 17552 4620 17604
rect 4672 17592 4678 17604
rect 4801 17595 4859 17601
rect 4801 17592 4813 17595
rect 4672 17564 4813 17592
rect 4672 17552 4678 17564
rect 4801 17561 4813 17564
rect 4847 17592 4859 17595
rect 12728 17592 12756 17688
rect 15948 17669 15976 17768
rect 17313 17765 17325 17799
rect 17359 17796 17371 17799
rect 18138 17796 18144 17808
rect 17359 17768 18144 17796
rect 17359 17765 17371 17768
rect 17313 17759 17371 17765
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 18049 17731 18107 17737
rect 18049 17697 18061 17731
rect 18095 17728 18107 17731
rect 18095 17700 18736 17728
rect 18095 17697 18107 17700
rect 18049 17691 18107 17697
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16022 17660 16028 17672
rect 15979 17632 16028 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 18064 17660 18092 17691
rect 16132 17632 18092 17660
rect 13633 17595 13691 17601
rect 13633 17592 13645 17595
rect 4847 17564 5304 17592
rect 4847 17561 4859 17564
rect 4801 17555 4859 17561
rect 5276 17536 5304 17564
rect 10612 17564 12434 17592
rect 12728 17564 13645 17592
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 5077 17527 5135 17533
rect 5077 17524 5089 17527
rect 4212 17496 5089 17524
rect 4212 17484 4218 17496
rect 5077 17493 5089 17496
rect 5123 17524 5135 17527
rect 5166 17524 5172 17536
rect 5123 17496 5172 17524
rect 5123 17493 5135 17496
rect 5077 17487 5135 17493
rect 5166 17484 5172 17496
rect 5224 17484 5230 17536
rect 5258 17484 5264 17536
rect 5316 17484 5322 17536
rect 10042 17484 10048 17536
rect 10100 17524 10106 17536
rect 10612 17533 10640 17564
rect 12406 17536 12434 17564
rect 13633 17561 13645 17564
rect 13679 17592 13691 17595
rect 16132 17592 16160 17632
rect 13679 17564 16160 17592
rect 16200 17595 16258 17601
rect 13679 17561 13691 17564
rect 13633 17555 13691 17561
rect 16200 17561 16212 17595
rect 16246 17592 16258 17595
rect 17494 17592 17500 17604
rect 16246 17564 17500 17592
rect 16246 17561 16258 17564
rect 16200 17555 16258 17561
rect 17494 17552 17500 17564
rect 17552 17552 17558 17604
rect 17773 17595 17831 17601
rect 17773 17561 17785 17595
rect 17819 17592 17831 17595
rect 18598 17592 18604 17604
rect 17819 17564 18604 17592
rect 17819 17561 17831 17564
rect 17773 17555 17831 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 10137 17527 10195 17533
rect 10137 17524 10149 17527
rect 10100 17496 10149 17524
rect 10100 17484 10106 17496
rect 10137 17493 10149 17496
rect 10183 17493 10195 17527
rect 10137 17487 10195 17493
rect 10597 17527 10655 17533
rect 10597 17493 10609 17527
rect 10643 17493 10655 17527
rect 10597 17487 10655 17493
rect 11054 17484 11060 17536
rect 11112 17484 11118 17536
rect 12406 17496 12440 17536
rect 12434 17484 12440 17496
rect 12492 17524 12498 17536
rect 12805 17527 12863 17533
rect 12805 17524 12817 17527
rect 12492 17496 12817 17524
rect 12492 17484 12498 17496
rect 12805 17493 12817 17496
rect 12851 17493 12863 17527
rect 12805 17487 12863 17493
rect 12894 17484 12900 17536
rect 12952 17484 12958 17536
rect 13262 17484 13268 17536
rect 13320 17484 13326 17536
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 14792 17496 14933 17524
rect 14792 17484 14798 17496
rect 14921 17493 14933 17496
rect 14967 17493 14979 17527
rect 14921 17487 14979 17493
rect 15470 17484 15476 17536
rect 15528 17484 15534 17536
rect 15565 17527 15623 17533
rect 15565 17493 15577 17527
rect 15611 17524 15623 17527
rect 16574 17524 16580 17536
rect 15611 17496 16580 17524
rect 15611 17493 15623 17496
rect 15565 17487 15623 17493
rect 16574 17484 16580 17496
rect 16632 17524 16638 17536
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 16632 17496 17877 17524
rect 16632 17484 16638 17496
rect 17865 17493 17877 17496
rect 17911 17493 17923 17527
rect 17865 17487 17923 17493
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 18708 17524 18736 17700
rect 20916 17660 20944 17824
rect 22097 17731 22155 17737
rect 22097 17697 22109 17731
rect 22143 17728 22155 17731
rect 22296 17728 22324 17836
rect 24673 17833 24685 17836
rect 24719 17864 24731 17867
rect 24946 17864 24952 17876
rect 24719 17836 24952 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 24946 17824 24952 17836
rect 25004 17824 25010 17876
rect 26326 17824 26332 17876
rect 26384 17824 26390 17876
rect 26786 17824 26792 17876
rect 26844 17864 26850 17876
rect 26844 17836 37320 17864
rect 26844 17824 26850 17836
rect 34701 17799 34759 17805
rect 34701 17796 34713 17799
rect 22388 17768 24348 17796
rect 22388 17737 22416 17768
rect 24320 17740 24348 17768
rect 34532 17768 34713 17796
rect 22143 17700 22324 17728
rect 22373 17731 22431 17737
rect 22143 17697 22155 17700
rect 22097 17691 22155 17697
rect 22373 17697 22385 17731
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22557 17731 22615 17737
rect 22557 17728 22569 17731
rect 22520 17700 22569 17728
rect 22520 17688 22526 17700
rect 22557 17697 22569 17700
rect 22603 17697 22615 17731
rect 22557 17691 22615 17697
rect 23477 17731 23535 17737
rect 23477 17697 23489 17731
rect 23523 17728 23535 17731
rect 23658 17728 23664 17740
rect 23523 17700 23664 17728
rect 23523 17697 23535 17700
rect 23477 17691 23535 17697
rect 23658 17688 23664 17700
rect 23716 17688 23722 17740
rect 24302 17688 24308 17740
rect 24360 17688 24366 17740
rect 26878 17688 26884 17740
rect 26936 17688 26942 17740
rect 27341 17731 27399 17737
rect 27341 17697 27353 17731
rect 27387 17728 27399 17731
rect 28166 17728 28172 17740
rect 27387 17700 28172 17728
rect 27387 17697 27399 17700
rect 27341 17691 27399 17697
rect 28166 17688 28172 17700
rect 28224 17688 28230 17740
rect 34532 17737 34560 17768
rect 34701 17765 34713 17768
rect 34747 17765 34759 17799
rect 36357 17799 36415 17805
rect 36357 17796 36369 17799
rect 34701 17759 34759 17765
rect 35176 17768 36369 17796
rect 34517 17731 34575 17737
rect 34517 17697 34529 17731
rect 34563 17697 34575 17731
rect 35176 17728 35204 17768
rect 36357 17765 36369 17768
rect 36403 17765 36415 17799
rect 37292 17796 37320 17836
rect 37366 17824 37372 17876
rect 37424 17824 37430 17876
rect 37826 17796 37832 17808
rect 37292 17768 37832 17796
rect 36357 17759 36415 17765
rect 37826 17756 37832 17768
rect 37884 17756 37890 17808
rect 34517 17691 34575 17697
rect 35084 17700 35204 17728
rect 20916 17632 25360 17660
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19613 17595 19671 17601
rect 19613 17592 19625 17595
rect 19484 17564 19625 17592
rect 19484 17552 19490 17564
rect 19613 17561 19625 17564
rect 19659 17561 19671 17595
rect 19613 17555 19671 17561
rect 21358 17552 21364 17604
rect 21416 17592 21422 17604
rect 21416 17564 22048 17592
rect 21416 17552 21422 17564
rect 18966 17524 18972 17536
rect 18555 17496 18972 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 21450 17484 21456 17536
rect 21508 17484 21514 17536
rect 21836 17533 21864 17564
rect 22020 17536 22048 17564
rect 22646 17552 22652 17604
rect 22704 17552 22710 17604
rect 24213 17595 24271 17601
rect 24213 17561 24225 17595
rect 24259 17592 24271 17595
rect 24486 17592 24492 17604
rect 24259 17564 24492 17592
rect 24259 17561 24271 17564
rect 24213 17555 24271 17561
rect 24486 17552 24492 17564
rect 24544 17592 24550 17604
rect 24949 17595 25007 17601
rect 24949 17592 24961 17595
rect 24544 17564 24961 17592
rect 24544 17552 24550 17564
rect 24949 17561 24961 17564
rect 24995 17561 25007 17595
rect 25332 17592 25360 17632
rect 25682 17620 25688 17672
rect 25740 17660 25746 17672
rect 27706 17660 27712 17672
rect 25740 17632 27712 17660
rect 25740 17620 25746 17632
rect 27706 17620 27712 17632
rect 27764 17660 27770 17672
rect 27985 17663 28043 17669
rect 27985 17660 27997 17663
rect 27764 17632 27997 17660
rect 27764 17620 27770 17632
rect 27985 17629 27997 17632
rect 28031 17660 28043 17663
rect 28258 17660 28264 17672
rect 28031 17632 28264 17660
rect 28031 17629 28043 17632
rect 27985 17623 28043 17629
rect 28258 17620 28264 17632
rect 28316 17620 28322 17672
rect 28626 17620 28632 17672
rect 28684 17620 28690 17672
rect 35084 17669 35112 17700
rect 35250 17688 35256 17740
rect 35308 17688 35314 17740
rect 35342 17688 35348 17740
rect 35400 17688 35406 17740
rect 35621 17731 35679 17737
rect 35621 17728 35633 17731
rect 35452 17700 35633 17728
rect 35069 17663 35127 17669
rect 35069 17629 35081 17663
rect 35115 17629 35127 17663
rect 35268 17660 35296 17688
rect 35452 17660 35480 17700
rect 35621 17697 35633 17700
rect 35667 17728 35679 17731
rect 36538 17728 36544 17740
rect 35667 17700 36544 17728
rect 35667 17697 35679 17700
rect 35621 17691 35679 17697
rect 36538 17688 36544 17700
rect 36596 17688 36602 17740
rect 37274 17688 37280 17740
rect 37332 17728 37338 17740
rect 37921 17731 37979 17737
rect 37921 17728 37933 17731
rect 37332 17700 37933 17728
rect 37332 17688 37338 17700
rect 37921 17697 37933 17700
rect 37967 17697 37979 17731
rect 37921 17691 37979 17697
rect 35268 17632 35480 17660
rect 35069 17623 35127 17629
rect 36170 17620 36176 17672
rect 36228 17660 36234 17672
rect 36446 17660 36452 17672
rect 36228 17632 36452 17660
rect 36228 17620 36234 17632
rect 36446 17620 36452 17632
rect 36504 17620 36510 17672
rect 36906 17620 36912 17672
rect 36964 17620 36970 17672
rect 28644 17592 28672 17620
rect 34974 17592 34980 17604
rect 25332 17564 28672 17592
rect 33336 17564 34980 17592
rect 24949 17555 25007 17561
rect 21821 17527 21879 17533
rect 21821 17493 21833 17527
rect 21867 17493 21879 17527
rect 21821 17487 21879 17493
rect 21910 17484 21916 17536
rect 21968 17484 21974 17536
rect 22002 17484 22008 17536
rect 22060 17484 22066 17536
rect 22738 17484 22744 17536
rect 22796 17524 22802 17536
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22796 17496 23029 17524
rect 22796 17484 22802 17496
rect 23017 17493 23029 17496
rect 23063 17493 23075 17527
rect 24964 17524 24992 17555
rect 33336 17536 33364 17564
rect 34974 17552 34980 17564
rect 35032 17552 35038 17604
rect 35805 17595 35863 17601
rect 35805 17561 35817 17595
rect 35851 17592 35863 17595
rect 36078 17592 36084 17604
rect 35851 17564 36084 17592
rect 35851 17561 35863 17564
rect 35805 17555 35863 17561
rect 36078 17552 36084 17564
rect 36136 17552 36142 17604
rect 36188 17564 36400 17592
rect 28994 17524 29000 17536
rect 24964 17496 29000 17524
rect 23017 17487 23075 17493
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 29178 17484 29184 17536
rect 29236 17524 29242 17536
rect 29730 17524 29736 17536
rect 29236 17496 29736 17524
rect 29236 17484 29242 17496
rect 29730 17484 29736 17496
rect 29788 17484 29794 17536
rect 33318 17484 33324 17536
rect 33376 17484 33382 17536
rect 33778 17484 33784 17536
rect 33836 17484 33842 17536
rect 33870 17484 33876 17536
rect 33928 17484 33934 17536
rect 34698 17484 34704 17536
rect 34756 17524 34762 17536
rect 35161 17527 35219 17533
rect 35161 17524 35173 17527
rect 34756 17496 35173 17524
rect 34756 17484 34762 17496
rect 35161 17493 35173 17496
rect 35207 17524 35219 17527
rect 35897 17527 35955 17533
rect 35897 17524 35909 17527
rect 35207 17496 35909 17524
rect 35207 17493 35219 17496
rect 35161 17487 35219 17493
rect 35897 17493 35909 17496
rect 35943 17524 35955 17527
rect 36188 17524 36216 17564
rect 35943 17496 36216 17524
rect 35943 17493 35955 17496
rect 35897 17487 35955 17493
rect 36262 17484 36268 17536
rect 36320 17484 36326 17536
rect 36372 17524 36400 17564
rect 37550 17524 37556 17536
rect 36372 17496 37556 17524
rect 37550 17484 37556 17496
rect 37608 17484 37614 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 4893 17323 4951 17329
rect 4893 17289 4905 17323
rect 4939 17320 4951 17323
rect 4982 17320 4988 17332
rect 4939 17292 4988 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 26786 17320 26792 17332
rect 6748 17292 26792 17320
rect 4614 17212 4620 17264
rect 4672 17252 4678 17264
rect 6748 17252 6776 17292
rect 26786 17280 26792 17292
rect 26844 17280 26850 17332
rect 28994 17280 29000 17332
rect 29052 17280 29058 17332
rect 29086 17280 29092 17332
rect 29144 17320 29150 17332
rect 29181 17323 29239 17329
rect 29181 17320 29193 17323
rect 29144 17292 29193 17320
rect 29144 17280 29150 17292
rect 29181 17289 29193 17292
rect 29227 17289 29239 17323
rect 29181 17283 29239 17289
rect 33870 17280 33876 17332
rect 33928 17280 33934 17332
rect 34701 17323 34759 17329
rect 34701 17289 34713 17323
rect 34747 17320 34759 17323
rect 36078 17320 36084 17332
rect 34747 17292 36084 17320
rect 34747 17289 34759 17292
rect 34701 17283 34759 17289
rect 36078 17280 36084 17292
rect 36136 17320 36142 17332
rect 36906 17320 36912 17332
rect 36136 17292 36912 17320
rect 36136 17280 36142 17292
rect 36906 17280 36912 17292
rect 36964 17280 36970 17332
rect 37642 17280 37648 17332
rect 37700 17280 37706 17332
rect 4672 17224 6776 17252
rect 4672 17212 4678 17224
rect 7834 17212 7840 17264
rect 7892 17252 7898 17264
rect 9493 17255 9551 17261
rect 9493 17252 9505 17255
rect 7892 17224 9505 17252
rect 7892 17212 7898 17224
rect 9493 17221 9505 17224
rect 9539 17252 9551 17255
rect 9539 17224 11008 17252
rect 9539 17221 9551 17224
rect 9493 17215 9551 17221
rect 4798 17144 4804 17196
rect 4856 17144 4862 17196
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10209 17187 10267 17193
rect 10209 17184 10221 17187
rect 10100 17156 10221 17184
rect 10100 17144 10106 17156
rect 10209 17153 10221 17156
rect 10255 17153 10267 17187
rect 10209 17147 10267 17153
rect 3418 17076 3424 17128
rect 3476 17076 3482 17128
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17116 4215 17119
rect 4706 17116 4712 17128
rect 4203 17088 4712 17116
rect 4203 17085 4215 17088
rect 4157 17079 4215 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17116 6239 17119
rect 7006 17116 7012 17128
rect 6227 17088 7012 17116
rect 6227 17085 6239 17088
rect 6181 17079 6239 17085
rect 7006 17076 7012 17088
rect 7064 17076 7070 17128
rect 7558 17076 7564 17128
rect 7616 17076 7622 17128
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 8386 17116 8392 17128
rect 8343 17088 8392 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 9953 17119 10011 17125
rect 9953 17085 9965 17119
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 6687 17020 8340 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 2774 16940 2780 16992
rect 2832 16940 2838 16992
rect 3142 16940 3148 16992
rect 3200 16980 3206 16992
rect 3513 16983 3571 16989
rect 3513 16980 3525 16983
rect 3200 16952 3525 16980
rect 3200 16940 3206 16952
rect 3513 16949 3525 16952
rect 3559 16949 3571 16983
rect 3513 16943 3571 16949
rect 5258 16940 5264 16992
rect 5316 16940 5322 16992
rect 5534 16940 5540 16992
rect 5592 16940 5598 16992
rect 6914 16940 6920 16992
rect 6972 16940 6978 16992
rect 7650 16940 7656 16992
rect 7708 16940 7714 16992
rect 8312 16980 8340 17020
rect 8478 17008 8484 17060
rect 8536 17048 8542 17060
rect 8662 17048 8668 17060
rect 8536 17020 8668 17048
rect 8536 17008 8542 17020
rect 8662 17008 8668 17020
rect 8720 17048 8726 17060
rect 9858 17048 9864 17060
rect 8720 17020 9864 17048
rect 8720 17008 8726 17020
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 9968 16992 9996 17079
rect 10980 17060 11008 17224
rect 13262 17212 13268 17264
rect 13320 17212 13326 17264
rect 15013 17255 15071 17261
rect 15013 17221 15025 17255
rect 15059 17252 15071 17255
rect 15470 17252 15476 17264
rect 15059 17224 15476 17252
rect 15059 17221 15071 17224
rect 15013 17215 15071 17221
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 18598 17212 18604 17264
rect 18656 17212 18662 17264
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 20901 17255 20959 17261
rect 20901 17252 20913 17255
rect 20772 17224 20913 17252
rect 20772 17212 20778 17224
rect 20901 17221 20913 17224
rect 20947 17221 20959 17255
rect 20901 17215 20959 17221
rect 21450 17212 21456 17264
rect 21508 17212 21514 17264
rect 21821 17255 21879 17261
rect 21821 17221 21833 17255
rect 21867 17252 21879 17255
rect 21910 17252 21916 17264
rect 21867 17224 21916 17252
rect 21867 17221 21879 17224
rect 21821 17215 21879 17221
rect 21910 17212 21916 17224
rect 21968 17212 21974 17264
rect 29012 17252 29040 17280
rect 33042 17252 33048 17264
rect 29012 17224 33048 17252
rect 33042 17212 33048 17224
rect 33100 17252 33106 17264
rect 33137 17255 33195 17261
rect 33137 17252 33149 17255
rect 33100 17224 33149 17252
rect 33100 17212 33106 17224
rect 33137 17221 33149 17224
rect 33183 17221 33195 17255
rect 33137 17215 33195 17221
rect 33588 17255 33646 17261
rect 33588 17221 33600 17255
rect 33634 17252 33646 17255
rect 33888 17252 33916 17280
rect 35250 17252 35256 17264
rect 33634 17224 33916 17252
rect 35084 17224 35256 17252
rect 33634 17221 33646 17224
rect 33588 17215 33646 17221
rect 13280 17184 13308 17212
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13280 17156 14013 17184
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 15194 17184 15200 17196
rect 14507 17156 15200 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15378 17193 15384 17196
rect 15372 17147 15384 17193
rect 15378 17144 15384 17147
rect 15436 17144 15442 17196
rect 17301 17144 17307 17196
rect 17359 17144 17365 17196
rect 18138 17144 18144 17196
rect 18196 17144 18202 17196
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 19153 17187 19211 17193
rect 19153 17184 19165 17187
rect 18380 17156 19165 17184
rect 18380 17144 18386 17156
rect 19153 17153 19165 17156
rect 19199 17153 19211 17187
rect 21468 17184 21496 17212
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 21468 17156 21557 17184
rect 19153 17147 19211 17153
rect 21545 17153 21557 17156
rect 21591 17153 21603 17187
rect 21545 17147 21603 17153
rect 22370 17144 22376 17196
rect 22428 17144 22434 17196
rect 29273 17187 29331 17193
rect 29273 17153 29285 17187
rect 29319 17184 29331 17187
rect 29914 17184 29920 17196
rect 29319 17156 29920 17184
rect 29319 17153 29331 17156
rect 29273 17147 29331 17153
rect 29914 17144 29920 17156
rect 29972 17144 29978 17196
rect 35084 17193 35112 17224
rect 35250 17212 35256 17224
rect 35308 17212 35314 17264
rect 35069 17187 35127 17193
rect 35069 17153 35081 17187
rect 35115 17153 35127 17187
rect 35069 17147 35127 17153
rect 36078 17144 36084 17196
rect 36136 17193 36142 17196
rect 36136 17187 36164 17193
rect 36152 17153 36164 17187
rect 36136 17147 36164 17153
rect 36909 17187 36967 17193
rect 36909 17153 36921 17187
rect 36955 17184 36967 17187
rect 37553 17187 37611 17193
rect 37553 17184 37565 17187
rect 36955 17156 37565 17184
rect 36955 17153 36967 17156
rect 36909 17147 36967 17153
rect 37553 17153 37565 17156
rect 37599 17153 37611 17187
rect 37553 17147 37611 17153
rect 36136 17144 36142 17147
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11112 17088 11529 17116
rect 11112 17076 11118 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11698 17076 11704 17128
rect 11756 17076 11762 17128
rect 12618 17125 12624 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12268 17088 12449 17116
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 12161 17051 12219 17057
rect 12161 17048 12173 17051
rect 11020 17020 12173 17048
rect 11020 17008 11026 17020
rect 12161 17017 12173 17020
rect 12207 17017 12219 17051
rect 12161 17011 12219 17017
rect 9306 16980 9312 16992
rect 8312 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16980 9370 16992
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 9364 16952 9781 16980
rect 9364 16940 9370 16952
rect 9769 16949 9781 16952
rect 9815 16949 9827 16983
rect 9769 16943 9827 16949
rect 9950 16940 9956 16992
rect 10008 16940 10014 16992
rect 11330 16940 11336 16992
rect 11388 16980 11394 16992
rect 12268 16980 12296 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12575 17119 12624 17125
rect 12575 17085 12587 17119
rect 12621 17085 12624 17119
rect 12575 17079 12624 17085
rect 12618 17076 12624 17079
rect 12676 17076 12682 17128
rect 12713 17119 12771 17125
rect 12713 17085 12725 17119
rect 12759 17116 12771 17119
rect 13078 17116 13084 17128
rect 12759 17088 13084 17116
rect 12759 17085 12771 17088
rect 12713 17079 12771 17085
rect 13078 17076 13084 17088
rect 13136 17116 13142 17128
rect 13136 17088 14228 17116
rect 13136 17076 13142 17088
rect 13262 17008 13268 17060
rect 13320 17048 13326 17060
rect 13449 17051 13507 17057
rect 13449 17048 13461 17051
rect 13320 17020 13461 17048
rect 13320 17008 13326 17020
rect 13449 17017 13461 17020
rect 13495 17017 13507 17051
rect 13449 17011 13507 17017
rect 11388 16952 12296 16980
rect 11388 16940 11394 16952
rect 13354 16940 13360 16992
rect 13412 16940 13418 16992
rect 14200 16980 14228 17088
rect 15102 17076 15108 17128
rect 15160 17076 15166 17128
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 17451 17119 17509 17125
rect 17451 17116 17463 17119
rect 16264 17088 17463 17116
rect 16264 17076 16270 17088
rect 17451 17085 17463 17088
rect 17497 17085 17509 17119
rect 17451 17079 17509 17085
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17116 17647 17119
rect 18156 17116 18184 17144
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 17635 17088 17816 17116
rect 18156 17088 18521 17116
rect 17635 17085 17647 17088
rect 17589 17079 17647 17085
rect 16482 17008 16488 17060
rect 16540 17048 16546 17060
rect 16540 17020 16988 17048
rect 16540 17008 16546 17020
rect 16298 16980 16304 16992
rect 14200 16952 16304 16980
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 16960 16980 16988 17020
rect 17788 16980 17816 17088
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 23201 17119 23259 17125
rect 23201 17085 23213 17119
rect 23247 17116 23259 17119
rect 23382 17116 23388 17128
rect 23247 17088 23388 17116
rect 23247 17085 23259 17088
rect 23201 17079 23259 17085
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 23842 17076 23848 17128
rect 23900 17076 23906 17128
rect 26510 17076 26516 17128
rect 26568 17116 26574 17128
rect 26789 17119 26847 17125
rect 26789 17116 26801 17119
rect 26568 17088 26801 17116
rect 26568 17076 26574 17088
rect 26789 17085 26801 17088
rect 26835 17116 26847 17119
rect 27430 17116 27436 17128
rect 26835 17088 27436 17116
rect 26835 17085 26847 17088
rect 26789 17079 26847 17085
rect 27430 17076 27436 17088
rect 27488 17076 27494 17128
rect 27614 17076 27620 17128
rect 27672 17076 27678 17128
rect 27890 17076 27896 17128
rect 27948 17116 27954 17128
rect 28261 17119 28319 17125
rect 28261 17116 28273 17119
rect 27948 17088 28273 17116
rect 27948 17076 27954 17088
rect 28261 17085 28273 17088
rect 28307 17085 28319 17119
rect 28261 17079 28319 17085
rect 33134 17076 33140 17128
rect 33192 17116 33198 17128
rect 33321 17119 33379 17125
rect 33321 17116 33333 17119
rect 33192 17088 33333 17116
rect 33192 17076 33198 17088
rect 33321 17085 33333 17088
rect 33367 17085 33379 17119
rect 33321 17079 33379 17085
rect 35253 17119 35311 17125
rect 35253 17085 35265 17119
rect 35299 17116 35311 17119
rect 35434 17116 35440 17128
rect 35299 17088 35440 17116
rect 35299 17085 35311 17088
rect 35253 17079 35311 17085
rect 35434 17076 35440 17088
rect 35492 17076 35498 17128
rect 35618 17076 35624 17128
rect 35676 17116 35682 17128
rect 35989 17119 36047 17125
rect 35989 17116 36001 17119
rect 35676 17088 36001 17116
rect 35676 17076 35682 17088
rect 35989 17085 36001 17088
rect 36035 17085 36047 17119
rect 35989 17079 36047 17085
rect 36265 17119 36323 17125
rect 36265 17085 36277 17119
rect 36311 17116 36323 17119
rect 36446 17116 36452 17128
rect 36311 17088 36452 17116
rect 36311 17085 36323 17088
rect 36265 17079 36323 17085
rect 36446 17076 36452 17088
rect 36504 17076 36510 17128
rect 37461 17119 37519 17125
rect 37461 17085 37473 17119
rect 37507 17116 37519 17119
rect 38102 17116 38108 17128
rect 37507 17088 38108 17116
rect 37507 17085 37519 17088
rect 37461 17079 37519 17085
rect 38102 17076 38108 17088
rect 38160 17116 38166 17128
rect 38289 17119 38347 17125
rect 38289 17116 38301 17119
rect 38160 17088 38301 17116
rect 38160 17076 38166 17088
rect 38289 17085 38301 17088
rect 38335 17085 38347 17119
rect 38289 17079 38347 17085
rect 17862 17008 17868 17060
rect 17920 17008 17926 17060
rect 24578 17008 24584 17060
rect 24636 17048 24642 17060
rect 32769 17051 32827 17057
rect 32769 17048 32781 17051
rect 24636 17020 32781 17048
rect 24636 17008 24642 17020
rect 32769 17017 32781 17020
rect 32815 17017 32827 17051
rect 32769 17011 32827 17017
rect 35713 17051 35771 17057
rect 35713 17017 35725 17051
rect 35759 17017 35771 17051
rect 35713 17011 35771 17017
rect 16960 16952 17816 16980
rect 22554 16940 22560 16992
rect 22612 16940 22618 16992
rect 23290 16940 23296 16992
rect 23348 16940 23354 16992
rect 24302 16940 24308 16992
rect 24360 16980 24366 16992
rect 25498 16980 25504 16992
rect 24360 16952 25504 16980
rect 24360 16940 24366 16952
rect 25498 16940 25504 16952
rect 25556 16940 25562 16992
rect 26234 16940 26240 16992
rect 26292 16980 26298 16992
rect 26329 16983 26387 16989
rect 26329 16980 26341 16983
rect 26292 16952 26341 16980
rect 26292 16940 26298 16952
rect 26329 16949 26341 16952
rect 26375 16949 26387 16983
rect 26329 16943 26387 16949
rect 26786 16940 26792 16992
rect 26844 16980 26850 16992
rect 26973 16983 27031 16989
rect 26973 16980 26985 16983
rect 26844 16952 26985 16980
rect 26844 16940 26850 16952
rect 26973 16949 26985 16952
rect 27019 16949 27031 16983
rect 26973 16943 27031 16949
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 27709 16983 27767 16989
rect 27709 16980 27721 16983
rect 27120 16952 27721 16980
rect 27120 16940 27126 16952
rect 27709 16949 27721 16952
rect 27755 16949 27767 16983
rect 27709 16943 27767 16949
rect 30377 16983 30435 16989
rect 30377 16949 30389 16983
rect 30423 16980 30435 16983
rect 30926 16980 30932 16992
rect 30423 16952 30932 16980
rect 30423 16949 30435 16952
rect 30377 16943 30435 16949
rect 30926 16940 30932 16952
rect 30984 16940 30990 16992
rect 32784 16980 32812 17011
rect 35728 16980 35756 17011
rect 36722 16980 36728 16992
rect 32784 16952 36728 16980
rect 36722 16940 36728 16952
rect 36780 16940 36786 16992
rect 38013 16983 38071 16989
rect 38013 16949 38025 16983
rect 38059 16980 38071 16983
rect 38194 16980 38200 16992
rect 38059 16952 38200 16980
rect 38059 16949 38071 16952
rect 38013 16943 38071 16949
rect 38194 16940 38200 16952
rect 38252 16940 38258 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 3142 16736 3148 16788
rect 3200 16736 3206 16788
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 3605 16779 3663 16785
rect 3605 16776 3617 16779
rect 3476 16748 3617 16776
rect 3476 16736 3482 16748
rect 3605 16745 3617 16748
rect 3651 16745 3663 16779
rect 3605 16739 3663 16745
rect 7006 16736 7012 16788
rect 7064 16736 7070 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7616 16748 7849 16776
rect 7616 16736 7622 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 12434 16776 12440 16788
rect 10008 16748 12440 16776
rect 10008 16736 10014 16748
rect 12434 16736 12440 16748
rect 12492 16776 12498 16788
rect 12492 16748 12848 16776
rect 12492 16736 12498 16748
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2958 16640 2964 16652
rect 2087 16612 2964 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3160 16649 3188 16736
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16609 3203 16643
rect 3145 16603 3203 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4522 16640 4528 16652
rect 4479 16612 4528 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 7098 16600 7104 16652
rect 7156 16640 7162 16652
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 7156 16612 7297 16640
rect 7156 16600 7162 16612
rect 7285 16609 7297 16612
rect 7331 16640 7343 16643
rect 8662 16640 8668 16652
rect 7331 16612 8668 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9968 16649 9996 16736
rect 11425 16711 11483 16717
rect 11425 16677 11437 16711
rect 11471 16677 11483 16711
rect 11425 16671 11483 16677
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 2130 16532 2136 16584
rect 2188 16532 2194 16584
rect 2976 16572 3004 16600
rect 3878 16572 3884 16584
rect 2976 16544 3884 16572
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 6178 16572 6184 16584
rect 5675 16544 6184 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 8478 16532 8484 16584
rect 8536 16532 8542 16584
rect 10220 16575 10278 16581
rect 10220 16541 10232 16575
rect 10266 16572 10278 16575
rect 10502 16572 10508 16584
rect 10266 16544 10508 16572
rect 10266 16541 10278 16544
rect 10220 16535 10278 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11440 16572 11468 16671
rect 12820 16649 12848 16748
rect 12894 16736 12900 16788
rect 12952 16736 12958 16788
rect 15102 16776 15108 16788
rect 14844 16748 15108 16776
rect 14844 16649 14872 16748
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 15194 16736 15200 16788
rect 15252 16776 15258 16788
rect 16206 16776 16212 16788
rect 15252 16748 16212 16776
rect 15252 16736 15258 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16577 16779 16635 16785
rect 16577 16776 16589 16779
rect 16356 16748 16589 16776
rect 16356 16736 16362 16748
rect 16577 16745 16589 16748
rect 16623 16776 16635 16779
rect 17310 16776 17316 16788
rect 16623 16748 17316 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 18049 16779 18107 16785
rect 18049 16745 18061 16779
rect 18095 16776 18107 16779
rect 18322 16776 18328 16788
rect 18095 16748 18328 16776
rect 18095 16745 18107 16748
rect 18049 16739 18107 16745
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 20162 16736 20168 16788
rect 20220 16776 20226 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 20220 16748 21189 16776
rect 20220 16736 20226 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 21177 16739 21235 16745
rect 23109 16779 23167 16785
rect 23109 16745 23121 16779
rect 23155 16776 23167 16779
rect 23842 16776 23848 16788
rect 23155 16748 23848 16776
rect 23155 16745 23167 16748
rect 23109 16739 23167 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 24673 16779 24731 16785
rect 24673 16745 24685 16779
rect 24719 16776 24731 16779
rect 24946 16776 24952 16788
rect 24719 16748 24952 16776
rect 24719 16745 24731 16748
rect 24673 16739 24731 16745
rect 22480 16680 24072 16708
rect 12805 16643 12863 16649
rect 12805 16609 12817 16643
rect 12851 16640 12863 16643
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 12851 16612 14841 16640
rect 12851 16609 12863 16612
rect 12805 16603 12863 16609
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 22480 16649 22508 16680
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16080 16612 16681 16640
rect 16080 16600 16086 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 24044 16649 24072 16680
rect 22649 16643 22707 16649
rect 22649 16640 22661 16643
rect 22612 16612 22661 16640
rect 22612 16600 22618 16612
rect 22649 16609 22661 16612
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 24029 16643 24087 16649
rect 24029 16609 24041 16643
rect 24075 16640 24087 16643
rect 24688 16640 24716 16739
rect 24946 16736 24952 16748
rect 25004 16736 25010 16788
rect 25961 16779 26019 16785
rect 25961 16745 25973 16779
rect 26007 16776 26019 16779
rect 26418 16776 26424 16788
rect 26007 16748 26424 16776
rect 26007 16745 26019 16748
rect 25961 16739 26019 16745
rect 24075 16612 26004 16640
rect 24075 16609 24087 16612
rect 24029 16603 24087 16609
rect 11698 16572 11704 16584
rect 11440 16544 11704 16572
rect 11698 16532 11704 16544
rect 11756 16572 11762 16584
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 11756 16544 13461 16572
rect 11756 16532 11762 16544
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 13630 16532 13636 16584
rect 13688 16532 13694 16584
rect 15102 16581 15108 16584
rect 15096 16535 15108 16581
rect 15160 16572 15166 16584
rect 16936 16575 16994 16581
rect 15160 16544 15196 16572
rect 15102 16532 15108 16535
rect 15160 16532 15166 16544
rect 16936 16541 16948 16575
rect 16982 16572 16994 16575
rect 17218 16572 17224 16584
rect 16982 16544 17224 16572
rect 16982 16541 16994 16544
rect 16936 16535 16994 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 18141 16575 18199 16581
rect 18141 16572 18153 16575
rect 17552 16544 18153 16572
rect 17552 16532 17558 16544
rect 18141 16541 18153 16544
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 18690 16532 18696 16584
rect 18748 16532 18754 16584
rect 22281 16575 22339 16581
rect 22281 16572 22293 16575
rect 18800 16544 22293 16572
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 3237 16507 3295 16513
rect 3237 16504 3249 16507
rect 2464 16476 3249 16504
rect 2464 16464 2470 16476
rect 3237 16473 3249 16476
rect 3283 16504 3295 16507
rect 4157 16507 4215 16513
rect 3283 16476 4108 16504
rect 3283 16473 3295 16476
rect 3237 16467 3295 16473
rect 2590 16396 2596 16448
rect 2648 16436 2654 16448
rect 2777 16439 2835 16445
rect 2777 16436 2789 16439
rect 2648 16408 2789 16436
rect 2648 16396 2654 16408
rect 2777 16405 2789 16408
rect 2823 16405 2835 16439
rect 2777 16399 2835 16405
rect 3786 16396 3792 16448
rect 3844 16396 3850 16448
rect 4080 16436 4108 16476
rect 4157 16473 4169 16507
rect 4203 16504 4215 16507
rect 4798 16504 4804 16516
rect 4203 16476 4804 16504
rect 4203 16473 4215 16476
rect 4157 16467 4215 16473
rect 4798 16464 4804 16476
rect 4856 16464 4862 16516
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16504 5595 16507
rect 5874 16507 5932 16513
rect 5874 16504 5886 16507
rect 5583 16476 5886 16504
rect 5583 16473 5595 16476
rect 5537 16467 5595 16473
rect 5874 16473 5886 16476
rect 5920 16473 5932 16507
rect 5874 16467 5932 16473
rect 7377 16507 7435 16513
rect 7377 16473 7389 16507
rect 7423 16504 7435 16507
rect 7929 16507 7987 16513
rect 7929 16504 7941 16507
rect 7423 16476 7941 16504
rect 7423 16473 7435 16476
rect 7377 16467 7435 16473
rect 7929 16473 7941 16476
rect 7975 16473 7987 16507
rect 12560 16507 12618 16513
rect 7929 16467 7987 16473
rect 11348 16476 12434 16504
rect 4249 16439 4307 16445
rect 4249 16436 4261 16439
rect 4080 16408 4261 16436
rect 4249 16405 4261 16408
rect 4295 16436 4307 16439
rect 5442 16436 5448 16448
rect 4295 16408 5448 16436
rect 4295 16405 4307 16408
rect 4249 16399 4307 16405
rect 5442 16396 5448 16408
rect 5500 16436 5506 16448
rect 7469 16439 7527 16445
rect 7469 16436 7481 16439
rect 5500 16408 7481 16436
rect 5500 16396 5506 16408
rect 7469 16405 7481 16408
rect 7515 16436 7527 16439
rect 7742 16436 7748 16448
rect 7515 16408 7748 16436
rect 7515 16405 7527 16408
rect 7469 16399 7527 16405
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 11348 16445 11376 16476
rect 11333 16439 11391 16445
rect 11333 16405 11345 16439
rect 11379 16405 11391 16439
rect 12406 16436 12434 16476
rect 12560 16473 12572 16507
rect 12606 16504 12618 16507
rect 13262 16504 13268 16516
rect 12606 16476 13268 16504
rect 12606 16473 12618 16476
rect 12560 16467 12618 16473
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 12710 16436 12716 16448
rect 12406 16408 12716 16436
rect 11333 16399 11391 16405
rect 12710 16396 12716 16408
rect 12768 16436 12774 16448
rect 13648 16436 13676 16532
rect 17586 16464 17592 16516
rect 17644 16504 17650 16516
rect 18800 16504 18828 16544
rect 22281 16541 22293 16544
rect 22327 16572 22339 16575
rect 23201 16575 23259 16581
rect 23201 16572 23213 16575
rect 22327 16544 23213 16572
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 23201 16541 23213 16544
rect 23247 16541 23259 16575
rect 23201 16535 23259 16541
rect 25038 16532 25044 16584
rect 25096 16532 25102 16584
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 17644 16476 18828 16504
rect 17644 16464 17650 16476
rect 21266 16464 21272 16516
rect 21324 16464 21330 16516
rect 12768 16408 13676 16436
rect 22741 16439 22799 16445
rect 12768 16396 12774 16408
rect 22741 16405 22753 16439
rect 22787 16436 22799 16439
rect 23566 16436 23572 16448
rect 22787 16408 23572 16436
rect 22787 16405 22799 16408
rect 22741 16399 22799 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 25056 16436 25084 16532
rect 25976 16504 26004 16612
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 26160 16649 26188 16748
rect 26418 16736 26424 16748
rect 26476 16736 26482 16788
rect 26789 16779 26847 16785
rect 26789 16745 26801 16779
rect 26835 16776 26847 16779
rect 26835 16748 30144 16776
rect 26835 16745 26847 16748
rect 26789 16739 26847 16745
rect 26234 16668 26240 16720
rect 26292 16708 26298 16720
rect 27982 16708 27988 16720
rect 26292 16680 27988 16708
rect 26292 16668 26298 16680
rect 27982 16668 27988 16680
rect 28040 16708 28046 16720
rect 29546 16708 29552 16720
rect 28040 16680 29552 16708
rect 28040 16668 28046 16680
rect 29546 16668 29552 16680
rect 29604 16668 29610 16720
rect 26145 16643 26203 16649
rect 26145 16640 26157 16643
rect 26108 16612 26157 16640
rect 26108 16600 26114 16612
rect 26145 16609 26157 16612
rect 26191 16609 26203 16643
rect 26145 16603 26203 16609
rect 26329 16643 26387 16649
rect 26329 16609 26341 16643
rect 26375 16640 26387 16643
rect 27062 16640 27068 16652
rect 26375 16612 27068 16640
rect 26375 16609 26387 16612
rect 26329 16603 26387 16609
rect 27062 16600 27068 16612
rect 27120 16600 27126 16652
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16609 27399 16643
rect 27341 16603 27399 16609
rect 27356 16572 27384 16603
rect 27430 16600 27436 16652
rect 27488 16600 27494 16652
rect 28169 16643 28227 16649
rect 28169 16640 28181 16643
rect 27540 16612 28181 16640
rect 27540 16572 27568 16612
rect 28169 16609 28181 16612
rect 28215 16609 28227 16643
rect 28169 16603 28227 16609
rect 28258 16600 28264 16652
rect 28316 16600 28322 16652
rect 28534 16600 28540 16652
rect 28592 16640 28598 16652
rect 30116 16649 30144 16748
rect 37737 16711 37795 16717
rect 37737 16677 37749 16711
rect 37783 16677 37795 16711
rect 37737 16671 37795 16677
rect 29089 16643 29147 16649
rect 29089 16640 29101 16643
rect 28592 16612 29101 16640
rect 28592 16600 28598 16612
rect 29089 16609 29101 16612
rect 29135 16609 29147 16643
rect 29089 16603 29147 16609
rect 30101 16643 30159 16649
rect 30101 16609 30113 16643
rect 30147 16609 30159 16643
rect 33134 16640 33140 16652
rect 30101 16603 30159 16609
rect 31496 16612 33140 16640
rect 26436 16544 27568 16572
rect 26326 16504 26332 16516
rect 25976 16476 26332 16504
rect 26326 16464 26332 16476
rect 26384 16464 26390 16516
rect 26436 16448 26464 16544
rect 30374 16532 30380 16584
rect 30432 16572 30438 16584
rect 30469 16575 30527 16581
rect 30469 16572 30481 16575
rect 30432 16544 30481 16572
rect 30432 16532 30438 16544
rect 30469 16541 30481 16544
rect 30515 16572 30527 16575
rect 31496 16572 31524 16612
rect 33134 16600 33140 16612
rect 33192 16600 33198 16652
rect 36081 16643 36139 16649
rect 36081 16609 36093 16643
rect 36127 16640 36139 16643
rect 36170 16640 36176 16652
rect 36127 16612 36176 16640
rect 36127 16609 36139 16612
rect 36081 16603 36139 16609
rect 36170 16600 36176 16612
rect 36228 16640 36234 16652
rect 36357 16643 36415 16649
rect 36357 16640 36369 16643
rect 36228 16612 36369 16640
rect 36228 16600 36234 16612
rect 36357 16609 36369 16612
rect 36403 16609 36415 16643
rect 36357 16603 36415 16609
rect 37752 16584 37780 16671
rect 30515 16544 31524 16572
rect 30515 16541 30527 16544
rect 30469 16535 30527 16541
rect 32582 16532 32588 16584
rect 32640 16532 32646 16584
rect 35434 16532 35440 16584
rect 35492 16572 35498 16584
rect 37734 16572 37740 16584
rect 35492 16544 37740 16572
rect 35492 16532 35498 16544
rect 37734 16532 37740 16544
rect 37792 16532 37798 16584
rect 38378 16532 38384 16584
rect 38436 16532 38442 16584
rect 27249 16507 27307 16513
rect 27249 16473 27261 16507
rect 27295 16504 27307 16507
rect 28537 16507 28595 16513
rect 28537 16504 28549 16507
rect 27295 16476 28549 16504
rect 27295 16473 27307 16476
rect 27249 16467 27307 16473
rect 28537 16473 28549 16476
rect 28583 16473 28595 16507
rect 28537 16467 28595 16473
rect 30736 16507 30794 16513
rect 30736 16473 30748 16507
rect 30782 16504 30794 16507
rect 31941 16507 31999 16513
rect 31941 16504 31953 16507
rect 30782 16476 31953 16504
rect 30782 16473 30794 16476
rect 30736 16467 30794 16473
rect 31941 16473 31953 16476
rect 31987 16473 31999 16507
rect 31941 16467 31999 16473
rect 33404 16507 33462 16513
rect 33404 16473 33416 16507
rect 33450 16504 33462 16507
rect 33870 16504 33876 16516
rect 33450 16476 33876 16504
rect 33450 16473 33462 16476
rect 33404 16467 33462 16473
rect 33870 16464 33876 16476
rect 33928 16464 33934 16516
rect 35618 16504 35624 16516
rect 34532 16476 35624 16504
rect 25133 16439 25191 16445
rect 25133 16436 25145 16439
rect 25056 16408 25145 16436
rect 25133 16405 25145 16408
rect 25179 16405 25191 16439
rect 25133 16399 25191 16405
rect 26418 16396 26424 16448
rect 26476 16396 26482 16448
rect 26881 16439 26939 16445
rect 26881 16405 26893 16439
rect 26927 16436 26939 16439
rect 27614 16436 27620 16448
rect 26927 16408 27620 16436
rect 26927 16405 26939 16408
rect 26881 16399 26939 16405
rect 27614 16396 27620 16408
rect 27672 16396 27678 16448
rect 27709 16439 27767 16445
rect 27709 16405 27721 16439
rect 27755 16436 27767 16439
rect 27982 16436 27988 16448
rect 27755 16408 27988 16436
rect 27755 16405 27767 16408
rect 27709 16399 27767 16405
rect 27982 16396 27988 16408
rect 28040 16396 28046 16448
rect 28074 16396 28080 16448
rect 28132 16396 28138 16448
rect 29086 16396 29092 16448
rect 29144 16436 29150 16448
rect 29549 16439 29607 16445
rect 29549 16436 29561 16439
rect 29144 16408 29561 16436
rect 29144 16396 29150 16408
rect 29549 16405 29561 16408
rect 29595 16405 29607 16439
rect 29549 16399 29607 16405
rect 31846 16396 31852 16448
rect 31904 16396 31910 16448
rect 34532 16445 34560 16476
rect 35618 16464 35624 16476
rect 35676 16464 35682 16516
rect 35836 16507 35894 16513
rect 35836 16473 35848 16507
rect 35882 16504 35894 16507
rect 36078 16504 36084 16516
rect 35882 16476 36084 16504
rect 35882 16473 35894 16476
rect 35836 16467 35894 16473
rect 36078 16464 36084 16476
rect 36136 16464 36142 16516
rect 36624 16507 36682 16513
rect 36624 16473 36636 16507
rect 36670 16504 36682 16507
rect 37829 16507 37887 16513
rect 37829 16504 37841 16507
rect 36670 16476 37841 16504
rect 36670 16473 36682 16476
rect 36624 16467 36682 16473
rect 37829 16473 37841 16476
rect 37875 16473 37887 16507
rect 37829 16467 37887 16473
rect 34517 16439 34575 16445
rect 34517 16405 34529 16439
rect 34563 16405 34575 16439
rect 34517 16399 34575 16405
rect 34701 16439 34759 16445
rect 34701 16405 34713 16439
rect 34747 16436 34759 16439
rect 35342 16436 35348 16448
rect 34747 16408 35348 16436
rect 34747 16405 34759 16408
rect 34701 16399 34759 16405
rect 35342 16396 35348 16408
rect 35400 16396 35406 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 3786 16192 3792 16244
rect 3844 16192 3850 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5445 16235 5503 16241
rect 5445 16232 5457 16235
rect 5040 16204 5457 16232
rect 5040 16192 5046 16204
rect 5445 16201 5457 16204
rect 5491 16201 5503 16235
rect 5445 16195 5503 16201
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5813 16235 5871 16241
rect 5813 16232 5825 16235
rect 5592 16204 5825 16232
rect 5592 16192 5598 16204
rect 5813 16201 5825 16204
rect 5859 16201 5871 16235
rect 5813 16195 5871 16201
rect 5920 16204 7604 16232
rect 2584 16167 2642 16173
rect 2584 16133 2596 16167
rect 2630 16164 2642 16167
rect 2774 16164 2780 16176
rect 2630 16136 2780 16164
rect 2630 16133 2642 16136
rect 2584 16127 2642 16133
rect 2774 16124 2780 16136
rect 2832 16124 2838 16176
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 3804 16096 3832 16192
rect 4522 16124 4528 16176
rect 4580 16164 4586 16176
rect 5258 16164 5264 16176
rect 4580 16136 5264 16164
rect 4580 16124 4586 16136
rect 5258 16124 5264 16136
rect 5316 16164 5322 16176
rect 5920 16164 5948 16204
rect 5316 16136 5948 16164
rect 6724 16167 6782 16173
rect 5316 16124 5322 16136
rect 6724 16133 6736 16167
rect 6770 16164 6782 16167
rect 6914 16164 6920 16176
rect 6770 16136 6920 16164
rect 6770 16133 6782 16136
rect 6724 16127 6782 16133
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 1719 16068 3832 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 2314 15988 2320 16040
rect 2372 15988 2378 16040
rect 4540 16037 4568 16124
rect 4614 16056 4620 16108
rect 4672 16096 4678 16108
rect 4709 16099 4767 16105
rect 4709 16096 4721 16099
rect 4672 16068 4721 16096
rect 4672 16056 4678 16068
rect 4709 16065 4721 16068
rect 4755 16096 4767 16099
rect 5350 16096 5356 16108
rect 4755 16068 5356 16096
rect 4755 16065 4767 16068
rect 4709 16059 4767 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 5905 16031 5963 16037
rect 5905 16028 5917 16031
rect 5500 16000 5917 16028
rect 5500 15988 5506 16000
rect 5905 15997 5917 16000
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 6089 16031 6147 16037
rect 6089 15997 6101 16031
rect 6135 15997 6147 16031
rect 6089 15991 6147 15997
rect 5353 15963 5411 15969
rect 5353 15929 5365 15963
rect 5399 15960 5411 15963
rect 5994 15960 6000 15972
rect 5399 15932 6000 15960
rect 5399 15929 5411 15932
rect 5353 15923 5411 15929
rect 5994 15920 6000 15932
rect 6052 15960 6058 15972
rect 6104 15960 6132 15991
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6457 16031 6515 16037
rect 6457 16028 6469 16031
rect 6236 16000 6469 16028
rect 6236 15988 6242 16000
rect 6457 15997 6469 16000
rect 6503 15997 6515 16031
rect 6457 15991 6515 15997
rect 6362 15960 6368 15972
rect 6052 15932 6368 15960
rect 6052 15920 6058 15932
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 2225 15895 2283 15901
rect 2225 15861 2237 15895
rect 2271 15892 2283 15895
rect 3050 15892 3056 15904
rect 2271 15864 3056 15892
rect 2271 15861 2283 15864
rect 2225 15855 2283 15861
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 3697 15895 3755 15901
rect 3697 15861 3709 15895
rect 3743 15892 3755 15895
rect 4706 15892 4712 15904
rect 3743 15864 4712 15892
rect 3743 15861 3755 15864
rect 3697 15855 3755 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 7576 15892 7604 16204
rect 7742 16192 7748 16244
rect 7800 16192 7806 16244
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16201 7895 16235
rect 7837 16195 7895 16201
rect 7929 16235 7987 16241
rect 7929 16201 7941 16235
rect 7975 16232 7987 16235
rect 8386 16232 8392 16244
rect 7975 16204 8392 16232
rect 7975 16201 7987 16204
rect 7929 16195 7987 16201
rect 7760 16028 7788 16192
rect 7852 16164 7880 16195
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8478 16192 8484 16244
rect 8536 16192 8542 16244
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 10505 16235 10563 16241
rect 10505 16232 10517 16235
rect 9916 16204 10517 16232
rect 9916 16192 9922 16204
rect 10505 16201 10517 16204
rect 10551 16201 10563 16235
rect 10505 16195 10563 16201
rect 8496 16164 8524 16192
rect 7852 16136 8524 16164
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 8343 16068 8769 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 8757 16065 8769 16068
rect 8803 16065 8815 16099
rect 8757 16059 8815 16065
rect 8386 16028 8392 16040
rect 7760 16000 8392 16028
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 9214 16028 9220 16040
rect 8619 16000 9220 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 15997 9367 16031
rect 10520 16028 10548 16195
rect 12250 16192 12256 16244
rect 12308 16232 12314 16244
rect 12345 16235 12403 16241
rect 12345 16232 12357 16235
rect 12308 16204 12357 16232
rect 12308 16192 12314 16204
rect 12345 16201 12357 16204
rect 12391 16201 12403 16235
rect 12345 16195 12403 16201
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 15896 16204 16221 16232
rect 15896 16192 15902 16204
rect 16209 16201 16221 16204
rect 16255 16201 16267 16235
rect 16209 16195 16267 16201
rect 16574 16192 16580 16244
rect 16632 16192 16638 16244
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16232 17463 16235
rect 18690 16232 18696 16244
rect 17451 16204 18696 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 18874 16192 18880 16244
rect 18932 16192 18938 16244
rect 23290 16232 23296 16244
rect 23216 16204 23296 16232
rect 16117 16167 16175 16173
rect 16117 16133 16129 16167
rect 16163 16164 16175 16167
rect 16592 16164 16620 16192
rect 16942 16164 16948 16176
rect 16163 16136 16948 16164
rect 16163 16133 16175 16136
rect 16117 16127 16175 16133
rect 16942 16124 16948 16136
rect 17000 16164 17006 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 17000 16136 17049 16164
rect 17000 16124 17006 16136
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17037 16127 17095 16133
rect 18414 16124 18420 16176
rect 18472 16164 18478 16176
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 18472 16136 18521 16164
rect 18472 16124 18478 16136
rect 18509 16133 18521 16136
rect 18555 16164 18567 16167
rect 18892 16164 18920 16192
rect 18555 16136 18920 16164
rect 23048 16167 23106 16173
rect 18555 16133 18567 16136
rect 18509 16127 18567 16133
rect 23048 16133 23060 16167
rect 23094 16164 23106 16167
rect 23216 16164 23244 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 26329 16235 26387 16241
rect 26329 16201 26341 16235
rect 26375 16201 26387 16235
rect 26329 16195 26387 16201
rect 26234 16164 26240 16176
rect 23094 16136 23244 16164
rect 23308 16136 26240 16164
rect 23094 16133 23106 16136
rect 23048 16127 23106 16133
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16096 10839 16099
rect 11054 16096 11060 16108
rect 10827 16068 11060 16096
rect 10827 16065 10839 16068
rect 10781 16059 10839 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16096 11391 16099
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 11379 16068 11897 16096
rect 11379 16065 11391 16068
rect 11333 16059 11391 16065
rect 11885 16065 11897 16068
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12526 16096 12532 16108
rect 12023 16068 12532 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 18138 16056 18144 16108
rect 18196 16056 18202 16108
rect 23198 16056 23204 16108
rect 23256 16096 23262 16108
rect 23308 16105 23336 16136
rect 24780 16105 24808 16136
rect 26234 16124 26240 16136
rect 26292 16164 26298 16176
rect 26344 16164 26372 16195
rect 29546 16192 29552 16244
rect 29604 16232 29610 16244
rect 29917 16235 29975 16241
rect 29917 16232 29929 16235
rect 29604 16204 29929 16232
rect 29604 16192 29610 16204
rect 29917 16201 29929 16204
rect 29963 16201 29975 16235
rect 29917 16195 29975 16201
rect 34698 16192 34704 16244
rect 34756 16192 34762 16244
rect 35986 16192 35992 16244
rect 36044 16192 36050 16244
rect 36078 16192 36084 16244
rect 36136 16192 36142 16244
rect 37093 16235 37151 16241
rect 37093 16201 37105 16235
rect 37139 16232 37151 16235
rect 37182 16232 37188 16244
rect 37139 16204 37188 16232
rect 37139 16201 37151 16204
rect 37093 16195 37151 16201
rect 37182 16192 37188 16204
rect 37240 16192 37246 16244
rect 38013 16235 38071 16241
rect 38013 16201 38025 16235
rect 38059 16232 38071 16235
rect 38378 16232 38384 16244
rect 38059 16204 38384 16232
rect 38059 16201 38071 16204
rect 38013 16195 38071 16201
rect 38378 16192 38384 16204
rect 38436 16192 38442 16244
rect 26292 16136 26372 16164
rect 26292 16124 26298 16136
rect 23293 16099 23351 16105
rect 23293 16096 23305 16099
rect 23256 16068 23305 16096
rect 23256 16056 23262 16068
rect 23293 16065 23305 16068
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 24509 16099 24567 16105
rect 24509 16065 24521 16099
rect 24555 16096 24567 16099
rect 24765 16099 24823 16105
rect 24555 16068 24716 16096
rect 24555 16065 24567 16068
rect 24509 16059 24567 16065
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 10520 16000 11713 16028
rect 9309 15991 9367 15997
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 16206 16028 16212 16040
rect 15335 16000 16212 16028
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 9324 15960 9352 15991
rect 8260 15932 9352 15960
rect 11716 15960 11744 15991
rect 16206 15988 16212 16000
rect 16264 16028 16270 16040
rect 16301 16031 16359 16037
rect 16301 16028 16313 16031
rect 16264 16000 16313 16028
rect 16264 15988 16270 16000
rect 16301 15997 16313 16000
rect 16347 15997 16359 16031
rect 16758 16028 16764 16040
rect 16301 15991 16359 15997
rect 16408 16000 16764 16028
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 11716 15932 15577 15960
rect 8260 15920 8266 15932
rect 15565 15929 15577 15932
rect 15611 15960 15623 15963
rect 16408 15960 16436 16000
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 16991 16000 17509 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 24688 16028 24716 16068
rect 24765 16065 24777 16099
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 26142 16096 26148 16108
rect 25096 16068 26148 16096
rect 25096 16056 25102 16068
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 26344 16096 26372 16136
rect 28626 16124 28632 16176
rect 28684 16124 28690 16176
rect 31846 16124 31852 16176
rect 31904 16164 31910 16176
rect 31904 16136 34192 16164
rect 31904 16124 31910 16136
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26344 16068 26985 16096
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27240 16099 27298 16105
rect 27240 16065 27252 16099
rect 27286 16096 27298 16099
rect 27706 16096 27712 16108
rect 27286 16068 27712 16096
rect 27286 16065 27298 16068
rect 27240 16059 27298 16065
rect 27706 16056 27712 16068
rect 27764 16056 27770 16108
rect 34164 16105 34192 16136
rect 30736 16099 30794 16105
rect 30736 16065 30748 16099
rect 30782 16096 30794 16099
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 30782 16068 32137 16096
rect 30782 16065 30794 16068
rect 30736 16059 30794 16065
rect 32125 16065 32137 16068
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 34149 16099 34207 16105
rect 34149 16065 34161 16099
rect 34195 16065 34207 16099
rect 34149 16059 34207 16065
rect 35342 16056 35348 16108
rect 35400 16056 35406 16108
rect 36262 16056 36268 16108
rect 36320 16096 36326 16108
rect 36633 16099 36691 16105
rect 36633 16096 36645 16099
rect 36320 16068 36645 16096
rect 36320 16056 36326 16068
rect 36633 16065 36645 16068
rect 36679 16065 36691 16099
rect 36633 16059 36691 16065
rect 24946 16028 24952 16040
rect 24688 16000 24952 16028
rect 17497 15991 17555 15997
rect 24946 15988 24952 16000
rect 25004 15988 25010 16040
rect 29730 15988 29736 16040
rect 29788 16028 29794 16040
rect 30374 16028 30380 16040
rect 29788 16000 30380 16028
rect 29788 15988 29794 16000
rect 30374 15988 30380 16000
rect 30432 16028 30438 16040
rect 30469 16031 30527 16037
rect 30469 16028 30481 16031
rect 30432 16000 30481 16028
rect 30432 15988 30438 16000
rect 30469 15997 30481 16000
rect 30515 15997 30527 16031
rect 30469 15991 30527 15997
rect 32398 15988 32404 16040
rect 32456 16028 32462 16040
rect 32677 16031 32735 16037
rect 32677 16028 32689 16031
rect 32456 16000 32689 16028
rect 32456 15988 32462 16000
rect 32677 15997 32689 16000
rect 32723 15997 32735 16031
rect 32677 15991 32735 15997
rect 33413 16031 33471 16037
rect 33413 15997 33425 16031
rect 33459 15997 33471 16031
rect 33413 15991 33471 15997
rect 15611 15932 16436 15960
rect 15611 15929 15623 15932
rect 15565 15923 15623 15929
rect 31570 15920 31576 15972
rect 31628 15960 31634 15972
rect 31849 15963 31907 15969
rect 31849 15960 31861 15963
rect 31628 15932 31861 15960
rect 31628 15920 31634 15932
rect 31849 15929 31861 15932
rect 31895 15960 31907 15963
rect 33428 15960 33456 15991
rect 34790 15988 34796 16040
rect 34848 15988 34854 16040
rect 34977 16031 35035 16037
rect 34977 15997 34989 16031
rect 35023 16028 35035 16031
rect 35710 16028 35716 16040
rect 35023 16000 35716 16028
rect 35023 15997 35035 16000
rect 34977 15991 35035 15997
rect 34992 15960 35020 15991
rect 35710 15988 35716 16000
rect 35768 15988 35774 16040
rect 37200 16028 37228 16192
rect 37642 16056 37648 16108
rect 37700 16056 37706 16108
rect 37366 16028 37372 16040
rect 37200 16000 37372 16028
rect 37366 15988 37372 16000
rect 37424 15988 37430 16040
rect 37550 15988 37556 16040
rect 37608 16028 37614 16040
rect 38378 16028 38384 16040
rect 37608 16000 38384 16028
rect 37608 15988 37614 16000
rect 38378 15988 38384 16000
rect 38436 15988 38442 16040
rect 31895 15932 33456 15960
rect 33520 15932 35020 15960
rect 31895 15929 31907 15932
rect 31849 15923 31907 15929
rect 8846 15892 8852 15904
rect 7576 15864 8852 15892
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 15746 15852 15752 15904
rect 15804 15852 15810 15904
rect 21913 15895 21971 15901
rect 21913 15861 21925 15895
rect 21959 15892 21971 15895
rect 23290 15892 23296 15904
rect 21959 15864 23296 15892
rect 21959 15861 21971 15864
rect 21913 15855 21971 15861
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 23382 15852 23388 15904
rect 23440 15852 23446 15904
rect 28353 15895 28411 15901
rect 28353 15861 28365 15895
rect 28399 15892 28411 15895
rect 28442 15892 28448 15904
rect 28399 15864 28448 15892
rect 28399 15861 28411 15864
rect 28353 15855 28411 15861
rect 28442 15852 28448 15864
rect 28500 15852 28506 15904
rect 32858 15852 32864 15904
rect 32916 15852 32922 15904
rect 32950 15852 32956 15904
rect 33008 15892 33014 15904
rect 33520 15892 33548 15932
rect 33008 15864 33548 15892
rect 33008 15852 33014 15864
rect 33594 15852 33600 15904
rect 33652 15852 33658 15904
rect 34330 15852 34336 15904
rect 34388 15852 34394 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 2130 15648 2136 15700
rect 2188 15648 2194 15700
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 4856 15660 5733 15688
rect 4856 15648 4862 15660
rect 5721 15657 5733 15660
rect 5767 15657 5779 15691
rect 5721 15651 5779 15657
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 9824 15660 10057 15688
rect 9824 15648 9830 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15565 15691 15623 15697
rect 15565 15688 15577 15691
rect 15436 15660 15577 15688
rect 15436 15648 15442 15660
rect 15565 15657 15577 15660
rect 15611 15657 15623 15691
rect 15565 15651 15623 15657
rect 15746 15648 15752 15700
rect 15804 15648 15810 15700
rect 17034 15688 17040 15700
rect 16592 15660 17040 15688
rect 3602 15580 3608 15632
rect 3660 15620 3666 15632
rect 7653 15623 7711 15629
rect 3660 15592 4568 15620
rect 3660 15580 3666 15592
rect 1578 15512 1584 15564
rect 1636 15512 1642 15564
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 4540 15552 4568 15592
rect 7653 15589 7665 15623
rect 7699 15620 7711 15623
rect 7834 15620 7840 15632
rect 7699 15592 7840 15620
rect 7699 15589 7711 15592
rect 7653 15583 7711 15589
rect 7834 15580 7840 15592
rect 7892 15580 7898 15632
rect 12069 15623 12127 15629
rect 12069 15589 12081 15623
rect 12115 15589 12127 15623
rect 12069 15583 12127 15589
rect 4826 15555 4884 15561
rect 4826 15552 4838 15555
rect 4540 15524 4838 15552
rect 4826 15521 4838 15524
rect 4872 15521 4884 15555
rect 4826 15515 4884 15521
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5031 15524 6592 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15484 2283 15487
rect 2314 15484 2320 15496
rect 2271 15456 2320 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2314 15444 2320 15456
rect 2372 15484 2378 15496
rect 2774 15484 2780 15496
rect 2372 15456 2780 15484
rect 2372 15444 2378 15456
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3620 15456 3801 15484
rect 2492 15419 2550 15425
rect 2492 15385 2504 15419
rect 2538 15416 2550 15419
rect 2590 15416 2596 15428
rect 2538 15388 2596 15416
rect 2538 15385 2550 15388
rect 2492 15379 2550 15385
rect 2590 15376 2596 15388
rect 2648 15376 2654 15428
rect 1670 15308 1676 15360
rect 1728 15308 1734 15360
rect 1765 15351 1823 15357
rect 1765 15317 1777 15351
rect 1811 15348 1823 15351
rect 2406 15348 2412 15360
rect 1811 15320 2412 15348
rect 1811 15317 1823 15320
rect 1765 15311 1823 15317
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 3326 15308 3332 15360
rect 3384 15348 3390 15360
rect 3620 15357 3648 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 3605 15351 3663 15357
rect 3605 15348 3617 15351
rect 3384 15320 3617 15348
rect 3384 15308 3390 15320
rect 3605 15317 3617 15320
rect 3651 15317 3663 15351
rect 3988 15348 4016 15447
rect 4706 15444 4712 15496
rect 4764 15444 4770 15496
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 6288 15416 6316 15447
rect 5460 15388 6316 15416
rect 4154 15348 4160 15360
rect 3988 15320 4160 15348
rect 3605 15311 3663 15317
rect 4154 15308 4160 15320
rect 4212 15348 4218 15360
rect 5460 15348 5488 15388
rect 4212 15320 5488 15348
rect 4212 15308 4218 15320
rect 5626 15308 5632 15360
rect 5684 15308 5690 15360
rect 6454 15308 6460 15360
rect 6512 15308 6518 15360
rect 6564 15348 6592 15524
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 8113 15555 8171 15561
rect 6972 15524 7282 15552
rect 6972 15512 6978 15524
rect 7098 15444 7104 15496
rect 7156 15444 7162 15496
rect 7254 15493 7282 15524
rect 8113 15521 8125 15555
rect 8159 15552 8171 15555
rect 8202 15552 8208 15564
rect 8159 15524 8208 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 8478 15552 8484 15564
rect 8343 15524 8484 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15552 12035 15555
rect 12084 15552 12112 15583
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 12023 15524 12112 15552
rect 12406 15524 12725 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 7239 15487 7297 15493
rect 7239 15453 7251 15487
rect 7285 15453 7297 15487
rect 7239 15447 7297 15453
rect 7374 15444 7380 15496
rect 7432 15444 7438 15496
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 12406 15484 12434 15524
rect 12713 15521 12725 15524
rect 12759 15552 12771 15555
rect 13814 15552 13820 15564
rect 12759 15524 13820 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 15764 15552 15792 15648
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 15764 15524 16129 15552
rect 16117 15521 16129 15524
rect 16163 15521 16175 15555
rect 16117 15515 16175 15521
rect 11296 15456 12434 15484
rect 11296 15444 11302 15456
rect 12526 15444 12532 15496
rect 12584 15444 12590 15496
rect 12894 15444 12900 15496
rect 12952 15484 12958 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 12952 15456 13461 15484
rect 12952 15444 12958 15456
rect 13449 15453 13461 15456
rect 13495 15484 13507 15487
rect 13538 15484 13544 15496
rect 13495 15456 13544 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 16592 15484 16620 15660
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 26234 15688 26240 15700
rect 26068 15660 26240 15688
rect 17494 15620 17500 15632
rect 16960 15592 17500 15620
rect 16960 15564 16988 15592
rect 17494 15580 17500 15592
rect 17552 15620 17558 15632
rect 17552 15592 18552 15620
rect 17552 15580 17558 15592
rect 16666 15512 16672 15564
rect 16724 15512 16730 15564
rect 16942 15512 16948 15564
rect 17000 15512 17006 15564
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 17865 15555 17923 15561
rect 17865 15521 17877 15555
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 18325 15555 18383 15561
rect 18325 15521 18337 15555
rect 18371 15552 18383 15555
rect 18414 15552 18420 15564
rect 18371 15524 18420 15552
rect 18371 15521 18383 15524
rect 18325 15515 18383 15521
rect 15028 15456 16620 15484
rect 16684 15484 16712 15512
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 16684 15456 17785 15484
rect 8665 15419 8723 15425
rect 8665 15385 8677 15419
rect 8711 15416 8723 15419
rect 9306 15416 9312 15428
rect 8711 15388 9312 15416
rect 8711 15385 8723 15388
rect 8665 15379 8723 15385
rect 7098 15348 7104 15360
rect 6564 15320 7104 15348
rect 7098 15308 7104 15320
rect 7156 15348 7162 15360
rect 8680 15348 8708 15379
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 9950 15376 9956 15428
rect 10008 15376 10014 15428
rect 12437 15419 12495 15425
rect 12437 15385 12449 15419
rect 12483 15416 12495 15419
rect 12544 15416 12572 15444
rect 12802 15416 12808 15428
rect 12483 15388 12808 15416
rect 12483 15385 12495 15388
rect 12437 15379 12495 15385
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 7156 15320 8708 15348
rect 7156 15308 7162 15320
rect 9214 15308 9220 15360
rect 9272 15348 9278 15360
rect 9674 15348 9680 15360
rect 9272 15320 9680 15348
rect 9272 15308 9278 15320
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11606 15348 11612 15360
rect 11379 15320 11612 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12575 15320 12909 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12897 15317 12909 15320
rect 12943 15317 12955 15351
rect 12897 15311 12955 15317
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 15028 15357 15056 15456
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 17880 15416 17908 15515
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 18524 15493 18552 15592
rect 22830 15512 22836 15564
rect 22888 15552 22894 15564
rect 23382 15552 23388 15564
rect 22888 15524 23388 15552
rect 22888 15512 22894 15524
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 23566 15512 23572 15564
rect 23624 15512 23630 15564
rect 23753 15555 23811 15561
rect 23753 15521 23765 15555
rect 23799 15552 23811 15555
rect 23799 15524 24992 15552
rect 23799 15521 23811 15524
rect 23753 15515 23811 15521
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 15528 15388 17908 15416
rect 18524 15416 18552 15447
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 23198 15484 23204 15496
rect 21692 15456 23204 15484
rect 21692 15444 21698 15456
rect 23198 15444 23204 15456
rect 23256 15444 23262 15496
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 24302 15484 24308 15496
rect 23523 15456 24308 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 24302 15444 24308 15456
rect 24360 15444 24366 15496
rect 24857 15487 24915 15493
rect 24857 15453 24869 15487
rect 24903 15453 24915 15487
rect 24857 15447 24915 15453
rect 20070 15416 20076 15428
rect 18524 15388 20076 15416
rect 15528 15376 15534 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 21910 15425 21916 15428
rect 21904 15379 21916 15425
rect 21910 15376 21916 15379
rect 21968 15376 21974 15428
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 23032 15388 23888 15416
rect 15013 15351 15071 15357
rect 15013 15348 15025 15351
rect 13964 15320 15025 15348
rect 13964 15308 13970 15320
rect 15013 15317 15025 15320
rect 15059 15317 15071 15351
rect 15013 15311 15071 15317
rect 16482 15308 16488 15360
rect 16540 15308 16546 15360
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 17310 15308 17316 15360
rect 17368 15308 17374 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 17460 15320 17693 15348
rect 17460 15308 17466 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 18414 15308 18420 15360
rect 18472 15308 18478 15360
rect 18877 15351 18935 15357
rect 18877 15317 18889 15351
rect 18923 15348 18935 15351
rect 19334 15348 19340 15360
rect 18923 15320 19340 15348
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 19334 15308 19340 15320
rect 19392 15308 19398 15360
rect 20438 15308 20444 15360
rect 20496 15348 20502 15360
rect 23032 15357 23060 15388
rect 23860 15360 23888 15388
rect 23952 15388 24685 15416
rect 23952 15360 23980 15388
rect 24673 15385 24685 15388
rect 24719 15416 24731 15419
rect 24872 15416 24900 15447
rect 24719 15388 24900 15416
rect 24719 15385 24731 15388
rect 24673 15379 24731 15385
rect 20533 15351 20591 15357
rect 20533 15348 20545 15351
rect 20496 15320 20545 15348
rect 20496 15308 20502 15320
rect 20533 15317 20545 15320
rect 20579 15317 20591 15351
rect 20533 15311 20591 15317
rect 23017 15351 23075 15357
rect 23017 15317 23029 15351
rect 23063 15317 23075 15351
rect 23017 15311 23075 15317
rect 23106 15308 23112 15360
rect 23164 15308 23170 15360
rect 23842 15308 23848 15360
rect 23900 15308 23906 15360
rect 23934 15308 23940 15360
rect 23992 15308 23998 15360
rect 24213 15351 24271 15357
rect 24213 15317 24225 15351
rect 24259 15348 24271 15351
rect 24964 15348 24992 15524
rect 25682 15512 25688 15564
rect 25740 15512 25746 15564
rect 26068 15561 26096 15660
rect 26234 15648 26240 15660
rect 26292 15648 26298 15700
rect 27433 15691 27491 15697
rect 27433 15657 27445 15691
rect 27479 15688 27491 15691
rect 27798 15688 27804 15700
rect 27479 15660 27804 15688
rect 27479 15657 27491 15660
rect 27433 15651 27491 15657
rect 27798 15648 27804 15660
rect 27856 15688 27862 15700
rect 28534 15688 28540 15700
rect 27856 15660 28540 15688
rect 27856 15648 27862 15660
rect 28534 15648 28540 15660
rect 28592 15648 28598 15700
rect 29086 15648 29092 15700
rect 29144 15648 29150 15700
rect 30098 15648 30104 15700
rect 30156 15688 30162 15700
rect 30156 15660 32352 15688
rect 30156 15648 30162 15660
rect 27525 15623 27583 15629
rect 27525 15589 27537 15623
rect 27571 15620 27583 15623
rect 27890 15620 27896 15632
rect 27571 15592 27896 15620
rect 27571 15589 27583 15592
rect 27525 15583 27583 15589
rect 27890 15580 27896 15592
rect 27948 15580 27954 15632
rect 26053 15555 26111 15561
rect 26053 15521 26065 15555
rect 26099 15521 26111 15555
rect 26053 15515 26111 15521
rect 26320 15487 26378 15493
rect 26320 15453 26332 15487
rect 26366 15484 26378 15487
rect 26786 15484 26792 15496
rect 26366 15456 26792 15484
rect 26366 15453 26378 15456
rect 26320 15447 26378 15453
rect 26786 15444 26792 15456
rect 26844 15444 26850 15496
rect 27908 15416 27936 15580
rect 29104 15552 29132 15648
rect 31846 15580 31852 15632
rect 31904 15580 31910 15632
rect 28828 15524 29132 15552
rect 29365 15555 29423 15561
rect 28649 15487 28707 15493
rect 28649 15453 28661 15487
rect 28695 15484 28707 15487
rect 28828 15484 28856 15524
rect 29365 15521 29377 15555
rect 29411 15552 29423 15555
rect 30282 15552 30288 15564
rect 29411 15524 30288 15552
rect 29411 15521 29423 15524
rect 29365 15515 29423 15521
rect 30282 15512 30288 15524
rect 30340 15512 30346 15564
rect 30926 15512 30932 15564
rect 30984 15552 30990 15564
rect 31113 15555 31171 15561
rect 31113 15552 31125 15555
rect 30984 15524 31125 15552
rect 30984 15512 30990 15524
rect 31113 15521 31125 15524
rect 31159 15521 31171 15555
rect 31113 15515 31171 15521
rect 31386 15512 31392 15564
rect 31444 15512 31450 15564
rect 31570 15512 31576 15564
rect 31628 15552 31634 15564
rect 31665 15555 31723 15561
rect 31665 15552 31677 15555
rect 31628 15524 31677 15552
rect 31628 15512 31634 15524
rect 31665 15521 31677 15524
rect 31711 15521 31723 15555
rect 31864 15552 31892 15580
rect 32125 15555 32183 15561
rect 32125 15552 32137 15555
rect 31864 15524 32137 15552
rect 31665 15515 31723 15521
rect 32125 15521 32137 15524
rect 32171 15521 32183 15555
rect 32324 15552 32352 15660
rect 33870 15648 33876 15700
rect 33928 15648 33934 15700
rect 34330 15648 34336 15700
rect 34388 15648 34394 15700
rect 34701 15691 34759 15697
rect 34701 15657 34713 15691
rect 34747 15688 34759 15691
rect 34790 15688 34796 15700
rect 34747 15660 34796 15688
rect 34747 15657 34759 15660
rect 34701 15651 34759 15657
rect 34790 15648 34796 15660
rect 34848 15648 34854 15700
rect 35618 15648 35624 15700
rect 35676 15648 35682 15700
rect 35710 15648 35716 15700
rect 35768 15648 35774 15700
rect 36354 15648 36360 15700
rect 36412 15648 36418 15700
rect 37642 15648 37648 15700
rect 37700 15688 37706 15700
rect 37737 15691 37795 15697
rect 37737 15688 37749 15691
rect 37700 15660 37749 15688
rect 37700 15648 37706 15660
rect 37737 15657 37749 15660
rect 37783 15657 37795 15691
rect 37737 15651 37795 15657
rect 32401 15623 32459 15629
rect 32401 15589 32413 15623
rect 32447 15620 32459 15623
rect 33134 15620 33140 15632
rect 32447 15592 33140 15620
rect 32447 15589 32459 15592
rect 32401 15583 32459 15589
rect 33134 15580 33140 15592
rect 33192 15580 33198 15632
rect 32324 15524 32536 15552
rect 32125 15515 32183 15521
rect 28695 15456 28856 15484
rect 28905 15487 28963 15493
rect 28695 15453 28707 15456
rect 28649 15447 28707 15453
rect 28905 15453 28917 15487
rect 28951 15484 28963 15487
rect 29730 15484 29736 15496
rect 28951 15456 29736 15484
rect 28951 15453 28963 15456
rect 28905 15447 28963 15453
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 31202 15444 31208 15496
rect 31260 15493 31266 15496
rect 31260 15487 31309 15493
rect 31260 15453 31263 15487
rect 31297 15453 31309 15487
rect 31260 15447 31309 15453
rect 31260 15444 31266 15447
rect 32306 15444 32312 15496
rect 32364 15444 32370 15496
rect 28810 15416 28816 15428
rect 27908 15388 28816 15416
rect 28810 15376 28816 15388
rect 28868 15376 28874 15428
rect 30009 15419 30067 15425
rect 30009 15385 30021 15419
rect 30055 15416 30067 15419
rect 30558 15416 30564 15428
rect 30055 15388 30564 15416
rect 30055 15385 30067 15388
rect 30009 15379 30067 15385
rect 30558 15376 30564 15388
rect 30616 15376 30622 15428
rect 32508 15360 32536 15524
rect 32674 15512 32680 15564
rect 32732 15552 32738 15564
rect 32953 15555 33011 15561
rect 32953 15552 32965 15555
rect 32732 15524 32965 15552
rect 32732 15512 32738 15524
rect 32953 15521 32965 15524
rect 32999 15552 33011 15555
rect 33318 15552 33324 15564
rect 32999 15524 33324 15552
rect 32999 15521 33011 15524
rect 32953 15515 33011 15521
rect 33318 15512 33324 15524
rect 33376 15552 33382 15564
rect 33413 15555 33471 15561
rect 33413 15552 33425 15555
rect 33376 15524 33425 15552
rect 33376 15512 33382 15524
rect 33413 15521 33425 15524
rect 33459 15521 33471 15555
rect 34348 15552 34376 15648
rect 34425 15555 34483 15561
rect 34425 15552 34437 15555
rect 34348 15524 34437 15552
rect 33413 15515 33471 15521
rect 34425 15521 34437 15524
rect 34471 15521 34483 15555
rect 34425 15515 34483 15521
rect 35345 15555 35403 15561
rect 35345 15521 35357 15555
rect 35391 15552 35403 15555
rect 35636 15552 35664 15648
rect 35391 15524 35664 15552
rect 35391 15521 35403 15524
rect 35345 15515 35403 15521
rect 37734 15512 37740 15564
rect 37792 15552 37798 15564
rect 38289 15555 38347 15561
rect 38289 15552 38301 15555
rect 37792 15524 38301 15552
rect 37792 15512 37798 15524
rect 38289 15521 38301 15524
rect 38335 15521 38347 15555
rect 38289 15515 38347 15521
rect 36446 15376 36452 15428
rect 36504 15376 36510 15428
rect 25222 15348 25228 15360
rect 24259 15320 25228 15348
rect 24259 15317 24271 15320
rect 24213 15311 24271 15317
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 29641 15351 29699 15357
rect 29641 15317 29653 15351
rect 29687 15348 29699 15351
rect 29914 15348 29920 15360
rect 29687 15320 29920 15348
rect 29687 15317 29699 15320
rect 29641 15311 29699 15317
rect 29914 15308 29920 15320
rect 29972 15308 29978 15360
rect 30098 15308 30104 15360
rect 30156 15308 30162 15360
rect 30469 15351 30527 15357
rect 30469 15317 30481 15351
rect 30515 15348 30527 15351
rect 32122 15348 32128 15360
rect 30515 15320 32128 15348
rect 30515 15317 30527 15320
rect 30469 15311 30527 15317
rect 32122 15308 32128 15320
rect 32180 15308 32186 15360
rect 32490 15308 32496 15360
rect 32548 15348 32554 15360
rect 32769 15351 32827 15357
rect 32769 15348 32781 15351
rect 32548 15320 32781 15348
rect 32548 15308 32554 15320
rect 32769 15317 32781 15320
rect 32815 15317 32827 15351
rect 32769 15311 32827 15317
rect 32861 15351 32919 15357
rect 32861 15317 32873 15351
rect 32907 15348 32919 15351
rect 33226 15348 33232 15360
rect 32907 15320 33232 15348
rect 32907 15317 32919 15320
rect 32861 15311 32919 15317
rect 33226 15308 33232 15320
rect 33284 15308 33290 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1596 15116 4108 15144
rect 1596 15088 1624 15116
rect 1578 15036 1584 15088
rect 1636 15036 1642 15088
rect 2406 15036 2412 15088
rect 2464 15036 2470 15088
rect 3050 15085 3056 15088
rect 3022 15079 3056 15085
rect 3022 15045 3034 15079
rect 3022 15039 3056 15045
rect 3050 15036 3056 15039
rect 3108 15036 3114 15088
rect 4080 15076 4108 15116
rect 4154 15104 4160 15156
rect 4212 15104 4218 15156
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 4488 15116 5580 15144
rect 4488 15104 4494 15116
rect 4890 15076 4896 15088
rect 4080 15048 4896 15076
rect 4890 15036 4896 15048
rect 4948 15076 4954 15088
rect 5552 15076 5580 15116
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5684 15116 5825 15144
rect 5684 15104 5690 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 5905 15147 5963 15153
rect 5905 15113 5917 15147
rect 5951 15144 5963 15147
rect 6454 15144 6460 15156
rect 5951 15116 6460 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 7834 15144 7840 15156
rect 6696 15116 7840 15144
rect 6696 15104 6702 15116
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 8113 15147 8171 15153
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 8573 15147 8631 15153
rect 8573 15144 8585 15147
rect 8444 15116 8585 15144
rect 8444 15104 8450 15116
rect 8573 15113 8585 15116
rect 8619 15113 8631 15147
rect 8573 15107 8631 15113
rect 10962 15104 10968 15156
rect 11020 15104 11026 15156
rect 11072 15116 12848 15144
rect 6656 15076 6684 15104
rect 4948 15048 5120 15076
rect 5552 15048 6684 15076
rect 7000 15079 7058 15085
rect 4948 15036 4954 15048
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 15008 2375 15011
rect 2866 15008 2872 15020
rect 2363 14980 2872 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 4430 14968 4436 15020
rect 4488 14968 4494 15020
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 2593 14903 2651 14909
rect 1857 14875 1915 14881
rect 1857 14841 1869 14875
rect 1903 14872 1915 14875
rect 2608 14872 2636 14903
rect 2774 14900 2780 14952
rect 2832 14900 2838 14952
rect 5092 14949 5120 15048
rect 7000 15045 7012 15079
rect 7046 15076 7058 15079
rect 7650 15076 7656 15088
rect 7046 15048 7656 15076
rect 7046 15045 7058 15048
rect 7000 15039 7058 15045
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 11072 15076 11100 15116
rect 12434 15076 12440 15088
rect 7760 15048 11100 15076
rect 11532 15048 12440 15076
rect 7760 15008 7788 15048
rect 6196 14980 7788 15008
rect 8404 14980 8616 15008
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5123 14912 5948 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 1903 14844 2636 14872
rect 1903 14841 1915 14844
rect 1857 14835 1915 14841
rect 1946 14764 1952 14816
rect 2004 14764 2010 14816
rect 2608 14804 2636 14844
rect 4246 14804 4252 14816
rect 2608 14776 4252 14804
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 5445 14807 5503 14813
rect 5445 14804 5457 14807
rect 4856 14776 5457 14804
rect 4856 14764 4862 14776
rect 5445 14773 5457 14776
rect 5491 14773 5503 14807
rect 5920 14804 5948 14912
rect 6086 14900 6092 14952
rect 6144 14940 6150 14952
rect 6196 14940 6224 14980
rect 8404 14949 8432 14980
rect 8588 14952 8616 14980
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 9364 14980 11284 15008
rect 9364 14968 9370 14980
rect 6144 14912 6224 14940
rect 6733 14943 6791 14949
rect 6144 14900 6150 14912
rect 6733 14909 6745 14943
rect 6779 14909 6791 14943
rect 6733 14903 6791 14909
rect 8389 14943 8447 14949
rect 8389 14909 8401 14943
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 6178 14832 6184 14884
rect 6236 14872 6242 14884
rect 6748 14872 6776 14903
rect 8478 14900 8484 14952
rect 8536 14900 8542 14952
rect 8570 14900 8576 14952
rect 8628 14900 8634 14952
rect 9585 14943 9643 14949
rect 9585 14940 9597 14943
rect 8956 14912 9597 14940
rect 8956 14881 8984 14912
rect 9585 14909 9597 14912
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 6236 14844 6776 14872
rect 8941 14875 8999 14881
rect 6236 14832 6242 14844
rect 8941 14841 8953 14875
rect 8987 14841 8999 14875
rect 11256 14872 11284 14980
rect 11330 14900 11336 14952
rect 11388 14940 11394 14952
rect 11532 14949 11560 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 12820 15076 12848 15116
rect 12894 15104 12900 15156
rect 12952 15104 12958 15156
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 13354 15144 13360 15156
rect 13311 15116 13360 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 14461 15147 14519 15153
rect 14461 15113 14473 15147
rect 14507 15144 14519 15147
rect 15470 15144 15476 15156
rect 14507 15116 15476 15144
rect 14507 15113 14519 15116
rect 14461 15107 14519 15113
rect 12820 15048 13216 15076
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11773 15011 11831 15017
rect 11773 15008 11785 15011
rect 11664 14980 11785 15008
rect 11664 14968 11670 14980
rect 11773 14977 11785 14980
rect 11819 14977 11831 15011
rect 11773 14971 11831 14977
rect 13188 14949 13216 15048
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11388 14912 11529 14940
rect 11388 14900 11394 14912
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 14476 14940 14504 15107
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 16669 15147 16727 15153
rect 16669 15113 16681 15147
rect 16715 15144 16727 15147
rect 16850 15144 16856 15156
rect 16715 15116 16856 15144
rect 16715 15113 16727 15116
rect 16669 15107 16727 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17402 15104 17408 15156
rect 17460 15104 17466 15156
rect 17954 15144 17960 15156
rect 17512 15116 17960 15144
rect 15749 15079 15807 15085
rect 15749 15045 15761 15079
rect 15795 15076 15807 15079
rect 17512 15076 17540 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 20070 15144 20076 15156
rect 19576 15116 20076 15144
rect 19576 15104 19582 15116
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 21821 15147 21879 15153
rect 21821 15113 21833 15147
rect 21867 15144 21879 15147
rect 21910 15144 21916 15156
rect 21867 15116 21916 15144
rect 21867 15113 21879 15116
rect 21821 15107 21879 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 23106 15144 23112 15156
rect 22480 15116 23112 15144
rect 15795 15048 17540 15076
rect 15795 15045 15807 15048
rect 15749 15039 15807 15045
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 16482 15008 16488 15020
rect 15979 14980 16488 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 18046 14968 18052 15020
rect 18104 14968 18110 15020
rect 18892 14980 19748 15008
rect 13219 14912 14504 14940
rect 17313 14943 17371 14949
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 17862 14940 17868 14952
rect 17359 14912 17868 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 17862 14900 17868 14912
rect 17920 14940 17926 14952
rect 18187 14943 18245 14949
rect 18187 14940 18199 14943
rect 17920 14912 18199 14940
rect 17920 14900 17926 14912
rect 18187 14909 18199 14912
rect 18233 14909 18245 14943
rect 18187 14903 18245 14909
rect 18325 14943 18383 14949
rect 18325 14909 18337 14943
rect 18371 14940 18383 14943
rect 18506 14940 18512 14952
rect 18371 14912 18512 14940
rect 18371 14909 18383 14912
rect 18325 14903 18383 14909
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 18598 14900 18604 14952
rect 18656 14900 18662 14952
rect 11256 14844 11376 14872
rect 8941 14835 8999 14841
rect 8202 14804 8208 14816
rect 5920 14776 8208 14804
rect 5445 14767 5503 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 9030 14764 9036 14816
rect 9088 14764 9094 14816
rect 11348 14813 11376 14844
rect 12986 14832 12992 14884
rect 13044 14872 13050 14884
rect 15289 14875 15347 14881
rect 15289 14872 15301 14875
rect 13044 14844 15301 14872
rect 13044 14832 13050 14844
rect 15289 14841 15301 14844
rect 15335 14872 15347 14875
rect 17402 14872 17408 14884
rect 15335 14844 17408 14872
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 17402 14832 17408 14844
rect 17460 14832 17466 14884
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 12250 14804 12256 14816
rect 11379 14776 12256 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 12250 14764 12256 14776
rect 12308 14804 12314 14816
rect 13078 14804 13084 14816
rect 12308 14776 13084 14804
rect 12308 14764 12314 14776
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13722 14764 13728 14816
rect 13780 14764 13786 14816
rect 14090 14764 14096 14816
rect 14148 14764 14154 14816
rect 16485 14807 16543 14813
rect 16485 14773 16497 14807
rect 16531 14804 16543 14807
rect 16666 14804 16672 14816
rect 16531 14776 16672 14804
rect 16531 14773 16543 14776
rect 16485 14767 16543 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 18892 14804 18920 14980
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14909 19119 14943
rect 19061 14903 19119 14909
rect 19076 14872 19104 14903
rect 19242 14900 19248 14952
rect 19300 14900 19306 14952
rect 19720 14872 19748 14980
rect 20438 14968 20444 15020
rect 20496 15017 20502 15020
rect 20496 15011 20519 15017
rect 20507 14977 20519 15011
rect 20496 14971 20519 14977
rect 20496 14968 20502 14971
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21634 15008 21640 15020
rect 20772 14980 21640 15008
rect 20772 14968 20778 14980
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 22480 15017 22508 15116
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 26605 15147 26663 15153
rect 26605 15144 26617 15147
rect 23808 15116 26617 15144
rect 23808 15104 23814 15116
rect 26605 15113 26617 15116
rect 26651 15113 26663 15147
rect 26605 15107 26663 15113
rect 26050 15036 26056 15088
rect 26108 15036 26114 15088
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 23750 14968 23756 15020
rect 23808 14968 23814 15020
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24320 14980 24501 15008
rect 22278 14900 22284 14952
rect 22336 14940 22342 14952
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 22336 14912 22569 14940
rect 22336 14900 22342 14912
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 22738 14900 22744 14952
rect 22796 14900 22802 14952
rect 23290 14900 23296 14952
rect 23348 14940 23354 14952
rect 23658 14949 23664 14952
rect 23477 14943 23535 14949
rect 23477 14940 23489 14943
rect 23348 14912 23489 14940
rect 23348 14900 23354 14912
rect 23477 14909 23489 14912
rect 23523 14909 23535 14943
rect 23477 14903 23535 14909
rect 23615 14943 23664 14949
rect 23615 14909 23627 14943
rect 23661 14909 23664 14943
rect 23615 14903 23664 14909
rect 23658 14900 23664 14903
rect 23716 14900 23722 14952
rect 19076 14844 19380 14872
rect 19720 14844 19840 14872
rect 19352 14813 19380 14844
rect 17092 14776 18920 14804
rect 19337 14807 19395 14813
rect 17092 14764 17098 14776
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 19702 14804 19708 14816
rect 19383 14776 19708 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 19812 14804 19840 14844
rect 22646 14832 22652 14884
rect 22704 14872 22710 14884
rect 23201 14875 23259 14881
rect 23201 14872 23213 14875
rect 22704 14844 23213 14872
rect 22704 14832 22710 14844
rect 23201 14841 23213 14844
rect 23247 14841 23259 14875
rect 23201 14835 23259 14841
rect 23750 14804 23756 14816
rect 19812 14776 23756 14804
rect 23750 14764 23756 14776
rect 23808 14804 23814 14816
rect 24320 14804 24348 14980
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 24762 14968 24768 15020
rect 24820 15008 24826 15020
rect 25961 15011 26019 15017
rect 25961 15008 25973 15011
rect 24820 14980 25973 15008
rect 24820 14968 24826 14980
rect 25961 14977 25973 14980
rect 26007 14977 26019 15011
rect 26068 15008 26096 15036
rect 26068 14980 26188 15008
rect 25961 14971 26019 14977
rect 25222 14900 25228 14952
rect 25280 14940 25286 14952
rect 25317 14943 25375 14949
rect 25317 14940 25329 14943
rect 25280 14912 25329 14940
rect 25280 14900 25286 14912
rect 25317 14909 25329 14912
rect 25363 14909 25375 14943
rect 25317 14903 25375 14909
rect 25332 14872 25360 14903
rect 26050 14900 26056 14952
rect 26108 14900 26114 14952
rect 26160 14949 26188 14980
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14909 26203 14943
rect 26620 14940 26648 15107
rect 26694 15104 26700 15156
rect 26752 15144 26758 15156
rect 28905 15147 28963 15153
rect 28905 15144 28917 15147
rect 26752 15116 28917 15144
rect 26752 15104 26758 15116
rect 28905 15113 28917 15116
rect 28951 15113 28963 15147
rect 28905 15107 28963 15113
rect 30282 15104 30288 15156
rect 30340 15144 30346 15156
rect 31478 15144 31484 15156
rect 30340 15116 31484 15144
rect 30340 15104 30346 15116
rect 31478 15104 31484 15116
rect 31536 15104 31542 15156
rect 32125 15147 32183 15153
rect 32125 15113 32137 15147
rect 32171 15144 32183 15147
rect 32398 15144 32404 15156
rect 32171 15116 32404 15144
rect 32171 15113 32183 15116
rect 32125 15107 32183 15113
rect 32398 15104 32404 15116
rect 32456 15104 32462 15156
rect 32585 15147 32643 15153
rect 32585 15113 32597 15147
rect 32631 15144 32643 15147
rect 32858 15144 32864 15156
rect 32631 15116 32864 15144
rect 32631 15113 32643 15116
rect 32585 15107 32643 15113
rect 32858 15104 32864 15116
rect 32916 15104 32922 15156
rect 33321 15147 33379 15153
rect 33321 15113 33333 15147
rect 33367 15144 33379 15147
rect 33594 15144 33600 15156
rect 33367 15116 33600 15144
rect 33367 15113 33379 15116
rect 33321 15107 33379 15113
rect 33594 15104 33600 15116
rect 33652 15104 33658 15156
rect 33965 15147 34023 15153
rect 33965 15113 33977 15147
rect 34011 15144 34023 15147
rect 34238 15144 34244 15156
rect 34011 15116 34244 15144
rect 34011 15113 34023 15116
rect 33965 15107 34023 15113
rect 34238 15104 34244 15116
rect 34296 15104 34302 15156
rect 34422 15104 34428 15156
rect 34480 15144 34486 15156
rect 37366 15144 37372 15156
rect 34480 15116 37372 15144
rect 34480 15104 34486 15116
rect 37366 15104 37372 15116
rect 37424 15104 37430 15156
rect 38286 15104 38292 15156
rect 38344 15144 38350 15156
rect 38562 15144 38568 15156
rect 38344 15116 38568 15144
rect 38344 15104 38350 15116
rect 38562 15104 38568 15116
rect 38620 15104 38626 15156
rect 29546 15036 29552 15088
rect 29604 15076 29610 15088
rect 30193 15079 30251 15085
rect 30193 15076 30205 15079
rect 29604 15048 30205 15076
rect 29604 15036 29610 15048
rect 30193 15045 30205 15048
rect 30239 15045 30251 15079
rect 30193 15039 30251 15045
rect 27798 15017 27804 15020
rect 27776 15011 27804 15017
rect 27776 14977 27788 15011
rect 27776 14971 27804 14977
rect 27798 14968 27804 14971
rect 27856 14968 27862 15020
rect 29457 15011 29515 15017
rect 29457 15008 29469 15011
rect 28552 14980 29469 15008
rect 27062 14940 27068 14952
rect 26620 14912 27068 14940
rect 26145 14903 26203 14909
rect 27062 14900 27068 14912
rect 27120 14940 27126 14952
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 27120 14912 27629 14940
rect 27120 14900 27126 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 27893 14943 27951 14949
rect 27893 14909 27905 14943
rect 27939 14940 27951 14943
rect 28442 14940 28448 14952
rect 27939 14912 28448 14940
rect 27939 14909 27951 14912
rect 27893 14903 27951 14909
rect 28442 14900 28448 14912
rect 28500 14940 28506 14952
rect 28552 14940 28580 14980
rect 29457 14977 29469 14980
rect 29503 14977 29515 15011
rect 29457 14971 29515 14977
rect 32398 14968 32404 15020
rect 32456 15008 32462 15020
rect 32493 15011 32551 15017
rect 32493 15008 32505 15011
rect 32456 14980 32505 15008
rect 32456 14968 32462 14980
rect 32493 14977 32505 14980
rect 32539 15008 32551 15011
rect 33413 15011 33471 15017
rect 33413 15008 33425 15011
rect 32539 14980 33425 15008
rect 32539 14977 32551 14980
rect 32493 14971 32551 14977
rect 33413 14977 33425 14980
rect 33459 14977 33471 15011
rect 33413 14971 33471 14977
rect 33870 14968 33876 15020
rect 33928 14968 33934 15020
rect 28500 14912 28580 14940
rect 28500 14900 28506 14912
rect 28626 14900 28632 14952
rect 28684 14900 28690 14952
rect 28810 14900 28816 14952
rect 28868 14900 28874 14952
rect 32677 14943 32735 14949
rect 32677 14909 32689 14943
rect 32723 14909 32735 14943
rect 32677 14903 32735 14909
rect 33597 14943 33655 14949
rect 33597 14909 33609 14943
rect 33643 14940 33655 14943
rect 34440 14940 34468 15104
rect 33643 14912 34468 14940
rect 33643 14909 33655 14912
rect 33597 14903 33655 14909
rect 27154 14872 27160 14884
rect 25332 14844 27160 14872
rect 27154 14832 27160 14844
rect 27212 14832 27218 14884
rect 28169 14875 28227 14881
rect 28169 14841 28181 14875
rect 28215 14872 28227 14875
rect 31570 14872 31576 14884
rect 28215 14844 28994 14872
rect 28215 14841 28227 14844
rect 28169 14835 28227 14841
rect 23808 14776 24348 14804
rect 23808 14764 23814 14776
rect 24394 14764 24400 14816
rect 24452 14764 24458 14816
rect 24670 14764 24676 14816
rect 24728 14804 24734 14816
rect 25593 14807 25651 14813
rect 25593 14804 25605 14807
rect 24728 14776 25605 14804
rect 24728 14764 24734 14776
rect 25593 14773 25605 14776
rect 25639 14773 25651 14807
rect 25593 14767 25651 14773
rect 26973 14807 27031 14813
rect 26973 14773 26985 14807
rect 27019 14804 27031 14807
rect 27614 14804 27620 14816
rect 27019 14776 27620 14804
rect 27019 14773 27031 14776
rect 26973 14767 27031 14773
rect 27614 14764 27620 14776
rect 27672 14764 27678 14816
rect 28966 14804 28994 14844
rect 30668 14844 31576 14872
rect 30668 14816 30696 14844
rect 31570 14832 31576 14844
rect 31628 14832 31634 14884
rect 32692 14872 32720 14903
rect 34790 14900 34796 14952
rect 34848 14940 34854 14952
rect 35069 14943 35127 14949
rect 35069 14940 35081 14943
rect 34848 14912 35081 14940
rect 34848 14900 34854 14912
rect 35069 14909 35081 14912
rect 35115 14909 35127 14943
rect 35069 14903 35127 14909
rect 35894 14900 35900 14952
rect 35952 14900 35958 14952
rect 36538 14900 36544 14952
rect 36596 14900 36602 14952
rect 37918 14900 37924 14952
rect 37976 14900 37982 14952
rect 32766 14872 32772 14884
rect 32692 14844 32772 14872
rect 32766 14832 32772 14844
rect 32824 14832 32830 14884
rect 30101 14807 30159 14813
rect 30101 14804 30113 14807
rect 28966 14776 30113 14804
rect 30101 14773 30113 14776
rect 30147 14804 30159 14807
rect 30650 14804 30656 14816
rect 30147 14776 30656 14804
rect 30147 14773 30159 14776
rect 30101 14767 30159 14773
rect 30650 14764 30656 14776
rect 30708 14764 30714 14816
rect 31018 14764 31024 14816
rect 31076 14804 31082 14816
rect 31481 14807 31539 14813
rect 31481 14804 31493 14807
rect 31076 14776 31493 14804
rect 31076 14764 31082 14776
rect 31481 14773 31493 14776
rect 31527 14773 31539 14807
rect 31481 14767 31539 14773
rect 32582 14764 32588 14816
rect 32640 14804 32646 14816
rect 32953 14807 33011 14813
rect 32953 14804 32965 14807
rect 32640 14776 32965 14804
rect 32640 14764 32646 14776
rect 32953 14773 32965 14776
rect 32999 14773 33011 14807
rect 32953 14767 33011 14773
rect 34514 14764 34520 14816
rect 34572 14764 34578 14816
rect 35253 14807 35311 14813
rect 35253 14773 35265 14807
rect 35299 14804 35311 14807
rect 35342 14804 35348 14816
rect 35299 14776 35348 14804
rect 35299 14773 35311 14776
rect 35253 14767 35311 14773
rect 35342 14764 35348 14776
rect 35400 14764 35406 14816
rect 37093 14807 37151 14813
rect 37093 14773 37105 14807
rect 37139 14804 37151 14807
rect 37182 14804 37188 14816
rect 37139 14776 37188 14804
rect 37139 14773 37151 14776
rect 37093 14767 37151 14773
rect 37182 14764 37188 14776
rect 37240 14764 37246 14816
rect 37274 14764 37280 14816
rect 37332 14764 37338 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1946 14560 1952 14612
rect 2004 14560 2010 14612
rect 3602 14560 3608 14612
rect 3660 14560 3666 14612
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 4614 14600 4620 14612
rect 4203 14572 4620 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 7432 14572 7573 14600
rect 7432 14560 7438 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 7561 14563 7619 14569
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 1964 14464 1992 14560
rect 1627 14436 1992 14464
rect 7576 14464 7604 14563
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 8757 14603 8815 14609
rect 8757 14600 8769 14603
rect 8536 14572 8769 14600
rect 8536 14560 8542 14572
rect 8757 14569 8769 14572
rect 8803 14569 8815 14603
rect 8757 14563 8815 14569
rect 9030 14560 9036 14612
rect 9088 14560 9094 14612
rect 11330 14600 11336 14612
rect 10336 14572 11336 14600
rect 8113 14467 8171 14473
rect 8113 14464 8125 14467
rect 7576 14436 8125 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 8113 14433 8125 14436
rect 8159 14433 8171 14467
rect 8113 14427 8171 14433
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2774 14396 2780 14408
rect 2271 14368 2780 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2774 14356 2780 14368
rect 2832 14396 2838 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 2832 14368 5825 14396
rect 2832 14356 2838 14368
rect 5813 14365 5825 14368
rect 5859 14396 5871 14399
rect 6178 14396 6184 14408
rect 5859 14368 6184 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 6448 14399 6506 14405
rect 6448 14365 6460 14399
rect 6494 14396 6506 14399
rect 9048 14396 9076 14560
rect 6494 14368 9076 14396
rect 6494 14365 6506 14368
rect 6448 14359 6506 14365
rect 10134 14356 10140 14408
rect 10192 14396 10198 14408
rect 10336 14405 10364 14572
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 11793 14603 11851 14609
rect 11793 14569 11805 14603
rect 11839 14600 11851 14603
rect 13354 14600 13360 14612
rect 11839 14572 13360 14600
rect 11839 14569 11851 14572
rect 11793 14563 11851 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 15286 14560 15292 14612
rect 15344 14560 15350 14612
rect 17681 14603 17739 14609
rect 16224 14572 17172 14600
rect 15197 14535 15255 14541
rect 15197 14501 15209 14535
rect 15243 14532 15255 14535
rect 15304 14532 15332 14560
rect 15243 14504 15332 14532
rect 15243 14501 15255 14504
rect 15197 14495 15255 14501
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12437 14467 12495 14473
rect 12437 14464 12449 14467
rect 12308 14436 12449 14464
rect 12308 14424 12314 14436
rect 12437 14433 12449 14436
rect 12483 14433 12495 14467
rect 12437 14427 12495 14433
rect 12710 14424 12716 14476
rect 12768 14424 12774 14476
rect 12986 14424 12992 14476
rect 13044 14424 13050 14476
rect 14090 14424 14096 14476
rect 14148 14464 14154 14476
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14148 14436 14749 14464
rect 14148 14424 14154 14436
rect 14737 14433 14749 14436
rect 14783 14464 14795 14467
rect 15562 14464 15568 14476
rect 14783 14436 15568 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 15562 14424 15568 14436
rect 15620 14464 15626 14476
rect 16224 14464 16252 14572
rect 17144 14532 17172 14572
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 18138 14600 18144 14612
rect 17727 14572 18144 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 18138 14560 18144 14572
rect 18196 14600 18202 14612
rect 19242 14600 19248 14612
rect 18196 14572 19248 14600
rect 18196 14560 18202 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 20070 14560 20076 14612
rect 20128 14600 20134 14612
rect 20128 14572 23704 14600
rect 20128 14560 20134 14572
rect 20714 14532 20720 14544
rect 17144 14504 17724 14532
rect 15620 14436 16252 14464
rect 15620 14424 15626 14436
rect 12618 14405 12624 14408
rect 10321 14399 10379 14405
rect 10321 14396 10333 14399
rect 10192 14368 10333 14396
rect 10192 14356 10198 14368
rect 10321 14365 10333 14368
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 12575 14399 12624 14405
rect 12575 14365 12587 14399
rect 12621 14365 12624 14399
rect 12575 14359 12624 14365
rect 12618 14356 12624 14359
rect 12676 14356 12682 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 13596 14368 13645 14396
rect 13596 14356 13602 14368
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 13633 14359 13691 14365
rect 13740 14368 14565 14396
rect 2133 14331 2191 14337
rect 2133 14297 2145 14331
rect 2179 14328 2191 14331
rect 2470 14331 2528 14337
rect 2470 14328 2482 14331
rect 2179 14300 2482 14328
rect 2179 14297 2191 14300
rect 2133 14291 2191 14297
rect 2470 14297 2482 14300
rect 2516 14297 2528 14331
rect 2470 14291 2528 14297
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 7006 14328 7012 14340
rect 4295 14300 7012 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 7006 14288 7012 14300
rect 7064 14288 7070 14340
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 9122 14328 9128 14340
rect 8628 14300 9128 14328
rect 8628 14288 8634 14300
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 10588 14331 10646 14337
rect 10588 14297 10600 14331
rect 10634 14328 10646 14331
rect 11422 14328 11428 14340
rect 10634 14300 11428 14328
rect 10634 14297 10646 14300
rect 10588 14291 10646 14297
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 13740 14328 13768 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16298 14396 16304 14408
rect 16255 14368 16304 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17586 14396 17592 14408
rect 17460 14368 17592 14396
rect 17460 14356 17466 14368
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 17696 14396 17724 14504
rect 19076 14504 20720 14532
rect 19076 14473 19104 14504
rect 20714 14492 20720 14504
rect 20772 14492 20778 14544
rect 23676 14532 23704 14572
rect 23750 14560 23756 14612
rect 23808 14600 23814 14612
rect 24121 14603 24179 14609
rect 24121 14600 24133 14603
rect 23808 14572 24133 14600
rect 23808 14560 23814 14572
rect 24121 14569 24133 14572
rect 24167 14569 24179 14603
rect 24121 14563 24179 14569
rect 24302 14560 24308 14612
rect 24360 14600 24366 14612
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 24360 14572 24409 14600
rect 24360 14560 24366 14572
rect 24397 14569 24409 14572
rect 24443 14569 24455 14603
rect 27893 14603 27951 14609
rect 24397 14563 24455 14569
rect 26528 14572 27844 14600
rect 26528 14532 26556 14572
rect 23676 14504 26556 14532
rect 19061 14467 19119 14473
rect 19061 14433 19073 14467
rect 19107 14433 19119 14467
rect 19061 14427 19119 14433
rect 19429 14467 19487 14473
rect 19429 14433 19441 14467
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 19444 14396 19472 14427
rect 19518 14424 19524 14476
rect 19576 14424 19582 14476
rect 19702 14424 19708 14476
rect 19760 14464 19766 14476
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 19760 14436 20637 14464
rect 19760 14424 19766 14436
rect 20625 14433 20637 14436
rect 20671 14433 20683 14467
rect 20625 14427 20683 14433
rect 23842 14424 23848 14476
rect 23900 14464 23906 14476
rect 24949 14467 25007 14473
rect 24949 14464 24961 14467
rect 23900 14436 24961 14464
rect 23900 14424 23906 14436
rect 24949 14433 24961 14436
rect 24995 14433 25007 14467
rect 24949 14427 25007 14433
rect 25682 14424 25688 14476
rect 25740 14464 25746 14476
rect 25777 14467 25835 14473
rect 25777 14464 25789 14467
rect 25740 14436 25789 14464
rect 25740 14424 25746 14436
rect 25777 14433 25789 14436
rect 25823 14433 25835 14467
rect 25777 14427 25835 14433
rect 26234 14424 26240 14476
rect 26292 14464 26298 14476
rect 26513 14467 26571 14473
rect 26513 14464 26525 14467
rect 26292 14436 26525 14464
rect 26292 14424 26298 14436
rect 26513 14433 26525 14436
rect 26559 14433 26571 14467
rect 26513 14427 26571 14433
rect 23661 14399 23719 14405
rect 23661 14396 23673 14399
rect 17696 14368 20208 14396
rect 13464 14300 13768 14328
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 11238 14260 11244 14272
rect 8260 14232 11244 14260
rect 8260 14220 8266 14232
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12710 14260 12716 14272
rect 11747 14232 12716 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13464 14260 13492 14300
rect 14182 14288 14188 14340
rect 14240 14328 14246 14340
rect 16482 14337 16488 14340
rect 15013 14331 15071 14337
rect 15013 14328 15025 14331
rect 14240 14300 15025 14328
rect 14240 14288 14246 14300
rect 15013 14297 15025 14300
rect 15059 14297 15071 14331
rect 15013 14291 15071 14297
rect 16476 14291 16488 14337
rect 16482 14288 16488 14291
rect 16540 14288 16546 14340
rect 18782 14288 18788 14340
rect 18840 14337 18846 14340
rect 18840 14291 18852 14337
rect 18840 14288 18846 14291
rect 20180 14272 20208 14368
rect 23308 14368 23673 14396
rect 23308 14340 23336 14368
rect 23661 14365 23673 14368
rect 23707 14365 23719 14399
rect 27522 14396 27528 14408
rect 23661 14359 23719 14365
rect 24136 14368 27528 14396
rect 23290 14288 23296 14340
rect 23348 14288 23354 14340
rect 23416 14331 23474 14337
rect 23416 14297 23428 14331
rect 23462 14328 23474 14331
rect 24026 14328 24032 14340
rect 23462 14300 24032 14328
rect 23462 14297 23474 14300
rect 23416 14291 23474 14297
rect 24026 14288 24032 14300
rect 24084 14288 24090 14340
rect 12860 14232 13492 14260
rect 12860 14220 12866 14232
rect 14090 14220 14096 14272
rect 14148 14220 14154 14272
rect 14458 14220 14464 14272
rect 14516 14220 14522 14272
rect 17589 14263 17647 14269
rect 17589 14229 17601 14263
rect 17635 14260 17647 14263
rect 18506 14260 18512 14272
rect 17635 14232 18512 14260
rect 17635 14229 17647 14232
rect 17589 14223 17647 14229
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19659 14232 20085 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 20073 14229 20085 14232
rect 20119 14229 20131 14263
rect 20073 14223 20131 14229
rect 20162 14220 20168 14272
rect 20220 14220 20226 14272
rect 22278 14220 22284 14272
rect 22336 14220 22342 14272
rect 22738 14220 22744 14272
rect 22796 14260 22802 14272
rect 24136 14260 24164 14368
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 27816 14396 27844 14572
rect 27893 14569 27905 14603
rect 27939 14569 27951 14603
rect 27893 14563 27951 14569
rect 27908 14532 27936 14563
rect 28074 14560 28080 14612
rect 28132 14600 28138 14612
rect 28721 14603 28779 14609
rect 28721 14600 28733 14603
rect 28132 14572 28733 14600
rect 28132 14560 28138 14572
rect 28721 14569 28733 14572
rect 28767 14569 28779 14603
rect 30742 14600 30748 14612
rect 28721 14563 28779 14569
rect 29472 14572 30748 14600
rect 28626 14532 28632 14544
rect 27908 14504 28632 14532
rect 28626 14492 28632 14504
rect 28684 14532 28690 14544
rect 28684 14504 29316 14532
rect 28684 14492 28690 14504
rect 27982 14424 27988 14476
rect 28040 14464 28046 14476
rect 29288 14473 29316 14504
rect 28537 14467 28595 14473
rect 28537 14464 28549 14467
rect 28040 14436 28549 14464
rect 28040 14424 28046 14436
rect 28537 14433 28549 14436
rect 28583 14433 28595 14467
rect 28537 14427 28595 14433
rect 29273 14467 29331 14473
rect 29273 14433 29285 14467
rect 29319 14433 29331 14467
rect 29273 14427 29331 14433
rect 29472 14396 29500 14572
rect 30742 14560 30748 14572
rect 30800 14560 30806 14612
rect 30929 14603 30987 14609
rect 30929 14569 30941 14603
rect 30975 14600 30987 14603
rect 31202 14600 31208 14612
rect 30975 14572 31208 14600
rect 30975 14569 30987 14572
rect 30929 14563 30987 14569
rect 31202 14560 31208 14572
rect 31260 14560 31266 14612
rect 32306 14560 32312 14612
rect 32364 14600 32370 14612
rect 32401 14603 32459 14609
rect 32401 14600 32413 14603
rect 32364 14572 32413 14600
rect 32364 14560 32370 14572
rect 32401 14569 32413 14572
rect 32447 14569 32459 14603
rect 32401 14563 32459 14569
rect 32416 14532 32444 14563
rect 33226 14560 33232 14612
rect 33284 14560 33290 14612
rect 34790 14560 34796 14612
rect 34848 14560 34854 14612
rect 35342 14560 35348 14612
rect 35400 14560 35406 14612
rect 36538 14560 36544 14612
rect 36596 14600 36602 14612
rect 37001 14603 37059 14609
rect 37001 14600 37013 14603
rect 36596 14572 37013 14600
rect 36596 14560 36602 14572
rect 37001 14569 37013 14572
rect 37047 14569 37059 14603
rect 37001 14563 37059 14569
rect 37274 14560 37280 14612
rect 37332 14560 37338 14612
rect 37366 14560 37372 14612
rect 37424 14560 37430 14612
rect 35360 14532 35388 14560
rect 37292 14532 37320 14560
rect 32416 14504 33824 14532
rect 33134 14424 33140 14476
rect 33192 14424 33198 14476
rect 33796 14473 33824 14504
rect 35176 14504 35388 14532
rect 36648 14504 37320 14532
rect 37384 14532 37412 14560
rect 38105 14535 38163 14541
rect 38105 14532 38117 14535
rect 37384 14504 38117 14532
rect 33781 14467 33839 14473
rect 33781 14433 33793 14467
rect 33827 14433 33839 14467
rect 33781 14427 33839 14433
rect 27816 14368 29500 14396
rect 29549 14399 29607 14405
rect 29549 14365 29561 14399
rect 29595 14396 29607 14399
rect 31018 14396 31024 14408
rect 29595 14368 31024 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 24762 14328 24768 14340
rect 24228 14300 24768 14328
rect 24228 14272 24256 14300
rect 24762 14288 24768 14300
rect 24820 14328 24826 14340
rect 25593 14331 25651 14337
rect 24820 14300 25360 14328
rect 24820 14288 24826 14300
rect 22796 14232 24164 14260
rect 22796 14220 22802 14232
rect 24210 14220 24216 14272
rect 24268 14220 24274 14272
rect 25222 14220 25228 14272
rect 25280 14220 25286 14272
rect 25332 14260 25360 14300
rect 25593 14297 25605 14331
rect 25639 14328 25651 14331
rect 26780 14331 26838 14337
rect 25639 14300 26740 14328
rect 25639 14297 25651 14300
rect 25593 14291 25651 14297
rect 25685 14263 25743 14269
rect 25685 14260 25697 14263
rect 25332 14232 25697 14260
rect 25685 14229 25697 14232
rect 25731 14229 25743 14263
rect 25685 14223 25743 14229
rect 26326 14220 26332 14272
rect 26384 14220 26390 14272
rect 26712 14260 26740 14300
rect 26780 14297 26792 14331
rect 26826 14328 26838 14331
rect 27985 14331 28043 14337
rect 27985 14328 27997 14331
rect 26826 14300 27997 14328
rect 26826 14297 26838 14300
rect 26780 14291 26838 14297
rect 27985 14297 27997 14300
rect 28031 14297 28043 14331
rect 27985 14291 28043 14297
rect 29748 14272 29776 14368
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 35176 14405 35204 14504
rect 35345 14467 35403 14473
rect 35345 14464 35357 14467
rect 35268 14436 35357 14464
rect 35161 14399 35219 14405
rect 35161 14365 35173 14399
rect 35207 14365 35219 14399
rect 35161 14359 35219 14365
rect 29816 14331 29874 14337
rect 29816 14297 29828 14331
rect 29862 14328 29874 14331
rect 30098 14328 30104 14340
rect 29862 14300 30104 14328
rect 29862 14297 29874 14300
rect 29816 14291 29874 14297
rect 30098 14288 30104 14300
rect 30156 14288 30162 14340
rect 31288 14331 31346 14337
rect 31288 14297 31300 14331
rect 31334 14328 31346 14331
rect 32493 14331 32551 14337
rect 32493 14328 32505 14331
rect 31334 14300 32505 14328
rect 31334 14297 31346 14300
rect 31288 14291 31346 14297
rect 32493 14297 32505 14300
rect 32539 14297 32551 14331
rect 35268 14328 35296 14436
rect 35345 14433 35357 14436
rect 35391 14433 35403 14467
rect 35345 14427 35403 14433
rect 35621 14399 35679 14405
rect 35621 14365 35633 14399
rect 35667 14396 35679 14399
rect 36170 14396 36176 14408
rect 35667 14368 36176 14396
rect 35667 14365 35679 14368
rect 35621 14359 35679 14365
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 32493 14291 32551 14297
rect 34440 14300 35296 14328
rect 35888 14331 35946 14337
rect 26970 14260 26976 14272
rect 26712 14232 26976 14260
rect 26970 14220 26976 14232
rect 27028 14220 27034 14272
rect 29730 14220 29736 14272
rect 29788 14220 29794 14272
rect 31478 14220 31484 14272
rect 31536 14260 31542 14272
rect 33778 14260 33784 14272
rect 31536 14232 33784 14260
rect 31536 14220 31542 14232
rect 33778 14220 33784 14232
rect 33836 14260 33842 14272
rect 34440 14269 34468 14300
rect 35888 14297 35900 14331
rect 35934 14328 35946 14331
rect 36648 14328 36676 14504
rect 37660 14473 37688 14504
rect 38105 14501 38117 14504
rect 38151 14532 38163 14535
rect 38286 14532 38292 14544
rect 38151 14504 38292 14532
rect 38151 14501 38163 14504
rect 38105 14495 38163 14501
rect 38286 14492 38292 14504
rect 38344 14492 38350 14544
rect 37645 14467 37703 14473
rect 37645 14433 37657 14467
rect 37691 14433 37703 14467
rect 37645 14427 37703 14433
rect 37461 14399 37519 14405
rect 37461 14365 37473 14399
rect 37507 14396 37519 14399
rect 37826 14396 37832 14408
rect 37507 14368 37832 14396
rect 37507 14365 37519 14368
rect 37461 14359 37519 14365
rect 37826 14356 37832 14368
rect 37884 14356 37890 14408
rect 37553 14331 37611 14337
rect 37553 14328 37565 14331
rect 35934 14300 36676 14328
rect 37016 14300 37565 14328
rect 35934 14297 35946 14300
rect 35888 14291 35946 14297
rect 34425 14263 34483 14269
rect 34425 14260 34437 14263
rect 33836 14232 34437 14260
rect 33836 14220 33842 14232
rect 34425 14229 34437 14232
rect 34471 14229 34483 14263
rect 34425 14223 34483 14229
rect 35253 14263 35311 14269
rect 35253 14229 35265 14263
rect 35299 14260 35311 14263
rect 37016 14260 37044 14300
rect 37553 14297 37565 14300
rect 37599 14328 37611 14331
rect 37642 14328 37648 14340
rect 37599 14300 37648 14328
rect 37599 14297 37611 14300
rect 37553 14291 37611 14297
rect 37642 14288 37648 14300
rect 37700 14288 37706 14340
rect 35299 14232 37044 14260
rect 37093 14263 37151 14269
rect 35299 14229 35311 14232
rect 35253 14223 35311 14229
rect 37093 14229 37105 14263
rect 37139 14260 37151 14263
rect 37366 14260 37372 14272
rect 37139 14232 37372 14260
rect 37139 14229 37151 14232
rect 37093 14223 37151 14229
rect 37366 14220 37372 14232
rect 37424 14220 37430 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 2685 14059 2743 14065
rect 2685 14056 2697 14059
rect 1728 14028 2697 14056
rect 1728 14016 1734 14028
rect 2685 14025 2697 14028
rect 2731 14025 2743 14059
rect 2685 14019 2743 14025
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6638 14056 6644 14068
rect 6052 14028 6644 14056
rect 6052 14016 6058 14028
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 9456 14028 11744 14056
rect 9456 14016 9462 14028
rect 1578 13948 1584 14000
rect 1636 13988 1642 14000
rect 2225 13991 2283 13997
rect 2225 13988 2237 13991
rect 1636 13960 2237 13988
rect 1636 13948 1642 13960
rect 2225 13957 2237 13960
rect 2271 13957 2283 13991
rect 2225 13951 2283 13957
rect 7006 13948 7012 14000
rect 7064 13988 7070 14000
rect 8294 13988 8300 14000
rect 7064 13960 8300 13988
rect 7064 13948 7070 13960
rect 8294 13948 8300 13960
rect 8352 13988 8358 14000
rect 11716 13988 11744 14028
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12526 14056 12532 14068
rect 12032 14028 12532 14056
rect 12032 14016 12038 14028
rect 12526 14016 12532 14028
rect 12584 14056 12590 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12584 14028 12909 14056
rect 12584 14016 12590 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 14090 14016 14096 14068
rect 14148 14016 14154 14068
rect 16666 14016 16672 14068
rect 16724 14016 16730 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 17920 14028 18061 14056
rect 17920 14016 17926 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 18138 14016 18144 14068
rect 18196 14016 18202 14068
rect 18782 14016 18788 14068
rect 18840 14056 18846 14068
rect 18877 14059 18935 14065
rect 18877 14056 18889 14059
rect 18840 14028 18889 14056
rect 18840 14016 18846 14028
rect 18877 14025 18889 14028
rect 18923 14025 18935 14059
rect 18877 14019 18935 14025
rect 20070 14016 20076 14068
rect 20128 14016 20134 14068
rect 20162 14016 20168 14068
rect 20220 14056 20226 14068
rect 23934 14056 23940 14068
rect 20220 14028 23940 14056
rect 20220 14016 20226 14028
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 24026 14016 24032 14068
rect 24084 14016 24090 14068
rect 24670 14016 24676 14068
rect 24728 14016 24734 14068
rect 24946 14016 24952 14068
rect 25004 14016 25010 14068
rect 25222 14016 25228 14068
rect 25280 14016 25286 14068
rect 25958 14016 25964 14068
rect 26016 14016 26022 14068
rect 26329 14059 26387 14065
rect 26329 14025 26341 14059
rect 26375 14056 26387 14059
rect 26694 14056 26700 14068
rect 26375 14028 26700 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 26694 14016 26700 14028
rect 26752 14016 26758 14068
rect 26789 14059 26847 14065
rect 26789 14025 26801 14059
rect 26835 14025 26847 14059
rect 26789 14019 26847 14025
rect 8352 13960 11652 13988
rect 11716 13960 14044 13988
rect 8352 13948 8358 13960
rect 3326 13880 3332 13932
rect 3384 13880 3390 13932
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3476 13892 3709 13920
rect 3476 13880 3482 13892
rect 3697 13889 3709 13892
rect 3743 13920 3755 13923
rect 3970 13920 3976 13932
rect 3743 13892 3976 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 8205 13923 8263 13929
rect 8205 13889 8217 13923
rect 8251 13920 8263 13923
rect 9769 13923 9827 13929
rect 8251 13892 9536 13920
rect 8251 13889 8263 13892
rect 8205 13883 8263 13889
rect 9508 13864 9536 13892
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10410 13920 10416 13932
rect 9815 13892 10416 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 3016 13824 4537 13852
rect 3016 13812 3022 13824
rect 4525 13821 4537 13824
rect 4571 13852 4583 13855
rect 4571 13824 6675 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4614 13744 4620 13796
rect 4672 13784 4678 13796
rect 5074 13784 5080 13796
rect 4672 13756 5080 13784
rect 4672 13744 4678 13756
rect 5074 13744 5080 13756
rect 5132 13744 5138 13796
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 6086 13716 6092 13728
rect 5684 13688 6092 13716
rect 5684 13676 5690 13688
rect 6086 13676 6092 13688
rect 6144 13716 6150 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6144 13688 6561 13716
rect 6144 13676 6150 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6647 13716 6675 13824
rect 7926 13812 7932 13864
rect 7984 13852 7990 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 7984 13824 8401 13852
rect 7984 13812 7990 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9490 13812 9496 13864
rect 9548 13812 9554 13864
rect 7834 13744 7840 13796
rect 7892 13784 7898 13796
rect 9784 13784 9812 13883
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 11624 13929 11652 13960
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10551 13892 10977 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 11609 13923 11667 13929
rect 11103 13892 11560 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 9999 13824 10364 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 7892 13756 9812 13784
rect 7892 13744 7898 13756
rect 9214 13716 9220 13728
rect 6647 13688 9220 13716
rect 6549 13679 6607 13685
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9398 13676 9404 13728
rect 9456 13676 9462 13728
rect 10336 13716 10364 13824
rect 10980 13824 11161 13852
rect 10980 13796 11008 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11532 13852 11560 13892
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 11790 13920 11796 13932
rect 11655 13892 11796 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 12802 13920 12808 13932
rect 12406 13892 12808 13920
rect 12406 13852 12434 13892
rect 12544 13864 12572 13892
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 11532 13824 12434 13852
rect 11149 13815 11207 13821
rect 12526 13812 12532 13864
rect 12584 13812 12590 13864
rect 14016 13852 14044 13960
rect 14108 13920 14136 14016
rect 14274 13948 14280 14000
rect 14332 13988 14338 14000
rect 14737 13991 14795 13997
rect 14737 13988 14749 13991
rect 14332 13960 14749 13988
rect 14332 13948 14338 13960
rect 14737 13957 14749 13960
rect 14783 13957 14795 13991
rect 16684 13988 16712 14016
rect 16914 13991 16972 13997
rect 16914 13988 16926 13991
rect 16684 13960 16926 13988
rect 14737 13951 14795 13957
rect 16914 13957 16926 13960
rect 16960 13957 16972 13991
rect 16914 13951 16972 13957
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 14108 13892 14197 13920
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 18156 13929 18184 14016
rect 20088 13988 20116 14016
rect 18248 13960 20116 13988
rect 18141 13923 18199 13929
rect 15028 13892 17724 13920
rect 15028 13852 15056 13892
rect 14016 13824 15056 13852
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 16666 13852 16672 13864
rect 16356 13824 16672 13852
rect 16356 13812 16362 13824
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 17696 13852 17724 13892
rect 18141 13889 18153 13923
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 18248 13852 18276 13960
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19392 13892 19441 13920
rect 19392 13880 19398 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20180 13920 20208 14016
rect 22186 13948 22192 14000
rect 22244 13948 22250 14000
rect 23477 13991 23535 13997
rect 23477 13957 23489 13991
rect 23523 13988 23535 13991
rect 23658 13988 23664 14000
rect 23523 13960 23664 13988
rect 23523 13957 23535 13960
rect 23477 13951 23535 13957
rect 23658 13948 23664 13960
rect 23716 13988 23722 14000
rect 24210 13988 24216 14000
rect 23716 13960 24216 13988
rect 23716 13948 23722 13960
rect 24210 13948 24216 13960
rect 24268 13948 24274 14000
rect 22097 13923 22155 13929
rect 22097 13920 22109 13923
rect 19935 13892 20208 13920
rect 21560 13892 22109 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 17696 13824 18276 13852
rect 18414 13812 18420 13864
rect 18472 13852 18478 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18472 13824 18797 13852
rect 18472 13812 18478 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 21560 13861 21588 13892
rect 22097 13889 22109 13892
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 21545 13855 21603 13861
rect 21545 13852 21557 13855
rect 20772 13824 21557 13852
rect 20772 13812 20778 13824
rect 21545 13821 21557 13824
rect 21591 13821 21603 13855
rect 21545 13815 21603 13821
rect 21726 13812 21732 13864
rect 21784 13852 21790 13864
rect 22204 13852 22232 13948
rect 23566 13880 23572 13932
rect 23624 13880 23630 13932
rect 24688 13929 24716 14016
rect 24673 13923 24731 13929
rect 24673 13889 24685 13923
rect 24719 13889 24731 13923
rect 25240 13920 25268 14016
rect 25501 13923 25559 13929
rect 25501 13920 25513 13923
rect 25240 13892 25513 13920
rect 24673 13883 24731 13889
rect 25501 13889 25513 13892
rect 25547 13889 25559 13923
rect 25501 13883 25559 13889
rect 26418 13880 26424 13932
rect 26476 13880 26482 13932
rect 26804 13920 26832 14019
rect 26970 14016 26976 14068
rect 27028 14016 27034 14068
rect 27706 14016 27712 14068
rect 27764 14016 27770 14068
rect 29546 14016 29552 14068
rect 29604 14016 29610 14068
rect 30098 14016 30104 14068
rect 30156 14056 30162 14068
rect 30377 14059 30435 14065
rect 30377 14056 30389 14059
rect 30156 14028 30389 14056
rect 30156 14016 30162 14028
rect 30377 14025 30389 14028
rect 30423 14025 30435 14059
rect 30377 14019 30435 14025
rect 30558 14016 30564 14068
rect 30616 14016 30622 14068
rect 32401 14059 32459 14065
rect 32401 14025 32413 14059
rect 32447 14056 32459 14059
rect 32766 14056 32772 14068
rect 32447 14028 32772 14056
rect 32447 14025 32459 14028
rect 32401 14019 32459 14025
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 35161 14059 35219 14065
rect 35161 14025 35173 14059
rect 35207 14056 35219 14059
rect 35894 14056 35900 14068
rect 35207 14028 35900 14056
rect 35207 14025 35219 14028
rect 35161 14019 35219 14025
rect 35894 14016 35900 14028
rect 35952 14016 35958 14068
rect 36538 14016 36544 14068
rect 36596 14056 36602 14068
rect 36596 14028 37136 14056
rect 36596 14016 36602 14028
rect 27430 13948 27436 14000
rect 27488 13988 27494 14000
rect 30282 13988 30288 14000
rect 27488 13960 30288 13988
rect 27488 13948 27494 13960
rect 30282 13948 30288 13960
rect 30340 13948 30346 14000
rect 33796 13960 34836 13988
rect 28261 13923 28319 13929
rect 28261 13920 28273 13923
rect 26804 13892 28273 13920
rect 28261 13889 28273 13892
rect 28307 13889 28319 13923
rect 28261 13883 28319 13889
rect 29825 13923 29883 13929
rect 29825 13889 29837 13923
rect 29871 13920 29883 13923
rect 29914 13920 29920 13932
rect 29871 13892 29920 13920
rect 29871 13889 29883 13892
rect 29825 13883 29883 13889
rect 29914 13880 29920 13892
rect 29972 13880 29978 13932
rect 31202 13880 31208 13932
rect 31260 13880 31266 13932
rect 33796 13929 33824 13960
rect 33781 13923 33839 13929
rect 33781 13889 33793 13923
rect 33827 13889 33839 13923
rect 33781 13883 33839 13889
rect 34048 13923 34106 13929
rect 34048 13889 34060 13923
rect 34094 13920 34106 13923
rect 34514 13920 34520 13932
rect 34094 13892 34520 13920
rect 34094 13889 34106 13892
rect 34048 13883 34106 13889
rect 34514 13880 34520 13892
rect 34572 13880 34578 13932
rect 22465 13855 22523 13861
rect 22465 13852 22477 13855
rect 21784 13824 22477 13852
rect 21784 13812 21790 13824
rect 22465 13821 22477 13824
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 23385 13855 23443 13861
rect 23385 13821 23397 13855
rect 23431 13821 23443 13855
rect 25682 13852 25688 13864
rect 23385 13815 23443 13821
rect 23952 13824 25688 13852
rect 10410 13744 10416 13796
rect 10468 13784 10474 13796
rect 10962 13784 10968 13796
rect 10468 13756 10968 13784
rect 10468 13744 10474 13756
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 23400 13784 23428 13815
rect 23474 13784 23480 13796
rect 23400 13756 23480 13784
rect 23474 13744 23480 13756
rect 23532 13784 23538 13796
rect 23842 13784 23848 13796
rect 23532 13756 23848 13784
rect 23532 13744 23538 13756
rect 23842 13744 23848 13756
rect 23900 13744 23906 13796
rect 23952 13793 23980 13824
rect 25682 13812 25688 13824
rect 25740 13812 25746 13864
rect 26237 13855 26295 13861
rect 26237 13821 26249 13855
rect 26283 13821 26295 13855
rect 26436 13852 26464 13880
rect 34808 13864 34836 13960
rect 35986 13880 35992 13932
rect 36044 13929 36050 13932
rect 37108 13929 37136 14028
rect 37182 14016 37188 14068
rect 37240 14056 37246 14068
rect 37553 14059 37611 14065
rect 37553 14056 37565 14059
rect 37240 14028 37565 14056
rect 37240 14016 37246 14028
rect 37553 14025 37565 14028
rect 37599 14025 37611 14059
rect 37553 14019 37611 14025
rect 37642 14016 37648 14068
rect 37700 14016 37706 14068
rect 37918 14016 37924 14068
rect 37976 14056 37982 14068
rect 38013 14059 38071 14065
rect 38013 14056 38025 14059
rect 37976 14028 38025 14056
rect 37976 14016 37982 14028
rect 38013 14025 38025 14028
rect 38059 14025 38071 14059
rect 38013 14019 38071 14025
rect 37660 13932 37688 14016
rect 36044 13923 36093 13929
rect 36044 13889 36047 13923
rect 36081 13889 36093 13923
rect 36044 13883 36093 13889
rect 37093 13923 37151 13929
rect 37093 13889 37105 13923
rect 37139 13889 37151 13923
rect 37093 13883 37151 13889
rect 36044 13880 36050 13883
rect 37642 13880 37648 13932
rect 37700 13880 37706 13932
rect 27430 13852 27436 13864
rect 26436 13824 27436 13852
rect 26237 13815 26295 13821
rect 23937 13787 23995 13793
rect 23937 13753 23949 13787
rect 23983 13753 23995 13787
rect 23937 13747 23995 13753
rect 24302 13744 24308 13796
rect 24360 13784 24366 13796
rect 24578 13784 24584 13796
rect 24360 13756 24584 13784
rect 24360 13744 24366 13756
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 26252 13784 26280 13815
rect 27430 13812 27436 13824
rect 27488 13812 27494 13864
rect 27522 13812 27528 13864
rect 27580 13812 27586 13864
rect 34790 13812 34796 13864
rect 34848 13812 34854 13864
rect 35897 13855 35955 13861
rect 35897 13852 35909 13855
rect 34900 13824 35909 13852
rect 26510 13784 26516 13796
rect 26252 13756 26516 13784
rect 26510 13744 26516 13756
rect 26568 13744 26574 13796
rect 10502 13716 10508 13728
rect 10336 13688 10508 13716
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 10594 13676 10600 13728
rect 10652 13676 10658 13728
rect 13630 13676 13636 13728
rect 13688 13676 13694 13728
rect 30466 13676 30472 13728
rect 30524 13716 30530 13728
rect 30926 13716 30932 13728
rect 30524 13688 30932 13716
rect 30524 13676 30530 13688
rect 30926 13676 30932 13688
rect 30984 13716 30990 13728
rect 33597 13719 33655 13725
rect 33597 13716 33609 13719
rect 30984 13688 33609 13716
rect 30984 13676 30990 13688
rect 33597 13685 33609 13688
rect 33643 13716 33655 13719
rect 34900 13716 34928 13824
rect 35897 13821 35909 13824
rect 35943 13821 35955 13855
rect 35897 13815 35955 13821
rect 36173 13855 36231 13861
rect 36173 13821 36185 13855
rect 36219 13852 36231 13855
rect 36354 13852 36360 13864
rect 36219 13824 36360 13852
rect 36219 13821 36231 13824
rect 36173 13815 36231 13821
rect 36354 13812 36360 13824
rect 36412 13812 36418 13864
rect 36909 13855 36967 13861
rect 36909 13821 36921 13855
rect 36955 13852 36967 13855
rect 37461 13855 37519 13861
rect 36955 13824 37320 13852
rect 36955 13821 36967 13824
rect 36909 13815 36967 13821
rect 36449 13787 36507 13793
rect 36449 13753 36461 13787
rect 36495 13784 36507 13787
rect 36998 13784 37004 13796
rect 36495 13756 37004 13784
rect 36495 13753 36507 13756
rect 36449 13747 36507 13753
rect 36998 13744 37004 13756
rect 37056 13744 37062 13796
rect 37292 13784 37320 13824
rect 37461 13821 37473 13855
rect 37507 13852 37519 13855
rect 37507 13824 38424 13852
rect 37507 13821 37519 13824
rect 37461 13815 37519 13821
rect 37734 13784 37740 13796
rect 37292 13756 37740 13784
rect 37734 13744 37740 13756
rect 37792 13744 37798 13796
rect 33643 13688 34928 13716
rect 35253 13719 35311 13725
rect 33643 13685 33655 13688
rect 33597 13679 33655 13685
rect 35253 13685 35265 13719
rect 35299 13716 35311 13719
rect 37458 13716 37464 13728
rect 35299 13688 37464 13716
rect 35299 13685 35311 13688
rect 35253 13679 35311 13685
rect 37458 13676 37464 13688
rect 37516 13676 37522 13728
rect 38396 13725 38424 13824
rect 38381 13719 38439 13725
rect 38381 13685 38393 13719
rect 38427 13716 38439 13719
rect 38746 13716 38752 13728
rect 38427 13688 38752 13716
rect 38427 13685 38439 13688
rect 38381 13679 38439 13685
rect 38746 13676 38752 13688
rect 38804 13676 38810 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 2961 13475 3019 13481
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 12618 13512 12624 13524
rect 10560 13484 12624 13512
rect 10560 13472 10566 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 13357 13515 13415 13521
rect 13357 13481 13369 13515
rect 13403 13512 13415 13515
rect 13446 13512 13452 13524
rect 13403 13484 13452 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14516 13484 14749 13512
rect 14516 13472 14522 13484
rect 14737 13481 14749 13484
rect 14783 13481 14795 13515
rect 14737 13475 14795 13481
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16482 13512 16488 13524
rect 16439 13484 16488 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 17236 13484 22094 13512
rect 3602 13336 3608 13388
rect 3660 13336 3666 13388
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 9309 13379 9367 13385
rect 9309 13376 9321 13379
rect 6604 13348 9321 13376
rect 6604 13336 6610 13348
rect 9309 13345 9321 13348
rect 9355 13376 9367 13379
rect 10226 13376 10232 13388
rect 9355 13348 10232 13376
rect 9355 13345 9367 13348
rect 9309 13339 9367 13345
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 13464 13376 13492 13472
rect 17129 13447 17187 13453
rect 17129 13413 17141 13447
rect 17175 13413 17187 13447
rect 17129 13407 17187 13413
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13464 13348 14105 13376
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 14093 13339 14151 13345
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 17144 13376 17172 13407
rect 17083 13348 17172 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 8754 13268 8760 13320
rect 8812 13268 8818 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 11885 13311 11943 13317
rect 9171 13280 11744 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 8021 13243 8079 13249
rect 8021 13240 8033 13243
rect 6972 13212 8033 13240
rect 6972 13200 6978 13212
rect 8021 13209 8033 13212
rect 8067 13240 8079 13243
rect 9140 13240 9168 13271
rect 8067 13212 9168 13240
rect 10336 13212 11100 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 10336 13184 10364 13212
rect 8110 13132 8116 13184
rect 8168 13132 8174 13184
rect 10318 13132 10324 13184
rect 10376 13132 10382 13184
rect 11072 13172 11100 13212
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 11618 13243 11676 13249
rect 11618 13240 11630 13243
rect 11388 13212 11630 13240
rect 11388 13200 11394 13212
rect 11618 13209 11630 13212
rect 11664 13209 11676 13243
rect 11716 13240 11744 13280
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 11974 13308 11980 13320
rect 11931 13280 11980 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12244 13311 12302 13317
rect 12244 13277 12256 13311
rect 12290 13308 12302 13311
rect 13630 13308 13636 13320
rect 12290 13280 13636 13308
rect 12290 13277 12302 13280
rect 12244 13271 12302 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 16298 13268 16304 13320
rect 16356 13268 16362 13320
rect 17236 13240 17264 13484
rect 22066 13444 22094 13484
rect 23290 13472 23296 13524
rect 23348 13512 23354 13524
rect 23477 13515 23535 13521
rect 23477 13512 23489 13515
rect 23348 13484 23489 13512
rect 23348 13472 23354 13484
rect 23477 13481 23489 13484
rect 23523 13481 23535 13515
rect 23477 13475 23535 13481
rect 23842 13472 23848 13524
rect 23900 13512 23906 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 23900 13484 24593 13512
rect 23900 13472 23906 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 25409 13515 25467 13521
rect 25409 13481 25421 13515
rect 25455 13512 25467 13515
rect 26050 13512 26056 13524
rect 25455 13484 26056 13512
rect 25455 13481 25467 13484
rect 25409 13475 25467 13481
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 26326 13472 26332 13524
rect 26384 13512 26390 13524
rect 26602 13512 26608 13524
rect 26384 13484 26608 13512
rect 26384 13472 26390 13484
rect 26602 13472 26608 13484
rect 26660 13472 26666 13524
rect 27062 13472 27068 13524
rect 27120 13472 27126 13524
rect 27985 13515 28043 13521
rect 27985 13481 27997 13515
rect 28031 13512 28043 13515
rect 28350 13512 28356 13524
rect 28031 13484 28356 13512
rect 28031 13481 28043 13484
rect 27985 13475 28043 13481
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 36170 13472 36176 13524
rect 36228 13512 36234 13524
rect 36265 13515 36323 13521
rect 36265 13512 36277 13515
rect 36228 13484 36277 13512
rect 36228 13472 36234 13484
rect 36265 13481 36277 13484
rect 36311 13481 36323 13515
rect 36265 13475 36323 13481
rect 28718 13444 28724 13456
rect 22066 13416 28724 13444
rect 28718 13404 28724 13416
rect 28776 13404 28782 13456
rect 17678 13336 17684 13388
rect 17736 13336 17742 13388
rect 18506 13336 18512 13388
rect 18564 13336 18570 13388
rect 21545 13379 21603 13385
rect 21545 13345 21557 13379
rect 21591 13376 21603 13379
rect 21591 13348 22094 13376
rect 21591 13345 21603 13348
rect 21545 13339 21603 13345
rect 22066 13320 22094 13348
rect 22278 13336 22284 13388
rect 22336 13376 22342 13388
rect 24765 13379 24823 13385
rect 24765 13376 24777 13379
rect 22336 13348 24777 13376
rect 22336 13336 22342 13348
rect 24765 13345 24777 13348
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 25774 13336 25780 13388
rect 25832 13376 25838 13388
rect 26053 13379 26111 13385
rect 26053 13376 26065 13379
rect 25832 13348 26065 13376
rect 25832 13336 25838 13348
rect 26053 13345 26065 13348
rect 26099 13376 26111 13379
rect 28166 13376 28172 13388
rect 26099 13348 28172 13376
rect 26099 13345 26111 13348
rect 26053 13339 26111 13345
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 34790 13336 34796 13388
rect 34848 13376 34854 13388
rect 36280 13376 36308 13475
rect 37734 13472 37740 13524
rect 37792 13512 37798 13524
rect 37918 13512 37924 13524
rect 37792 13484 37924 13512
rect 37792 13472 37798 13484
rect 37918 13472 37924 13484
rect 37976 13512 37982 13524
rect 38197 13515 38255 13521
rect 38197 13512 38209 13515
rect 37976 13484 38209 13512
rect 37976 13472 37982 13484
rect 38197 13481 38209 13484
rect 38243 13481 38255 13515
rect 38197 13475 38255 13481
rect 36817 13379 36875 13385
rect 36817 13376 36829 13379
rect 34848 13348 36829 13376
rect 34848 13336 34854 13348
rect 36817 13345 36829 13348
rect 36863 13345 36875 13379
rect 36817 13339 36875 13345
rect 17494 13268 17500 13320
rect 17552 13268 17558 13320
rect 22066 13280 22100 13320
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22189 13311 22247 13317
rect 22189 13277 22201 13311
rect 22235 13308 22247 13311
rect 22235 13280 23152 13308
rect 22235 13277 22247 13280
rect 22189 13271 22247 13277
rect 23124 13240 23152 13280
rect 23198 13268 23204 13320
rect 23256 13308 23262 13320
rect 27706 13308 27712 13320
rect 23256 13280 27712 13308
rect 23256 13268 23262 13280
rect 27706 13268 27712 13280
rect 27764 13308 27770 13320
rect 28445 13311 28503 13317
rect 28445 13308 28457 13311
rect 27764 13280 28457 13308
rect 27764 13268 27770 13280
rect 28445 13277 28457 13280
rect 28491 13277 28503 13311
rect 28445 13271 28503 13277
rect 30650 13268 30656 13320
rect 30708 13268 30714 13320
rect 31938 13268 31944 13320
rect 31996 13268 32002 13320
rect 32030 13268 32036 13320
rect 32088 13308 32094 13320
rect 32493 13311 32551 13317
rect 32493 13308 32505 13311
rect 32088 13280 32505 13308
rect 32088 13268 32094 13280
rect 32493 13277 32505 13280
rect 32539 13277 32551 13311
rect 32493 13271 32551 13277
rect 25038 13240 25044 13252
rect 11716 13212 17264 13240
rect 17328 13212 22232 13240
rect 23124 13212 25044 13240
rect 11618 13203 11676 13209
rect 17328 13172 17356 13212
rect 11072 13144 17356 13172
rect 17589 13175 17647 13181
rect 17589 13141 17601 13175
rect 17635 13172 17647 13175
rect 17957 13175 18015 13181
rect 17957 13172 17969 13175
rect 17635 13144 17969 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 17957 13141 17969 13144
rect 18003 13141 18015 13175
rect 17957 13135 18015 13141
rect 22094 13132 22100 13184
rect 22152 13132 22158 13184
rect 22204 13172 22232 13212
rect 25038 13200 25044 13212
rect 25096 13240 25102 13252
rect 25685 13243 25743 13249
rect 25685 13240 25697 13243
rect 25096 13212 25697 13240
rect 25096 13200 25102 13212
rect 25685 13209 25697 13212
rect 25731 13209 25743 13243
rect 28077 13243 28135 13249
rect 25685 13203 25743 13209
rect 25976 13212 28028 13240
rect 25976 13172 26004 13212
rect 22204 13144 26004 13172
rect 26510 13132 26516 13184
rect 26568 13172 26574 13184
rect 26786 13172 26792 13184
rect 26568 13144 26792 13172
rect 26568 13132 26574 13144
rect 26786 13132 26792 13144
rect 26844 13172 26850 13184
rect 27338 13172 27344 13184
rect 26844 13144 27344 13172
rect 26844 13132 26850 13144
rect 27338 13132 27344 13144
rect 27396 13132 27402 13184
rect 27522 13132 27528 13184
rect 27580 13172 27586 13184
rect 27709 13175 27767 13181
rect 27709 13172 27721 13175
rect 27580 13144 27721 13172
rect 27580 13132 27586 13144
rect 27709 13141 27721 13144
rect 27755 13141 27767 13175
rect 28000 13172 28028 13212
rect 28077 13209 28089 13243
rect 28123 13240 28135 13243
rect 28626 13240 28632 13252
rect 28123 13212 28632 13240
rect 28123 13209 28135 13212
rect 28077 13203 28135 13209
rect 28626 13200 28632 13212
rect 28684 13200 28690 13252
rect 29730 13200 29736 13252
rect 29788 13240 29794 13252
rect 30469 13243 30527 13249
rect 30469 13240 30481 13243
rect 29788 13212 30481 13240
rect 29788 13200 29794 13212
rect 30469 13209 30481 13212
rect 30515 13240 30527 13243
rect 30558 13240 30564 13252
rect 30515 13212 30564 13240
rect 30515 13209 30527 13212
rect 30469 13203 30527 13209
rect 30558 13200 30564 13212
rect 30616 13240 30622 13252
rect 34149 13243 34207 13249
rect 30616 13212 33824 13240
rect 30616 13200 30622 13212
rect 33796 13184 33824 13212
rect 34149 13209 34161 13243
rect 34195 13240 34207 13243
rect 34330 13240 34336 13252
rect 34195 13212 34336 13240
rect 34195 13209 34207 13212
rect 34149 13203 34207 13209
rect 34330 13200 34336 13212
rect 34388 13240 34394 13252
rect 34977 13243 35035 13249
rect 34977 13240 34989 13243
rect 34388 13212 34989 13240
rect 34388 13200 34394 13212
rect 34977 13209 34989 13212
rect 35023 13209 35035 13243
rect 34977 13203 35035 13209
rect 37084 13243 37142 13249
rect 37084 13209 37096 13243
rect 37130 13240 37142 13243
rect 37274 13240 37280 13252
rect 37130 13212 37280 13240
rect 37130 13209 37142 13212
rect 37084 13203 37142 13209
rect 37274 13200 37280 13212
rect 37332 13200 37338 13252
rect 29270 13172 29276 13184
rect 28000 13144 29276 13172
rect 27709 13135 27767 13141
rect 29270 13132 29276 13144
rect 29328 13132 29334 13184
rect 31202 13132 31208 13184
rect 31260 13132 31266 13184
rect 31294 13132 31300 13184
rect 31352 13132 31358 13184
rect 33778 13132 33784 13184
rect 33836 13172 33842 13184
rect 34517 13175 34575 13181
rect 34517 13172 34529 13175
rect 33836 13144 34529 13172
rect 33836 13132 33842 13144
rect 34517 13141 34529 13144
rect 34563 13172 34575 13175
rect 36998 13172 37004 13184
rect 34563 13144 37004 13172
rect 34563 13141 34575 13144
rect 34517 13135 34575 13141
rect 36998 13132 37004 13144
rect 37056 13132 37062 13184
rect 37458 13132 37464 13184
rect 37516 13172 37522 13184
rect 37734 13172 37740 13184
rect 37516 13144 37740 13172
rect 37516 13132 37522 13144
rect 37734 13132 37740 13144
rect 37792 13132 37798 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7926 12928 7932 12980
rect 7984 12928 7990 12980
rect 11330 12928 11336 12980
rect 11388 12928 11394 12980
rect 17037 12971 17095 12977
rect 17037 12937 17049 12971
rect 17083 12968 17095 12971
rect 17678 12968 17684 12980
rect 17083 12940 17684 12968
rect 17083 12937 17095 12940
rect 17037 12931 17095 12937
rect 2777 12903 2835 12909
rect 2777 12900 2789 12903
rect 1964 12872 2789 12900
rect 1964 12844 1992 12872
rect 2777 12869 2789 12872
rect 2823 12900 2835 12903
rect 4157 12903 4215 12909
rect 4157 12900 4169 12903
rect 2823 12872 4169 12900
rect 2823 12869 2835 12872
rect 2777 12863 2835 12869
rect 4157 12869 4169 12872
rect 4203 12869 4215 12903
rect 4157 12863 4215 12869
rect 6380 12872 9168 12900
rect 6380 12844 6408 12872
rect 1946 12792 1952 12844
rect 2004 12792 2010 12844
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3142 12832 3148 12844
rect 3007 12804 3148 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 2700 12764 2728 12795
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3789 12835 3847 12841
rect 3789 12832 3801 12835
rect 3292 12804 3801 12832
rect 3292 12792 3298 12804
rect 3789 12801 3801 12804
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 6362 12792 6368 12844
rect 6420 12792 6426 12844
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 9042 12835 9100 12841
rect 9042 12832 9054 12835
rect 8352 12804 9054 12832
rect 8352 12792 8358 12804
rect 9042 12801 9054 12804
rect 9088 12801 9100 12835
rect 9140 12832 9168 12872
rect 9214 12860 9220 12912
rect 9272 12900 9278 12912
rect 9272 12872 12434 12900
rect 9272 12860 9278 12872
rect 9398 12832 9404 12844
rect 9140 12804 9404 12832
rect 9042 12795 9100 12801
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 9916 12804 10241 12832
rect 9916 12792 9922 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10594 12792 10600 12844
rect 10652 12832 10658 12844
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10652 12804 10701 12832
rect 10652 12792 10658 12804
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 12406 12776 12434 12872
rect 12526 12860 12532 12912
rect 12584 12860 12590 12912
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 12768 12872 13584 12900
rect 12768 12860 12774 12872
rect 13556 12841 13584 12872
rect 13722 12860 13728 12912
rect 13780 12900 13786 12912
rect 15654 12900 15660 12912
rect 13780 12872 15660 12900
rect 13780 12860 13786 12872
rect 15654 12860 15660 12872
rect 15712 12900 15718 12912
rect 17052 12900 17080 12931
rect 17678 12928 17684 12940
rect 17736 12928 17742 12980
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 24397 12971 24455 12977
rect 24397 12968 24409 12971
rect 23624 12940 24409 12968
rect 23624 12928 23630 12940
rect 24397 12937 24409 12940
rect 24443 12937 24455 12971
rect 24397 12931 24455 12937
rect 27338 12928 27344 12980
rect 27396 12968 27402 12980
rect 27396 12940 30604 12968
rect 27396 12928 27402 12940
rect 15712 12872 17080 12900
rect 17589 12903 17647 12909
rect 15712 12860 15718 12872
rect 17589 12869 17601 12903
rect 17635 12900 17647 12903
rect 18230 12900 18236 12912
rect 17635 12872 18236 12900
rect 17635 12869 17647 12872
rect 17589 12863 17647 12869
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 22094 12909 22100 12912
rect 18693 12903 18751 12909
rect 18693 12900 18705 12903
rect 18380 12872 18705 12900
rect 18380 12860 18386 12872
rect 18693 12869 18705 12872
rect 18739 12869 18751 12903
rect 22088 12900 22100 12909
rect 22055 12872 22100 12900
rect 18693 12863 18751 12869
rect 22088 12863 22100 12872
rect 22094 12860 22100 12863
rect 22152 12860 22158 12912
rect 23014 12860 23020 12912
rect 23072 12900 23078 12912
rect 25133 12903 25191 12909
rect 25133 12900 25145 12903
rect 23072 12872 25145 12900
rect 23072 12860 23078 12872
rect 25133 12869 25145 12872
rect 25179 12869 25191 12903
rect 27433 12903 27491 12909
rect 25133 12863 25191 12869
rect 25608 12872 27292 12900
rect 12621 12835 12679 12841
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12667 12804 13001 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 2866 12764 2872 12776
rect 2700 12736 2872 12764
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 2961 12699 3019 12705
rect 2961 12665 2973 12699
rect 3007 12696 3019 12699
rect 3620 12696 3648 12727
rect 7282 12724 7288 12776
rect 7340 12724 7346 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 10134 12764 10140 12776
rect 9355 12736 10140 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 12406 12736 12440 12776
rect 12434 12724 12440 12736
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12764 12863 12767
rect 13740 12764 13768 12860
rect 17494 12792 17500 12844
rect 17552 12792 17558 12844
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12832 18935 12835
rect 19334 12832 19340 12844
rect 18923 12804 19340 12832
rect 18923 12801 18935 12804
rect 18877 12795 18935 12801
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12832 21879 12835
rect 21910 12832 21916 12844
rect 21867 12804 21916 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 23198 12792 23204 12844
rect 23256 12832 23262 12844
rect 23293 12835 23351 12841
rect 23293 12832 23305 12835
rect 23256 12804 23305 12832
rect 23256 12792 23262 12804
rect 23293 12801 23305 12804
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 24118 12792 24124 12844
rect 24176 12832 24182 12844
rect 24762 12832 24768 12844
rect 24176 12804 24768 12832
rect 24176 12792 24182 12804
rect 24762 12792 24768 12804
rect 24820 12832 24826 12844
rect 25608 12832 25636 12872
rect 24820 12804 25636 12832
rect 24820 12792 24826 12804
rect 25682 12792 25688 12844
rect 25740 12792 25746 12844
rect 12851 12736 13768 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 14274 12724 14280 12776
rect 14332 12724 14338 12776
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 3007 12668 3648 12696
rect 3007 12665 3019 12668
rect 2961 12659 3019 12665
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 15948 12696 15976 12727
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 17681 12767 17739 12773
rect 17681 12764 17693 12767
rect 16816 12736 17693 12764
rect 16816 12724 16822 12736
rect 17681 12733 17693 12736
rect 17727 12764 17739 12767
rect 18141 12767 18199 12773
rect 18141 12764 18153 12767
rect 17727 12736 18153 12764
rect 17727 12733 17739 12736
rect 17681 12727 17739 12733
rect 18141 12733 18153 12736
rect 18187 12733 18199 12767
rect 18141 12727 18199 12733
rect 20898 12724 20904 12776
rect 20956 12724 20962 12776
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12733 25007 12767
rect 24949 12727 25007 12733
rect 26789 12767 26847 12773
rect 26789 12733 26801 12767
rect 26835 12733 26847 12767
rect 26789 12727 26847 12733
rect 17129 12699 17187 12705
rect 17129 12696 17141 12699
rect 11848 12668 15884 12696
rect 15948 12668 17141 12696
rect 11848 12656 11854 12668
rect 15856 12640 15884 12668
rect 17129 12665 17141 12668
rect 17175 12665 17187 12699
rect 24964 12696 24992 12727
rect 17129 12659 17187 12665
rect 22756 12668 24992 12696
rect 26804 12696 26832 12727
rect 26973 12699 27031 12705
rect 26973 12696 26985 12699
rect 26804 12668 26985 12696
rect 3050 12588 3056 12640
rect 3108 12588 3114 12640
rect 7650 12588 7656 12640
rect 7708 12628 7714 12640
rect 7837 12631 7895 12637
rect 7837 12628 7849 12631
rect 7708 12600 7849 12628
rect 7708 12588 7714 12600
rect 7837 12597 7849 12600
rect 7883 12597 7895 12631
rect 7837 12591 7895 12597
rect 12158 12588 12164 12640
rect 12216 12588 12222 12640
rect 13722 12588 13728 12640
rect 13780 12588 13786 12640
rect 15838 12588 15844 12640
rect 15896 12588 15902 12640
rect 16485 12631 16543 12637
rect 16485 12597 16497 12631
rect 16531 12628 16543 12631
rect 16850 12628 16856 12640
rect 16531 12600 16856 12628
rect 16531 12597 16543 12600
rect 16485 12591 16543 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 21542 12588 21548 12640
rect 21600 12588 21606 12640
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 22756 12628 22784 12668
rect 26973 12665 26985 12668
rect 27019 12665 27031 12699
rect 27264 12696 27292 12872
rect 27433 12869 27445 12903
rect 27479 12900 27491 12903
rect 28442 12900 28448 12912
rect 27479 12872 28448 12900
rect 27479 12869 27491 12872
rect 27433 12863 27491 12869
rect 28442 12860 28448 12872
rect 28500 12860 28506 12912
rect 29825 12903 29883 12909
rect 29825 12869 29837 12903
rect 29871 12900 29883 12903
rect 30466 12900 30472 12912
rect 29871 12872 30472 12900
rect 29871 12869 29883 12872
rect 29825 12863 29883 12869
rect 30466 12860 30472 12872
rect 30524 12860 30530 12912
rect 27341 12835 27399 12841
rect 27341 12801 27353 12835
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27356 12764 27384 12795
rect 30576 12776 30604 12940
rect 30650 12928 30656 12980
rect 30708 12928 30714 12980
rect 31113 12971 31171 12977
rect 31113 12937 31125 12971
rect 31159 12968 31171 12971
rect 31294 12968 31300 12980
rect 31159 12940 31300 12968
rect 31159 12937 31171 12940
rect 31113 12931 31171 12937
rect 31294 12928 31300 12940
rect 31352 12928 31358 12980
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 32401 12971 32459 12977
rect 32401 12968 32413 12971
rect 32180 12940 32413 12968
rect 32180 12928 32186 12940
rect 32401 12937 32413 12940
rect 32447 12937 32459 12971
rect 32401 12931 32459 12937
rect 36081 12971 36139 12977
rect 36081 12937 36093 12971
rect 36127 12968 36139 12971
rect 36354 12968 36360 12980
rect 36127 12940 36360 12968
rect 36127 12937 36139 12940
rect 36081 12931 36139 12937
rect 36354 12928 36360 12940
rect 36412 12928 36418 12980
rect 37274 12928 37280 12980
rect 37332 12928 37338 12980
rect 38286 12928 38292 12980
rect 38344 12928 38350 12980
rect 33686 12860 33692 12912
rect 33744 12900 33750 12912
rect 34514 12900 34520 12912
rect 33744 12872 34520 12900
rect 33744 12860 33750 12872
rect 34514 12860 34520 12872
rect 34572 12860 34578 12912
rect 37550 12860 37556 12912
rect 37608 12900 37614 12912
rect 38102 12900 38108 12912
rect 37608 12872 38108 12900
rect 37608 12860 37614 12872
rect 38102 12860 38108 12872
rect 38160 12860 38166 12912
rect 31018 12792 31024 12844
rect 31076 12792 31082 12844
rect 32490 12792 32496 12844
rect 32548 12792 32554 12844
rect 34701 12835 34759 12841
rect 34701 12801 34713 12835
rect 34747 12832 34759 12835
rect 34790 12832 34796 12844
rect 34747 12804 34796 12832
rect 34747 12801 34759 12804
rect 34701 12795 34759 12801
rect 34790 12792 34796 12804
rect 34848 12792 34854 12844
rect 34968 12835 35026 12841
rect 34968 12801 34980 12835
rect 35014 12832 35026 12835
rect 36173 12835 36231 12841
rect 36173 12832 36185 12835
rect 35014 12804 36185 12832
rect 35014 12801 35026 12804
rect 34968 12795 35026 12801
rect 36173 12801 36185 12804
rect 36219 12801 36231 12835
rect 36173 12795 36231 12801
rect 37366 12792 37372 12844
rect 37424 12832 37430 12844
rect 37829 12835 37887 12841
rect 37829 12832 37841 12835
rect 37424 12804 37841 12832
rect 37424 12792 37430 12804
rect 37829 12801 37841 12804
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 27430 12764 27436 12776
rect 27356 12736 27436 12764
rect 27430 12724 27436 12736
rect 27488 12724 27494 12776
rect 27522 12724 27528 12776
rect 27580 12724 27586 12776
rect 28350 12724 28356 12776
rect 28408 12724 28414 12776
rect 28810 12724 28816 12776
rect 28868 12764 28874 12776
rect 29089 12767 29147 12773
rect 29089 12764 29101 12767
rect 28868 12736 29101 12764
rect 28868 12724 28874 12736
rect 29089 12733 29101 12736
rect 29135 12733 29147 12767
rect 29089 12727 29147 12733
rect 30466 12724 30472 12776
rect 30524 12724 30530 12776
rect 30558 12724 30564 12776
rect 30616 12764 30622 12776
rect 31205 12767 31263 12773
rect 31205 12764 31217 12767
rect 30616 12736 31217 12764
rect 30616 12724 30622 12736
rect 31205 12733 31217 12736
rect 31251 12733 31263 12767
rect 31205 12727 31263 12733
rect 31941 12767 31999 12773
rect 31941 12733 31953 12767
rect 31987 12764 31999 12767
rect 32122 12764 32128 12776
rect 31987 12736 32128 12764
rect 31987 12733 31999 12736
rect 31941 12727 31999 12733
rect 32122 12724 32128 12736
rect 32180 12764 32186 12776
rect 32217 12767 32275 12773
rect 32217 12764 32229 12767
rect 32180 12736 32229 12764
rect 32180 12724 32186 12736
rect 32217 12733 32229 12736
rect 32263 12733 32275 12767
rect 32217 12727 32275 12733
rect 33134 12724 33140 12776
rect 33192 12764 33198 12776
rect 33505 12767 33563 12773
rect 33505 12764 33517 12767
rect 33192 12736 33517 12764
rect 33192 12724 33198 12736
rect 33505 12733 33517 12736
rect 33551 12733 33563 12767
rect 33505 12727 33563 12733
rect 36722 12724 36728 12776
rect 36780 12724 36786 12776
rect 27540 12696 27568 12724
rect 32766 12696 32772 12708
rect 27264 12668 32772 12696
rect 26973 12659 27031 12665
rect 32766 12656 32772 12668
rect 32824 12656 32830 12708
rect 34238 12696 34244 12708
rect 32876 12668 34244 12696
rect 22612 12600 22784 12628
rect 22612 12588 22618 12600
rect 22830 12588 22836 12640
rect 22888 12628 22894 12640
rect 23201 12631 23259 12637
rect 23201 12628 23213 12631
rect 22888 12600 23213 12628
rect 22888 12588 22894 12600
rect 23201 12597 23213 12600
rect 23247 12628 23259 12631
rect 24946 12628 24952 12640
rect 23247 12600 24952 12628
rect 23247 12597 23259 12600
rect 23201 12591 23259 12597
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 26145 12631 26203 12637
rect 26145 12597 26157 12631
rect 26191 12628 26203 12631
rect 26326 12628 26332 12640
rect 26191 12600 26332 12628
rect 26191 12597 26203 12600
rect 26145 12591 26203 12597
rect 26326 12588 26332 12600
rect 26384 12588 26390 12640
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27801 12631 27859 12637
rect 27801 12628 27813 12631
rect 26752 12600 27813 12628
rect 26752 12588 26758 12600
rect 27801 12597 27813 12600
rect 27847 12597 27859 12631
rect 27801 12591 27859 12597
rect 28534 12588 28540 12640
rect 28592 12588 28598 12640
rect 29914 12588 29920 12640
rect 29972 12588 29978 12640
rect 32876 12637 32904 12668
rect 34238 12656 34244 12668
rect 34296 12656 34302 12708
rect 32861 12631 32919 12637
rect 32861 12597 32873 12631
rect 32907 12597 32919 12631
rect 32861 12591 32919 12597
rect 32950 12588 32956 12640
rect 33008 12588 33014 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 2866 12384 2872 12436
rect 2924 12384 2930 12436
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 3970 12424 3976 12436
rect 3007 12396 3976 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2976 12356 3004 12387
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4614 12424 4620 12436
rect 4295 12396 4620 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5902 12384 5908 12436
rect 5960 12424 5966 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 5960 12396 6377 12424
rect 5960 12384 5966 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 7285 12427 7343 12433
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 8294 12424 8300 12436
rect 7331 12396 8300 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 8754 12384 8760 12436
rect 8812 12384 8818 12436
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12492 12396 12541 12424
rect 12492 12384 12498 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 15804 12396 15945 12424
rect 15804 12384 15810 12396
rect 15933 12393 15945 12396
rect 15979 12393 15991 12427
rect 15933 12387 15991 12393
rect 18230 12384 18236 12436
rect 18288 12384 18294 12436
rect 20533 12427 20591 12433
rect 20533 12393 20545 12427
rect 20579 12424 20591 12427
rect 20579 12396 22784 12424
rect 20579 12393 20591 12396
rect 20533 12387 20591 12393
rect 2556 12328 3004 12356
rect 2556 12316 2562 12328
rect 3510 12316 3516 12368
rect 3568 12356 3574 12368
rect 4798 12356 4804 12368
rect 3568 12328 4804 12356
rect 3568 12316 3574 12328
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 18141 12359 18199 12365
rect 18141 12325 18153 12359
rect 18187 12356 18199 12359
rect 18598 12356 18604 12368
rect 18187 12328 18604 12356
rect 18187 12325 18199 12328
rect 18141 12319 18199 12325
rect 18598 12316 18604 12328
rect 18656 12356 18662 12368
rect 18656 12328 18828 12356
rect 18656 12316 18662 12328
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 6236 12260 7389 12288
rect 6236 12248 6242 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12288 12127 12291
rect 12158 12288 12164 12300
rect 12115 12260 12164 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 13906 12288 13912 12300
rect 13403 12260 13912 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 14792 12260 15117 12288
rect 14792 12248 14798 12260
rect 15105 12257 15117 12260
rect 15151 12288 15163 12291
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 15151 12260 16497 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 2314 12180 2320 12232
rect 2372 12180 2378 12232
rect 3602 12180 3608 12232
rect 3660 12180 3666 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 7650 12229 7656 12232
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 4856 12192 5365 12220
rect 4856 12180 4862 12192
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 7644 12183 7656 12229
rect 4157 12155 4215 12161
rect 2746 12124 3096 12152
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 2746 12084 2774 12124
rect 2464 12056 2774 12084
rect 3068 12084 3096 12124
rect 4157 12121 4169 12155
rect 4203 12152 4215 12155
rect 4982 12152 4988 12164
rect 4203 12124 4988 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 4982 12112 4988 12124
rect 5040 12112 5046 12164
rect 4801 12087 4859 12093
rect 4801 12084 4813 12087
rect 3068 12056 4813 12084
rect 2464 12044 2470 12056
rect 4801 12053 4813 12056
rect 4847 12053 4859 12087
rect 6564 12084 6592 12183
rect 6748 12152 6776 12183
rect 7650 12180 7656 12183
rect 7708 12180 7714 12232
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8444 12192 9137 12220
rect 8444 12180 8450 12192
rect 9125 12189 9137 12192
rect 9171 12220 9183 12223
rect 9582 12220 9588 12232
rect 9171 12192 9588 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 14645 12223 14703 12229
rect 14645 12220 14657 12223
rect 13504 12192 14657 12220
rect 13504 12180 13510 12192
rect 14645 12189 14657 12192
rect 14691 12189 14703 12223
rect 14645 12183 14703 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 8478 12152 8484 12164
rect 6748 12124 8484 12152
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 9214 12112 9220 12164
rect 9272 12152 9278 12164
rect 11057 12155 11115 12161
rect 11057 12152 11069 12155
rect 9272 12124 11069 12152
rect 9272 12112 9278 12124
rect 11057 12121 11069 12124
rect 11103 12152 11115 12155
rect 12158 12152 12164 12164
rect 11103 12124 12164 12152
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 15304 12096 15332 12183
rect 15841 12155 15899 12161
rect 15841 12121 15853 12155
rect 15887 12152 15899 12155
rect 16301 12155 16359 12161
rect 16301 12152 16313 12155
rect 15887 12124 16313 12152
rect 15887 12121 15899 12124
rect 15841 12115 15899 12121
rect 16301 12121 16313 12124
rect 16347 12121 16359 12155
rect 16500 12152 16528 12251
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 18800 12297 18828 12328
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16724 12260 16773 12288
rect 16724 12248 16730 12260
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 18785 12291 18843 12297
rect 18785 12257 18797 12291
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 20548 12288 20576 12387
rect 19935 12260 20576 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 20714 12248 20720 12300
rect 20772 12248 20778 12300
rect 22189 12291 22247 12297
rect 22189 12257 22201 12291
rect 22235 12288 22247 12291
rect 22554 12288 22560 12300
rect 22235 12260 22560 12288
rect 22235 12257 22247 12260
rect 22189 12251 22247 12257
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 22646 12248 22652 12300
rect 22704 12248 22710 12300
rect 22756 12288 22784 12396
rect 28350 12384 28356 12436
rect 28408 12384 28414 12436
rect 28442 12384 28448 12436
rect 28500 12384 28506 12436
rect 30745 12427 30803 12433
rect 30745 12393 30757 12427
rect 30791 12424 30803 12427
rect 32490 12424 32496 12436
rect 30791 12396 32496 12424
rect 30791 12393 30803 12396
rect 30745 12387 30803 12393
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 32766 12384 32772 12436
rect 32824 12424 32830 12436
rect 34885 12427 34943 12433
rect 34885 12424 34897 12427
rect 32824 12396 34897 12424
rect 32824 12384 32830 12396
rect 34885 12393 34897 12396
rect 34931 12393 34943 12427
rect 34885 12387 34943 12393
rect 35805 12427 35863 12433
rect 35805 12393 35817 12427
rect 35851 12424 35863 12427
rect 36722 12424 36728 12436
rect 35851 12396 36728 12424
rect 35851 12393 35863 12396
rect 35805 12387 35863 12393
rect 27525 12359 27583 12365
rect 27525 12325 27537 12359
rect 27571 12356 27583 12359
rect 28810 12356 28816 12368
rect 27571 12328 28816 12356
rect 27571 12325 27583 12328
rect 27525 12319 27583 12325
rect 28810 12316 28816 12328
rect 28868 12316 28874 12368
rect 30926 12316 30932 12368
rect 30984 12316 30990 12368
rect 31941 12359 31999 12365
rect 31941 12325 31953 12359
rect 31987 12356 31999 12359
rect 33413 12359 33471 12365
rect 31987 12328 33272 12356
rect 31987 12325 31999 12328
rect 31941 12319 31999 12325
rect 23042 12291 23100 12297
rect 23042 12288 23054 12291
rect 22756 12260 23054 12288
rect 23042 12257 23054 12260
rect 23088 12257 23100 12291
rect 23042 12251 23100 12257
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12288 23259 12291
rect 24210 12288 24216 12300
rect 23247 12260 24216 12288
rect 23247 12257 23259 12260
rect 23201 12251 23259 12257
rect 24210 12248 24216 12260
rect 24268 12248 24274 12300
rect 24762 12248 24768 12300
rect 24820 12288 24826 12300
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 24820 12260 25053 12288
rect 24820 12248 24826 12260
rect 25041 12257 25053 12260
rect 25087 12288 25099 12291
rect 25222 12288 25228 12300
rect 25087 12260 25228 12288
rect 25087 12257 25099 12260
rect 25041 12251 25099 12257
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 25409 12291 25467 12297
rect 25409 12257 25421 12291
rect 25455 12288 25467 12291
rect 25498 12288 25504 12300
rect 25455 12260 25504 12288
rect 25455 12257 25467 12260
rect 25409 12251 25467 12257
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 26145 12291 26203 12297
rect 26145 12257 26157 12291
rect 26191 12257 26203 12291
rect 26145 12251 26203 12257
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17017 12223 17075 12229
rect 17017 12220 17029 12223
rect 16908 12192 17029 12220
rect 16908 12180 16914 12192
rect 17017 12189 17029 12192
rect 17063 12189 17075 12223
rect 17017 12183 17075 12189
rect 20732 12152 20760 12248
rect 21634 12180 21640 12232
rect 21692 12229 21698 12232
rect 21692 12183 21704 12229
rect 21692 12180 21698 12183
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21876 12192 21925 12220
rect 21876 12180 21882 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 22005 12223 22063 12229
rect 22005 12189 22017 12223
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 16500 12124 20760 12152
rect 16301 12115 16359 12121
rect 8202 12084 8208 12096
rect 6564 12056 8208 12084
rect 4801 12047 4859 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 12710 12044 12716 12096
rect 12768 12044 12774 12096
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 13170 12044 13176 12096
rect 13228 12044 13234 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 13909 12087 13967 12093
rect 13909 12084 13921 12087
rect 13872 12056 13921 12084
rect 13872 12044 13878 12056
rect 13909 12053 13921 12056
rect 13955 12084 13967 12087
rect 13998 12084 14004 12096
rect 13955 12056 14004 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 14090 12044 14096 12096
rect 14148 12044 14154 12096
rect 15286 12044 15292 12096
rect 15344 12044 15350 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 15436 12056 16405 12084
rect 15436 12044 15442 12056
rect 16393 12053 16405 12056
rect 16439 12084 16451 12087
rect 17494 12084 17500 12096
rect 16439 12056 17500 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 20438 12044 20444 12096
rect 20496 12044 20502 12096
rect 22020 12084 22048 12183
rect 22922 12180 22928 12232
rect 22980 12180 22986 12232
rect 24394 12180 24400 12232
rect 24452 12220 24458 12232
rect 25593 12223 25651 12229
rect 25593 12220 25605 12223
rect 24452 12192 25605 12220
rect 24452 12180 24458 12192
rect 25593 12189 25605 12192
rect 25639 12189 25651 12223
rect 26160 12220 26188 12251
rect 27706 12248 27712 12300
rect 27764 12248 27770 12300
rect 27893 12291 27951 12297
rect 27893 12257 27905 12291
rect 27939 12288 27951 12291
rect 28534 12288 28540 12300
rect 27939 12260 28540 12288
rect 27939 12257 27951 12260
rect 27893 12251 27951 12257
rect 28534 12248 28540 12260
rect 28592 12248 28598 12300
rect 30944 12288 30972 12316
rect 31389 12291 31447 12297
rect 31389 12288 31401 12291
rect 28644 12260 31401 12288
rect 26234 12220 26240 12232
rect 26160 12192 26240 12220
rect 25593 12183 25651 12189
rect 26234 12180 26240 12192
rect 26292 12180 26298 12232
rect 28644 12220 28672 12260
rect 31389 12257 31401 12260
rect 31435 12257 31447 12291
rect 31389 12251 31447 12257
rect 31548 12291 31606 12297
rect 31548 12257 31560 12291
rect 31594 12288 31606 12291
rect 31846 12288 31852 12300
rect 31594 12260 31852 12288
rect 31594 12257 31606 12260
rect 31548 12251 31606 12257
rect 31846 12248 31852 12260
rect 31904 12248 31910 12300
rect 32030 12248 32036 12300
rect 32088 12288 32094 12300
rect 32769 12291 32827 12297
rect 32769 12288 32781 12291
rect 32088 12260 32781 12288
rect 32088 12248 32094 12260
rect 32769 12257 32781 12260
rect 32815 12257 32827 12291
rect 32769 12251 32827 12257
rect 32950 12248 32956 12300
rect 33008 12248 33014 12300
rect 33134 12248 33140 12300
rect 33192 12248 33198 12300
rect 27847 12192 28672 12220
rect 28997 12223 29055 12229
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 25501 12155 25559 12161
rect 25501 12152 25513 12155
rect 23891 12124 25513 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 25501 12121 25513 12124
rect 25547 12121 25559 12155
rect 25501 12115 25559 12121
rect 26412 12155 26470 12161
rect 26412 12121 26424 12155
rect 26458 12152 26470 12155
rect 26694 12152 26700 12164
rect 26458 12124 26700 12152
rect 26458 12121 26470 12124
rect 26412 12115 26470 12121
rect 26694 12112 26700 12124
rect 26752 12112 26758 12164
rect 27062 12112 27068 12164
rect 27120 12152 27126 12164
rect 27847 12152 27875 12192
rect 28997 12189 29009 12223
rect 29043 12189 29055 12223
rect 28997 12183 29055 12189
rect 27120 12124 27875 12152
rect 27120 12112 27126 12124
rect 28442 12112 28448 12164
rect 28500 12152 28506 12164
rect 29012 12152 29040 12183
rect 30098 12180 30104 12232
rect 30156 12180 30162 12232
rect 31662 12180 31668 12232
rect 31720 12180 31726 12232
rect 32401 12223 32459 12229
rect 32401 12189 32413 12223
rect 32447 12189 32459 12223
rect 32401 12183 32459 12189
rect 32585 12223 32643 12229
rect 32585 12189 32597 12223
rect 32631 12220 32643 12223
rect 33152 12220 33180 12248
rect 32631 12192 33180 12220
rect 33244 12220 33272 12328
rect 33413 12325 33425 12359
rect 33459 12325 33471 12359
rect 33413 12319 33471 12325
rect 33428 12288 33456 12319
rect 34057 12291 34115 12297
rect 34057 12288 34069 12291
rect 33428 12260 34069 12288
rect 34057 12257 34069 12260
rect 34103 12257 34115 12291
rect 34900 12288 34928 12387
rect 36722 12384 36728 12396
rect 36780 12384 36786 12436
rect 37458 12384 37464 12436
rect 37516 12384 37522 12436
rect 37826 12384 37832 12436
rect 37884 12384 37890 12436
rect 35161 12291 35219 12297
rect 35161 12288 35173 12291
rect 34900 12260 35173 12288
rect 34057 12251 34115 12257
rect 35161 12257 35173 12260
rect 35207 12257 35219 12291
rect 35161 12251 35219 12257
rect 36446 12248 36452 12300
rect 36504 12248 36510 12300
rect 37918 12248 37924 12300
rect 37976 12288 37982 12300
rect 38381 12291 38439 12297
rect 38381 12288 38393 12291
rect 37976 12260 38393 12288
rect 37976 12248 37982 12260
rect 38381 12257 38393 12260
rect 38427 12257 38439 12291
rect 38381 12251 38439 12257
rect 33778 12220 33784 12232
rect 33244 12192 33784 12220
rect 32631 12189 32643 12192
rect 32585 12183 32643 12189
rect 28500 12124 29040 12152
rect 28500 12112 28506 12124
rect 32416 12096 32444 12183
rect 33778 12180 33784 12192
rect 33836 12180 33842 12232
rect 35345 12155 35403 12161
rect 35345 12121 35357 12155
rect 35391 12152 35403 12155
rect 35897 12155 35955 12161
rect 35897 12152 35909 12155
rect 35391 12124 35909 12152
rect 35391 12121 35403 12124
rect 35345 12115 35403 12121
rect 35897 12121 35909 12124
rect 35943 12121 35955 12155
rect 35897 12115 35955 12121
rect 37553 12155 37611 12161
rect 37553 12121 37565 12155
rect 37599 12152 37611 12155
rect 38010 12152 38016 12164
rect 37599 12124 38016 12152
rect 37599 12121 37611 12124
rect 37553 12115 37611 12121
rect 38010 12112 38016 12124
rect 38068 12112 38074 12164
rect 22830 12084 22836 12096
rect 22020 12056 22836 12084
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 23198 12044 23204 12096
rect 23256 12084 23262 12096
rect 24121 12087 24179 12093
rect 24121 12084 24133 12087
rect 23256 12056 24133 12084
rect 23256 12044 23262 12056
rect 24121 12053 24133 12056
rect 24167 12053 24179 12087
rect 24121 12047 24179 12053
rect 24394 12044 24400 12096
rect 24452 12044 24458 12096
rect 24762 12044 24768 12096
rect 24820 12044 24826 12096
rect 24854 12044 24860 12096
rect 24912 12044 24918 12096
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 25961 12087 26019 12093
rect 25961 12084 25973 12087
rect 25832 12056 25973 12084
rect 25832 12044 25838 12056
rect 25961 12053 25973 12056
rect 26007 12053 26019 12087
rect 25961 12047 26019 12053
rect 27430 12044 27436 12096
rect 27488 12084 27494 12096
rect 27982 12084 27988 12096
rect 27488 12056 27988 12084
rect 27488 12044 27494 12056
rect 27982 12044 27988 12056
rect 28040 12044 28046 12096
rect 29086 12044 29092 12096
rect 29144 12084 29150 12096
rect 29549 12087 29607 12093
rect 29549 12084 29561 12087
rect 29144 12056 29561 12084
rect 29144 12044 29150 12056
rect 29549 12053 29561 12056
rect 29595 12053 29607 12087
rect 29549 12047 29607 12053
rect 30558 12044 30564 12096
rect 30616 12044 30622 12096
rect 31110 12044 31116 12096
rect 31168 12084 31174 12096
rect 31662 12084 31668 12096
rect 31168 12056 31668 12084
rect 31168 12044 31174 12056
rect 31662 12044 31668 12056
rect 31720 12084 31726 12096
rect 31938 12084 31944 12096
rect 31720 12056 31944 12084
rect 31720 12044 31726 12056
rect 31938 12044 31944 12056
rect 31996 12044 32002 12096
rect 32398 12044 32404 12096
rect 32456 12044 32462 12096
rect 32490 12044 32496 12096
rect 32548 12084 32554 12096
rect 33045 12087 33103 12093
rect 33045 12084 33057 12087
rect 32548 12056 33057 12084
rect 32548 12044 32554 12056
rect 33045 12053 33057 12056
rect 33091 12053 33103 12087
rect 33045 12047 33103 12053
rect 33226 12044 33232 12096
rect 33284 12084 33290 12096
rect 33505 12087 33563 12093
rect 33505 12084 33517 12087
rect 33284 12056 33517 12084
rect 33284 12044 33290 12056
rect 33505 12053 33517 12056
rect 33551 12053 33563 12087
rect 33505 12047 33563 12053
rect 34514 12044 34520 12096
rect 34572 12044 34578 12096
rect 35437 12087 35495 12093
rect 35437 12053 35449 12087
rect 35483 12084 35495 12087
rect 36078 12084 36084 12096
rect 35483 12056 36084 12084
rect 35483 12053 35495 12056
rect 35437 12047 35495 12053
rect 36078 12044 36084 12056
rect 36136 12044 36142 12096
rect 37182 12044 37188 12096
rect 37240 12044 37246 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 2314 11840 2320 11892
rect 2372 11880 2378 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2372 11852 2421 11880
rect 2372 11840 2378 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3660 11852 3985 11880
rect 3660 11840 3666 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 5258 11880 5264 11892
rect 3973 11843 4031 11849
rect 4264 11852 5264 11880
rect 1762 11772 1768 11824
rect 1820 11772 1826 11824
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 1965 11815 2023 11821
rect 1965 11812 1977 11815
rect 1912 11784 1977 11812
rect 1912 11772 1918 11784
rect 1965 11781 1977 11784
rect 2011 11781 2023 11815
rect 1965 11775 2023 11781
rect 2860 11815 2918 11821
rect 2860 11781 2872 11815
rect 2906 11812 2918 11815
rect 3050 11812 3056 11824
rect 2906 11784 3056 11812
rect 2906 11781 2918 11784
rect 2860 11775 2918 11781
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3988 11812 4016 11843
rect 4264 11821 4292 11852
rect 5258 11840 5264 11852
rect 5316 11880 5322 11892
rect 5362 11883 5420 11889
rect 5362 11880 5374 11883
rect 5316 11852 5374 11880
rect 5316 11840 5322 11852
rect 5362 11849 5374 11852
rect 5408 11849 5420 11883
rect 5362 11843 5420 11849
rect 6454 11840 6460 11892
rect 6512 11880 6518 11892
rect 6730 11880 6736 11892
rect 6512 11852 6736 11880
rect 6512 11840 6518 11852
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 7340 11852 7389 11880
rect 7340 11840 7346 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 7377 11843 7435 11849
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11880 7895 11883
rect 8110 11880 8116 11892
rect 7883 11852 8116 11880
rect 7883 11849 7895 11852
rect 7837 11843 7895 11849
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9732 11852 10640 11880
rect 9732 11840 9738 11852
rect 4249 11815 4307 11821
rect 4249 11812 4261 11815
rect 3988 11784 4261 11812
rect 4249 11781 4261 11784
rect 4295 11781 4307 11815
rect 4249 11775 4307 11781
rect 4663 11815 4721 11821
rect 4663 11781 4675 11815
rect 4709 11812 4721 11815
rect 5166 11812 5172 11824
rect 4709 11784 5172 11812
rect 4709 11781 4721 11784
rect 4663 11775 4721 11781
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 8386 11812 8392 11824
rect 5644 11784 8392 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2332 11620 2360 11707
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 5644 11753 5672 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 2314 11608 2320 11620
rect 1964 11580 2320 11608
rect 1964 11549 1992 11580
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 1949 11543 2007 11549
rect 1949 11509 1961 11543
rect 1995 11509 2007 11543
rect 1949 11503 2007 11509
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 2498 11540 2504 11552
rect 2179 11512 2504 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 2608 11540 2636 11639
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 5000 11676 5028 11707
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7009 11747 7067 11753
rect 7009 11713 7021 11747
rect 7055 11744 7067 11747
rect 7742 11744 7748 11756
rect 7055 11716 7748 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 8018 11704 8024 11756
rect 8076 11744 8082 11756
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 8076 11716 8217 11744
rect 8076 11704 8082 11716
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10612 11744 10640 11852
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11020 11852 11897 11880
rect 11020 11840 11026 11852
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 10612 11716 11161 11744
rect 6730 11676 6736 11688
rect 4856 11648 5028 11676
rect 5092 11648 6736 11676
rect 4856 11636 4862 11648
rect 4816 11608 4844 11636
rect 4632 11580 4844 11608
rect 2774 11540 2780 11552
rect 2608 11512 2780 11540
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 4632 11549 4660 11580
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 5092 11540 5120 11648
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 6181 11611 6239 11617
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 6638 11608 6644 11620
rect 6227 11580 6644 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 7116 11608 7144 11639
rect 6696 11580 7144 11608
rect 6696 11568 6702 11580
rect 7944 11552 7972 11639
rect 8386 11636 8392 11688
rect 8444 11636 8450 11688
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 8812 11648 9137 11676
rect 8812 11636 8818 11648
rect 9125 11645 9137 11648
rect 9171 11645 9183 11679
rect 9125 11639 9183 11645
rect 9214 11636 9220 11688
rect 9272 11685 9278 11688
rect 9272 11679 9300 11685
rect 9288 11645 9300 11679
rect 9272 11639 9300 11645
rect 9272 11636 9278 11639
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 10704 11685 10732 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 9640 11648 10609 11676
rect 9640 11636 9646 11648
rect 10597 11645 10609 11648
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11645 10747 11679
rect 10689 11639 10747 11645
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 8849 11611 8907 11617
rect 8849 11608 8861 11611
rect 8628 11580 8861 11608
rect 8628 11568 8634 11580
rect 8849 11577 8861 11580
rect 8895 11577 8907 11611
rect 8849 11571 8907 11577
rect 10045 11611 10103 11617
rect 10045 11577 10057 11611
rect 10091 11608 10103 11611
rect 10318 11608 10324 11620
rect 10091 11580 10324 11608
rect 10091 11577 10103 11580
rect 10045 11571 10103 11577
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 4847 11512 5120 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5224 11512 5365 11540
rect 5224 11500 5230 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 6546 11500 6552 11552
rect 6604 11500 6610 11552
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 9122 11540 9128 11552
rect 7984 11512 9128 11540
rect 7984 11500 7990 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10134 11500 10140 11552
rect 10192 11500 10198 11552
rect 11900 11540 11928 11843
rect 13446 11840 13452 11892
rect 13504 11840 13510 11892
rect 13817 11883 13875 11889
rect 13817 11849 13829 11883
rect 13863 11880 13875 11883
rect 14090 11880 14096 11892
rect 13863 11852 14096 11880
rect 13863 11849 13875 11852
rect 13817 11843 13875 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14274 11840 14280 11892
rect 14332 11840 14338 11892
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 17402 11880 17408 11892
rect 17184 11852 17408 11880
rect 17184 11840 17190 11852
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17552 11852 18552 11880
rect 17552 11840 17558 11852
rect 12336 11815 12394 11821
rect 12336 11781 12348 11815
rect 12382 11812 12394 11815
rect 13722 11812 13728 11824
rect 12382 11784 13728 11812
rect 12382 11781 12394 11784
rect 12336 11775 12394 11781
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 16206 11772 16212 11824
rect 16264 11821 16270 11824
rect 16264 11815 16298 11821
rect 16286 11781 16298 11815
rect 16264 11775 16298 11781
rect 16264 11772 16270 11775
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 12032 11716 12081 11744
rect 12032 11704 12038 11716
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13228 11716 13921 11744
rect 13228 11704 13234 11716
rect 13909 11713 13921 11716
rect 13955 11744 13967 11747
rect 15378 11744 15384 11756
rect 13955 11716 15384 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16666 11744 16672 11756
rect 16531 11716 16672 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 14918 11636 14924 11688
rect 14976 11636 14982 11688
rect 17543 11679 17601 11685
rect 17543 11676 17555 11679
rect 16776 11648 17555 11676
rect 16776 11608 16804 11648
rect 17543 11645 17555 11648
rect 17589 11645 17601 11679
rect 17543 11639 17601 11645
rect 17681 11679 17739 11685
rect 17681 11645 17693 11679
rect 17727 11676 17739 11679
rect 18046 11676 18052 11688
rect 17727 11648 18052 11676
rect 17727 11645 17739 11648
rect 17681 11639 17739 11645
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18414 11676 18420 11688
rect 18340 11648 18420 11676
rect 16500 11580 16804 11608
rect 17957 11611 18015 11617
rect 13906 11540 13912 11552
rect 11900 11512 13912 11540
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14369 11543 14427 11549
rect 14369 11540 14381 11543
rect 14148 11512 14381 11540
rect 14148 11500 14154 11512
rect 14369 11509 14381 11512
rect 14415 11509 14427 11543
rect 14369 11503 14427 11509
rect 15105 11543 15163 11549
rect 15105 11509 15117 11543
rect 15151 11540 15163 11543
rect 15286 11540 15292 11552
rect 15151 11512 15292 11540
rect 15151 11509 15163 11512
rect 15105 11503 15163 11509
rect 15286 11500 15292 11512
rect 15344 11540 15350 11552
rect 16500 11540 16528 11580
rect 17957 11577 17969 11611
rect 18003 11577 18015 11611
rect 17957 11571 18015 11577
rect 15344 11512 16528 11540
rect 15344 11500 15350 11512
rect 16758 11500 16764 11552
rect 16816 11500 16822 11552
rect 17586 11500 17592 11552
rect 17644 11540 17650 11552
rect 17972 11540 18000 11571
rect 17644 11512 18000 11540
rect 18340 11540 18368 11648
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 18524 11676 18552 11852
rect 18598 11840 18604 11892
rect 18656 11840 18662 11892
rect 20438 11840 20444 11892
rect 20496 11840 20502 11892
rect 20898 11840 20904 11892
rect 20956 11840 20962 11892
rect 21361 11883 21419 11889
rect 21361 11849 21373 11883
rect 21407 11880 21419 11883
rect 21407 11852 22094 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 18616 11753 18644 11840
rect 20456 11812 20484 11840
rect 21269 11815 21327 11821
rect 21269 11812 21281 11815
rect 20456 11784 21281 11812
rect 21269 11781 21281 11784
rect 21315 11781 21327 11815
rect 22066 11812 22094 11852
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 23198 11880 23204 11892
rect 22336 11852 23204 11880
rect 22336 11840 22342 11852
rect 23198 11840 23204 11852
rect 23256 11840 23262 11892
rect 26789 11883 26847 11889
rect 26789 11849 26801 11883
rect 26835 11880 26847 11883
rect 27706 11880 27712 11892
rect 26835 11852 27712 11880
rect 26835 11849 26847 11852
rect 26789 11843 26847 11849
rect 27706 11840 27712 11852
rect 27764 11840 27770 11892
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 29181 11883 29239 11889
rect 29181 11880 29193 11883
rect 28040 11852 29193 11880
rect 28040 11840 28046 11852
rect 29181 11849 29193 11852
rect 29227 11849 29239 11883
rect 29181 11843 29239 11849
rect 29641 11883 29699 11889
rect 29641 11849 29653 11883
rect 29687 11880 29699 11883
rect 30098 11880 30104 11892
rect 29687 11852 30104 11880
rect 29687 11849 29699 11852
rect 29641 11843 29699 11849
rect 30098 11840 30104 11852
rect 30156 11840 30162 11892
rect 32125 11883 32183 11889
rect 32125 11849 32137 11883
rect 32171 11880 32183 11883
rect 33134 11880 33140 11892
rect 32171 11852 33140 11880
rect 32171 11849 32183 11852
rect 32125 11843 32183 11849
rect 33134 11840 33140 11852
rect 33192 11840 33198 11892
rect 38286 11880 38292 11892
rect 33244 11852 38292 11880
rect 22370 11812 22376 11824
rect 22066 11784 22376 11812
rect 21269 11775 21327 11781
rect 22370 11772 22376 11784
rect 22428 11772 22434 11824
rect 22646 11812 22652 11824
rect 22480 11784 22652 11812
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11744 19119 11747
rect 19521 11747 19579 11753
rect 19521 11744 19533 11747
rect 19107 11716 19533 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 19521 11713 19533 11716
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 22088 11747 22146 11753
rect 22088 11713 22100 11747
rect 22134 11744 22146 11747
rect 22480 11744 22508 11784
rect 22646 11772 22652 11784
rect 22704 11772 22710 11824
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 24762 11812 24768 11824
rect 23624 11784 24768 11812
rect 23624 11772 23630 11784
rect 24762 11772 24768 11784
rect 24820 11772 24826 11824
rect 27062 11772 27068 11824
rect 27120 11772 27126 11824
rect 29914 11772 29920 11824
rect 29972 11812 29978 11824
rect 30184 11815 30242 11821
rect 30184 11812 30196 11815
rect 29972 11784 30196 11812
rect 29972 11772 29978 11784
rect 30184 11781 30196 11784
rect 30230 11781 30242 11815
rect 30184 11775 30242 11781
rect 32030 11772 32036 11824
rect 32088 11812 32094 11824
rect 33244 11812 33272 11852
rect 38286 11840 38292 11852
rect 38344 11840 38350 11892
rect 32088 11784 33272 11812
rect 34517 11815 34575 11821
rect 32088 11772 32094 11784
rect 34517 11781 34529 11815
rect 34563 11812 34575 11815
rect 35774 11815 35832 11821
rect 35774 11812 35786 11815
rect 34563 11784 35786 11812
rect 34563 11781 34575 11784
rect 34517 11775 34575 11781
rect 35774 11781 35786 11784
rect 35820 11781 35832 11815
rect 35774 11775 35832 11781
rect 37645 11815 37703 11821
rect 37645 11781 37657 11815
rect 37691 11812 37703 11815
rect 37734 11812 37740 11824
rect 37691 11784 37740 11812
rect 37691 11781 37703 11784
rect 37645 11775 37703 11781
rect 37734 11772 37740 11784
rect 37792 11772 37798 11824
rect 22134 11716 22508 11744
rect 22134 11713 22146 11716
rect 22088 11707 22146 11713
rect 23382 11704 23388 11756
rect 23440 11704 23446 11756
rect 24946 11704 24952 11756
rect 25004 11704 25010 11756
rect 25676 11747 25734 11753
rect 25676 11713 25688 11747
rect 25722 11744 25734 11747
rect 26142 11744 26148 11756
rect 25722 11716 26148 11744
rect 25722 11713 25734 11716
rect 25676 11707 25734 11713
rect 26142 11704 26148 11716
rect 26200 11704 26206 11756
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 18524 11648 19165 11676
rect 19153 11645 19165 11648
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 19242 11636 19248 11688
rect 19300 11636 19306 11688
rect 20073 11679 20131 11685
rect 20073 11645 20085 11679
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 21545 11679 21603 11685
rect 21545 11645 21557 11679
rect 21591 11676 21603 11679
rect 21726 11676 21732 11688
rect 21591 11648 21732 11676
rect 21591 11645 21603 11648
rect 21545 11639 21603 11645
rect 20088 11608 20116 11639
rect 21726 11636 21732 11648
rect 21784 11636 21790 11688
rect 21818 11636 21824 11688
rect 21876 11636 21882 11688
rect 23290 11636 23296 11688
rect 23348 11636 23354 11688
rect 23842 11636 23848 11688
rect 23900 11676 23906 11688
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 23900 11648 24133 11676
rect 23900 11636 23906 11648
rect 24121 11645 24133 11648
rect 24167 11676 24179 11679
rect 24578 11676 24584 11688
rect 24167 11648 24584 11676
rect 24167 11645 24179 11648
rect 24121 11639 24179 11645
rect 24578 11636 24584 11648
rect 24636 11636 24642 11688
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11645 25467 11679
rect 27080 11676 27108 11772
rect 27798 11753 27804 11756
rect 27776 11747 27804 11753
rect 27776 11713 27788 11747
rect 27776 11707 27804 11713
rect 27798 11704 27804 11707
rect 27856 11704 27862 11756
rect 28442 11704 28448 11756
rect 28500 11704 28506 11756
rect 28810 11704 28816 11756
rect 28868 11704 28874 11756
rect 29270 11704 29276 11756
rect 29328 11704 29334 11756
rect 33226 11704 33232 11756
rect 33284 11753 33290 11756
rect 33284 11744 33296 11753
rect 33284 11716 33329 11744
rect 33284 11707 33296 11716
rect 33284 11704 33290 11707
rect 33502 11704 33508 11756
rect 33560 11744 33566 11756
rect 33560 11716 34836 11744
rect 33560 11704 33566 11716
rect 27617 11679 27675 11685
rect 27617 11676 27629 11679
rect 27080 11648 27629 11676
rect 25409 11639 25467 11645
rect 27617 11645 27629 11648
rect 27663 11645 27675 11679
rect 27617 11639 27675 11645
rect 18616 11580 20116 11608
rect 18616 11540 18644 11580
rect 18340 11512 18644 11540
rect 17644 11500 17650 11512
rect 18690 11500 18696 11552
rect 18748 11500 18754 11552
rect 21836 11540 21864 11636
rect 23308 11608 23336 11636
rect 22756 11580 23336 11608
rect 22756 11540 22784 11580
rect 21836 11512 22784 11540
rect 22922 11500 22928 11552
rect 22980 11540 22986 11552
rect 23198 11540 23204 11552
rect 22980 11512 23204 11540
rect 22980 11500 22986 11512
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 24397 11543 24455 11549
rect 24397 11540 24409 11543
rect 23532 11512 24409 11540
rect 23532 11500 23538 11512
rect 24397 11509 24409 11512
rect 24443 11509 24455 11543
rect 25424 11540 25452 11639
rect 27890 11636 27896 11688
rect 27948 11676 27954 11688
rect 28460 11676 28488 11704
rect 34808 11688 34836 11716
rect 37200 11716 37872 11744
rect 37200 11688 37228 11716
rect 27948 11648 28488 11676
rect 28629 11679 28687 11685
rect 27948 11636 27954 11648
rect 28629 11645 28641 11679
rect 28675 11676 28687 11679
rect 28718 11676 28724 11688
rect 28675 11648 28724 11676
rect 28675 11645 28687 11648
rect 28629 11639 28687 11645
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 28994 11636 29000 11688
rect 29052 11636 29058 11688
rect 29822 11636 29828 11688
rect 29880 11676 29886 11688
rect 29917 11679 29975 11685
rect 29917 11676 29929 11679
rect 29880 11648 29929 11676
rect 29880 11636 29886 11648
rect 29917 11645 29929 11648
rect 29963 11645 29975 11679
rect 29917 11639 29975 11645
rect 33965 11679 34023 11685
rect 33965 11645 33977 11679
rect 34011 11645 34023 11679
rect 33965 11639 34023 11645
rect 28074 11568 28080 11620
rect 28132 11608 28138 11620
rect 28169 11611 28227 11617
rect 28169 11608 28181 11611
rect 28132 11580 28181 11608
rect 28132 11568 28138 11580
rect 28169 11577 28181 11580
rect 28215 11608 28227 11611
rect 29730 11608 29736 11620
rect 28215 11580 29736 11608
rect 28215 11577 28227 11580
rect 28169 11571 28227 11577
rect 29730 11568 29736 11580
rect 29788 11568 29794 11620
rect 33980 11608 34008 11639
rect 34698 11636 34704 11688
rect 34756 11636 34762 11688
rect 34790 11636 34796 11688
rect 34848 11676 34854 11688
rect 35526 11676 35532 11688
rect 34848 11648 35532 11676
rect 34848 11636 34854 11648
rect 35526 11636 35532 11648
rect 35584 11636 35590 11688
rect 37182 11636 37188 11688
rect 37240 11636 37246 11688
rect 37458 11636 37464 11688
rect 37516 11676 37522 11688
rect 37844 11685 37872 11716
rect 37737 11679 37795 11685
rect 37737 11676 37749 11679
rect 37516 11648 37749 11676
rect 37516 11636 37522 11648
rect 37737 11645 37749 11648
rect 37783 11645 37795 11679
rect 37737 11639 37795 11645
rect 37829 11679 37887 11685
rect 37829 11645 37841 11679
rect 37875 11645 37887 11679
rect 37829 11639 37887 11645
rect 36909 11611 36967 11617
rect 33980 11580 35572 11608
rect 25590 11540 25596 11552
rect 25424 11512 25596 11540
rect 24397 11503 24455 11509
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 26973 11543 27031 11549
rect 26973 11509 26985 11543
rect 27019 11540 27031 11543
rect 28258 11540 28264 11552
rect 27019 11512 28264 11540
rect 27019 11509 27031 11512
rect 26973 11503 27031 11509
rect 28258 11500 28264 11512
rect 28316 11500 28322 11552
rect 31297 11543 31355 11549
rect 31297 11509 31309 11543
rect 31343 11540 31355 11543
rect 31846 11540 31852 11552
rect 31343 11512 31852 11540
rect 31343 11509 31355 11512
rect 31297 11503 31355 11509
rect 31846 11500 31852 11512
rect 31904 11500 31910 11552
rect 35253 11543 35311 11549
rect 35253 11509 35265 11543
rect 35299 11540 35311 11543
rect 35342 11540 35348 11552
rect 35299 11512 35348 11540
rect 35299 11509 35311 11512
rect 35253 11503 35311 11509
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 35544 11540 35572 11580
rect 36909 11577 36921 11611
rect 36955 11608 36967 11611
rect 37366 11608 37372 11620
rect 36955 11580 37372 11608
rect 36955 11577 36967 11580
rect 36909 11571 36967 11577
rect 37366 11568 37372 11580
rect 37424 11568 37430 11620
rect 37752 11608 37780 11639
rect 37918 11636 37924 11688
rect 37976 11636 37982 11688
rect 37936 11608 37964 11636
rect 37752 11580 37964 11608
rect 37090 11540 37096 11552
rect 35544 11512 37096 11540
rect 37090 11500 37096 11512
rect 37148 11500 37154 11552
rect 37277 11543 37335 11549
rect 37277 11509 37289 11543
rect 37323 11540 37335 11543
rect 37826 11540 37832 11552
rect 37323 11512 37832 11540
rect 37323 11509 37335 11512
rect 37277 11503 37335 11509
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1489 11339 1547 11345
rect 1489 11305 1501 11339
rect 1535 11336 1547 11339
rect 1854 11336 1860 11348
rect 1535 11308 1860 11336
rect 1535 11305 1547 11308
rect 1489 11299 1547 11305
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 4948 11308 5825 11336
rect 4948 11296 4954 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 6181 11339 6239 11345
rect 6181 11305 6193 11339
rect 6227 11336 6239 11339
rect 6362 11336 6368 11348
rect 6227 11308 6368 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6546 11296 6552 11348
rect 6604 11296 6610 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 8294 11336 8300 11348
rect 6788 11308 8300 11336
rect 6788 11296 6794 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 8754 11296 8760 11348
rect 8812 11336 8818 11348
rect 9214 11336 9220 11348
rect 8812 11308 9220 11336
rect 8812 11296 8818 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 9456 11308 10609 11336
rect 9456 11296 9462 11308
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 11974 11336 11980 11348
rect 10597 11299 10655 11305
rect 11072 11308 11980 11336
rect 5258 11228 5264 11280
rect 5316 11268 5322 11280
rect 5353 11271 5411 11277
rect 5353 11268 5365 11271
rect 5316 11240 5365 11268
rect 5316 11228 5322 11240
rect 5353 11237 5365 11240
rect 5399 11237 5411 11271
rect 5353 11231 5411 11237
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 5721 11271 5779 11277
rect 5721 11268 5733 11271
rect 5592 11240 5733 11268
rect 5592 11228 5598 11240
rect 5721 11237 5733 11240
rect 5767 11237 5779 11271
rect 5721 11231 5779 11237
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 6564 11200 6592 11296
rect 8404 11268 8432 11296
rect 8938 11268 8944 11280
rect 8404 11240 8944 11268
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 11072 11209 11100 11308
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 12986 11336 12992 11348
rect 12575 11308 12992 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 12986 11296 12992 11308
rect 13044 11336 13050 11348
rect 14829 11339 14887 11345
rect 13044 11308 14320 11336
rect 13044 11296 13050 11308
rect 14090 11268 14096 11280
rect 13924 11240 14096 11268
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6564 11172 6653 11200
rect 5905 11163 5963 11169
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10367 11172 11069 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 13924 11200 13952 11240
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 11057 11163 11115 11169
rect 13832 11172 13952 11200
rect 2038 11092 2044 11144
rect 2096 11092 2102 11144
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2774 11132 2780 11144
rect 2271 11104 2780 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2774 11092 2780 11104
rect 2832 11132 2838 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 2832 11104 3801 11132
rect 2832 11092 2838 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 2492 11067 2550 11073
rect 2492 11033 2504 11067
rect 2538 11064 2550 11067
rect 2590 11064 2596 11076
rect 2538 11036 2596 11064
rect 2538 11033 2550 11036
rect 2492 11027 2550 11033
rect 2590 11024 2596 11036
rect 2648 11024 2654 11076
rect 3326 11024 3332 11076
rect 3384 11064 3390 11076
rect 4034 11067 4092 11073
rect 4034 11064 4046 11067
rect 3384 11036 4046 11064
rect 3384 11024 3390 11036
rect 4034 11033 4046 11036
rect 4080 11033 4092 11067
rect 5920 11064 5948 11163
rect 7190 11092 7196 11144
rect 7248 11132 7254 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7248 11104 7389 11132
rect 7248 11092 7254 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 13653 11135 13711 11141
rect 13653 11101 13665 11135
rect 13699 11132 13711 11135
rect 13832 11132 13860 11172
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 14056 11172 14197 11200
rect 14056 11160 14062 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14292 11200 14320 11308
rect 14829 11305 14841 11339
rect 14875 11336 14887 11339
rect 14918 11336 14924 11348
rect 14875 11308 14924 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15160 11308 15945 11336
rect 15160 11296 15166 11308
rect 15933 11305 15945 11308
rect 15979 11336 15991 11339
rect 16574 11336 16580 11348
rect 15979 11308 16580 11336
rect 15979 11305 15991 11308
rect 15933 11299 15991 11305
rect 16574 11296 16580 11308
rect 16632 11336 16638 11348
rect 17126 11336 17132 11348
rect 16632 11308 17132 11336
rect 16632 11296 16638 11308
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21726 11336 21732 11348
rect 21232 11308 21732 11336
rect 21232 11296 21238 11308
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 21913 11339 21971 11345
rect 21913 11305 21925 11339
rect 21959 11336 21971 11339
rect 22554 11336 22560 11348
rect 21959 11308 22560 11336
rect 21959 11305 21971 11308
rect 21913 11299 21971 11305
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 24912 11308 25053 11336
rect 24912 11296 24918 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 27433 11339 27491 11345
rect 27433 11305 27445 11339
rect 27479 11336 27491 11339
rect 28810 11336 28816 11348
rect 27479 11308 28816 11336
rect 27479 11305 27491 11308
rect 27433 11299 27491 11305
rect 28810 11296 28816 11308
rect 28868 11296 28874 11348
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29089 11339 29147 11345
rect 29089 11336 29101 11339
rect 29052 11308 29101 11336
rect 29052 11296 29058 11308
rect 29089 11305 29101 11308
rect 29135 11305 29147 11339
rect 29089 11299 29147 11305
rect 30101 11339 30159 11345
rect 30101 11305 30113 11339
rect 30147 11336 30159 11339
rect 31110 11336 31116 11348
rect 30147 11308 31116 11336
rect 30147 11305 30159 11308
rect 30101 11299 30159 11305
rect 31110 11296 31116 11308
rect 31168 11296 31174 11348
rect 31294 11296 31300 11348
rect 31352 11336 31358 11348
rect 32766 11336 32772 11348
rect 31352 11308 32772 11336
rect 31352 11296 31358 11308
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 33502 11296 33508 11348
rect 33560 11296 33566 11348
rect 34698 11296 34704 11348
rect 34756 11296 34762 11348
rect 35529 11339 35587 11345
rect 35529 11305 35541 11339
rect 35575 11336 35587 11339
rect 37642 11336 37648 11348
rect 35575 11308 37648 11336
rect 35575 11305 35587 11308
rect 35529 11299 35587 11305
rect 37642 11296 37648 11308
rect 37700 11296 37706 11348
rect 38286 11296 38292 11348
rect 38344 11296 38350 11348
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 19521 11271 19579 11277
rect 19521 11268 19533 11271
rect 16264 11240 19533 11268
rect 16264 11228 16270 11240
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 14292 11172 15485 11200
rect 14185 11163 14243 11169
rect 15473 11169 15485 11172
rect 15519 11169 15531 11203
rect 15473 11163 15531 11169
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 18064 11209 18092 11240
rect 19521 11237 19533 11240
rect 19567 11268 19579 11271
rect 22278 11268 22284 11280
rect 19567 11240 22284 11268
rect 19567 11237 19579 11240
rect 19521 11231 19579 11237
rect 22278 11228 22284 11240
rect 22336 11228 22342 11280
rect 27341 11271 27399 11277
rect 27341 11237 27353 11271
rect 27387 11268 27399 11271
rect 27798 11268 27804 11280
rect 27387 11240 27804 11268
rect 27387 11237 27399 11240
rect 27341 11231 27399 11237
rect 27798 11228 27804 11240
rect 27856 11228 27862 11280
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 16724 11172 17601 11200
rect 16724 11160 16730 11172
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 23290 11160 23296 11212
rect 23348 11200 23354 11212
rect 25590 11200 25596 11212
rect 23348 11172 25596 11200
rect 23348 11160 23354 11172
rect 25590 11160 25596 11172
rect 25648 11200 25654 11212
rect 25961 11203 26019 11209
rect 25961 11200 25973 11203
rect 25648 11172 25973 11200
rect 25648 11160 25654 11172
rect 25961 11169 25973 11172
rect 26007 11169 26019 11203
rect 25961 11163 26019 11169
rect 28813 11203 28871 11209
rect 28813 11169 28825 11203
rect 28859 11200 28871 11203
rect 29822 11200 29828 11212
rect 28859 11172 29828 11200
rect 28859 11169 28871 11172
rect 28813 11163 28871 11169
rect 29822 11160 29828 11172
rect 29880 11160 29886 11212
rect 32953 11203 33011 11209
rect 32953 11169 32965 11203
rect 32999 11200 33011 11203
rect 33520 11200 33548 11296
rect 34238 11228 34244 11280
rect 34296 11268 34302 11280
rect 35710 11268 35716 11280
rect 34296 11240 35716 11268
rect 34296 11228 34302 11240
rect 35710 11228 35716 11240
rect 35768 11228 35774 11280
rect 36725 11271 36783 11277
rect 36725 11237 36737 11271
rect 36771 11268 36783 11271
rect 36771 11240 36952 11268
rect 36771 11237 36783 11240
rect 36725 11231 36783 11237
rect 32999 11172 33548 11200
rect 33873 11203 33931 11209
rect 32999 11169 33011 11172
rect 32953 11163 33011 11169
rect 33873 11169 33885 11203
rect 33919 11200 33931 11203
rect 33962 11200 33968 11212
rect 33919 11172 33968 11200
rect 33919 11169 33931 11172
rect 33873 11163 33931 11169
rect 33962 11160 33968 11172
rect 34020 11160 34026 11212
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 35253 11203 35311 11209
rect 35253 11200 35265 11203
rect 34572 11172 35265 11200
rect 34572 11160 34578 11172
rect 35253 11169 35265 11172
rect 35299 11169 35311 11203
rect 35253 11163 35311 11169
rect 36187 11203 36245 11209
rect 36187 11169 36199 11203
rect 36233 11200 36245 11203
rect 36814 11200 36820 11212
rect 36233 11172 36820 11200
rect 36233 11169 36245 11172
rect 36187 11163 36245 11169
rect 36814 11160 36820 11172
rect 36872 11160 36878 11212
rect 36924 11200 36952 11240
rect 37090 11228 37096 11280
rect 37148 11268 37154 11280
rect 37461 11271 37519 11277
rect 37461 11268 37473 11271
rect 37148 11240 37473 11268
rect 37148 11228 37154 11240
rect 37461 11237 37473 11240
rect 37507 11237 37519 11271
rect 37461 11231 37519 11237
rect 36998 11200 37004 11212
rect 36924 11172 37004 11200
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 37366 11160 37372 11212
rect 37424 11160 37430 11212
rect 38105 11203 38163 11209
rect 38105 11169 38117 11203
rect 38151 11200 38163 11203
rect 38304 11200 38332 11296
rect 38151 11172 38332 11200
rect 38151 11169 38163 11172
rect 38105 11163 38163 11169
rect 13699 11104 13860 11132
rect 13909 11135 13967 11141
rect 13699 11101 13711 11104
rect 13653 11095 13711 11101
rect 13909 11101 13921 11135
rect 13955 11132 13967 11135
rect 14274 11132 14280 11144
rect 13955 11104 14280 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14507 11104 15424 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 15396 11076 15424 11104
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17552 11104 18245 11132
rect 17552 11092 17558 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 19260 11104 21956 11132
rect 19260 11076 19288 11104
rect 4034 11027 4092 11033
rect 5184 11036 5948 11064
rect 7285 11067 7343 11073
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 3418 10996 3424 11008
rect 1728 10968 3424 10996
rect 1728 10956 1734 10968
rect 3418 10956 3424 10968
rect 3476 10956 3482 11008
rect 3602 10956 3608 11008
rect 3660 10956 3666 11008
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 5184 11005 5212 11036
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 7622 11067 7680 11073
rect 7622 11064 7634 11067
rect 7331 11036 7634 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 7622 11033 7634 11036
rect 7668 11033 7680 11067
rect 7622 11027 7680 11033
rect 10042 11024 10048 11076
rect 10100 11073 10106 11076
rect 10100 11027 10112 11073
rect 11324 11067 11382 11073
rect 11324 11033 11336 11067
rect 11370 11064 11382 11067
rect 11514 11064 11520 11076
rect 11370 11036 11520 11064
rect 11370 11033 11382 11036
rect 11324 11027 11382 11033
rect 10100 11024 10106 11027
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13814 11064 13820 11076
rect 13504 11036 13820 11064
rect 13504 11024 13510 11036
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14369 11067 14427 11073
rect 14369 11033 14381 11067
rect 14415 11064 14427 11067
rect 14921 11067 14979 11073
rect 14921 11064 14933 11067
rect 14415 11036 14933 11064
rect 14415 11033 14427 11036
rect 14369 11027 14427 11033
rect 14921 11033 14933 11036
rect 14967 11033 14979 11067
rect 14921 11027 14979 11033
rect 15378 11024 15384 11076
rect 15436 11024 15442 11076
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16025 11067 16083 11073
rect 16025 11064 16037 11067
rect 15896 11036 16037 11064
rect 15896 11024 15902 11036
rect 16025 11033 16037 11036
rect 16071 11033 16083 11067
rect 16025 11027 16083 11033
rect 18874 11024 18880 11076
rect 18932 11064 18938 11076
rect 19242 11064 19248 11076
rect 18932 11036 19248 11064
rect 18932 11024 18938 11036
rect 19242 11024 19248 11036
rect 19300 11024 19306 11076
rect 21928 11064 21956 11104
rect 22002 11092 22008 11144
rect 22060 11132 22066 11144
rect 22060 11104 22968 11132
rect 22060 11092 22066 11104
rect 22940 11064 22968 11104
rect 23014 11092 23020 11144
rect 23072 11141 23078 11144
rect 23072 11095 23084 11141
rect 23072 11092 23078 11095
rect 23198 11092 23204 11144
rect 23256 11132 23262 11144
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 23256 11104 24409 11132
rect 23256 11092 23262 11104
rect 24397 11101 24409 11104
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 25498 11092 25504 11144
rect 25556 11132 25562 11144
rect 25777 11135 25835 11141
rect 25777 11132 25789 11135
rect 25556 11104 25789 11132
rect 25556 11092 25562 11104
rect 25777 11101 25789 11104
rect 25823 11132 25835 11135
rect 26050 11132 26056 11144
rect 25823 11104 26056 11132
rect 25823 11101 25835 11104
rect 25777 11095 25835 11101
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 26234 11141 26240 11144
rect 26228 11095 26240 11141
rect 26234 11092 26240 11095
rect 26292 11092 26298 11144
rect 28557 11135 28615 11141
rect 28557 11101 28569 11135
rect 28603 11132 28615 11135
rect 29086 11132 29092 11144
rect 28603 11104 29092 11132
rect 28603 11101 28615 11104
rect 28557 11095 28615 11101
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 31202 11092 31208 11144
rect 31260 11141 31266 11144
rect 31260 11132 31272 11141
rect 31481 11135 31539 11141
rect 31260 11104 31305 11132
rect 31260 11095 31272 11104
rect 31481 11101 31493 11135
rect 31527 11132 31539 11135
rect 31938 11132 31944 11144
rect 31527 11104 31944 11132
rect 31527 11101 31539 11104
rect 31481 11095 31539 11101
rect 31260 11092 31266 11095
rect 31938 11092 31944 11104
rect 31996 11092 32002 11144
rect 32398 11132 32404 11144
rect 32048 11104 32404 11132
rect 21928 11036 22876 11064
rect 22940 11036 23888 11064
rect 5169 10999 5227 11005
rect 5169 10996 5181 10999
rect 4856 10968 5181 10996
rect 4856 10956 4862 10968
rect 5169 10965 5181 10968
rect 5215 10965 5227 10999
rect 5169 10959 5227 10965
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 14090 10996 14096 11008
rect 12492 10968 14096 10996
rect 12492 10956 12498 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 18138 10956 18144 11008
rect 18196 10956 18202 11008
rect 18598 10956 18604 11008
rect 18656 10956 18662 11008
rect 22848 10996 22876 11036
rect 23382 10996 23388 11008
rect 22848 10968 23388 10996
rect 23382 10956 23388 10968
rect 23440 10996 23446 11008
rect 23860 11005 23888 11036
rect 23934 11024 23940 11076
rect 23992 11024 23998 11076
rect 25222 11024 25228 11076
rect 25280 11064 25286 11076
rect 25317 11067 25375 11073
rect 25317 11064 25329 11067
rect 25280 11036 25329 11064
rect 25280 11024 25286 11036
rect 25317 11033 25329 11036
rect 25363 11033 25375 11067
rect 28074 11064 28080 11076
rect 25317 11027 25375 11033
rect 26804 11036 28080 11064
rect 26804 11008 26832 11036
rect 28074 11024 28080 11036
rect 28132 11024 28138 11076
rect 32048 11064 32076 11104
rect 32398 11092 32404 11104
rect 32456 11132 32462 11144
rect 36354 11141 36360 11144
rect 33597 11135 33655 11141
rect 33597 11132 33609 11135
rect 32456 11104 33609 11132
rect 32456 11092 32462 11104
rect 33597 11101 33609 11104
rect 33643 11101 33655 11135
rect 33597 11095 33655 11101
rect 36311 11135 36360 11141
rect 36311 11101 36323 11135
rect 36357 11101 36360 11135
rect 36311 11095 36360 11101
rect 36354 11092 36360 11095
rect 36412 11092 36418 11144
rect 36446 11092 36452 11144
rect 36504 11092 36510 11144
rect 37185 11135 37243 11141
rect 37185 11101 37197 11135
rect 37231 11132 37243 11135
rect 37458 11132 37464 11144
rect 37231 11104 37464 11132
rect 37231 11101 37243 11104
rect 37185 11095 37243 11101
rect 37458 11092 37464 11104
rect 37516 11092 37522 11144
rect 37918 11092 37924 11144
rect 37976 11092 37982 11144
rect 31588 11036 32076 11064
rect 32708 11067 32766 11073
rect 23569 10999 23627 11005
rect 23569 10996 23581 10999
rect 23440 10968 23581 10996
rect 23440 10956 23446 10968
rect 23569 10965 23581 10968
rect 23615 10965 23627 10999
rect 23569 10959 23627 10965
rect 23845 10999 23903 11005
rect 23845 10965 23857 10999
rect 23891 10965 23903 10999
rect 23845 10959 23903 10965
rect 26786 10956 26792 11008
rect 26844 10956 26850 11008
rect 31588 11005 31616 11036
rect 32708 11033 32720 11067
rect 32754 11064 32766 11067
rect 32950 11064 32956 11076
rect 32754 11036 32956 11064
rect 32754 11033 32766 11036
rect 32708 11027 32766 11033
rect 32950 11024 32956 11036
rect 33008 11024 33014 11076
rect 34517 11067 34575 11073
rect 34517 11033 34529 11067
rect 34563 11064 34575 11067
rect 35069 11067 35127 11073
rect 35069 11064 35081 11067
rect 34563 11036 35081 11064
rect 34563 11033 34575 11036
rect 34517 11027 34575 11033
rect 35069 11033 35081 11036
rect 35115 11033 35127 11067
rect 35069 11027 35127 11033
rect 35161 11067 35219 11073
rect 35161 11033 35173 11067
rect 35207 11064 35219 11067
rect 37829 11067 37887 11073
rect 37829 11064 37841 11067
rect 35207 11036 35756 11064
rect 35207 11033 35219 11036
rect 35161 11027 35219 11033
rect 31573 10999 31631 11005
rect 31573 10965 31585 10999
rect 31619 10965 31631 10999
rect 31573 10959 31631 10965
rect 33042 10956 33048 11008
rect 33100 10956 33106 11008
rect 35728 10996 35756 11036
rect 37200 11036 37841 11064
rect 36078 10996 36084 11008
rect 35728 10968 36084 10996
rect 36078 10956 36084 10968
rect 36136 10996 36142 11008
rect 37200 10996 37228 11036
rect 37829 11033 37841 11036
rect 37875 11064 37887 11067
rect 37936 11064 37964 11092
rect 38654 11064 38660 11076
rect 37875 11036 38660 11064
rect 37875 11033 37887 11036
rect 37829 11027 37887 11033
rect 38654 11024 38660 11036
rect 38712 11024 38718 11076
rect 36136 10968 37228 10996
rect 36136 10956 36142 10968
rect 37918 10956 37924 11008
rect 37976 10956 37982 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1670 10752 1676 10804
rect 1728 10752 1734 10804
rect 2038 10752 2044 10804
rect 2096 10752 2102 10804
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 3234 10792 3240 10804
rect 2372 10764 3240 10792
rect 2372 10752 2378 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 3326 10752 3332 10804
rect 3384 10752 3390 10804
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4706 10792 4712 10804
rect 4111 10764 4712 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5074 10792 5080 10804
rect 4816 10764 5080 10792
rect 1946 10684 1952 10736
rect 2004 10684 2010 10736
rect 3418 10684 3424 10736
rect 3476 10724 3482 10736
rect 4816 10724 4844 10764
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5258 10752 5264 10804
rect 5316 10752 5322 10804
rect 5350 10752 5356 10804
rect 5408 10752 5414 10804
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6822 10792 6828 10804
rect 6043 10764 6828 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 6972 10764 7757 10792
rect 6972 10752 6978 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 7926 10752 7932 10804
rect 7984 10752 7990 10804
rect 8478 10752 8484 10804
rect 8536 10752 8542 10804
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 9030 10792 9036 10804
rect 8987 10764 9036 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10100 10764 10149 10792
rect 10100 10752 10106 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 11514 10752 11520 10804
rect 11572 10752 11578 10804
rect 12897 10795 12955 10801
rect 12897 10761 12909 10795
rect 12943 10792 12955 10795
rect 13078 10792 13084 10804
rect 12943 10764 13084 10792
rect 12943 10761 12955 10764
rect 12897 10755 12955 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 16945 10795 17003 10801
rect 13188 10764 16344 10792
rect 5276 10724 5304 10752
rect 5629 10727 5687 10733
rect 5629 10724 5641 10727
rect 3476 10696 4844 10724
rect 5092 10696 5641 10724
rect 3476 10684 3482 10696
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 3142 10656 3148 10668
rect 1811 10628 3148 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3568 10659 3626 10665
rect 3568 10656 3580 10659
rect 3200 10628 3580 10656
rect 3200 10616 3206 10628
rect 3568 10625 3580 10628
rect 3614 10656 3626 10659
rect 3614 10625 3648 10656
rect 3568 10619 3648 10625
rect 2222 10548 2228 10600
rect 2280 10548 2286 10600
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10557 2375 10591
rect 2317 10551 2375 10557
rect 2332 10520 2360 10551
rect 2406 10548 2412 10600
rect 2464 10548 2470 10600
rect 2498 10548 2504 10600
rect 2556 10548 2562 10600
rect 2682 10548 2688 10600
rect 2740 10548 2746 10600
rect 2866 10520 2872 10532
rect 2332 10492 2872 10520
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 3620 10452 3648 10619
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 3752 10628 3832 10656
rect 3752 10616 3758 10628
rect 3804 10597 3832 10628
rect 4798 10616 4804 10668
rect 4856 10616 4862 10668
rect 5092 10665 5120 10696
rect 5629 10693 5641 10696
rect 5675 10693 5687 10727
rect 5629 10687 5687 10693
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10693 5871 10727
rect 5813 10687 5871 10693
rect 7653 10727 7711 10733
rect 7653 10693 7665 10727
rect 7699 10724 7711 10727
rect 7944 10724 7972 10752
rect 7699 10696 7972 10724
rect 7699 10693 7711 10696
rect 7653 10687 7711 10693
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5077 10619 5135 10625
rect 5184 10628 5549 10656
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10557 3847 10591
rect 3789 10551 3847 10557
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4706 10520 4712 10532
rect 3743 10492 4712 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 4706 10480 4712 10492
rect 4764 10520 4770 10532
rect 4816 10520 4844 10616
rect 5184 10600 5212 10628
rect 5537 10625 5549 10628
rect 5583 10656 5595 10659
rect 5828 10656 5856 10687
rect 5583 10628 5856 10656
rect 8389 10659 8447 10665
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8754 10656 8760 10668
rect 8435 10628 8760 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 8849 10619 8907 10625
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 8864 10588 8892 10619
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9401 10659 9459 10665
rect 9401 10656 9413 10659
rect 8996 10628 9413 10656
rect 8996 10616 9002 10628
rect 9401 10625 9413 10628
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10192 10628 10701 10656
rect 10192 10616 10198 10628
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10656 12403 10659
rect 12434 10656 12440 10668
rect 12391 10628 12440 10656
rect 12391 10625 12403 10628
rect 12345 10619 12403 10625
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13188 10600 13216 10764
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 16316 10665 16344 10764
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17586 10792 17592 10804
rect 16991 10764 17592 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 18414 10752 18420 10804
rect 18472 10752 18478 10804
rect 22186 10752 22192 10804
rect 22244 10752 22250 10804
rect 22646 10752 22652 10804
rect 22704 10792 22710 10804
rect 23293 10795 23351 10801
rect 23293 10792 23305 10795
rect 22704 10764 23305 10792
rect 22704 10752 22710 10764
rect 23293 10761 23305 10764
rect 23339 10761 23351 10795
rect 23293 10755 23351 10761
rect 23474 10752 23480 10804
rect 23532 10752 23538 10804
rect 23842 10752 23848 10804
rect 23900 10792 23906 10804
rect 24210 10792 24216 10804
rect 23900 10764 24216 10792
rect 23900 10752 23906 10764
rect 24210 10752 24216 10764
rect 24268 10752 24274 10804
rect 26142 10752 26148 10804
rect 26200 10752 26206 10804
rect 27614 10752 27620 10804
rect 27672 10792 27678 10804
rect 28169 10795 28227 10801
rect 28169 10792 28181 10795
rect 27672 10764 28181 10792
rect 27672 10752 27678 10764
rect 28169 10761 28181 10764
rect 28215 10761 28227 10795
rect 28169 10755 28227 10761
rect 28258 10752 28264 10804
rect 28316 10752 28322 10804
rect 29270 10752 29276 10804
rect 29328 10752 29334 10804
rect 29825 10795 29883 10801
rect 29825 10761 29837 10795
rect 29871 10792 29883 10795
rect 30190 10792 30196 10804
rect 29871 10764 30196 10792
rect 29871 10761 29883 10764
rect 29825 10755 29883 10761
rect 30190 10752 30196 10764
rect 30248 10752 30254 10804
rect 30466 10752 30472 10804
rect 30524 10752 30530 10804
rect 30929 10795 30987 10801
rect 30929 10761 30941 10795
rect 30975 10792 30987 10795
rect 31018 10792 31024 10804
rect 30975 10764 31024 10792
rect 30975 10761 30987 10764
rect 30929 10755 30987 10761
rect 31018 10752 31024 10764
rect 31076 10752 31082 10804
rect 32493 10795 32551 10801
rect 32493 10761 32505 10795
rect 32539 10792 32551 10795
rect 33042 10792 33048 10804
rect 32539 10764 33048 10792
rect 32539 10761 32551 10764
rect 32493 10755 32551 10761
rect 33042 10752 33048 10764
rect 33100 10752 33106 10804
rect 33962 10752 33968 10804
rect 34020 10792 34026 10804
rect 34241 10795 34299 10801
rect 34241 10792 34253 10795
rect 34020 10764 34253 10792
rect 34020 10752 34026 10764
rect 34241 10761 34253 10764
rect 34287 10761 34299 10795
rect 34241 10755 34299 10761
rect 34624 10764 35572 10792
rect 22370 10684 22376 10736
rect 22428 10724 22434 10736
rect 22557 10727 22615 10733
rect 22557 10724 22569 10727
rect 22428 10696 22569 10724
rect 22428 10684 22434 10696
rect 22557 10693 22569 10696
rect 22603 10724 22615 10727
rect 23382 10724 23388 10736
rect 22603 10696 23388 10724
rect 22603 10693 22615 10696
rect 22557 10687 22615 10693
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15335 10628 15761 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16666 10616 16672 10668
rect 16724 10656 16730 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16724 10628 17049 10656
rect 16724 10616 16730 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17304 10659 17362 10665
rect 17304 10625 17316 10659
rect 17350 10656 17362 10659
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 17350 10628 18521 10656
rect 17350 10625 17362 10628
rect 17304 10619 17362 10625
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 18690 10616 18696 10668
rect 18748 10656 18754 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 18748 10628 19073 10656
rect 18748 10616 18754 10628
rect 19061 10625 19073 10628
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 23492 10656 23520 10752
rect 29917 10727 29975 10733
rect 29917 10693 29929 10727
rect 29963 10724 29975 10727
rect 32306 10724 32312 10736
rect 29963 10696 32312 10724
rect 29963 10693 29975 10696
rect 29917 10687 29975 10693
rect 32306 10684 32312 10696
rect 32364 10684 32370 10736
rect 32950 10684 32956 10736
rect 33008 10684 33014 10736
rect 22695 10628 23520 10656
rect 23937 10659 23995 10665
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 23937 10625 23949 10659
rect 23983 10656 23995 10659
rect 24394 10656 24400 10668
rect 23983 10628 24400 10656
rect 23983 10625 23995 10628
rect 23937 10619 23995 10625
rect 24394 10616 24400 10628
rect 24452 10616 24458 10668
rect 27338 10616 27344 10668
rect 27396 10616 27402 10668
rect 27430 10616 27436 10668
rect 27488 10656 27494 10668
rect 27488 10628 28304 10656
rect 27488 10616 27494 10628
rect 9125 10591 9183 10597
rect 8864 10560 9076 10588
rect 9048 10520 9076 10560
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9858 10588 9864 10600
rect 9171 10560 9864 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 10502 10588 10508 10600
rect 10091 10560 10508 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10557 12219 10591
rect 12710 10588 12716 10600
rect 12161 10551 12219 10557
rect 12406 10560 12716 10588
rect 9582 10520 9588 10532
rect 4764 10492 5856 10520
rect 4764 10480 4770 10492
rect 4798 10452 4804 10464
rect 3620 10424 4804 10452
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5828 10461 5856 10492
rect 9048 10492 9588 10520
rect 9048 10464 9076 10492
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 12176 10520 12204 10551
rect 12406 10520 12434 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 12986 10548 12992 10600
rect 13044 10548 13050 10600
rect 13170 10548 13176 10600
rect 13228 10548 13234 10600
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14090 10597 14096 10600
rect 14047 10591 14096 10597
rect 14047 10557 14059 10591
rect 14093 10557 14096 10591
rect 14047 10551 14096 10557
rect 14090 10548 14096 10551
rect 14148 10548 14154 10600
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 15120 10588 15148 10616
rect 28276 10600 28304 10628
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 30837 10659 30895 10665
rect 30837 10625 30849 10659
rect 30883 10656 30895 10659
rect 31297 10659 31355 10665
rect 31297 10656 31309 10659
rect 30883 10628 31309 10656
rect 30883 10625 30895 10628
rect 30837 10619 30895 10625
rect 31297 10625 31309 10628
rect 31343 10625 31355 10659
rect 31297 10619 31355 10625
rect 31846 10616 31852 10668
rect 31904 10616 31910 10668
rect 34057 10659 34115 10665
rect 34057 10656 34069 10659
rect 32140 10628 34069 10656
rect 14240 10560 15148 10588
rect 14240 10548 14246 10560
rect 15378 10548 15384 10600
rect 15436 10548 15442 10600
rect 15562 10548 15568 10600
rect 15620 10548 15626 10600
rect 22833 10591 22891 10597
rect 22833 10557 22845 10591
rect 22879 10588 22891 10591
rect 23014 10588 23020 10600
rect 22879 10560 23020 10588
rect 22879 10557 22891 10560
rect 22833 10551 22891 10557
rect 23014 10548 23020 10560
rect 23072 10548 23078 10600
rect 26789 10591 26847 10597
rect 26789 10557 26801 10591
rect 26835 10557 26847 10591
rect 27525 10591 27583 10597
rect 27525 10588 27537 10591
rect 26789 10551 26847 10557
rect 27080 10560 27537 10588
rect 12176 10492 12434 10520
rect 12802 10480 12808 10532
rect 12860 10520 12866 10532
rect 13633 10523 13691 10529
rect 13633 10520 13645 10523
rect 12860 10492 13645 10520
rect 12860 10480 12866 10492
rect 13633 10489 13645 10492
rect 13679 10489 13691 10523
rect 13633 10483 13691 10489
rect 14829 10523 14887 10529
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 16022 10520 16028 10532
rect 14875 10492 16028 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 26804 10520 26832 10551
rect 26973 10523 27031 10529
rect 26973 10520 26985 10523
rect 26804 10492 26985 10520
rect 26973 10489 26985 10492
rect 27019 10489 27031 10523
rect 26973 10483 27031 10489
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10421 5871 10455
rect 5813 10415 5871 10421
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6822 10452 6828 10464
rect 6052 10424 6828 10452
rect 6052 10412 6058 10424
rect 6822 10412 6828 10424
rect 6880 10452 6886 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 6880 10424 7205 10452
rect 6880 10412 6886 10424
rect 7193 10421 7205 10424
rect 7239 10452 7251 10455
rect 8570 10452 8576 10464
rect 7239 10424 8576 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9030 10412 9036 10464
rect 9088 10412 9094 10464
rect 14918 10412 14924 10464
rect 14976 10412 14982 10464
rect 24670 10412 24676 10464
rect 24728 10412 24734 10464
rect 25038 10412 25044 10464
rect 25096 10452 25102 10464
rect 25961 10455 26019 10461
rect 25961 10452 25973 10455
rect 25096 10424 25973 10452
rect 25096 10412 25102 10424
rect 25961 10421 25973 10424
rect 26007 10452 26019 10455
rect 27080 10452 27108 10560
rect 27525 10557 27537 10560
rect 27571 10557 27583 10591
rect 27525 10551 27583 10557
rect 27540 10520 27568 10551
rect 28258 10548 28264 10600
rect 28316 10548 28322 10600
rect 28350 10548 28356 10600
rect 28408 10548 28414 10600
rect 31021 10591 31079 10597
rect 31021 10588 31033 10591
rect 30576 10560 31033 10588
rect 30466 10520 30472 10532
rect 27540 10492 30472 10520
rect 30466 10480 30472 10492
rect 30524 10480 30530 10532
rect 26007 10424 27108 10452
rect 26007 10421 26019 10424
rect 25961 10415 26019 10421
rect 27798 10412 27804 10464
rect 27856 10412 27862 10464
rect 29362 10412 29368 10464
rect 29420 10452 29426 10464
rect 30282 10452 30288 10464
rect 29420 10424 30288 10452
rect 29420 10412 29426 10424
rect 30282 10412 30288 10424
rect 30340 10452 30346 10464
rect 30377 10455 30435 10461
rect 30377 10452 30389 10455
rect 30340 10424 30389 10452
rect 30340 10412 30346 10424
rect 30377 10421 30389 10424
rect 30423 10452 30435 10455
rect 30576 10452 30604 10560
rect 31021 10557 31033 10560
rect 31067 10588 31079 10591
rect 32140 10588 32168 10628
rect 34057 10625 34069 10628
rect 34103 10656 34115 10659
rect 34514 10656 34520 10668
rect 34103 10628 34520 10656
rect 34103 10625 34115 10628
rect 34057 10619 34115 10625
rect 34514 10616 34520 10628
rect 34572 10616 34578 10668
rect 31067 10560 32168 10588
rect 31067 10557 31079 10560
rect 31021 10551 31079 10557
rect 32214 10548 32220 10600
rect 32272 10548 32278 10600
rect 32398 10548 32404 10600
rect 32456 10548 32462 10600
rect 33505 10591 33563 10597
rect 33505 10588 33517 10591
rect 32876 10560 33517 10588
rect 32416 10520 32444 10548
rect 32876 10529 32904 10560
rect 33505 10557 33517 10560
rect 33551 10557 33563 10591
rect 34624 10588 34652 10764
rect 35342 10684 35348 10736
rect 35400 10733 35406 10736
rect 35400 10724 35412 10733
rect 35544 10724 35572 10764
rect 36078 10752 36084 10804
rect 36136 10752 36142 10804
rect 36817 10795 36875 10801
rect 36817 10761 36829 10795
rect 36863 10792 36875 10795
rect 36998 10792 37004 10804
rect 36863 10764 37004 10792
rect 36863 10761 36875 10764
rect 36817 10755 36875 10761
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 37550 10752 37556 10804
rect 37608 10752 37614 10804
rect 37642 10752 37648 10804
rect 37700 10752 37706 10804
rect 37182 10724 37188 10736
rect 35400 10696 35445 10724
rect 35544 10696 37188 10724
rect 35400 10687 35412 10696
rect 35400 10684 35406 10687
rect 37182 10684 37188 10696
rect 37240 10684 37246 10736
rect 35526 10616 35532 10668
rect 35584 10656 35590 10668
rect 35621 10659 35679 10665
rect 35621 10656 35633 10659
rect 35584 10628 35633 10656
rect 35584 10616 35590 10628
rect 35621 10625 35633 10628
rect 35667 10625 35679 10659
rect 35621 10619 35679 10625
rect 38105 10659 38163 10665
rect 38105 10625 38117 10659
rect 38151 10625 38163 10659
rect 38105 10619 38163 10625
rect 33505 10551 33563 10557
rect 33612 10560 34652 10588
rect 31036 10492 32444 10520
rect 32861 10523 32919 10529
rect 31036 10464 31064 10492
rect 32861 10489 32873 10523
rect 32907 10489 32919 10523
rect 32861 10483 32919 10489
rect 33042 10480 33048 10532
rect 33100 10520 33106 10532
rect 33612 10520 33640 10560
rect 36170 10548 36176 10600
rect 36228 10548 36234 10600
rect 36262 10548 36268 10600
rect 36320 10548 36326 10600
rect 37274 10548 37280 10600
rect 37332 10588 37338 10600
rect 37369 10591 37427 10597
rect 37369 10588 37381 10591
rect 37332 10560 37381 10588
rect 37332 10548 37338 10560
rect 37369 10557 37381 10560
rect 37415 10588 37427 10591
rect 37642 10588 37648 10600
rect 37415 10560 37648 10588
rect 37415 10557 37427 10560
rect 37369 10551 37427 10557
rect 37642 10548 37648 10560
rect 37700 10548 37706 10600
rect 38120 10520 38148 10619
rect 38470 10520 38476 10532
rect 33100 10492 33640 10520
rect 33980 10492 34192 10520
rect 33100 10480 33106 10492
rect 30423 10424 30604 10452
rect 30423 10421 30435 10424
rect 30377 10415 30435 10421
rect 31018 10412 31024 10464
rect 31076 10412 31082 10464
rect 31386 10412 31392 10464
rect 31444 10452 31450 10464
rect 33980 10452 34008 10492
rect 31444 10424 34008 10452
rect 34164 10452 34192 10492
rect 35636 10492 38148 10520
rect 38212 10492 38476 10520
rect 35636 10452 35664 10492
rect 34164 10424 35664 10452
rect 35713 10455 35771 10461
rect 31444 10412 31450 10424
rect 35713 10421 35725 10455
rect 35759 10452 35771 10455
rect 35894 10452 35900 10464
rect 35759 10424 35900 10452
rect 35759 10421 35771 10424
rect 35713 10415 35771 10421
rect 35894 10412 35900 10424
rect 35952 10412 35958 10464
rect 38013 10455 38071 10461
rect 38013 10421 38025 10455
rect 38059 10452 38071 10455
rect 38212 10452 38240 10492
rect 38470 10480 38476 10492
rect 38528 10480 38534 10532
rect 38059 10424 38240 10452
rect 38059 10421 38071 10424
rect 38013 10415 38071 10421
rect 38286 10412 38292 10464
rect 38344 10412 38350 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10217 2375 10251
rect 2317 10211 2375 10217
rect 2332 10044 2360 10211
rect 2590 10208 2596 10260
rect 2648 10208 2654 10260
rect 5258 10248 5264 10260
rect 4632 10220 5264 10248
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10180 2559 10183
rect 2547 10152 2774 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 2746 10112 2774 10152
rect 3602 10140 3608 10192
rect 3660 10140 3666 10192
rect 3145 10115 3203 10121
rect 3145 10112 3157 10115
rect 2746 10084 3157 10112
rect 3145 10081 3157 10084
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 3418 10044 3424 10056
rect 2332 10016 3424 10044
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 3620 10044 3648 10140
rect 4632 10121 4660 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5445 10251 5503 10257
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 10226 10248 10232 10260
rect 5491 10220 10232 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 13170 10248 13176 10260
rect 13004 10220 13176 10248
rect 4706 10140 4712 10192
rect 4764 10140 4770 10192
rect 5074 10140 5080 10192
rect 5132 10180 5138 10192
rect 5534 10180 5540 10192
rect 5132 10152 5540 10180
rect 5132 10140 5138 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 7469 10183 7527 10189
rect 7469 10149 7481 10183
rect 7515 10180 7527 10183
rect 7650 10180 7656 10192
rect 7515 10152 7656 10180
rect 7515 10149 7527 10152
rect 7469 10143 7527 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 7834 10140 7840 10192
rect 7892 10140 7898 10192
rect 9858 10140 9864 10192
rect 9916 10140 9922 10192
rect 12529 10183 12587 10189
rect 12529 10149 12541 10183
rect 12575 10180 12587 10183
rect 13004 10180 13032 10220
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 14182 10208 14188 10260
rect 14240 10208 14246 10260
rect 14918 10208 14924 10260
rect 14976 10208 14982 10260
rect 15838 10208 15844 10260
rect 15896 10208 15902 10260
rect 18046 10208 18052 10260
rect 18104 10208 18110 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 18196 10220 18245 10248
rect 18196 10208 18202 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18233 10211 18291 10217
rect 27062 10208 27068 10260
rect 27120 10208 27126 10260
rect 27157 10251 27215 10257
rect 27157 10217 27169 10251
rect 27203 10248 27215 10251
rect 27338 10248 27344 10260
rect 27203 10220 27344 10248
rect 27203 10217 27215 10220
rect 27157 10211 27215 10217
rect 27338 10208 27344 10220
rect 27396 10208 27402 10260
rect 30377 10251 30435 10257
rect 30377 10217 30389 10251
rect 30423 10248 30435 10251
rect 30926 10248 30932 10260
rect 30423 10220 30932 10248
rect 30423 10217 30435 10220
rect 30377 10211 30435 10217
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 31294 10208 31300 10260
rect 31352 10208 31358 10260
rect 31662 10208 31668 10260
rect 31720 10248 31726 10260
rect 34149 10251 34207 10257
rect 34149 10248 34161 10251
rect 31720 10220 34161 10248
rect 31720 10208 31726 10220
rect 34149 10217 34161 10220
rect 34195 10248 34207 10251
rect 36262 10248 36268 10260
rect 34195 10220 36268 10248
rect 34195 10217 34207 10220
rect 34149 10211 34207 10217
rect 36262 10208 36268 10220
rect 36320 10208 36326 10260
rect 37458 10208 37464 10260
rect 37516 10248 37522 10260
rect 37645 10251 37703 10257
rect 37645 10248 37657 10251
rect 37516 10220 37657 10248
rect 37516 10208 37522 10220
rect 37645 10217 37657 10220
rect 37691 10217 37703 10251
rect 37645 10211 37703 10217
rect 37918 10208 37924 10260
rect 37976 10248 37982 10260
rect 38381 10251 38439 10257
rect 38381 10248 38393 10251
rect 37976 10220 38393 10248
rect 37976 10208 37982 10220
rect 38381 10217 38393 10220
rect 38427 10217 38439 10251
rect 38381 10211 38439 10217
rect 12575 10152 13032 10180
rect 12575 10149 12587 10152
rect 12529 10143 12587 10149
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10081 4675 10115
rect 4617 10075 4675 10081
rect 4724 10053 4752 10140
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 4856 10084 5181 10112
rect 4856 10072 4862 10084
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 7668 10112 7696 10140
rect 8662 10112 8668 10124
rect 7668 10084 8668 10112
rect 5169 10075 5227 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 9876 10112 9904 10140
rect 12894 10112 12900 10124
rect 9876 10084 12900 10112
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 14200 10112 14228 10208
rect 14936 10121 14964 10208
rect 13832 10084 14228 10112
rect 14921 10115 14979 10121
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 3620 10016 4261 10044
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 8018 10004 8024 10056
rect 8076 10004 8082 10056
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8904 10016 8953 10044
rect 8904 10004 8910 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 13832 10044 13860 10084
rect 14921 10081 14933 10115
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 16666 10072 16672 10124
rect 16724 10072 16730 10124
rect 18064 10112 18092 10208
rect 27080 10180 27108 10208
rect 27522 10180 27528 10192
rect 27080 10152 27528 10180
rect 27522 10140 27528 10152
rect 27580 10140 27586 10192
rect 28169 10183 28227 10189
rect 28169 10149 28181 10183
rect 28215 10180 28227 10183
rect 28350 10180 28356 10192
rect 28215 10152 28356 10180
rect 28215 10149 28227 10152
rect 28169 10143 28227 10149
rect 28350 10140 28356 10152
rect 28408 10180 28414 10192
rect 29178 10180 29184 10192
rect 28408 10152 29184 10180
rect 28408 10140 28414 10152
rect 29178 10140 29184 10152
rect 29236 10180 29242 10192
rect 30009 10183 30067 10189
rect 30009 10180 30021 10183
rect 29236 10152 30021 10180
rect 29236 10140 29242 10152
rect 30009 10149 30021 10152
rect 30055 10180 30067 10183
rect 31846 10180 31852 10192
rect 30055 10152 31852 10180
rect 30055 10149 30067 10152
rect 30009 10143 30067 10149
rect 31846 10140 31852 10152
rect 31904 10180 31910 10192
rect 32122 10180 32128 10192
rect 31904 10152 32128 10180
rect 31904 10140 31910 10152
rect 32122 10140 32128 10152
rect 32180 10140 32186 10192
rect 32401 10183 32459 10189
rect 32401 10149 32413 10183
rect 32447 10180 32459 10183
rect 34330 10180 34336 10192
rect 32447 10152 34336 10180
rect 32447 10149 32459 10152
rect 32401 10143 32459 10149
rect 18785 10115 18843 10121
rect 18785 10112 18797 10115
rect 18064 10084 18797 10112
rect 18785 10081 18797 10084
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 27706 10072 27712 10124
rect 27764 10072 27770 10124
rect 29822 10072 29828 10124
rect 29880 10112 29886 10124
rect 32416 10112 32444 10143
rect 34330 10140 34336 10152
rect 34388 10140 34394 10192
rect 29880 10084 32444 10112
rect 29880 10072 29886 10084
rect 33042 10072 33048 10124
rect 33100 10072 33106 10124
rect 33778 10072 33784 10124
rect 33836 10072 33842 10124
rect 37366 10072 37372 10124
rect 37424 10112 37430 10124
rect 37737 10115 37795 10121
rect 37737 10112 37749 10115
rect 37424 10084 37749 10112
rect 37424 10072 37430 10084
rect 37737 10081 37749 10084
rect 37783 10081 37795 10115
rect 37737 10075 37795 10081
rect 12483 10016 13860 10044
rect 13909 10047 13967 10053
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 13909 10013 13921 10047
rect 13955 10044 13967 10047
rect 14274 10044 14280 10056
rect 13955 10016 14280 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 14274 10004 14280 10016
rect 14332 10044 14338 10056
rect 15102 10044 15108 10056
rect 14332 10016 15108 10044
rect 14332 10004 14338 10016
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 30926 10004 30932 10056
rect 30984 10044 30990 10056
rect 31570 10044 31576 10056
rect 30984 10016 31576 10044
rect 30984 10004 30990 10016
rect 31570 10004 31576 10016
rect 31628 10044 31634 10056
rect 32033 10047 32091 10053
rect 31628 10016 31984 10044
rect 31628 10004 31634 10016
rect 1762 9936 1768 9988
rect 1820 9976 1826 9988
rect 2133 9979 2191 9985
rect 2133 9976 2145 9979
rect 1820 9948 2145 9976
rect 1820 9936 1826 9948
rect 2133 9945 2145 9948
rect 2179 9976 2191 9979
rect 3694 9976 3700 9988
rect 2179 9948 3700 9976
rect 2179 9945 2191 9948
rect 2133 9939 2191 9945
rect 3694 9936 3700 9948
rect 3752 9936 3758 9988
rect 12802 9976 12808 9988
rect 12406 9948 12808 9976
rect 2343 9911 2401 9917
rect 2343 9877 2355 9911
rect 2389 9908 2401 9911
rect 3050 9908 3056 9920
rect 2389 9880 3056 9908
rect 2389 9877 2401 9880
rect 2343 9871 2401 9877
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 4433 9911 4491 9917
rect 4433 9877 4445 9911
rect 4479 9908 4491 9911
rect 4706 9908 4712 9920
rect 4479 9880 4712 9908
rect 4479 9877 4491 9880
rect 4433 9871 4491 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8536 9880 8585 9908
rect 8536 9868 8542 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 8573 9871 8631 9877
rect 9582 9868 9588 9920
rect 9640 9868 9646 9920
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 12406 9908 12434 9948
rect 12802 9936 12808 9948
rect 12860 9936 12866 9988
rect 13664 9979 13722 9985
rect 13664 9945 13676 9979
rect 13710 9976 13722 9979
rect 14369 9979 14427 9985
rect 14369 9976 14381 9979
rect 13710 9948 14381 9976
rect 13710 9945 13722 9948
rect 13664 9939 13722 9945
rect 14369 9945 14381 9948
rect 14415 9945 14427 9979
rect 14369 9939 14427 9945
rect 16936 9979 16994 9985
rect 16936 9945 16948 9979
rect 16982 9976 16994 9979
rect 17678 9976 17684 9988
rect 16982 9948 17684 9976
rect 16982 9945 16994 9948
rect 16936 9939 16994 9945
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 31956 9976 31984 10016
rect 32033 10013 32045 10047
rect 32079 10044 32091 10047
rect 32214 10044 32220 10056
rect 32079 10016 32220 10044
rect 32079 10013 32091 10016
rect 32033 10007 32091 10013
rect 32214 10004 32220 10016
rect 32272 10044 32278 10056
rect 33060 10044 33088 10072
rect 32272 10016 33088 10044
rect 32272 10004 32278 10016
rect 34514 10004 34520 10056
rect 34572 10044 34578 10056
rect 34701 10047 34759 10053
rect 34701 10044 34713 10047
rect 34572 10016 34713 10044
rect 34572 10004 34578 10016
rect 34701 10013 34713 10016
rect 34747 10044 34759 10047
rect 36265 10047 36323 10053
rect 36265 10044 36277 10047
rect 34747 10016 36277 10044
rect 34747 10013 34759 10016
rect 34701 10007 34759 10013
rect 36265 10013 36277 10016
rect 36311 10013 36323 10047
rect 36814 10044 36820 10056
rect 36265 10007 36323 10013
rect 36464 10016 36820 10044
rect 34425 9979 34483 9985
rect 34425 9976 34437 9979
rect 31726 9948 31892 9976
rect 31956 9948 34437 9976
rect 12124 9880 12434 9908
rect 15381 9911 15439 9917
rect 12124 9868 12130 9880
rect 15381 9877 15393 9911
rect 15427 9908 15439 9911
rect 15562 9908 15568 9920
rect 15427 9880 15568 9908
rect 15427 9877 15439 9880
rect 15381 9871 15439 9877
rect 15562 9868 15568 9880
rect 15620 9908 15626 9920
rect 16850 9908 16856 9920
rect 15620 9880 16856 9908
rect 15620 9868 15626 9880
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 23014 9868 23020 9920
rect 23072 9868 23078 9920
rect 26697 9911 26755 9917
rect 26697 9877 26709 9911
rect 26743 9908 26755 9911
rect 26786 9908 26792 9920
rect 26743 9880 26792 9908
rect 26743 9877 26755 9880
rect 26697 9871 26755 9877
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 30742 9868 30748 9920
rect 30800 9908 30806 9920
rect 31726 9908 31754 9948
rect 30800 9880 31754 9908
rect 31864 9908 31892 9948
rect 34425 9945 34437 9948
rect 34471 9945 34483 9979
rect 34425 9939 34483 9945
rect 34968 9979 35026 9985
rect 34968 9945 34980 9979
rect 35014 9976 35026 9979
rect 35342 9976 35348 9988
rect 35014 9948 35348 9976
rect 35014 9945 35026 9948
rect 34968 9939 35026 9945
rect 32030 9908 32036 9920
rect 31864 9880 32036 9908
rect 30800 9868 30806 9880
rect 32030 9868 32036 9880
rect 32088 9868 32094 9920
rect 32122 9868 32128 9920
rect 32180 9908 32186 9920
rect 32677 9911 32735 9917
rect 32677 9908 32689 9911
rect 32180 9880 32689 9908
rect 32180 9868 32186 9880
rect 32677 9877 32689 9880
rect 32723 9877 32735 9911
rect 34440 9908 34468 9939
rect 35342 9936 35348 9948
rect 35400 9936 35406 9988
rect 36464 9976 36492 10016
rect 36814 10004 36820 10016
rect 36872 10004 36878 10056
rect 36004 9948 36492 9976
rect 36532 9979 36590 9985
rect 36004 9908 36032 9948
rect 36532 9945 36544 9979
rect 36578 9976 36590 9979
rect 37274 9976 37280 9988
rect 36578 9948 37280 9976
rect 36578 9945 36590 9948
rect 36532 9939 36590 9945
rect 37274 9936 37280 9948
rect 37332 9936 37338 9988
rect 34440 9880 36032 9908
rect 36081 9911 36139 9917
rect 32677 9871 32735 9877
rect 36081 9877 36093 9911
rect 36127 9908 36139 9911
rect 36446 9908 36452 9920
rect 36127 9880 36452 9908
rect 36127 9877 36139 9880
rect 36081 9871 36139 9877
rect 36446 9868 36452 9880
rect 36504 9908 36510 9920
rect 36814 9908 36820 9920
rect 36504 9880 36820 9908
rect 36504 9868 36510 9880
rect 36814 9868 36820 9880
rect 36872 9868 36878 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 2777 9707 2835 9713
rect 2777 9704 2789 9707
rect 2464 9676 2789 9704
rect 2464 9664 2470 9676
rect 2777 9673 2789 9676
rect 2823 9704 2835 9707
rect 2823 9676 2877 9704
rect 2823 9673 2835 9676
rect 2777 9667 2835 9673
rect 2792 9636 2820 9667
rect 3050 9664 3056 9716
rect 3108 9664 3114 9716
rect 3602 9664 3608 9716
rect 3660 9664 3666 9716
rect 4433 9707 4491 9713
rect 4433 9673 4445 9707
rect 4479 9704 4491 9707
rect 5166 9704 5172 9716
rect 4479 9676 5172 9704
rect 4479 9673 4491 9676
rect 4433 9667 4491 9673
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 8113 9707 8171 9713
rect 8113 9704 8125 9707
rect 8076 9676 8125 9704
rect 8076 9664 8082 9676
rect 8113 9673 8125 9676
rect 8159 9673 8171 9707
rect 8113 9667 8171 9673
rect 16022 9664 16028 9716
rect 16080 9664 16086 9716
rect 17678 9664 17684 9716
rect 17736 9664 17742 9716
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 25038 9704 25044 9716
rect 21232 9676 25044 9704
rect 21232 9664 21238 9676
rect 25038 9664 25044 9676
rect 25096 9664 25102 9716
rect 27617 9707 27675 9713
rect 27617 9673 27629 9707
rect 27663 9704 27675 9707
rect 28350 9704 28356 9716
rect 27663 9676 28356 9704
rect 27663 9673 27675 9676
rect 27617 9667 27675 9673
rect 28350 9664 28356 9676
rect 28408 9664 28414 9716
rect 31496 9676 31708 9704
rect 2792 9608 3464 9636
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2556 9540 2605 9568
rect 2556 9528 2562 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 2682 9500 2688 9512
rect 2280 9472 2688 9500
rect 2280 9460 2286 9472
rect 2682 9460 2688 9472
rect 2740 9500 2746 9512
rect 2976 9500 3004 9531
rect 3436 9512 3464 9608
rect 3620 9568 3648 9664
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 5442 9636 5448 9648
rect 4847 9608 5448 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 7800 9608 8493 9636
rect 7800 9596 7806 9608
rect 8481 9605 8493 9608
rect 8527 9636 8539 9639
rect 8527 9608 9076 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 9048 9580 9076 9608
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12805 9639 12863 9645
rect 12805 9636 12817 9639
rect 12584 9608 12817 9636
rect 12584 9596 12590 9608
rect 12805 9605 12817 9608
rect 12851 9605 12863 9639
rect 12805 9599 12863 9605
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 3620 9540 3801 9568
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 4274 9571 4332 9577
rect 4274 9568 4286 9571
rect 3789 9531 3847 9537
rect 3988 9540 4286 9568
rect 2740 9472 3004 9500
rect 2740 9460 2746 9472
rect 2869 9435 2927 9441
rect 2869 9401 2881 9435
rect 2915 9401 2927 9435
rect 2976 9432 3004 9472
rect 3418 9460 3424 9512
rect 3476 9460 3482 9512
rect 3602 9460 3608 9512
rect 3660 9460 3666 9512
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 3988 9500 4016 9540
rect 4274 9537 4286 9540
rect 4320 9537 4332 9571
rect 4274 9531 4332 9537
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8619 9540 8953 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9030 9528 9036 9580
rect 9088 9528 9094 9580
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 16040 9568 16068 9664
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 16816 9608 17141 9636
rect 16816 9596 16822 9608
rect 17129 9605 17141 9608
rect 17175 9605 17187 9639
rect 17129 9599 17187 9605
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 25409 9639 25467 9645
rect 25409 9636 25421 9639
rect 24728 9608 25421 9636
rect 24728 9596 24734 9608
rect 25409 9605 25421 9608
rect 25455 9636 25467 9639
rect 26786 9636 26792 9648
rect 25455 9608 26792 9636
rect 25455 9605 25467 9608
rect 25409 9599 25467 9605
rect 26786 9596 26792 9608
rect 26844 9596 26850 9648
rect 31496 9636 31524 9676
rect 31680 9674 31708 9676
rect 34256 9676 34560 9704
rect 31680 9646 31800 9674
rect 29104 9608 31524 9636
rect 31772 9636 31800 9646
rect 32214 9636 32220 9648
rect 31772 9608 32220 9636
rect 29104 9580 29132 9608
rect 32214 9596 32220 9608
rect 32272 9596 32278 9648
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 16040 9540 17233 9568
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 18598 9568 18604 9580
rect 18371 9540 18604 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 21637 9571 21695 9577
rect 21637 9568 21649 9571
rect 20772 9540 21649 9568
rect 20772 9528 20778 9540
rect 21637 9537 21649 9540
rect 21683 9568 21695 9571
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 21683 9540 22109 9568
rect 21683 9537 21695 9540
rect 21637 9531 21695 9537
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 29086 9528 29092 9580
rect 29144 9528 29150 9580
rect 30466 9528 30472 9580
rect 30524 9568 30530 9580
rect 31478 9568 31484 9580
rect 30524 9540 31484 9568
rect 30524 9528 30530 9540
rect 31478 9528 31484 9540
rect 31536 9528 31542 9580
rect 32674 9528 32680 9580
rect 32732 9568 32738 9580
rect 33042 9568 33048 9580
rect 32732 9540 33048 9568
rect 32732 9528 32738 9540
rect 33042 9528 33048 9540
rect 33100 9568 33106 9580
rect 34256 9568 34284 9676
rect 34330 9596 34336 9648
rect 34388 9636 34394 9648
rect 34425 9639 34483 9645
rect 34425 9636 34437 9639
rect 34388 9608 34437 9636
rect 34388 9596 34394 9608
rect 34425 9605 34437 9608
rect 34471 9605 34483 9639
rect 34532 9636 34560 9676
rect 36170 9664 36176 9716
rect 36228 9704 36234 9716
rect 36265 9707 36323 9713
rect 36265 9704 36277 9707
rect 36228 9676 36277 9704
rect 36228 9664 36234 9676
rect 36265 9673 36277 9676
rect 36311 9673 36323 9707
rect 36265 9667 36323 9673
rect 37274 9664 37280 9716
rect 37332 9664 37338 9716
rect 36078 9636 36084 9648
rect 34532 9608 36084 9636
rect 34425 9599 34483 9605
rect 36078 9596 36084 9608
rect 36136 9636 36142 9648
rect 38746 9636 38752 9648
rect 36136 9608 38752 9636
rect 36136 9596 36142 9608
rect 38746 9596 38752 9608
rect 38804 9596 38810 9648
rect 38473 9571 38531 9577
rect 38473 9568 38485 9571
rect 33100 9540 34284 9568
rect 34348 9540 38485 9568
rect 33100 9528 33106 9540
rect 3752 9472 4016 9500
rect 3752 9460 3758 9472
rect 4062 9460 4068 9512
rect 4120 9460 4126 9512
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 3970 9432 3976 9444
rect 2976 9404 3976 9432
rect 2869 9395 2927 9401
rect 2884 9364 2912 9395
rect 3970 9392 3976 9404
rect 4028 9432 4034 9444
rect 4172 9432 4200 9463
rect 4028 9404 4200 9432
rect 6656 9432 6684 9463
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8386 9500 8392 9512
rect 7892 9472 8392 9500
rect 7892 9460 7898 9472
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8662 9460 8668 9512
rect 8720 9460 8726 9512
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 8772 9472 9505 9500
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 6656 9404 7297 9432
rect 4028 9392 4034 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7285 9395 7343 9401
rect 3234 9364 3240 9376
rect 2884 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 7193 9367 7251 9373
rect 7193 9333 7205 9367
rect 7239 9364 7251 9367
rect 7466 9364 7472 9376
rect 7239 9336 7472 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8772 9364 8800 9472
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 10410 9460 10416 9512
rect 10468 9500 10474 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 10468 9472 16405 9500
rect 10468 9460 10474 9472
rect 16393 9469 16405 9472
rect 16439 9500 16451 9503
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16439 9472 16957 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 18966 9460 18972 9512
rect 19024 9460 19030 9512
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23014 9500 23020 9512
rect 22971 9472 23020 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23014 9460 23020 9472
rect 23072 9460 23078 9512
rect 23750 9460 23756 9512
rect 23808 9460 23814 9512
rect 26145 9503 26203 9509
rect 26145 9469 26157 9503
rect 26191 9500 26203 9503
rect 26326 9500 26332 9512
rect 26191 9472 26332 9500
rect 26191 9469 26203 9472
rect 26145 9463 26203 9469
rect 26326 9460 26332 9472
rect 26384 9460 26390 9512
rect 29914 9460 29920 9512
rect 29972 9460 29978 9512
rect 30558 9460 30564 9512
rect 30616 9460 30622 9512
rect 31202 9460 31208 9512
rect 31260 9460 31266 9512
rect 31294 9460 31300 9512
rect 31352 9500 31358 9512
rect 34348 9509 34376 9540
rect 38473 9537 38485 9540
rect 38519 9537 38531 9571
rect 38473 9531 38531 9537
rect 32309 9503 32367 9509
rect 32309 9500 32321 9503
rect 31352 9472 32321 9500
rect 31352 9460 31358 9472
rect 32309 9469 32321 9472
rect 32355 9469 32367 9503
rect 32309 9463 32367 9469
rect 33781 9503 33839 9509
rect 33781 9469 33793 9503
rect 33827 9469 33839 9503
rect 33781 9463 33839 9469
rect 34333 9503 34391 9509
rect 34333 9469 34345 9503
rect 34379 9469 34391 9503
rect 34333 9463 34391 9469
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 16666 9432 16672 9444
rect 15160 9404 16672 9432
rect 15160 9392 15166 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 17589 9435 17647 9441
rect 17589 9401 17601 9435
rect 17635 9432 17647 9435
rect 18506 9432 18512 9444
rect 17635 9404 18512 9432
rect 17635 9401 17647 9404
rect 17589 9395 17647 9401
rect 18506 9392 18512 9404
rect 18564 9392 18570 9444
rect 29089 9435 29147 9441
rect 29089 9401 29101 9435
rect 29135 9432 29147 9435
rect 29825 9435 29883 9441
rect 29825 9432 29837 9435
rect 29135 9404 29837 9432
rect 29135 9401 29147 9404
rect 29089 9395 29147 9401
rect 29825 9401 29837 9404
rect 29871 9432 29883 9435
rect 30576 9432 30604 9460
rect 31662 9432 31668 9444
rect 29871 9404 31668 9432
rect 29871 9401 29883 9404
rect 29825 9395 29883 9401
rect 31036 9376 31064 9404
rect 31662 9392 31668 9404
rect 31720 9392 31726 9444
rect 33796 9432 33824 9463
rect 36814 9460 36820 9512
rect 36872 9460 36878 9512
rect 37826 9460 37832 9512
rect 37884 9460 37890 9512
rect 38010 9460 38016 9512
rect 38068 9500 38074 9512
rect 38068 9472 38332 9500
rect 38068 9460 38074 9472
rect 38304 9441 38332 9472
rect 38289 9435 38347 9441
rect 33796 9404 38240 9432
rect 8168 9336 8800 9364
rect 8168 9324 8174 9336
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 8996 9336 9873 9364
rect 8996 9324 9002 9336
rect 9861 9333 9873 9336
rect 9907 9364 9919 9367
rect 11238 9364 11244 9376
rect 9907 9336 11244 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12158 9364 12164 9376
rect 12023 9336 12164 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 18414 9324 18420 9376
rect 18472 9324 18478 9376
rect 23198 9324 23204 9376
rect 23256 9324 23262 9376
rect 25498 9324 25504 9376
rect 25556 9324 25562 9376
rect 27154 9324 27160 9376
rect 27212 9324 27218 9376
rect 28994 9324 29000 9376
rect 29052 9364 29058 9376
rect 29365 9367 29423 9373
rect 29365 9364 29377 9367
rect 29052 9336 29377 9364
rect 29052 9324 29058 9336
rect 29365 9333 29377 9336
rect 29411 9333 29423 9367
rect 29365 9327 29423 9333
rect 30558 9324 30564 9376
rect 30616 9324 30622 9376
rect 30650 9324 30656 9376
rect 30708 9324 30714 9376
rect 31018 9324 31024 9376
rect 31076 9324 31082 9376
rect 31478 9324 31484 9376
rect 31536 9364 31542 9376
rect 31573 9367 31631 9373
rect 31573 9364 31585 9367
rect 31536 9336 31585 9364
rect 31536 9324 31542 9336
rect 31573 9333 31585 9336
rect 31619 9333 31631 9367
rect 31573 9327 31631 9333
rect 32950 9324 32956 9376
rect 33008 9324 33014 9376
rect 33318 9324 33324 9376
rect 33376 9324 33382 9376
rect 34514 9324 34520 9376
rect 34572 9364 34578 9376
rect 35713 9367 35771 9373
rect 35713 9364 35725 9367
rect 34572 9336 35725 9364
rect 34572 9324 34578 9336
rect 35713 9333 35725 9336
rect 35759 9333 35771 9367
rect 38212 9364 38240 9404
rect 38289 9401 38301 9435
rect 38335 9401 38347 9435
rect 38289 9395 38347 9401
rect 38930 9364 38936 9376
rect 38212 9336 38936 9364
rect 35713 9327 35771 9333
rect 38930 9324 38936 9336
rect 38988 9324 38994 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 658 9120 664 9172
rect 716 9160 722 9172
rect 19426 9160 19432 9172
rect 716 9132 19432 9160
rect 716 9120 722 9132
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 22738 9120 22744 9172
rect 22796 9160 22802 9172
rect 23290 9160 23296 9172
rect 22796 9132 23296 9160
rect 22796 9120 22802 9132
rect 23290 9120 23296 9132
rect 23348 9160 23354 9172
rect 24670 9160 24676 9172
rect 23348 9132 24676 9160
rect 23348 9120 23354 9132
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 30834 9120 30840 9172
rect 30892 9160 30898 9172
rect 31205 9163 31263 9169
rect 31205 9160 31217 9163
rect 30892 9132 31217 9160
rect 30892 9120 30898 9132
rect 31205 9129 31217 9132
rect 31251 9160 31263 9163
rect 31294 9160 31300 9172
rect 31251 9132 31300 9160
rect 31251 9129 31263 9132
rect 31205 9123 31263 9129
rect 31294 9120 31300 9132
rect 31352 9120 31358 9172
rect 34330 9120 34336 9172
rect 34388 9120 34394 9172
rect 35342 9120 35348 9172
rect 35400 9120 35406 9172
rect 37734 9120 37740 9172
rect 37792 9120 37798 9172
rect 3602 9052 3608 9104
rect 3660 9052 3666 9104
rect 4706 9092 4712 9104
rect 4448 9064 4712 9092
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 2740 8996 3188 9024
rect 2740 8984 2746 8996
rect 3160 8965 3188 8996
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4448 8965 4476 9064
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 7285 9095 7343 9101
rect 7285 9061 7297 9095
rect 7331 9092 7343 9095
rect 7650 9092 7656 9104
rect 7331 9064 7656 9092
rect 7331 9061 7343 9064
rect 7285 9055 7343 9061
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 9677 9095 9735 9101
rect 9677 9061 9689 9095
rect 9723 9061 9735 9095
rect 9677 9055 9735 9061
rect 12069 9095 12127 9101
rect 12069 9061 12081 9095
rect 12115 9061 12127 9095
rect 12069 9055 12127 9061
rect 26421 9095 26479 9101
rect 26421 9061 26433 9095
rect 26467 9092 26479 9095
rect 26602 9092 26608 9104
rect 26467 9064 26608 9092
rect 26467 9061 26479 9064
rect 26421 9055 26479 9061
rect 8938 8984 8944 9036
rect 8996 9024 9002 9036
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8996 8996 9045 9024
rect 8996 8984 9002 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9692 9024 9720 9055
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9692 8996 10333 9024
rect 9033 8987 9091 8993
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 12084 9024 12112 9055
rect 26602 9052 26608 9064
rect 26660 9052 26666 9104
rect 12023 8996 12112 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12713 9027 12771 9033
rect 12713 9024 12725 9027
rect 12216 8996 12725 9024
rect 12216 8984 12222 8996
rect 12713 8993 12725 8996
rect 12759 9024 12771 9027
rect 16206 9024 16212 9036
rect 12759 8996 16212 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 16666 8984 16672 9036
rect 16724 8984 16730 9036
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 34514 9024 34520 9036
rect 16807 8996 16988 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4264 8928 4445 8956
rect 3436 8888 3464 8916
rect 4264 8888 4292 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 4798 8956 4804 8968
rect 4580 8928 4804 8956
rect 4580 8916 4586 8928
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 6779 8928 8432 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 3436 8860 4292 8888
rect 4341 8891 4399 8897
rect 4341 8857 4353 8891
rect 4387 8888 4399 8891
rect 5074 8888 5080 8900
rect 4387 8860 5080 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 8110 8888 8116 8900
rect 7392 8860 8116 8888
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 3234 8820 3240 8832
rect 2924 8792 3240 8820
rect 2924 8780 2930 8792
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 7392 8829 7420 8860
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 4617 8823 4675 8829
rect 4617 8820 4629 8823
rect 3752 8792 4629 8820
rect 3752 8780 3758 8792
rect 4617 8789 4629 8792
rect 4663 8789 4675 8823
rect 4617 8783 4675 8789
rect 7377 8823 7435 8829
rect 7377 8789 7389 8823
rect 7423 8789 7435 8823
rect 8404 8820 8432 8928
rect 8478 8916 8484 8968
rect 8536 8965 8542 8968
rect 8536 8956 8548 8965
rect 8536 8928 8581 8956
rect 8536 8919 8548 8928
rect 8536 8916 8542 8919
rect 8754 8916 8760 8968
rect 8812 8916 8818 8968
rect 13446 8916 13452 8968
rect 13504 8916 13510 8968
rect 15930 8916 15936 8968
rect 15988 8916 15994 8968
rect 16684 8956 16712 8984
rect 16960 8968 16988 8996
rect 32600 8996 34520 9024
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16684 8928 16865 8956
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 16942 8916 16948 8968
rect 17000 8916 17006 8968
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 17552 8928 18613 8956
rect 17552 8916 17558 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 21082 8916 21088 8968
rect 21140 8916 21146 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 22204 8928 22569 8956
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 10502 8888 10508 8900
rect 8720 8860 10508 8888
rect 8720 8848 8726 8860
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 17120 8891 17178 8897
rect 17120 8857 17132 8891
rect 17166 8888 17178 8891
rect 18046 8888 18052 8900
rect 17166 8860 18052 8888
rect 17166 8857 17178 8860
rect 17120 8851 17178 8857
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 18417 8891 18475 8897
rect 18417 8857 18429 8891
rect 18463 8888 18475 8891
rect 18782 8888 18788 8900
rect 18463 8860 18788 8888
rect 18463 8857 18475 8860
rect 18417 8851 18475 8857
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 22204 8832 22232 8928
rect 22557 8925 22569 8928
rect 22603 8956 22615 8959
rect 24029 8959 24087 8965
rect 24029 8956 24041 8959
rect 22603 8928 24041 8956
rect 22603 8925 22615 8928
rect 22557 8919 22615 8925
rect 24029 8925 24041 8928
rect 24075 8956 24087 8959
rect 24670 8956 24676 8968
rect 24075 8928 24676 8956
rect 24075 8925 24087 8928
rect 24029 8919 24087 8925
rect 24670 8916 24676 8928
rect 24728 8956 24734 8968
rect 25041 8959 25099 8965
rect 25041 8956 25053 8959
rect 24728 8928 25053 8956
rect 24728 8916 24734 8928
rect 25041 8925 25053 8928
rect 25087 8925 25099 8959
rect 25041 8919 25099 8925
rect 27062 8916 27068 8968
rect 27120 8916 27126 8968
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 27801 8959 27859 8965
rect 27801 8956 27813 8959
rect 27672 8928 27813 8956
rect 27672 8916 27678 8928
rect 27801 8925 27813 8928
rect 27847 8925 27859 8959
rect 27801 8919 27859 8925
rect 29730 8916 29736 8968
rect 29788 8916 29794 8968
rect 30000 8959 30058 8965
rect 30000 8925 30012 8959
rect 30046 8956 30058 8959
rect 30558 8956 30564 8968
rect 30046 8928 30564 8956
rect 30046 8925 30058 8928
rect 30000 8919 30058 8925
rect 30558 8916 30564 8928
rect 30616 8916 30622 8968
rect 31938 8916 31944 8968
rect 31996 8956 32002 8968
rect 32600 8965 32628 8996
rect 34514 8984 34520 8996
rect 34572 8984 34578 9036
rect 35894 8984 35900 9036
rect 35952 8984 35958 9036
rect 37458 8984 37464 9036
rect 37516 9024 37522 9036
rect 38289 9027 38347 9033
rect 38289 9024 38301 9027
rect 37516 8996 38301 9024
rect 37516 8984 37522 8996
rect 38289 8993 38301 8996
rect 38335 8993 38347 9027
rect 38289 8987 38347 8993
rect 32585 8959 32643 8965
rect 32585 8956 32597 8959
rect 31996 8928 32597 8956
rect 31996 8916 32002 8928
rect 32585 8925 32597 8928
rect 32631 8925 32643 8959
rect 32585 8919 32643 8925
rect 32766 8916 32772 8968
rect 32824 8956 32830 8968
rect 33229 8959 33287 8965
rect 33229 8956 33241 8959
rect 32824 8928 33241 8956
rect 32824 8916 32830 8928
rect 33229 8925 33241 8928
rect 33275 8925 33287 8959
rect 33229 8919 33287 8925
rect 33962 8916 33968 8968
rect 34020 8916 34026 8968
rect 36630 8916 36636 8968
rect 36688 8916 36694 8968
rect 37366 8916 37372 8968
rect 37424 8916 37430 8968
rect 22312 8891 22370 8897
rect 22312 8857 22324 8891
rect 22358 8888 22370 8891
rect 23198 8888 23204 8900
rect 22358 8860 23204 8888
rect 22358 8857 22370 8860
rect 22312 8851 22370 8857
rect 23198 8848 23204 8860
rect 23256 8848 23262 8900
rect 23784 8891 23842 8897
rect 23784 8857 23796 8891
rect 23830 8888 23842 8891
rect 24394 8888 24400 8900
rect 23830 8860 24400 8888
rect 23830 8857 23842 8860
rect 23784 8851 23842 8857
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 25308 8891 25366 8897
rect 25308 8857 25320 8891
rect 25354 8888 25366 8891
rect 25498 8888 25504 8900
rect 25354 8860 25504 8888
rect 25354 8857 25366 8860
rect 25308 8851 25366 8857
rect 25498 8848 25504 8860
rect 25556 8848 25562 8900
rect 28166 8848 28172 8900
rect 28224 8888 28230 8900
rect 28261 8891 28319 8897
rect 28261 8888 28273 8891
rect 28224 8860 28273 8888
rect 28224 8848 28230 8860
rect 28261 8857 28273 8860
rect 28307 8888 28319 8891
rect 28997 8891 29055 8897
rect 28307 8860 28672 8888
rect 28307 8857 28319 8860
rect 28261 8851 28319 8857
rect 8938 8820 8944 8832
rect 8404 8792 8944 8820
rect 7377 8783 7435 8789
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 9088 8792 9229 8820
rect 9088 8780 9094 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 9306 8780 9312 8832
rect 9364 8780 9370 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 9732 8792 9781 8820
rect 9732 8780 9738 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 11330 8780 11336 8832
rect 11388 8780 11394 8832
rect 12434 8780 12440 8832
rect 12492 8780 12498 8832
rect 12529 8823 12587 8829
rect 12529 8789 12541 8823
rect 12575 8820 12587 8823
rect 12897 8823 12955 8829
rect 12897 8820 12909 8823
rect 12575 8792 12909 8820
rect 12575 8789 12587 8792
rect 12529 8783 12587 8789
rect 12897 8789 12909 8792
rect 12943 8789 12955 8823
rect 12897 8783 12955 8789
rect 15378 8780 15384 8832
rect 15436 8780 15442 8832
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 18230 8780 18236 8832
rect 18288 8780 18294 8832
rect 20441 8823 20499 8829
rect 20441 8789 20453 8823
rect 20487 8820 20499 8823
rect 20898 8820 20904 8832
rect 20487 8792 20904 8820
rect 20487 8789 20499 8792
rect 20441 8783 20499 8789
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 21177 8823 21235 8829
rect 21177 8789 21189 8823
rect 21223 8820 21235 8823
rect 21726 8820 21732 8832
rect 21223 8792 21732 8820
rect 21223 8789 21235 8792
rect 21177 8783 21235 8789
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 22186 8780 22192 8832
rect 22244 8780 22250 8832
rect 22462 8780 22468 8832
rect 22520 8820 22526 8832
rect 22649 8823 22707 8829
rect 22649 8820 22661 8823
rect 22520 8792 22661 8820
rect 22520 8780 22526 8792
rect 22649 8789 22661 8792
rect 22695 8820 22707 8823
rect 22738 8820 22744 8832
rect 22695 8792 22744 8820
rect 22695 8789 22707 8792
rect 22649 8783 22707 8789
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 26510 8780 26516 8832
rect 26568 8780 26574 8832
rect 27246 8780 27252 8832
rect 27304 8780 27310 8832
rect 27522 8780 27528 8832
rect 27580 8820 27586 8832
rect 27982 8820 27988 8832
rect 27580 8792 27988 8820
rect 27580 8780 27586 8792
rect 27982 8780 27988 8792
rect 28040 8820 28046 8832
rect 28537 8823 28595 8829
rect 28537 8820 28549 8823
rect 28040 8792 28549 8820
rect 28040 8780 28046 8792
rect 28537 8789 28549 8792
rect 28583 8789 28595 8823
rect 28644 8820 28672 8860
rect 28997 8857 29009 8891
rect 29043 8888 29055 8891
rect 30742 8888 30748 8900
rect 29043 8860 30748 8888
rect 29043 8857 29055 8860
rect 28997 8851 29055 8857
rect 29564 8832 29592 8860
rect 30742 8848 30748 8860
rect 30800 8848 30806 8900
rect 32340 8891 32398 8897
rect 32340 8857 32352 8891
rect 32386 8888 32398 8891
rect 33413 8891 33471 8897
rect 33413 8888 33425 8891
rect 32386 8860 33425 8888
rect 32386 8857 32398 8860
rect 32340 8851 32398 8857
rect 33413 8857 33425 8860
rect 33459 8857 33471 8891
rect 33413 8851 33471 8857
rect 29086 8820 29092 8832
rect 28644 8792 29092 8820
rect 28537 8783 28595 8789
rect 29086 8780 29092 8792
rect 29144 8780 29150 8832
rect 29362 8780 29368 8832
rect 29420 8780 29426 8832
rect 29546 8780 29552 8832
rect 29604 8780 29610 8832
rect 31110 8780 31116 8832
rect 31168 8780 31174 8832
rect 32674 8780 32680 8832
rect 32732 8780 32738 8832
rect 34146 8780 34152 8832
rect 34204 8820 34210 8832
rect 34885 8823 34943 8829
rect 34885 8820 34897 8823
rect 34204 8792 34897 8820
rect 34204 8780 34210 8792
rect 34885 8789 34897 8792
rect 34931 8789 34943 8823
rect 34885 8783 34943 8789
rect 35894 8780 35900 8832
rect 35952 8820 35958 8832
rect 36081 8823 36139 8829
rect 36081 8820 36093 8823
rect 35952 8792 36093 8820
rect 35952 8780 35958 8792
rect 36081 8789 36093 8792
rect 36127 8789 36139 8823
rect 36081 8783 36139 8789
rect 36814 8780 36820 8832
rect 36872 8780 36878 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 4154 8616 4160 8628
rect 3292 8588 4160 8616
rect 3292 8576 3298 8588
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 10318 8576 10324 8628
rect 10376 8576 10382 8628
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 12989 8619 13047 8625
rect 12989 8616 13001 8619
rect 12952 8588 13001 8616
rect 12952 8576 12958 8588
rect 12989 8585 13001 8588
rect 13035 8616 13047 8619
rect 13446 8616 13452 8628
rect 13035 8588 13452 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 16853 8619 16911 8625
rect 16853 8616 16865 8619
rect 16632 8588 16865 8616
rect 16632 8576 16638 8588
rect 16853 8585 16865 8588
rect 16899 8616 16911 8619
rect 17678 8616 17684 8628
rect 16899 8588 17684 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 18414 8576 18420 8628
rect 18472 8576 18478 8628
rect 22186 8616 22192 8628
rect 20272 8588 22192 8616
rect 6472 8520 7236 8548
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 4522 8480 4528 8492
rect 2924 8452 4528 8480
rect 2924 8440 2930 8452
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 6472 8489 6500 8520
rect 7208 8492 7236 8520
rect 6730 8489 6736 8492
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 6724 8443 6736 8489
rect 6730 8440 6736 8443
rect 6788 8440 6794 8492
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8128 8480 8156 8576
rect 11348 8548 11376 8576
rect 11854 8551 11912 8557
rect 11854 8548 11866 8551
rect 11348 8520 11866 8548
rect 11854 8517 11866 8520
rect 11900 8517 11912 8551
rect 11854 8511 11912 8517
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 13541 8551 13599 8557
rect 13541 8548 13553 8551
rect 12492 8520 13553 8548
rect 12492 8508 12498 8520
rect 13541 8517 13553 8520
rect 13587 8548 13599 8551
rect 14366 8548 14372 8560
rect 13587 8520 14372 8548
rect 13587 8517 13599 8520
rect 13541 8511 13599 8517
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 17396 8551 17454 8557
rect 17396 8517 17408 8551
rect 17442 8548 17454 8551
rect 18432 8548 18460 8576
rect 17442 8520 18460 8548
rect 17442 8517 17454 8520
rect 17396 8511 17454 8517
rect 7975 8452 8156 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 8938 8440 8944 8492
rect 8996 8489 9002 8492
rect 8996 8483 9024 8489
rect 9012 8449 9024 8483
rect 8996 8443 9024 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 10229 8483 10287 8489
rect 10229 8480 10241 8483
rect 9815 8452 10241 8480
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 10229 8449 10241 8452
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 13449 8483 13507 8489
rect 11379 8452 13124 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 8996 8440 9002 8443
rect 8110 8372 8116 8424
rect 8168 8372 8174 8424
rect 8864 8412 8892 8440
rect 8496 8384 8892 8412
rect 9125 8415 9183 8421
rect 6178 8304 6184 8356
rect 6236 8344 6242 8356
rect 7837 8347 7895 8353
rect 6236 8316 6500 8344
rect 6236 8304 6242 8316
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 5994 8276 6000 8288
rect 3752 8248 6000 8276
rect 3752 8236 3758 8248
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 6472 8276 6500 8316
rect 7837 8313 7849 8347
rect 7883 8344 7895 8347
rect 8496 8344 8524 8384
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9490 8412 9496 8424
rect 9171 8384 9496 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 10410 8372 10416 8424
rect 10468 8372 10474 8424
rect 11606 8372 11612 8424
rect 11664 8372 11670 8424
rect 7883 8316 8524 8344
rect 8573 8347 8631 8353
rect 7883 8313 7895 8316
rect 7837 8307 7895 8313
rect 8573 8313 8585 8347
rect 8619 8344 8631 8347
rect 8662 8344 8668 8356
rect 8619 8316 8668 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 6822 8276 6828 8288
rect 6472 8248 6828 8276
rect 6822 8236 6828 8248
rect 6880 8276 6886 8288
rect 8588 8276 8616 8307
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 13096 8353 13124 8452
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13495 8452 13921 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 15378 8489 15384 8492
rect 15372 8480 15384 8489
rect 15339 8452 15384 8480
rect 15372 8443 15384 8452
rect 15378 8440 15384 8443
rect 15436 8440 15442 8492
rect 16666 8440 16672 8492
rect 16724 8480 16730 8492
rect 20272 8489 20300 8588
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 22370 8576 22376 8628
rect 22428 8616 22434 8628
rect 26053 8619 26111 8625
rect 22428 8588 24440 8616
rect 22428 8576 22434 8588
rect 21082 8508 21088 8560
rect 21140 8508 21146 8560
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 16724 8452 17141 8480
rect 16724 8440 16730 8452
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20513 8483 20571 8489
rect 20513 8480 20525 8483
rect 20257 8443 20315 8449
rect 20364 8452 20525 8480
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 18690 8412 18696 8424
rect 18524 8384 18696 8412
rect 18524 8353 18552 8384
rect 18690 8372 18696 8384
rect 18748 8412 18754 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18748 8384 19165 8412
rect 18748 8372 18754 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19153 8375 19211 8381
rect 19610 8372 19616 8424
rect 19668 8372 19674 8424
rect 20165 8415 20223 8421
rect 20165 8381 20177 8415
rect 20211 8412 20223 8415
rect 20364 8412 20392 8452
rect 20513 8449 20525 8452
rect 20559 8449 20571 8483
rect 21100 8480 21128 8508
rect 21100 8452 22232 8480
rect 20513 8443 20571 8449
rect 20211 8384 20392 8412
rect 20211 8381 20223 8384
rect 20165 8375 20223 8381
rect 21652 8353 21680 8452
rect 21726 8372 21732 8424
rect 21784 8412 21790 8424
rect 21821 8415 21879 8421
rect 21821 8412 21833 8415
rect 21784 8384 21833 8412
rect 21784 8372 21790 8384
rect 21821 8381 21833 8384
rect 21867 8381 21879 8415
rect 21821 8375 21879 8381
rect 21910 8372 21916 8424
rect 21968 8412 21974 8424
rect 22005 8415 22063 8421
rect 22005 8412 22017 8415
rect 21968 8384 22017 8412
rect 21968 8372 21974 8384
rect 22005 8381 22017 8384
rect 22051 8381 22063 8415
rect 22204 8412 22232 8452
rect 22738 8440 22744 8492
rect 22796 8440 22802 8492
rect 24412 8489 24440 8588
rect 26053 8585 26065 8619
rect 26099 8616 26111 8619
rect 26418 8616 26424 8628
rect 26099 8588 26424 8616
rect 26099 8585 26111 8588
rect 26053 8579 26111 8585
rect 26418 8576 26424 8588
rect 26476 8616 26482 8628
rect 27062 8616 27068 8628
rect 26476 8588 27068 8616
rect 26476 8576 26482 8588
rect 27062 8576 27068 8588
rect 27120 8576 27126 8628
rect 30650 8576 30656 8628
rect 30708 8576 30714 8628
rect 30837 8619 30895 8625
rect 30837 8585 30849 8619
rect 30883 8585 30895 8619
rect 30837 8579 30895 8585
rect 30929 8619 30987 8625
rect 30929 8585 30941 8619
rect 30975 8616 30987 8619
rect 31202 8616 31208 8628
rect 30975 8588 31208 8616
rect 30975 8585 30987 8588
rect 30929 8579 30987 8585
rect 29724 8551 29782 8557
rect 24596 8520 26832 8548
rect 22858 8483 22916 8489
rect 22858 8480 22870 8483
rect 22848 8449 22870 8480
rect 22904 8449 22916 8483
rect 22848 8443 22916 8449
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8449 24455 8483
rect 24397 8443 24455 8449
rect 22848 8412 22876 8443
rect 24596 8424 24624 8520
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 24940 8483 24998 8489
rect 24940 8449 24952 8483
rect 24986 8480 24998 8483
rect 26145 8483 26203 8489
rect 26145 8480 26157 8483
rect 24986 8452 26157 8480
rect 24986 8449 24998 8452
rect 24940 8443 24998 8449
rect 26145 8449 26157 8452
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 22204 8384 22876 8412
rect 23017 8415 23075 8421
rect 22005 8375 22063 8381
rect 23017 8381 23029 8415
rect 23063 8412 23075 8415
rect 23842 8412 23848 8424
rect 23063 8384 23848 8412
rect 23063 8381 23075 8384
rect 23017 8375 23075 8381
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 26234 8372 26240 8424
rect 26292 8412 26298 8424
rect 26697 8415 26755 8421
rect 26697 8412 26709 8415
rect 26292 8384 26709 8412
rect 26292 8372 26298 8384
rect 26697 8381 26709 8384
rect 26743 8381 26755 8415
rect 26804 8412 26832 8520
rect 29724 8517 29736 8551
rect 29770 8548 29782 8551
rect 30668 8548 30696 8576
rect 29770 8520 30696 8548
rect 30852 8548 30880 8579
rect 31202 8576 31208 8588
rect 31260 8576 31266 8628
rect 31297 8619 31355 8625
rect 31297 8585 31309 8619
rect 31343 8616 31355 8619
rect 32674 8616 32680 8628
rect 31343 8588 32680 8616
rect 31343 8585 31355 8588
rect 31297 8579 31355 8585
rect 32674 8576 32680 8588
rect 32732 8576 32738 8628
rect 32766 8576 32772 8628
rect 32824 8576 32830 8628
rect 32950 8576 32956 8628
rect 33008 8616 33014 8628
rect 33321 8619 33379 8625
rect 33321 8616 33333 8619
rect 33008 8588 33333 8616
rect 33008 8576 33014 8588
rect 33321 8585 33333 8588
rect 33367 8585 33379 8619
rect 33321 8579 33379 8585
rect 33689 8619 33747 8625
rect 33689 8585 33701 8619
rect 33735 8616 33747 8619
rect 33962 8616 33968 8628
rect 33735 8588 33968 8616
rect 33735 8585 33747 8588
rect 33689 8579 33747 8585
rect 33962 8576 33968 8588
rect 34020 8576 34026 8628
rect 34422 8576 34428 8628
rect 34480 8576 34486 8628
rect 35805 8619 35863 8625
rect 35805 8585 35817 8619
rect 35851 8616 35863 8619
rect 36170 8616 36176 8628
rect 35851 8588 36176 8616
rect 35851 8585 35863 8588
rect 35805 8579 35863 8585
rect 36170 8576 36176 8588
rect 36228 8616 36234 8628
rect 36630 8616 36636 8628
rect 36228 8588 36636 8616
rect 36228 8576 36234 8588
rect 36630 8576 36636 8588
rect 36688 8576 36694 8628
rect 36725 8619 36783 8625
rect 36725 8585 36737 8619
rect 36771 8616 36783 8619
rect 37366 8616 37372 8628
rect 36771 8588 37372 8616
rect 36771 8585 36783 8588
rect 36725 8579 36783 8585
rect 37366 8576 37372 8588
rect 37424 8576 37430 8628
rect 38378 8576 38384 8628
rect 38436 8576 38442 8628
rect 31662 8548 31668 8560
rect 30852 8520 31668 8548
rect 29770 8517 29782 8520
rect 29724 8511 29782 8517
rect 31662 8508 31668 8520
rect 31720 8548 31726 8560
rect 32784 8548 32812 8576
rect 31720 8520 32812 8548
rect 31720 8508 31726 8520
rect 33042 8508 33048 8560
rect 33100 8548 33106 8560
rect 34057 8551 34115 8557
rect 34057 8548 34069 8551
rect 33100 8520 34069 8548
rect 33100 8508 33106 8520
rect 34057 8517 34069 8520
rect 34103 8517 34115 8551
rect 34440 8548 34468 8576
rect 34057 8511 34115 8517
rect 34256 8520 34836 8548
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8480 27399 8483
rect 27801 8483 27859 8489
rect 27801 8480 27813 8483
rect 27387 8452 27813 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 27801 8449 27813 8452
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 31389 8483 31447 8489
rect 31389 8449 31401 8483
rect 31435 8480 31447 8483
rect 32493 8483 32551 8489
rect 32493 8480 32505 8483
rect 31435 8452 32505 8480
rect 31435 8449 31447 8452
rect 31389 8443 31447 8449
rect 32493 8449 32505 8452
rect 32539 8480 32551 8483
rect 33229 8483 33287 8489
rect 33229 8480 33241 8483
rect 32539 8452 33241 8480
rect 32539 8449 32551 8452
rect 32493 8443 32551 8449
rect 33229 8449 33241 8452
rect 33275 8449 33287 8483
rect 33229 8443 33287 8449
rect 27065 8415 27123 8421
rect 27065 8412 27077 8415
rect 26804 8384 27077 8412
rect 26697 8375 26755 8381
rect 27065 8381 27077 8384
rect 27111 8412 27123 8415
rect 27154 8412 27160 8424
rect 27111 8384 27160 8412
rect 27111 8381 27123 8384
rect 27065 8375 27123 8381
rect 27154 8372 27160 8384
rect 27212 8372 27218 8424
rect 27249 8415 27307 8421
rect 27249 8381 27261 8415
rect 27295 8381 27307 8415
rect 27249 8375 27307 8381
rect 13081 8347 13139 8353
rect 13081 8313 13093 8347
rect 13127 8313 13139 8347
rect 13081 8307 13139 8313
rect 16485 8347 16543 8353
rect 16485 8313 16497 8347
rect 16531 8344 16543 8347
rect 18509 8347 18567 8353
rect 16531 8316 16988 8344
rect 16531 8313 16543 8316
rect 16485 8307 16543 8313
rect 16960 8288 16988 8316
rect 18509 8313 18521 8347
rect 18555 8313 18567 8347
rect 18509 8307 18567 8313
rect 21637 8347 21695 8353
rect 21637 8313 21649 8347
rect 21683 8313 21695 8347
rect 21744 8344 21772 8372
rect 22370 8344 22376 8356
rect 21744 8316 22376 8344
rect 21637 8307 21695 8313
rect 22370 8304 22376 8316
rect 22428 8304 22434 8356
rect 22465 8347 22523 8353
rect 22465 8313 22477 8347
rect 22511 8313 22523 8347
rect 22465 8307 22523 8313
rect 6880 8248 8616 8276
rect 6880 8236 6886 8248
rect 9858 8236 9864 8288
rect 9916 8236 9922 8288
rect 10686 8236 10692 8288
rect 10744 8236 10750 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 13262 8276 13268 8288
rect 11848 8248 13268 8276
rect 11848 8236 11854 8248
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 16942 8236 16948 8288
rect 17000 8236 17006 8288
rect 17126 8236 17132 8288
rect 17184 8276 17190 8288
rect 17770 8276 17776 8288
rect 17184 8248 17776 8276
rect 17184 8236 17190 8248
rect 17770 8236 17776 8248
rect 17828 8276 17834 8288
rect 18322 8276 18328 8288
rect 17828 8248 18328 8276
rect 17828 8236 17834 8248
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 18598 8236 18604 8288
rect 18656 8236 18662 8288
rect 22480 8276 22508 8307
rect 23658 8304 23664 8356
rect 23716 8304 23722 8356
rect 23198 8276 23204 8288
rect 22480 8248 23204 8276
rect 23198 8236 23204 8248
rect 23256 8236 23262 8288
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 23753 8279 23811 8285
rect 23753 8276 23765 8279
rect 23532 8248 23765 8276
rect 23532 8236 23538 8248
rect 23753 8245 23765 8248
rect 23799 8245 23811 8279
rect 27264 8276 27292 8375
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 28537 8415 28595 8421
rect 28537 8381 28549 8415
rect 28583 8381 28595 8415
rect 28537 8375 28595 8381
rect 27709 8347 27767 8353
rect 27709 8313 27721 8347
rect 27755 8344 27767 8347
rect 28552 8344 28580 8375
rect 29454 8372 29460 8424
rect 29512 8372 29518 8424
rect 31404 8344 31432 8443
rect 31478 8372 31484 8424
rect 31536 8412 31542 8424
rect 31573 8415 31631 8421
rect 31573 8412 31585 8415
rect 31536 8384 31585 8412
rect 31536 8372 31542 8384
rect 31573 8381 31585 8384
rect 31619 8381 31631 8415
rect 31573 8375 31631 8381
rect 27755 8316 28580 8344
rect 30392 8316 31432 8344
rect 31588 8344 31616 8375
rect 32582 8372 32588 8424
rect 32640 8372 32646 8424
rect 32769 8415 32827 8421
rect 32769 8381 32781 8415
rect 32815 8412 32827 8415
rect 33042 8412 33048 8424
rect 32815 8384 33048 8412
rect 32815 8381 32827 8384
rect 32769 8375 32827 8381
rect 33042 8372 33048 8384
rect 33100 8372 33106 8424
rect 33137 8415 33195 8421
rect 33137 8381 33149 8415
rect 33183 8412 33195 8415
rect 33318 8412 33324 8424
rect 33183 8384 33324 8412
rect 33183 8381 33195 8384
rect 33137 8375 33195 8381
rect 33318 8372 33324 8384
rect 33376 8412 33382 8424
rect 34256 8412 34284 8520
rect 34330 8440 34336 8492
rect 34388 8440 34394 8492
rect 34425 8483 34483 8489
rect 34425 8449 34437 8483
rect 34471 8480 34483 8483
rect 34514 8480 34520 8492
rect 34471 8452 34520 8480
rect 34471 8449 34483 8452
rect 34425 8443 34483 8449
rect 34514 8440 34520 8452
rect 34572 8440 34578 8492
rect 34698 8489 34704 8492
rect 34692 8443 34704 8489
rect 34698 8440 34704 8443
rect 34756 8440 34762 8492
rect 34808 8480 34836 8520
rect 35986 8508 35992 8560
rect 36044 8548 36050 8560
rect 36357 8551 36415 8557
rect 36357 8548 36369 8551
rect 36044 8520 36369 8548
rect 36044 8508 36050 8520
rect 36357 8517 36369 8520
rect 36403 8548 36415 8551
rect 36403 8520 37228 8548
rect 36403 8517 36415 8520
rect 36357 8511 36415 8517
rect 37200 8492 37228 8520
rect 34808 8452 36400 8480
rect 33376 8384 34284 8412
rect 33376 8372 33382 8384
rect 36078 8372 36084 8424
rect 36136 8372 36142 8424
rect 36265 8415 36323 8421
rect 36265 8381 36277 8415
rect 36311 8381 36323 8415
rect 36372 8412 36400 8452
rect 36446 8440 36452 8492
rect 36504 8480 36510 8492
rect 37001 8483 37059 8489
rect 37001 8480 37013 8483
rect 36504 8452 37013 8480
rect 36504 8440 36510 8452
rect 37001 8449 37013 8452
rect 37047 8449 37059 8483
rect 37001 8443 37059 8449
rect 37182 8440 37188 8492
rect 37240 8440 37246 8492
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 38197 8483 38255 8489
rect 38197 8449 38209 8483
rect 38243 8480 38255 8483
rect 38286 8480 38292 8492
rect 38243 8452 38292 8480
rect 38243 8449 38255 8452
rect 38197 8443 38255 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 36372 8384 38332 8412
rect 36265 8375 36323 8381
rect 31588 8316 32812 8344
rect 27755 8313 27767 8316
rect 27709 8307 27767 8313
rect 27338 8276 27344 8288
rect 27264 8248 27344 8276
rect 23753 8239 23811 8245
rect 27338 8236 27344 8248
rect 27396 8236 27402 8288
rect 29178 8236 29184 8288
rect 29236 8236 29242 8288
rect 30190 8236 30196 8288
rect 30248 8276 30254 8288
rect 30392 8276 30420 8316
rect 30248 8248 30420 8276
rect 30248 8236 30254 8248
rect 31570 8236 31576 8288
rect 31628 8276 31634 8288
rect 31846 8276 31852 8288
rect 31628 8248 31852 8276
rect 31628 8236 31634 8248
rect 31846 8236 31852 8248
rect 31904 8236 31910 8288
rect 32125 8279 32183 8285
rect 32125 8245 32137 8279
rect 32171 8276 32183 8279
rect 32674 8276 32680 8288
rect 32171 8248 32680 8276
rect 32171 8245 32183 8248
rect 32125 8239 32183 8245
rect 32674 8236 32680 8248
rect 32732 8236 32738 8288
rect 32784 8276 32812 8316
rect 34054 8304 34060 8356
rect 34112 8344 34118 8356
rect 34149 8347 34207 8353
rect 34149 8344 34161 8347
rect 34112 8316 34161 8344
rect 34112 8304 34118 8316
rect 34149 8313 34161 8316
rect 34195 8313 34207 8347
rect 34149 8307 34207 8313
rect 34238 8304 34244 8356
rect 34296 8304 34302 8356
rect 36280 8344 36308 8375
rect 38304 8356 38332 8384
rect 37274 8344 37280 8356
rect 36280 8316 37280 8344
rect 37274 8304 37280 8316
rect 37332 8304 37338 8356
rect 37461 8347 37519 8353
rect 37461 8313 37473 8347
rect 37507 8344 37519 8347
rect 37642 8344 37648 8356
rect 37507 8316 37648 8344
rect 37507 8313 37519 8316
rect 37461 8307 37519 8313
rect 37642 8304 37648 8316
rect 37700 8304 37706 8356
rect 37734 8304 37740 8356
rect 37792 8304 37798 8356
rect 38286 8304 38292 8356
rect 38344 8304 38350 8356
rect 34256 8276 34284 8304
rect 32784 8248 34284 8276
rect 36538 8236 36544 8288
rect 36596 8276 36602 8288
rect 36817 8279 36875 8285
rect 36817 8276 36829 8279
rect 36596 8248 36829 8276
rect 36596 8236 36602 8248
rect 36817 8245 36829 8248
rect 36863 8245 36875 8279
rect 36817 8239 36875 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 3878 8032 3884 8084
rect 3936 8032 3942 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4028 8044 4629 8072
rect 4028 8032 4034 8044
rect 4617 8041 4629 8044
rect 4663 8072 4675 8075
rect 5442 8072 5448 8084
rect 4663 8044 5448 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 6730 8072 6736 8084
rect 6687 8044 6736 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12066 8072 12072 8084
rect 11112 8044 12072 8072
rect 11112 8032 11118 8044
rect 12066 8032 12072 8044
rect 12124 8072 12130 8084
rect 13633 8075 13691 8081
rect 12124 8044 13216 8072
rect 12124 8032 12130 8044
rect 4172 7976 4384 8004
rect 4172 7945 4200 7976
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 4157 7939 4215 7945
rect 2915 7908 4016 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 2590 7828 2596 7880
rect 2648 7868 2654 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2648 7840 2697 7868
rect 2648 7828 2654 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2823 7840 2912 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2884 7744 2912 7840
rect 3145 7803 3203 7809
rect 3145 7769 3157 7803
rect 3191 7800 3203 7803
rect 3878 7800 3884 7812
rect 3191 7772 3884 7800
rect 3191 7769 3203 7772
rect 3145 7763 3203 7769
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 3988 7800 4016 7908
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4356 7936 4384 7976
rect 9490 7964 9496 8016
rect 9548 8004 9554 8016
rect 10042 8004 10048 8016
rect 9548 7976 10048 8004
rect 9548 7964 9554 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 5258 7936 5264 7948
rect 4356 7908 5264 7936
rect 4157 7899 4215 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 8812 7908 10456 7936
rect 8812 7896 8818 7908
rect 4062 7828 4068 7880
rect 4120 7877 4126 7880
rect 4120 7871 4137 7877
rect 4125 7837 4137 7871
rect 5902 7868 5908 7880
rect 4120 7831 4137 7837
rect 4172 7840 5908 7868
rect 4120 7828 4126 7831
rect 4172 7800 4200 7840
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8312 7840 8953 7868
rect 8312 7812 8340 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 9398 7868 9404 7880
rect 8987 7840 9404 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9674 7828 9680 7880
rect 9732 7828 9738 7880
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10428 7877 10456 7908
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 13188 7936 13216 8044
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13722 8072 13728 8084
rect 13679 8044 13728 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13722 8032 13728 8044
rect 13780 8072 13786 8084
rect 14734 8072 14740 8084
rect 13780 8044 14740 8072
rect 13780 8032 13786 8044
rect 14734 8032 14740 8044
rect 14792 8072 14798 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14792 8044 14841 8072
rect 14792 8032 14798 8044
rect 14829 8041 14841 8044
rect 14875 8041 14887 8075
rect 14829 8035 14887 8041
rect 15381 8075 15439 8081
rect 15381 8041 15393 8075
rect 15427 8072 15439 8075
rect 15930 8072 15936 8084
rect 15427 8044 15936 8072
rect 15427 8041 15439 8044
rect 15381 8035 15439 8041
rect 13265 8007 13323 8013
rect 13265 7973 13277 8007
rect 13311 8004 13323 8007
rect 13814 8004 13820 8016
rect 13311 7976 13820 8004
rect 13311 7973 13323 7976
rect 13265 7967 13323 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 13906 7964 13912 8016
rect 13964 7964 13970 8016
rect 13924 7936 13952 7964
rect 13188 7908 13952 7936
rect 14844 7936 14872 8035
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 17037 8075 17095 8081
rect 17037 8041 17049 8075
rect 17083 8072 17095 8075
rect 18138 8072 18144 8084
rect 17083 8044 18144 8072
rect 17083 8041 17095 8044
rect 17037 8035 17095 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18230 8032 18236 8084
rect 18288 8032 18294 8084
rect 19610 8032 19616 8084
rect 19668 8072 19674 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 19668 8044 20545 8072
rect 19668 8032 19674 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 20533 8035 20591 8041
rect 23569 8075 23627 8081
rect 23569 8041 23581 8075
rect 23615 8072 23627 8075
rect 23750 8072 23756 8084
rect 23615 8044 23756 8072
rect 23615 8041 23627 8044
rect 23569 8035 23627 8041
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 23842 8032 23848 8084
rect 23900 8072 23906 8084
rect 24581 8075 24639 8081
rect 24581 8072 24593 8075
rect 23900 8044 24593 8072
rect 23900 8032 23906 8044
rect 24581 8041 24593 8044
rect 24627 8041 24639 8075
rect 24581 8035 24639 8041
rect 25593 8075 25651 8081
rect 25593 8041 25605 8075
rect 25639 8072 25651 8075
rect 26234 8072 26240 8084
rect 25639 8044 26240 8072
rect 25639 8041 25651 8044
rect 25593 8035 25651 8041
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 15289 8007 15347 8013
rect 15289 8004 15301 8007
rect 15160 7976 15301 8004
rect 15160 7964 15166 7976
rect 15289 7973 15301 7976
rect 15335 8004 15347 8007
rect 17126 8004 17132 8016
rect 15335 7976 17132 8004
rect 15335 7973 15347 7976
rect 15289 7967 15347 7973
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 18248 8004 18276 8032
rect 24596 8004 24624 8035
rect 26234 8032 26240 8044
rect 26292 8032 26298 8084
rect 27617 8075 27675 8081
rect 27617 8072 27629 8075
rect 27356 8044 27629 8072
rect 18248 7976 18920 8004
rect 24596 7976 26004 8004
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 14844 7908 15945 7936
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 16264 7908 16313 7936
rect 16264 7896 16270 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17819 7939 17877 7945
rect 17819 7936 17831 7939
rect 17000 7908 17831 7936
rect 17000 7896 17006 7908
rect 17819 7905 17831 7908
rect 17865 7905 17877 7939
rect 17819 7899 17877 7905
rect 18233 7939 18291 7945
rect 18233 7905 18245 7939
rect 18279 7936 18291 7939
rect 18322 7936 18328 7948
rect 18279 7908 18328 7936
rect 18279 7905 18291 7908
rect 18233 7899 18291 7905
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 18690 7896 18696 7948
rect 18748 7896 18754 7948
rect 18892 7945 18920 7976
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 19797 7939 19855 7945
rect 19797 7936 19809 7939
rect 18923 7908 19809 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 19797 7905 19809 7908
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 21174 7896 21180 7948
rect 21232 7896 21238 7948
rect 23014 7896 23020 7948
rect 23072 7896 23078 7948
rect 23109 7939 23167 7945
rect 23109 7905 23121 7939
rect 23155 7936 23167 7939
rect 23474 7936 23480 7948
rect 23155 7908 23480 7936
rect 23155 7905 23167 7908
rect 23109 7899 23167 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 25038 7896 25044 7948
rect 25096 7896 25102 7948
rect 25976 7936 26004 7976
rect 26142 7936 26148 7948
rect 25976 7908 26148 7936
rect 26142 7896 26148 7908
rect 26200 7936 26206 7948
rect 26329 7939 26387 7945
rect 26329 7936 26341 7939
rect 26200 7908 26341 7936
rect 26200 7896 26206 7908
rect 26329 7905 26341 7908
rect 26375 7905 26387 7939
rect 26329 7899 26387 7905
rect 26418 7896 26424 7948
rect 26476 7945 26482 7948
rect 26476 7939 26525 7945
rect 26476 7905 26479 7939
rect 26513 7905 26525 7939
rect 26476 7899 26525 7905
rect 26476 7896 26482 7899
rect 26602 7896 26608 7948
rect 26660 7896 26666 7948
rect 26786 7896 26792 7948
rect 26844 7936 26850 7948
rect 27356 7945 27384 8044
rect 27617 8041 27629 8044
rect 27663 8072 27675 8075
rect 28350 8072 28356 8084
rect 27663 8044 28356 8072
rect 27663 8041 27675 8044
rect 27617 8035 27675 8041
rect 28350 8032 28356 8044
rect 28408 8032 28414 8084
rect 29825 8075 29883 8081
rect 29825 8041 29837 8075
rect 29871 8072 29883 8075
rect 29914 8072 29920 8084
rect 29871 8044 29920 8072
rect 29871 8041 29883 8044
rect 29825 8035 29883 8041
rect 29914 8032 29920 8044
rect 29972 8032 29978 8084
rect 30668 8044 32260 8072
rect 30668 7948 30696 8044
rect 31110 7964 31116 8016
rect 31168 8004 31174 8016
rect 31168 7976 31432 8004
rect 31168 7964 31174 7976
rect 26881 7939 26939 7945
rect 26881 7936 26893 7939
rect 26844 7908 26893 7936
rect 26844 7896 26850 7908
rect 26881 7905 26893 7908
rect 26927 7936 26939 7939
rect 27341 7939 27399 7945
rect 26927 7908 27200 7936
rect 26927 7905 26939 7908
rect 26881 7899 26939 7905
rect 10413 7871 10471 7877
rect 9824 7840 10180 7868
rect 9824 7828 9830 7840
rect 3988 7772 4200 7800
rect 4264 7772 4568 7800
rect 2866 7692 2872 7744
rect 2924 7692 2930 7744
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3510 7732 3516 7744
rect 3108 7704 3516 7732
rect 3108 7692 3114 7704
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 4264 7732 4292 7772
rect 3660 7704 4292 7732
rect 3660 7692 3666 7704
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 4540 7732 4568 7772
rect 4706 7760 4712 7812
rect 4764 7800 4770 7812
rect 4801 7803 4859 7809
rect 4801 7800 4813 7803
rect 4764 7772 4813 7800
rect 4764 7760 4770 7772
rect 4801 7769 4813 7772
rect 4847 7769 4859 7803
rect 4801 7763 4859 7769
rect 8294 7760 8300 7812
rect 8352 7760 8358 7812
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8512 7803 8570 7809
rect 8512 7769 8524 7803
rect 8558 7800 8570 7803
rect 9692 7800 9720 7828
rect 10152 7812 10180 7840
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 11624 7868 11652 7896
rect 10459 7840 11652 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7868 15807 7871
rect 16114 7868 16120 7880
rect 15795 7840 16120 7868
rect 15795 7837 15807 7840
rect 15749 7831 15807 7837
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 17678 7828 17684 7880
rect 17736 7828 17742 7880
rect 17954 7828 17960 7880
rect 18012 7828 18018 7880
rect 20898 7828 20904 7880
rect 20956 7828 20962 7880
rect 20993 7871 21051 7877
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 21039 7840 22094 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 8558 7772 9720 7800
rect 8558 7769 8570 7772
rect 8512 7763 8570 7769
rect 10134 7760 10140 7812
rect 10192 7760 10198 7812
rect 10686 7809 10692 7812
rect 10680 7800 10692 7809
rect 10647 7772 10692 7800
rect 10680 7763 10692 7772
rect 10686 7760 10692 7763
rect 10744 7760 10750 7812
rect 12158 7809 12164 7812
rect 12152 7763 12164 7809
rect 12158 7760 12164 7763
rect 12216 7760 12222 7812
rect 12802 7800 12808 7812
rect 12406 7772 12808 7800
rect 4596 7735 4654 7741
rect 4596 7732 4608 7735
rect 4540 7704 4608 7732
rect 4596 7701 4608 7704
rect 4642 7732 4654 7735
rect 4890 7732 4896 7744
rect 4642 7704 4896 7732
rect 4642 7701 4654 7704
rect 4596 7695 4654 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 7377 7735 7435 7741
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 8110 7732 8116 7744
rect 7423 7704 8116 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8404 7732 8432 7760
rect 9674 7732 9680 7744
rect 8404 7704 9680 7732
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 10100 7704 10333 7732
rect 10100 7692 10106 7704
rect 10321 7701 10333 7704
rect 10367 7732 10379 7735
rect 10962 7732 10968 7744
rect 10367 7704 10968 7732
rect 10367 7701 10379 7704
rect 10321 7695 10379 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11793 7735 11851 7741
rect 11793 7701 11805 7735
rect 11839 7732 11851 7735
rect 12406 7732 12434 7772
rect 12802 7760 12808 7772
rect 12860 7800 12866 7812
rect 14458 7800 14464 7812
rect 12860 7772 14464 7800
rect 12860 7760 12866 7772
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 16485 7803 16543 7809
rect 16485 7769 16497 7803
rect 16531 7800 16543 7803
rect 16531 7772 17264 7800
rect 16531 7769 16543 7772
rect 16485 7763 16543 7769
rect 11839 7704 12434 7732
rect 15841 7735 15899 7741
rect 11839 7701 11851 7704
rect 11793 7695 11851 7701
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 16206 7732 16212 7744
rect 15887 7704 16212 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 16206 7692 16212 7704
rect 16264 7732 16270 7744
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 16264 7704 16589 7732
rect 16264 7692 16270 7704
rect 16577 7701 16589 7704
rect 16623 7701 16635 7735
rect 16577 7695 16635 7701
rect 16942 7692 16948 7744
rect 17000 7692 17006 7744
rect 17236 7732 17264 7772
rect 18138 7732 18144 7744
rect 17236 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 18472 7704 19257 7732
rect 18472 7692 18478 7704
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19245 7695 19303 7701
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21910 7732 21916 7744
rect 21416 7704 21916 7732
rect 21416 7692 21422 7704
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22066 7732 22094 7840
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22741 7871 22799 7877
rect 22741 7868 22753 7871
rect 22244 7840 22753 7868
rect 22244 7828 22250 7840
rect 22741 7837 22753 7840
rect 22787 7837 22799 7871
rect 23032 7868 23060 7896
rect 27172 7868 27200 7908
rect 27341 7905 27353 7939
rect 27387 7905 27399 7939
rect 27341 7899 27399 7905
rect 27525 7939 27583 7945
rect 27525 7905 27537 7939
rect 27571 7936 27583 7939
rect 27614 7936 27620 7948
rect 27571 7908 27620 7936
rect 27571 7905 27583 7908
rect 27525 7899 27583 7905
rect 27614 7896 27620 7908
rect 27672 7896 27678 7948
rect 29365 7939 29423 7945
rect 29365 7905 29377 7939
rect 29411 7936 29423 7939
rect 30282 7936 30288 7948
rect 29411 7908 30288 7936
rect 29411 7905 29423 7908
rect 29365 7899 29423 7905
rect 30282 7896 30288 7908
rect 30340 7936 30346 7948
rect 30377 7939 30435 7945
rect 30377 7936 30389 7939
rect 30340 7908 30389 7936
rect 30340 7896 30346 7908
rect 30377 7905 30389 7908
rect 30423 7905 30435 7939
rect 30377 7899 30435 7905
rect 30650 7896 30656 7948
rect 30708 7896 30714 7948
rect 30834 7896 30840 7948
rect 30892 7896 30898 7948
rect 31202 7896 31208 7948
rect 31260 7936 31266 7948
rect 31297 7939 31355 7945
rect 31297 7936 31309 7939
rect 31260 7908 31309 7936
rect 31260 7896 31266 7908
rect 31297 7905 31309 7908
rect 31343 7905 31355 7939
rect 31404 7936 31432 7976
rect 31573 7939 31631 7945
rect 31573 7936 31585 7939
rect 31404 7908 31585 7936
rect 31297 7899 31355 7905
rect 31573 7905 31585 7908
rect 31619 7905 31631 7939
rect 31573 7899 31631 7905
rect 31662 7896 31668 7948
rect 31720 7945 31726 7948
rect 31720 7939 31748 7945
rect 31736 7905 31748 7939
rect 31720 7899 31748 7905
rect 31720 7896 31726 7899
rect 31846 7896 31852 7948
rect 31904 7896 31910 7948
rect 32232 7936 32260 8044
rect 32582 8032 32588 8084
rect 32640 8032 32646 8084
rect 33597 8075 33655 8081
rect 33597 8041 33609 8075
rect 33643 8072 33655 8075
rect 33870 8072 33876 8084
rect 33643 8044 33876 8072
rect 33643 8041 33655 8044
rect 33597 8035 33655 8041
rect 33870 8032 33876 8044
rect 33928 8032 33934 8084
rect 36078 8072 36084 8084
rect 34440 8044 36084 8072
rect 33137 7939 33195 7945
rect 33137 7936 33149 7939
rect 32232 7908 33149 7936
rect 33137 7905 33149 7908
rect 33183 7905 33195 7939
rect 33137 7899 33195 7905
rect 33965 7939 34023 7945
rect 33965 7905 33977 7939
rect 34011 7936 34023 7939
rect 34146 7936 34152 7948
rect 34011 7908 34152 7936
rect 34011 7905 34023 7908
rect 33965 7899 34023 7905
rect 34146 7896 34152 7908
rect 34204 7896 34210 7948
rect 34440 7880 34468 8044
rect 36078 8032 36084 8044
rect 36136 8032 36142 8084
rect 34514 7896 34520 7948
rect 34572 7936 34578 7948
rect 34701 7939 34759 7945
rect 34701 7936 34713 7939
rect 34572 7908 34713 7936
rect 34572 7896 34578 7908
rect 34701 7905 34713 7908
rect 34747 7905 34759 7939
rect 34701 7899 34759 7905
rect 28997 7871 29055 7877
rect 23032 7840 23980 7868
rect 27172 7840 27384 7868
rect 22741 7831 22799 7837
rect 22496 7803 22554 7809
rect 22496 7769 22508 7803
rect 22542 7800 22554 7803
rect 23474 7800 23480 7812
rect 22542 7772 23480 7800
rect 22542 7769 22554 7772
rect 22496 7763 22554 7769
rect 23474 7760 23480 7772
rect 23532 7760 23538 7812
rect 22922 7732 22928 7744
rect 22066 7704 22928 7732
rect 22922 7692 22928 7704
rect 22980 7732 22986 7744
rect 23952 7741 23980 7840
rect 25225 7803 25283 7809
rect 25225 7769 25237 7803
rect 25271 7800 25283 7803
rect 25271 7772 25912 7800
rect 25271 7769 25283 7772
rect 25225 7763 25283 7769
rect 23201 7735 23259 7741
rect 23201 7732 23213 7735
rect 22980 7704 23213 7732
rect 22980 7692 22986 7704
rect 23201 7701 23213 7704
rect 23247 7701 23259 7735
rect 23201 7695 23259 7701
rect 23937 7735 23995 7741
rect 23937 7701 23949 7735
rect 23983 7732 23995 7735
rect 24210 7732 24216 7744
rect 23983 7704 24216 7732
rect 23983 7701 23995 7704
rect 23937 7695 23995 7701
rect 24210 7692 24216 7704
rect 24268 7692 24274 7744
rect 25130 7692 25136 7744
rect 25188 7692 25194 7744
rect 25682 7692 25688 7744
rect 25740 7692 25746 7744
rect 25884 7732 25912 7772
rect 26510 7732 26516 7744
rect 25884 7704 26516 7732
rect 26510 7692 26516 7704
rect 26568 7692 26574 7744
rect 27356 7732 27384 7840
rect 28997 7837 29009 7871
rect 29043 7868 29055 7871
rect 29454 7868 29460 7880
rect 29043 7840 29460 7868
rect 29043 7837 29055 7840
rect 28997 7831 29055 7837
rect 29454 7828 29460 7840
rect 29512 7828 29518 7880
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 30190 7868 30196 7880
rect 29972 7840 30196 7868
rect 29972 7828 29978 7840
rect 30190 7828 30196 7840
rect 30248 7828 30254 7880
rect 33413 7871 33471 7877
rect 33413 7837 33425 7871
rect 33459 7837 33471 7871
rect 33413 7831 33471 7837
rect 34057 7871 34115 7877
rect 34057 7837 34069 7871
rect 34103 7868 34115 7871
rect 34238 7868 34244 7880
rect 34103 7840 34244 7868
rect 34103 7837 34115 7840
rect 34057 7831 34115 7837
rect 28752 7803 28810 7809
rect 28752 7769 28764 7803
rect 28798 7800 28810 7803
rect 29178 7800 29184 7812
rect 28798 7772 29184 7800
rect 28798 7769 28810 7772
rect 28752 7763 28810 7769
rect 29178 7760 29184 7772
rect 29236 7760 29242 7812
rect 33428 7800 33456 7831
rect 34238 7828 34244 7840
rect 34296 7828 34302 7880
rect 34422 7828 34428 7880
rect 34480 7828 34486 7880
rect 34716 7868 34744 7899
rect 37182 7896 37188 7948
rect 37240 7936 37246 7948
rect 38105 7939 38163 7945
rect 38105 7936 38117 7939
rect 37240 7908 38117 7936
rect 37240 7896 37246 7908
rect 38105 7905 38117 7908
rect 38151 7905 38163 7939
rect 38105 7899 38163 7905
rect 38286 7896 38292 7948
rect 38344 7896 38350 7948
rect 36173 7871 36231 7877
rect 36173 7868 36185 7871
rect 34716 7840 36185 7868
rect 36173 7837 36185 7840
rect 36219 7837 36231 7871
rect 36173 7831 36231 7837
rect 36440 7871 36498 7877
rect 36440 7837 36452 7871
rect 36486 7868 36498 7871
rect 36814 7868 36820 7880
rect 36486 7840 36820 7868
rect 36486 7837 36498 7840
rect 36440 7831 36498 7837
rect 36814 7828 36820 7840
rect 36872 7828 36878 7880
rect 34968 7803 35026 7809
rect 33428 7772 34928 7800
rect 28994 7732 29000 7744
rect 27356 7704 29000 7732
rect 28994 7692 29000 7704
rect 29052 7692 29058 7744
rect 30285 7735 30343 7741
rect 30285 7701 30297 7735
rect 30331 7732 30343 7735
rect 30742 7732 30748 7744
rect 30331 7704 30748 7732
rect 30331 7701 30343 7704
rect 30285 7695 30343 7701
rect 30742 7692 30748 7704
rect 30800 7692 30806 7744
rect 32490 7692 32496 7744
rect 32548 7692 32554 7744
rect 34146 7692 34152 7744
rect 34204 7692 34210 7744
rect 34514 7692 34520 7744
rect 34572 7692 34578 7744
rect 34900 7732 34928 7772
rect 34968 7769 34980 7803
rect 35014 7800 35026 7803
rect 35158 7800 35164 7812
rect 35014 7772 35164 7800
rect 35014 7769 35026 7772
rect 34968 7763 35026 7769
rect 35158 7760 35164 7772
rect 35216 7760 35222 7812
rect 36722 7800 36728 7812
rect 36004 7772 36728 7800
rect 36004 7732 36032 7772
rect 36722 7760 36728 7772
rect 36780 7760 36786 7812
rect 34900 7704 36032 7732
rect 37550 7692 37556 7744
rect 37608 7692 37614 7744
rect 37645 7735 37703 7741
rect 37645 7701 37657 7735
rect 37691 7732 37703 7735
rect 37918 7732 37924 7744
rect 37691 7704 37924 7732
rect 37691 7701 37703 7704
rect 37645 7695 37703 7701
rect 37918 7692 37924 7704
rect 37976 7692 37982 7744
rect 38010 7692 38016 7744
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2648 7500 3096 7528
rect 2648 7488 2654 7500
rect 3068 7401 3096 7500
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 3384 7500 4384 7528
rect 3384 7488 3390 7500
rect 3510 7420 3516 7472
rect 3568 7460 3574 7472
rect 3568 7432 4108 7460
rect 3568 7420 3574 7432
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7361 3111 7395
rect 3053 7355 3111 7361
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3752 7364 3801 7392
rect 3752 7352 3758 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 4080 7401 4108 7432
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4154 7352 4160 7404
rect 4212 7352 4218 7404
rect 4356 7392 4384 7500
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4706 7528 4712 7540
rect 4488 7500 4712 7528
rect 4488 7488 4494 7500
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 4948 7500 5580 7528
rect 4948 7488 4954 7500
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 5261 7463 5319 7469
rect 5261 7460 5273 7463
rect 4856 7432 5273 7460
rect 4856 7420 4862 7432
rect 5261 7429 5273 7432
rect 5307 7429 5319 7463
rect 5261 7423 5319 7429
rect 5442 7420 5448 7472
rect 5500 7420 5506 7472
rect 5552 7401 5580 7500
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 8665 7531 8723 7537
rect 8665 7528 8677 7531
rect 7340 7500 8677 7528
rect 7340 7488 7346 7500
rect 8665 7497 8677 7500
rect 8711 7497 8723 7531
rect 8665 7491 8723 7497
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9582 7528 9588 7540
rect 9171 7500 9588 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 14366 7488 14372 7540
rect 14424 7488 14430 7540
rect 15102 7488 15108 7540
rect 15160 7488 15166 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15749 7531 15807 7537
rect 15749 7528 15761 7531
rect 15528 7500 15761 7528
rect 15528 7488 15534 7500
rect 15749 7497 15761 7500
rect 15795 7497 15807 7531
rect 15749 7491 15807 7497
rect 17678 7488 17684 7540
rect 17736 7528 17742 7540
rect 18417 7531 18475 7537
rect 18417 7528 18429 7531
rect 17736 7500 18429 7528
rect 17736 7488 17742 7500
rect 18417 7497 18429 7500
rect 18463 7497 18475 7531
rect 18417 7491 18475 7497
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 18598 7528 18604 7540
rect 18555 7500 18604 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7528 18935 7531
rect 18966 7528 18972 7540
rect 18923 7500 18972 7528
rect 18923 7497 18935 7500
rect 18877 7491 18935 7497
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 21174 7488 21180 7540
rect 21232 7528 21238 7540
rect 21361 7531 21419 7537
rect 21361 7528 21373 7531
rect 21232 7500 21373 7528
rect 21232 7488 21238 7500
rect 21361 7497 21373 7500
rect 21407 7497 21419 7531
rect 21361 7491 21419 7497
rect 24394 7488 24400 7540
rect 24452 7488 24458 7540
rect 27246 7488 27252 7540
rect 27304 7488 27310 7540
rect 28258 7488 28264 7540
rect 28316 7488 28322 7540
rect 30285 7531 30343 7537
rect 30285 7497 30297 7531
rect 30331 7528 30343 7531
rect 30650 7528 30656 7540
rect 30331 7500 30656 7528
rect 30331 7497 30343 7500
rect 30285 7491 30343 7497
rect 30650 7488 30656 7500
rect 30708 7488 30714 7540
rect 31202 7488 31208 7540
rect 31260 7488 31266 7540
rect 31846 7488 31852 7540
rect 31904 7528 31910 7540
rect 32582 7528 32588 7540
rect 31904 7500 32588 7528
rect 31904 7488 31910 7500
rect 32582 7488 32588 7500
rect 32640 7528 32646 7540
rect 33045 7531 33103 7537
rect 33045 7528 33057 7531
rect 32640 7500 33057 7528
rect 32640 7488 32646 7500
rect 33045 7497 33057 7500
rect 33091 7497 33103 7531
rect 33045 7491 33103 7497
rect 33781 7531 33839 7537
rect 33781 7497 33793 7531
rect 33827 7528 33839 7531
rect 34146 7528 34152 7540
rect 33827 7500 34152 7528
rect 33827 7497 33839 7500
rect 33781 7491 33839 7497
rect 9398 7420 9404 7472
rect 9456 7460 9462 7472
rect 10045 7463 10103 7469
rect 10045 7460 10057 7463
rect 9456 7432 10057 7460
rect 9456 7420 9462 7432
rect 10045 7429 10057 7432
rect 10091 7429 10103 7463
rect 13906 7460 13912 7472
rect 10045 7423 10103 7429
rect 13648 7432 13912 7460
rect 7466 7401 7472 7404
rect 5537 7395 5595 7401
rect 4356 7364 5028 7392
rect 2682 7284 2688 7336
rect 2740 7284 2746 7336
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 3142 7324 3148 7336
rect 3007 7296 3148 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 2130 7216 2136 7268
rect 2188 7256 2194 7268
rect 4632 7256 4660 7287
rect 2188 7228 4660 7256
rect 2188 7216 2194 7228
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3568 7160 3709 7188
rect 3568 7148 3574 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 3697 7151 3755 7157
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4890 7188 4896 7200
rect 4479 7160 4896 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 5000 7188 5028 7364
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 7460 7392 7472 7401
rect 7427 7364 7472 7392
rect 5537 7355 5595 7361
rect 7460 7355 7472 7364
rect 7466 7352 7472 7355
rect 7524 7352 7530 7404
rect 9030 7352 9036 7404
rect 9088 7352 9094 7404
rect 12802 7401 12808 7404
rect 12780 7395 12808 7401
rect 12780 7361 12792 7395
rect 12780 7355 12808 7361
rect 12802 7352 12808 7355
rect 12860 7352 12866 7404
rect 12894 7352 12900 7404
rect 12952 7352 12958 7404
rect 13648 7392 13676 7432
rect 13906 7420 13912 7432
rect 13964 7460 13970 7472
rect 14550 7460 14556 7472
rect 13964 7432 14556 7460
rect 13964 7420 13970 7432
rect 14550 7420 14556 7432
rect 14608 7460 14614 7472
rect 15120 7460 15148 7488
rect 16393 7463 16451 7469
rect 16393 7460 16405 7463
rect 14608 7432 15148 7460
rect 15212 7432 16405 7460
rect 14608 7420 14614 7432
rect 13556 7364 13676 7392
rect 7190 7284 7196 7336
rect 7248 7284 7254 7336
rect 8938 7284 8944 7336
rect 8996 7284 9002 7336
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11020 7296 11897 7324
rect 11020 7284 11026 7296
rect 11885 7293 11897 7296
rect 11931 7324 11943 7327
rect 12250 7324 12256 7336
rect 11931 7296 12256 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 12250 7284 12256 7296
rect 12308 7324 12314 7336
rect 12621 7327 12679 7333
rect 12621 7324 12633 7327
rect 12308 7296 12633 7324
rect 12308 7284 12314 7296
rect 12621 7293 12633 7296
rect 12667 7293 12679 7327
rect 12621 7287 12679 7293
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7324 13231 7327
rect 13556 7324 13584 7364
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 14323 7364 14749 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 13722 7333 13728 7336
rect 13219 7296 13584 7324
rect 13679 7327 13728 7333
rect 13219 7293 13231 7296
rect 13173 7287 13231 7293
rect 13679 7293 13691 7327
rect 13725 7293 13728 7327
rect 13679 7287 13728 7293
rect 13722 7284 13728 7287
rect 13780 7324 13786 7336
rect 13780 7296 14228 7324
rect 13780 7284 13786 7296
rect 5169 7259 5227 7265
rect 5169 7225 5181 7259
rect 5215 7256 5227 7259
rect 5534 7256 5540 7268
rect 5215 7228 5540 7256
rect 5215 7225 5227 7228
rect 5169 7219 5227 7225
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8956 7256 8984 7284
rect 8619 7228 8984 7256
rect 14200 7256 14228 7296
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 15212 7324 15240 7432
rect 16393 7429 16405 7432
rect 16439 7460 16451 7463
rect 16439 7432 17816 7460
rect 16439 7429 16451 7432
rect 16393 7423 16451 7429
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15436 7364 15669 7392
rect 15436 7352 15442 7364
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16925 7395 16983 7401
rect 16925 7392 16937 7395
rect 16816 7364 16937 7392
rect 16816 7352 16822 7364
rect 16925 7361 16937 7364
rect 16971 7361 16983 7395
rect 16925 7355 16983 7361
rect 14516 7296 15240 7324
rect 15289 7327 15347 7333
rect 14516 7284 14522 7296
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 17788 7324 17816 7432
rect 18046 7420 18052 7472
rect 18104 7420 18110 7472
rect 26234 7460 26240 7472
rect 25424 7432 26240 7460
rect 18064 7392 18092 7420
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18064 7364 18981 7392
rect 18969 7361 18981 7364
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 25314 7392 25320 7404
rect 22603 7364 25320 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 25314 7352 25320 7364
rect 25372 7352 25378 7404
rect 25424 7401 25452 7432
rect 26234 7420 26240 7432
rect 26292 7460 26298 7472
rect 30193 7463 30251 7469
rect 26292 7432 29776 7460
rect 26292 7420 26298 7432
rect 29748 7404 29776 7432
rect 30193 7429 30205 7463
rect 30239 7460 30251 7463
rect 31220 7460 31248 7488
rect 30239 7432 31248 7460
rect 31420 7463 31478 7469
rect 30239 7429 30251 7432
rect 30193 7423 30251 7429
rect 31420 7429 31432 7463
rect 31466 7460 31478 7463
rect 32125 7463 32183 7469
rect 32125 7460 32137 7463
rect 31466 7432 32137 7460
rect 31466 7429 31478 7432
rect 31420 7423 31478 7429
rect 32125 7429 32137 7432
rect 32171 7429 32183 7463
rect 32125 7423 32183 7429
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25676 7395 25734 7401
rect 25676 7361 25688 7395
rect 25722 7392 25734 7395
rect 27154 7392 27160 7404
rect 25722 7364 27160 7392
rect 25722 7361 25734 7364
rect 25676 7355 25734 7361
rect 27154 7352 27160 7364
rect 27212 7352 27218 7404
rect 27246 7352 27252 7404
rect 27304 7392 27310 7404
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 27304 7364 27353 7392
rect 27304 7352 27310 7364
rect 27341 7361 27353 7364
rect 27387 7361 27399 7395
rect 27341 7355 27399 7361
rect 28353 7395 28411 7401
rect 28353 7361 28365 7395
rect 28399 7392 28411 7395
rect 29638 7392 29644 7404
rect 28399 7364 29644 7392
rect 28399 7361 28411 7364
rect 28353 7355 28411 7361
rect 29638 7352 29644 7364
rect 29696 7352 29702 7404
rect 29730 7352 29736 7404
rect 29788 7352 29794 7404
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 17788 7296 18245 7324
rect 15289 7287 15347 7293
rect 18233 7293 18245 7296
rect 18279 7324 18291 7327
rect 18874 7324 18880 7336
rect 18279 7296 18880 7324
rect 18279 7293 18291 7296
rect 18233 7287 18291 7293
rect 15304 7256 15332 7287
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 19518 7284 19524 7336
rect 19576 7284 19582 7336
rect 23750 7284 23756 7336
rect 23808 7324 23814 7336
rect 24949 7327 25007 7333
rect 24949 7324 24961 7327
rect 23808 7296 24961 7324
rect 23808 7284 23814 7296
rect 24949 7293 24961 7296
rect 24995 7293 25007 7327
rect 24949 7287 25007 7293
rect 27062 7284 27068 7336
rect 27120 7324 27126 7336
rect 28721 7327 28779 7333
rect 28721 7324 28733 7327
rect 27120 7296 28733 7324
rect 27120 7284 27126 7296
rect 28721 7293 28733 7296
rect 28767 7293 28779 7327
rect 28721 7287 28779 7293
rect 28994 7284 29000 7336
rect 29052 7324 29058 7336
rect 30208 7324 30236 7423
rect 32674 7352 32680 7404
rect 32732 7352 32738 7404
rect 29052 7296 30236 7324
rect 31665 7327 31723 7333
rect 29052 7284 29058 7296
rect 31665 7293 31677 7327
rect 31711 7324 31723 7327
rect 31938 7324 31944 7336
rect 31711 7296 31944 7324
rect 31711 7293 31723 7296
rect 31665 7287 31723 7293
rect 31938 7284 31944 7296
rect 31996 7284 32002 7336
rect 33060 7324 33088 7491
rect 34146 7488 34152 7500
rect 34204 7488 34210 7540
rect 35158 7488 35164 7540
rect 35216 7488 35222 7540
rect 36262 7528 36268 7540
rect 35452 7500 36268 7528
rect 33413 7463 33471 7469
rect 33413 7429 33425 7463
rect 33459 7460 33471 7463
rect 35452 7460 35480 7500
rect 36262 7488 36268 7500
rect 36320 7488 36326 7540
rect 37274 7488 37280 7540
rect 37332 7488 37338 7540
rect 37550 7488 37556 7540
rect 37608 7488 37614 7540
rect 33459 7432 35480 7460
rect 33459 7429 33471 7432
rect 33413 7423 33471 7429
rect 34333 7395 34391 7401
rect 34333 7361 34345 7395
rect 34379 7392 34391 7395
rect 34422 7392 34428 7404
rect 34379 7364 34428 7392
rect 34379 7361 34391 7364
rect 34333 7355 34391 7361
rect 34422 7352 34428 7364
rect 34480 7352 34486 7404
rect 34514 7352 34520 7404
rect 34572 7352 34578 7404
rect 36078 7401 36084 7404
rect 36056 7395 36084 7401
rect 36056 7361 36068 7395
rect 36056 7355 36084 7361
rect 36078 7352 36084 7355
rect 36136 7352 36142 7404
rect 36170 7352 36176 7404
rect 36228 7352 36234 7404
rect 37093 7395 37151 7401
rect 37093 7361 37105 7395
rect 37139 7392 37151 7395
rect 37568 7392 37596 7488
rect 37829 7395 37887 7401
rect 37829 7392 37841 7395
rect 37139 7364 37841 7392
rect 37139 7361 37151 7364
rect 37093 7355 37151 7361
rect 37829 7361 37841 7364
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 38102 7352 38108 7404
rect 38160 7392 38166 7404
rect 38197 7395 38255 7401
rect 38197 7392 38209 7395
rect 38160 7364 38209 7392
rect 38160 7352 38166 7364
rect 38197 7361 38209 7364
rect 38243 7361 38255 7395
rect 38197 7355 38255 7361
rect 35897 7327 35955 7333
rect 35897 7324 35909 7327
rect 33060 7296 35909 7324
rect 35897 7293 35909 7296
rect 35943 7293 35955 7327
rect 35897 7287 35955 7293
rect 36909 7327 36967 7333
rect 36909 7293 36921 7327
rect 36955 7324 36967 7327
rect 36998 7324 37004 7336
rect 36955 7296 37004 7324
rect 36955 7293 36967 7296
rect 36909 7287 36967 7293
rect 36998 7284 37004 7296
rect 37056 7284 37062 7336
rect 38286 7284 38292 7336
rect 38344 7324 38350 7336
rect 38381 7327 38439 7333
rect 38381 7324 38393 7327
rect 38344 7296 38393 7324
rect 38344 7284 38350 7296
rect 38381 7293 38393 7296
rect 38427 7293 38439 7327
rect 38381 7287 38439 7293
rect 14200 7228 15332 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 22186 7216 22192 7268
rect 22244 7256 22250 7268
rect 23845 7259 23903 7265
rect 23845 7256 23857 7259
rect 22244 7228 23857 7256
rect 22244 7216 22250 7228
rect 23845 7225 23857 7228
rect 23891 7225 23903 7259
rect 27982 7256 27988 7268
rect 23845 7219 23903 7225
rect 26712 7228 27988 7256
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 5000 7160 5273 7188
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5261 7151 5319 7157
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10410 7188 10416 7200
rect 9732 7160 10416 7188
rect 9732 7148 9738 7160
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11241 7191 11299 7197
rect 11241 7188 11253 7191
rect 11112 7160 11253 7188
rect 11112 7148 11118 7160
rect 11241 7157 11253 7160
rect 11287 7157 11299 7191
rect 11241 7151 11299 7157
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 13078 7188 13084 7200
rect 12023 7160 13084 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 13906 7148 13912 7200
rect 13964 7148 13970 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 18012 7160 18061 7188
rect 18012 7148 18018 7160
rect 18049 7157 18061 7160
rect 18095 7188 18107 7191
rect 18690 7188 18696 7200
rect 18095 7160 18696 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 21821 7191 21879 7197
rect 21821 7157 21833 7191
rect 21867 7188 21879 7191
rect 22094 7188 22100 7200
rect 21867 7160 22100 7188
rect 21867 7157 21879 7160
rect 21821 7151 21879 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 26142 7148 26148 7200
rect 26200 7188 26206 7200
rect 26712 7188 26740 7228
rect 27982 7216 27988 7228
rect 28040 7256 28046 7268
rect 28077 7259 28135 7265
rect 28077 7256 28089 7259
rect 28040 7228 28089 7256
rect 28040 7216 28046 7228
rect 28077 7225 28089 7228
rect 28123 7225 28135 7259
rect 28077 7219 28135 7225
rect 29181 7259 29239 7265
rect 29181 7225 29193 7259
rect 29227 7256 29239 7259
rect 29362 7256 29368 7268
rect 29227 7228 29368 7256
rect 29227 7225 29239 7228
rect 29181 7219 29239 7225
rect 29362 7216 29368 7228
rect 29420 7216 29426 7268
rect 36449 7259 36507 7265
rect 36449 7225 36461 7259
rect 36495 7256 36507 7259
rect 36538 7256 36544 7268
rect 36495 7228 36544 7256
rect 36495 7225 36507 7228
rect 36449 7219 36507 7225
rect 36538 7216 36544 7228
rect 36596 7216 36602 7268
rect 26200 7160 26740 7188
rect 26789 7191 26847 7197
rect 26200 7148 26206 7160
rect 26789 7157 26801 7191
rect 26835 7188 26847 7191
rect 27614 7188 27620 7200
rect 26835 7160 27620 7188
rect 26835 7157 26847 7160
rect 26789 7151 26847 7157
rect 27614 7148 27620 7160
rect 27672 7148 27678 7200
rect 27706 7148 27712 7200
rect 27764 7148 27770 7200
rect 29270 7148 29276 7200
rect 29328 7188 29334 7200
rect 29457 7191 29515 7197
rect 29457 7188 29469 7191
rect 29328 7160 29469 7188
rect 29328 7148 29334 7160
rect 29457 7157 29469 7160
rect 29503 7188 29515 7191
rect 29822 7188 29828 7200
rect 29503 7160 29828 7188
rect 29503 7157 29515 7160
rect 29457 7151 29515 7157
rect 29822 7148 29828 7160
rect 29880 7148 29886 7200
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 33321 7191 33379 7197
rect 33321 7188 33333 7191
rect 32456 7160 33333 7188
rect 32456 7148 32462 7160
rect 33321 7157 33333 7160
rect 33367 7157 33379 7191
rect 33321 7151 33379 7157
rect 35253 7191 35311 7197
rect 35253 7157 35265 7191
rect 35299 7188 35311 7191
rect 35802 7188 35808 7200
rect 35299 7160 35808 7188
rect 35299 7157 35311 7160
rect 35253 7151 35311 7157
rect 35802 7148 35808 7160
rect 35860 7148 35866 7200
rect 38013 7191 38071 7197
rect 38013 7157 38025 7191
rect 38059 7188 38071 7191
rect 38838 7188 38844 7200
rect 38059 7160 38844 7188
rect 38059 7157 38071 7160
rect 38013 7151 38071 7157
rect 38838 7148 38844 7160
rect 38896 7148 38902 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 2225 6987 2283 6993
rect 2225 6953 2237 6987
rect 2271 6984 2283 6987
rect 3694 6984 3700 6996
rect 2271 6956 3700 6984
rect 2271 6953 2283 6956
rect 2225 6947 2283 6953
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 5258 6944 5264 6996
rect 5316 6984 5322 6996
rect 5353 6987 5411 6993
rect 5353 6984 5365 6987
rect 5316 6956 5365 6984
rect 5316 6944 5322 6956
rect 5353 6953 5365 6956
rect 5399 6953 5411 6987
rect 5353 6947 5411 6953
rect 5902 6944 5908 6996
rect 5960 6944 5966 6996
rect 10962 6944 10968 6996
rect 11020 6944 11026 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12158 6984 12164 6996
rect 12115 6956 12164 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 13541 6987 13599 6993
rect 13541 6953 13553 6987
rect 13587 6984 13599 6987
rect 13722 6984 13728 6996
rect 13587 6956 13728 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 13909 6987 13967 6993
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 14458 6984 14464 6996
rect 13955 6956 14464 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 16117 6987 16175 6993
rect 16117 6953 16129 6987
rect 16163 6984 16175 6987
rect 16298 6984 16304 6996
rect 16163 6956 16304 6984
rect 16163 6953 16175 6956
rect 16117 6947 16175 6953
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 16577 6987 16635 6993
rect 16577 6953 16589 6987
rect 16623 6984 16635 6987
rect 16758 6984 16764 6996
rect 16623 6956 16764 6984
rect 16623 6953 16635 6956
rect 16577 6947 16635 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 18138 6944 18144 6996
rect 18196 6944 18202 6996
rect 23290 6984 23296 6996
rect 22756 6956 23296 6984
rect 21928 6888 22232 6916
rect 3605 6851 3663 6857
rect 3605 6817 3617 6851
rect 3651 6817 3663 6851
rect 3605 6811 3663 6817
rect 3338 6783 3396 6789
rect 3338 6749 3350 6783
rect 3384 6780 3396 6783
rect 3384 6776 3464 6780
rect 3510 6776 3516 6792
rect 3384 6752 3516 6776
rect 3384 6749 3396 6752
rect 3338 6743 3396 6749
rect 3436 6748 3516 6752
rect 3510 6740 3516 6748
rect 3568 6740 3574 6792
rect 2682 6672 2688 6724
rect 2740 6712 2746 6724
rect 3050 6712 3056 6724
rect 2740 6684 3056 6712
rect 2740 6672 2746 6684
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3620 6712 3648 6811
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 3936 6820 5549 6848
rect 3936 6808 3942 6820
rect 5537 6817 5549 6820
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8168 6820 8953 6848
rect 8168 6808 8174 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9364 6820 9597 6848
rect 9364 6808 9370 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 11238 6808 11244 6860
rect 11296 6808 11302 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 11940 6820 12173 6848
rect 11940 6808 11946 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 3694 6740 3700 6792
rect 3752 6776 3758 6792
rect 3789 6783 3847 6789
rect 3789 6776 3801 6783
rect 3752 6749 3801 6776
rect 3835 6749 3847 6783
rect 4430 6780 4436 6792
rect 3752 6748 3847 6749
rect 3752 6740 3758 6748
rect 3789 6743 3847 6748
rect 3896 6752 4436 6780
rect 3896 6712 3924 6752
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 5166 6740 5172 6792
rect 5224 6740 5230 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 5644 6712 5672 6743
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5868 6752 5917 6780
rect 5868 6740 5874 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6104 6712 6132 6743
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 9214 6780 9220 6792
rect 8628 6752 9220 6780
rect 8628 6740 8634 6752
rect 9214 6740 9220 6752
rect 9272 6780 9278 6792
rect 10410 6780 10416 6792
rect 9272 6752 10416 6780
rect 9272 6740 9278 6752
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 3620 6684 3924 6712
rect 3988 6684 6132 6712
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3988 6653 4016 6684
rect 3973 6647 4031 6653
rect 3973 6644 3985 6647
rect 3752 6616 3985 6644
rect 3752 6604 3758 6616
rect 3973 6613 3985 6616
rect 4019 6613 4031 6647
rect 3973 6607 4031 6613
rect 4522 6604 4528 6656
rect 4580 6604 4586 6656
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8754 6644 8760 6656
rect 8352 6616 8760 6644
rect 8352 6604 8358 6616
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 11054 6644 11060 6656
rect 10008 6616 11060 6644
rect 10008 6604 10014 6616
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11256 6644 11284 6808
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 12176 6780 12204 6811
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 13872 6820 14657 6848
rect 13872 6808 13878 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 15654 6808 15660 6860
rect 15712 6808 15718 6860
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 17000 6820 17141 6848
rect 17000 6808 17006 6820
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17497 6851 17555 6857
rect 17497 6817 17509 6851
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 18414 6848 18420 6860
rect 17635 6820 18420 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 12894 6780 12900 6792
rect 12176 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 13044 6752 16405 6780
rect 13044 6740 13050 6752
rect 16393 6749 16405 6752
rect 16439 6780 16451 6783
rect 17512 6780 17540 6811
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18690 6808 18696 6860
rect 18748 6808 18754 6860
rect 20714 6848 20720 6860
rect 18800 6820 20720 6848
rect 18800 6780 18828 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 21928 6848 21956 6888
rect 21039 6820 21956 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 22002 6808 22008 6860
rect 22060 6808 22066 6860
rect 22094 6808 22100 6860
rect 22152 6808 22158 6860
rect 22204 6848 22232 6888
rect 22756 6848 22784 6956
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 23474 6944 23480 6996
rect 23532 6944 23538 6996
rect 23750 6944 23756 6996
rect 23808 6944 23814 6996
rect 25038 6944 25044 6996
rect 25096 6944 25102 6996
rect 25314 6944 25320 6996
rect 25372 6944 25378 6996
rect 25700 6956 26556 6984
rect 23566 6916 23572 6928
rect 22848 6888 23572 6916
rect 22848 6857 22876 6888
rect 23566 6876 23572 6888
rect 23624 6876 23630 6928
rect 22204 6820 22784 6848
rect 22833 6851 22891 6857
rect 22833 6817 22845 6851
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 22922 6808 22928 6860
rect 22980 6808 22986 6860
rect 23768 6848 23796 6944
rect 23308 6820 23796 6848
rect 16439 6752 18828 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 19518 6740 19524 6792
rect 19576 6740 19582 6792
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6780 22247 6783
rect 22278 6780 22284 6792
rect 22235 6752 22284 6780
rect 22235 6749 22247 6752
rect 22189 6743 22247 6749
rect 22278 6740 22284 6752
rect 22336 6780 22342 6792
rect 22940 6780 22968 6808
rect 22336 6752 22968 6780
rect 22336 6740 22342 6752
rect 12428 6715 12486 6721
rect 12428 6681 12440 6715
rect 12474 6712 12486 6715
rect 13170 6712 13176 6724
rect 12474 6684 13176 6712
rect 12474 6681 12486 6684
rect 12428 6675 12486 6681
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 15470 6672 15476 6724
rect 15528 6712 15534 6724
rect 17218 6712 17224 6724
rect 15528 6684 17224 6712
rect 15528 6672 15534 6684
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 19536 6712 19564 6740
rect 23308 6712 23336 6820
rect 25038 6808 25044 6860
rect 25096 6848 25102 6860
rect 25222 6848 25228 6860
rect 25096 6820 25228 6848
rect 25096 6808 25102 6820
rect 25222 6808 25228 6820
rect 25280 6848 25286 6860
rect 25700 6857 25728 6956
rect 26528 6916 26556 6956
rect 27154 6944 27160 6996
rect 27212 6944 27218 6996
rect 27982 6944 27988 6996
rect 28040 6984 28046 6996
rect 28813 6987 28871 6993
rect 28813 6984 28825 6987
rect 28040 6956 28825 6984
rect 28040 6944 28046 6956
rect 28813 6953 28825 6956
rect 28859 6953 28871 6987
rect 30282 6984 30288 6996
rect 28813 6947 28871 6953
rect 29012 6956 30288 6984
rect 28077 6919 28135 6925
rect 28077 6916 28089 6919
rect 26528 6888 28089 6916
rect 28077 6885 28089 6888
rect 28123 6885 28135 6919
rect 28077 6879 28135 6885
rect 25685 6851 25743 6857
rect 25685 6848 25697 6851
rect 25280 6820 25697 6848
rect 25280 6808 25286 6820
rect 25685 6817 25697 6820
rect 25731 6817 25743 6851
rect 25685 6811 25743 6817
rect 26602 6808 26608 6860
rect 26660 6848 26666 6860
rect 26973 6851 27031 6857
rect 26973 6848 26985 6851
rect 26660 6820 26985 6848
rect 26660 6808 26666 6820
rect 26973 6817 26985 6820
rect 27019 6817 27031 6851
rect 26973 6811 27031 6817
rect 27706 6808 27712 6860
rect 27764 6808 27770 6860
rect 28092 6848 28120 6879
rect 29012 6848 29040 6956
rect 30282 6944 30288 6956
rect 30340 6944 30346 6996
rect 33962 6944 33968 6996
rect 34020 6984 34026 6996
rect 34701 6987 34759 6993
rect 34701 6984 34713 6987
rect 34020 6956 34713 6984
rect 34020 6944 34026 6956
rect 34701 6953 34713 6956
rect 34747 6953 34759 6987
rect 34701 6947 34759 6953
rect 35897 6987 35955 6993
rect 35897 6953 35909 6987
rect 35943 6984 35955 6987
rect 36078 6984 36084 6996
rect 35943 6956 36084 6984
rect 35943 6953 35955 6956
rect 35897 6947 35955 6953
rect 36078 6944 36084 6956
rect 36136 6944 36142 6996
rect 29181 6919 29239 6925
rect 29181 6885 29193 6919
rect 29227 6885 29239 6919
rect 29181 6879 29239 6885
rect 28092 6820 29040 6848
rect 29196 6848 29224 6879
rect 29454 6876 29460 6928
rect 29512 6916 29518 6928
rect 29512 6888 31754 6916
rect 29512 6876 29518 6888
rect 29914 6848 29920 6860
rect 29196 6820 29920 6848
rect 29914 6808 29920 6820
rect 29972 6808 29978 6860
rect 30742 6808 30748 6860
rect 30800 6808 30806 6860
rect 31110 6808 31116 6860
rect 31168 6848 31174 6860
rect 31297 6851 31355 6857
rect 31297 6848 31309 6851
rect 31168 6820 31309 6848
rect 31168 6808 31174 6820
rect 31297 6817 31309 6820
rect 31343 6817 31355 6851
rect 31297 6811 31355 6817
rect 31386 6808 31392 6860
rect 31444 6808 31450 6860
rect 31726 6848 31754 6888
rect 33704 6888 36032 6916
rect 31938 6848 31944 6860
rect 31726 6820 31944 6848
rect 31938 6808 31944 6820
rect 31996 6808 32002 6860
rect 32309 6851 32367 6857
rect 32309 6817 32321 6851
rect 32355 6848 32367 6851
rect 33704 6848 33732 6888
rect 32355 6820 33732 6848
rect 33781 6851 33839 6857
rect 32355 6817 32367 6820
rect 32309 6811 32367 6817
rect 33781 6817 33793 6851
rect 33827 6848 33839 6851
rect 33827 6820 35388 6848
rect 33827 6817 33839 6820
rect 33781 6811 33839 6817
rect 24029 6783 24087 6789
rect 24029 6780 24041 6783
rect 18064 6684 19564 6712
rect 22572 6684 23336 6712
rect 23400 6752 24041 6780
rect 12250 6644 12256 6656
rect 11256 6616 12256 6644
rect 12250 6604 12256 6616
rect 12308 6644 12314 6656
rect 13722 6644 13728 6656
rect 12308 6616 13728 6644
rect 12308 6604 12314 6616
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 15378 6644 15384 6656
rect 14516 6616 15384 6644
rect 14516 6604 14522 6616
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 17678 6644 17684 6656
rect 16264 6616 17684 6644
rect 16264 6604 16270 6616
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 18064 6653 18092 6684
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 20622 6604 20628 6656
rect 20680 6604 20686 6656
rect 21266 6604 21272 6656
rect 21324 6604 21330 6656
rect 21634 6604 21640 6656
rect 21692 6604 21698 6656
rect 22572 6653 22600 6684
rect 22557 6647 22615 6653
rect 22557 6613 22569 6647
rect 22603 6613 22615 6647
rect 22557 6607 22615 6613
rect 23014 6604 23020 6656
rect 23072 6604 23078 6656
rect 23400 6653 23428 6752
rect 24029 6749 24041 6752
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25961 6783 26019 6789
rect 25961 6780 25973 6783
rect 25188 6752 25973 6780
rect 25188 6740 25194 6752
rect 25961 6749 25973 6752
rect 26007 6780 26019 6783
rect 26142 6780 26148 6792
rect 26007 6752 26148 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26142 6740 26148 6752
rect 26200 6740 26206 6792
rect 28442 6740 28448 6792
rect 28500 6780 28506 6792
rect 28994 6780 29000 6792
rect 28500 6752 29000 6780
rect 28500 6740 28506 6752
rect 28994 6740 29000 6752
rect 29052 6740 29058 6792
rect 29365 6783 29423 6789
rect 29365 6749 29377 6783
rect 29411 6749 29423 6783
rect 29365 6743 29423 6749
rect 23566 6672 23572 6724
rect 23624 6712 23630 6724
rect 24578 6712 24584 6724
rect 23624 6684 24584 6712
rect 23624 6672 23630 6684
rect 24578 6672 24584 6684
rect 24636 6672 24642 6724
rect 25869 6715 25927 6721
rect 25869 6681 25881 6715
rect 25915 6712 25927 6715
rect 26421 6715 26479 6721
rect 26421 6712 26433 6715
rect 25915 6684 26433 6712
rect 25915 6681 25927 6684
rect 25869 6675 25927 6681
rect 26421 6681 26433 6684
rect 26467 6681 26479 6715
rect 29380 6712 29408 6743
rect 30098 6740 30104 6792
rect 30156 6740 30162 6792
rect 30653 6783 30711 6789
rect 30653 6749 30665 6783
rect 30699 6780 30711 6783
rect 31404 6780 31432 6808
rect 30699 6752 31432 6780
rect 31757 6783 31815 6789
rect 30699 6749 30711 6752
rect 30653 6743 30711 6749
rect 31757 6749 31769 6783
rect 31803 6780 31815 6783
rect 32398 6780 32404 6792
rect 31803 6752 32404 6780
rect 31803 6749 31815 6752
rect 31757 6743 31815 6749
rect 32398 6740 32404 6752
rect 32456 6740 32462 6792
rect 32493 6783 32551 6789
rect 32493 6749 32505 6783
rect 32539 6749 32551 6783
rect 32493 6743 32551 6749
rect 30374 6712 30380 6724
rect 29380 6684 30380 6712
rect 26421 6675 26479 6681
rect 30374 6672 30380 6684
rect 30432 6672 30438 6724
rect 32508 6712 32536 6743
rect 33226 6740 33232 6792
rect 33284 6740 33290 6792
rect 33965 6783 34023 6789
rect 33965 6749 33977 6783
rect 34011 6780 34023 6783
rect 34054 6780 34060 6792
rect 34011 6752 34060 6780
rect 34011 6749 34023 6752
rect 33965 6743 34023 6749
rect 34054 6740 34060 6752
rect 34112 6740 34118 6792
rect 34517 6783 34575 6789
rect 34517 6749 34529 6783
rect 34563 6780 34575 6783
rect 34885 6783 34943 6789
rect 34563 6752 34836 6780
rect 34563 6749 34575 6752
rect 34517 6743 34575 6749
rect 34808 6724 34836 6752
rect 34885 6749 34897 6783
rect 34931 6780 34943 6783
rect 35158 6780 35164 6792
rect 34931 6752 35164 6780
rect 34931 6749 34943 6752
rect 34885 6743 34943 6749
rect 35158 6740 35164 6752
rect 35216 6740 35222 6792
rect 33502 6712 33508 6724
rect 32508 6684 33508 6712
rect 33502 6672 33508 6684
rect 33560 6672 33566 6724
rect 34790 6672 34796 6724
rect 34848 6672 34854 6724
rect 35360 6712 35388 6820
rect 35526 6808 35532 6860
rect 35584 6808 35590 6860
rect 35894 6808 35900 6860
rect 35952 6808 35958 6860
rect 36004 6848 36032 6888
rect 36446 6848 36452 6860
rect 36004 6820 36452 6848
rect 36446 6808 36452 6820
rect 36504 6808 36510 6860
rect 37921 6851 37979 6857
rect 37921 6817 37933 6851
rect 37967 6848 37979 6851
rect 38654 6848 38660 6860
rect 37967 6820 38660 6848
rect 37967 6817 37979 6820
rect 37921 6811 37979 6817
rect 38654 6808 38660 6820
rect 38712 6808 38718 6860
rect 38746 6808 38752 6860
rect 38804 6808 38810 6860
rect 35437 6783 35495 6789
rect 35437 6749 35449 6783
rect 35483 6780 35495 6783
rect 35912 6780 35940 6808
rect 35483 6752 35940 6780
rect 36081 6783 36139 6789
rect 35483 6749 35495 6752
rect 35437 6743 35495 6749
rect 36081 6749 36093 6783
rect 36127 6780 36139 6783
rect 36127 6752 37412 6780
rect 36127 6749 36139 6752
rect 36081 6743 36139 6749
rect 36814 6712 36820 6724
rect 34900 6684 35296 6712
rect 35360 6684 36820 6712
rect 23385 6647 23443 6653
rect 23385 6613 23397 6647
rect 23431 6613 23443 6647
rect 23385 6607 23443 6613
rect 23750 6604 23756 6656
rect 23808 6644 23814 6656
rect 25958 6644 25964 6656
rect 23808 6616 25964 6644
rect 23808 6604 23814 6616
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 26326 6604 26332 6656
rect 26384 6604 26390 6656
rect 28994 6604 29000 6656
rect 29052 6644 29058 6656
rect 29733 6647 29791 6653
rect 29733 6644 29745 6647
rect 29052 6616 29745 6644
rect 29052 6604 29058 6616
rect 29733 6613 29745 6616
rect 29779 6613 29791 6647
rect 29733 6607 29791 6613
rect 33042 6604 33048 6656
rect 33100 6604 33106 6656
rect 34054 6604 34060 6656
rect 34112 6644 34118 6656
rect 34238 6644 34244 6656
rect 34112 6616 34244 6644
rect 34112 6604 34118 6616
rect 34238 6604 34244 6616
rect 34296 6644 34302 6656
rect 34900 6644 34928 6684
rect 34296 6616 34928 6644
rect 34296 6604 34302 6616
rect 34974 6604 34980 6656
rect 35032 6604 35038 6656
rect 35268 6644 35296 6684
rect 36814 6672 36820 6684
rect 36872 6672 36878 6724
rect 36998 6672 37004 6724
rect 37056 6672 37062 6724
rect 37274 6672 37280 6724
rect 37332 6721 37338 6724
rect 37332 6675 37344 6721
rect 37332 6672 37338 6675
rect 35345 6647 35403 6653
rect 35345 6644 35357 6647
rect 35268 6616 35357 6644
rect 35345 6613 35357 6616
rect 35391 6644 35403 6647
rect 35986 6644 35992 6656
rect 35391 6616 35992 6644
rect 35391 6613 35403 6616
rect 35345 6607 35403 6613
rect 35986 6604 35992 6616
rect 36044 6604 36050 6656
rect 36173 6647 36231 6653
rect 36173 6613 36185 6647
rect 36219 6644 36231 6647
rect 37016 6644 37044 6672
rect 36219 6616 37044 6644
rect 37384 6644 37412 6752
rect 37458 6740 37464 6792
rect 37516 6780 37522 6792
rect 37553 6783 37611 6789
rect 37553 6780 37565 6783
rect 37516 6752 37565 6780
rect 37516 6740 37522 6752
rect 37553 6749 37565 6752
rect 37599 6749 37611 6783
rect 37553 6743 37611 6749
rect 37642 6740 37648 6792
rect 37700 6780 37706 6792
rect 37737 6783 37795 6789
rect 37737 6780 37749 6783
rect 37700 6752 37749 6780
rect 37700 6740 37706 6752
rect 37737 6749 37749 6752
rect 37783 6749 37795 6783
rect 37737 6743 37795 6749
rect 38289 6783 38347 6789
rect 38289 6749 38301 6783
rect 38335 6780 38347 6783
rect 38764 6780 38792 6808
rect 38335 6752 38792 6780
rect 38335 6749 38347 6752
rect 38289 6743 38347 6749
rect 37642 6644 37648 6656
rect 37384 6616 37648 6644
rect 36219 6613 36231 6616
rect 36173 6607 36231 6613
rect 37642 6604 37648 6616
rect 37700 6604 37706 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2130 6400 2136 6452
rect 2188 6400 2194 6452
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 4522 6400 4528 6452
rect 4580 6400 4586 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5224 6412 5457 6440
rect 5224 6400 5230 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 7064 6412 8861 6440
rect 7064 6400 7070 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 2774 6372 2780 6384
rect 2148 6344 2780 6372
rect 2148 6313 2176 6344
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 3878 6372 3884 6384
rect 2976 6344 3884 6372
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2133 6307 2191 6313
rect 2133 6273 2145 6307
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 1964 6236 1992 6267
rect 2590 6264 2596 6316
rect 2648 6264 2654 6316
rect 2406 6236 2412 6248
rect 1964 6208 2412 6236
rect 2406 6196 2412 6208
rect 2464 6236 2470 6248
rect 2608 6236 2636 6264
rect 2464 6208 2636 6236
rect 2685 6239 2743 6245
rect 2464 6196 2470 6208
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 2976 6236 3004 6344
rect 3878 6332 3884 6344
rect 3936 6332 3942 6384
rect 4280 6375 4338 6381
rect 4280 6341 4292 6375
rect 4326 6372 4338 6375
rect 4540 6372 4568 6400
rect 4326 6344 4568 6372
rect 5552 6372 5580 6400
rect 7285 6375 7343 6381
rect 5552 6344 5948 6372
rect 4326 6341 4338 6344
rect 4280 6335 4338 6341
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3694 6304 3700 6316
rect 3099 6276 3700 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 4488 6276 4568 6304
rect 4488 6264 4494 6276
rect 3234 6236 3240 6248
rect 2731 6208 3240 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 4540 6245 4568 6276
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 4948 6276 5273 6304
rect 4948 6264 4954 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5408 6276 5733 6304
rect 5408 6264 5414 6276
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 5920 6313 5948 6344
rect 7285 6341 7297 6375
rect 7331 6372 7343 6375
rect 7374 6372 7380 6384
rect 7331 6344 7380 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 8570 6332 8576 6384
rect 8628 6332 8634 6384
rect 8864 6372 8892 6403
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9309 6443 9367 6449
rect 9309 6440 9321 6443
rect 9088 6412 9321 6440
rect 9088 6400 9094 6412
rect 9309 6409 9321 6412
rect 9355 6409 9367 6443
rect 9309 6403 9367 6409
rect 10502 6400 10508 6452
rect 10560 6440 10566 6452
rect 11422 6440 11428 6452
rect 10560 6412 11428 6440
rect 10560 6400 10566 6412
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 11572 6412 12357 6440
rect 11572 6400 11578 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12713 6443 12771 6449
rect 12713 6440 12725 6443
rect 12492 6412 12725 6440
rect 12492 6400 12498 6412
rect 12713 6409 12725 6412
rect 12759 6409 12771 6443
rect 12713 6403 12771 6409
rect 13170 6400 13176 6452
rect 13228 6400 13234 6452
rect 14090 6400 14096 6452
rect 14148 6400 14154 6452
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 15378 6440 15384 6452
rect 14875 6412 15384 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 15378 6400 15384 6412
rect 15436 6440 15442 6452
rect 15838 6440 15844 6452
rect 15436 6412 15844 6440
rect 15436 6400 15442 6412
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 22925 6443 22983 6449
rect 20680 6412 22876 6440
rect 20680 6400 20686 6412
rect 12805 6375 12863 6381
rect 8864 6344 12434 6372
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6089 6307 6147 6313
rect 6089 6304 6101 6307
rect 6052 6276 6101 6304
rect 6052 6264 6058 6276
rect 6089 6273 6101 6276
rect 6135 6304 6147 6307
rect 6362 6304 6368 6316
rect 6135 6276 6368 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 9214 6264 9220 6316
rect 9272 6264 9278 6316
rect 4525 6239 4583 6245
rect 4525 6205 4537 6239
rect 4571 6236 4583 6239
rect 5166 6236 5172 6248
rect 4571 6208 5172 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5828 6168 5856 6264
rect 9692 6208 11192 6236
rect 9692 6180 9720 6208
rect 2700 6140 3648 6168
rect 2700 6112 2728 6140
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2682 6100 2688 6112
rect 2363 6072 2688 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 2774 6060 2780 6112
rect 2832 6060 2838 6112
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 3050 6100 3056 6112
rect 2915 6072 3056 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 3620 6100 3648 6140
rect 4632 6140 5856 6168
rect 8205 6171 8263 6177
rect 4632 6100 4660 6140
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 8251 6140 8708 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 8680 6112 8708 6140
rect 9674 6128 9680 6180
rect 9732 6128 9738 6180
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 10192 6140 10241 6168
rect 10192 6128 10198 6140
rect 10229 6137 10241 6140
rect 10275 6168 10287 6171
rect 10870 6168 10876 6180
rect 10275 6140 10876 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 3620 6072 4660 6100
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 4890 6100 4896 6112
rect 4755 6072 4896 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7524 6072 7757 6100
rect 7524 6060 7530 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 8662 6060 8668 6112
rect 8720 6060 8726 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 8812 6072 9781 6100
rect 8812 6060 8818 6072
rect 9769 6069 9781 6072
rect 9815 6100 9827 6103
rect 9950 6100 9956 6112
rect 9815 6072 9956 6100
rect 9815 6069 9827 6072
rect 9769 6063 9827 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 10962 6100 10968 6112
rect 10735 6072 10968 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11164 6100 11192 6208
rect 11238 6196 11244 6248
rect 11296 6196 11302 6248
rect 11514 6196 11520 6248
rect 11572 6196 11578 6248
rect 12158 6196 12164 6248
rect 12216 6196 12222 6248
rect 12406 6168 12434 6344
rect 12805 6341 12817 6375
rect 12851 6372 12863 6375
rect 14108 6372 14136 6400
rect 12851 6344 14136 6372
rect 12851 6341 12863 6344
rect 12805 6335 12863 6341
rect 14642 6332 14648 6384
rect 14700 6372 14706 6384
rect 19242 6372 19248 6384
rect 14700 6344 19248 6372
rect 14700 6332 14706 6344
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 13906 6304 13912 6316
rect 13863 6276 13912 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 15580 6313 15608 6344
rect 19242 6332 19248 6344
rect 19300 6332 19306 6384
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 19306 6276 21312 6304
rect 12986 6196 12992 6248
rect 13044 6196 13050 6248
rect 15838 6196 15844 6248
rect 15896 6196 15902 6248
rect 17586 6196 17592 6248
rect 17644 6196 17650 6248
rect 18230 6196 18236 6248
rect 18288 6196 18294 6248
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18656 6208 18705 6236
rect 18656 6196 18662 6208
rect 18693 6205 18705 6208
rect 18739 6236 18751 6239
rect 19306 6236 19334 6276
rect 18739 6208 19334 6236
rect 18739 6205 18751 6208
rect 18693 6199 18751 6205
rect 20806 6196 20812 6248
rect 20864 6196 20870 6248
rect 21284 6236 21312 6276
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 21416 6276 22293 6304
rect 21416 6264 21422 6276
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 22848 6304 22876 6412
rect 22925 6409 22937 6443
rect 22971 6440 22983 6443
rect 23014 6440 23020 6452
rect 22971 6412 23020 6440
rect 22971 6409 22983 6412
rect 22925 6403 22983 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 23106 6400 23112 6452
rect 23164 6440 23170 6452
rect 24486 6440 24492 6452
rect 23164 6412 24492 6440
rect 23164 6400 23170 6412
rect 24486 6400 24492 6412
rect 24544 6400 24550 6452
rect 25958 6400 25964 6452
rect 26016 6440 26022 6452
rect 26016 6412 27752 6440
rect 26016 6400 26022 6412
rect 23382 6332 23388 6384
rect 23440 6332 23446 6384
rect 24118 6372 24124 6384
rect 23492 6344 24124 6372
rect 23492 6304 23520 6344
rect 24118 6332 24124 6344
rect 24176 6332 24182 6384
rect 24857 6375 24915 6381
rect 24857 6341 24869 6375
rect 24903 6372 24915 6375
rect 27246 6372 27252 6384
rect 24903 6344 27252 6372
rect 24903 6341 24915 6344
rect 24857 6335 24915 6341
rect 27246 6332 27252 6344
rect 27304 6332 27310 6384
rect 22848 6276 23520 6304
rect 23569 6307 23627 6313
rect 22281 6267 22339 6273
rect 23569 6273 23581 6307
rect 23615 6273 23627 6307
rect 23569 6267 23627 6273
rect 23845 6307 23903 6313
rect 23845 6273 23857 6307
rect 23891 6304 23903 6307
rect 23891 6276 24624 6304
rect 23891 6273 23903 6276
rect 23845 6267 23903 6273
rect 21726 6236 21732 6248
rect 21284 6208 21732 6236
rect 21726 6196 21732 6208
rect 21784 6236 21790 6248
rect 22005 6239 22063 6245
rect 22005 6236 22017 6239
rect 21784 6208 22017 6236
rect 21784 6196 21790 6208
rect 22005 6205 22017 6208
rect 22051 6205 22063 6239
rect 23584 6236 23612 6267
rect 24596 6248 24624 6276
rect 24670 6264 24676 6316
rect 24728 6264 24734 6316
rect 25777 6307 25835 6313
rect 25777 6273 25789 6307
rect 25823 6304 25835 6307
rect 26050 6304 26056 6316
rect 25823 6276 26056 6304
rect 25823 6273 25835 6276
rect 25777 6267 25835 6273
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 26237 6307 26295 6313
rect 26237 6273 26249 6307
rect 26283 6304 26295 6307
rect 26326 6304 26332 6316
rect 26283 6276 26332 6304
rect 26283 6273 26295 6276
rect 26237 6267 26295 6273
rect 26326 6264 26332 6276
rect 26384 6304 26390 6316
rect 27154 6304 27160 6316
rect 26384 6276 27160 6304
rect 26384 6264 26390 6276
rect 27154 6264 27160 6276
rect 27212 6264 27218 6316
rect 24394 6236 24400 6248
rect 23584 6208 24400 6236
rect 22005 6199 22063 6205
rect 24394 6196 24400 6208
rect 24452 6196 24458 6248
rect 24489 6239 24547 6245
rect 24489 6205 24501 6239
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 14461 6171 14519 6177
rect 14461 6168 14473 6171
rect 12406 6140 14473 6168
rect 14461 6137 14473 6140
rect 14507 6168 14519 6171
rect 14507 6140 15240 6168
rect 14507 6137 14519 6140
rect 14461 6131 14519 6137
rect 15212 6112 15240 6140
rect 19426 6128 19432 6180
rect 19484 6128 19490 6180
rect 20257 6171 20315 6177
rect 20257 6137 20269 6171
rect 20303 6168 20315 6171
rect 22370 6168 22376 6180
rect 20303 6140 22376 6168
rect 20303 6137 20315 6140
rect 20257 6131 20315 6137
rect 22370 6128 22376 6140
rect 22428 6128 22434 6180
rect 24121 6171 24179 6177
rect 24121 6137 24133 6171
rect 24167 6168 24179 6171
rect 24504 6168 24532 6199
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 25866 6236 25872 6248
rect 24636 6208 25872 6236
rect 24636 6196 24642 6208
rect 25866 6196 25872 6208
rect 25924 6196 25930 6248
rect 25958 6196 25964 6248
rect 26016 6196 26022 6248
rect 26145 6239 26203 6245
rect 26145 6205 26157 6239
rect 26191 6236 26203 6239
rect 26973 6239 27031 6245
rect 26973 6236 26985 6239
rect 26191 6208 26985 6236
rect 26191 6205 26203 6208
rect 26145 6199 26203 6205
rect 26973 6205 26985 6208
rect 27019 6205 27031 6239
rect 26973 6199 27031 6205
rect 27522 6196 27528 6248
rect 27580 6196 27586 6248
rect 27724 6236 27752 6412
rect 27798 6400 27804 6452
rect 27856 6400 27862 6452
rect 28537 6443 28595 6449
rect 28537 6409 28549 6443
rect 28583 6440 28595 6443
rect 28626 6440 28632 6452
rect 28583 6412 28632 6440
rect 28583 6409 28595 6412
rect 28537 6403 28595 6409
rect 28626 6400 28632 6412
rect 28684 6400 28690 6452
rect 30190 6400 30196 6452
rect 30248 6400 30254 6452
rect 32306 6400 32312 6452
rect 32364 6440 32370 6452
rect 32953 6443 33011 6449
rect 32953 6440 32965 6443
rect 32364 6412 32965 6440
rect 32364 6400 32370 6412
rect 32953 6409 32965 6412
rect 32999 6409 33011 6443
rect 32953 6403 33011 6409
rect 33042 6400 33048 6452
rect 33100 6400 33106 6452
rect 34057 6443 34115 6449
rect 34057 6409 34069 6443
rect 34103 6440 34115 6443
rect 34330 6440 34336 6452
rect 34103 6412 34336 6440
rect 34103 6409 34115 6412
rect 34057 6403 34115 6409
rect 34330 6400 34336 6412
rect 34388 6400 34394 6452
rect 34698 6400 34704 6452
rect 34756 6440 34762 6452
rect 34885 6443 34943 6449
rect 34885 6440 34897 6443
rect 34756 6412 34897 6440
rect 34756 6400 34762 6412
rect 34885 6409 34897 6412
rect 34931 6409 34943 6443
rect 34885 6403 34943 6409
rect 34974 6400 34980 6452
rect 35032 6400 35038 6452
rect 35894 6400 35900 6452
rect 35952 6440 35958 6452
rect 36078 6440 36084 6452
rect 35952 6412 36084 6440
rect 35952 6400 35958 6412
rect 36078 6400 36084 6412
rect 36136 6400 36142 6452
rect 37921 6443 37979 6449
rect 37921 6409 37933 6443
rect 37967 6440 37979 6443
rect 38010 6440 38016 6452
rect 37967 6412 38016 6440
rect 37967 6409 37979 6412
rect 37921 6403 37979 6409
rect 38010 6400 38016 6412
rect 38068 6400 38074 6452
rect 27816 6304 27844 6400
rect 29546 6372 29552 6384
rect 28368 6344 29552 6372
rect 28368 6313 28396 6344
rect 29546 6332 29552 6344
rect 29604 6372 29610 6384
rect 30650 6372 30656 6384
rect 29604 6344 30656 6372
rect 29604 6332 29610 6344
rect 30650 6332 30656 6344
rect 30708 6332 30714 6384
rect 33060 6372 33088 6400
rect 33060 6344 34928 6372
rect 27893 6307 27951 6313
rect 27893 6304 27905 6307
rect 27816 6276 27905 6304
rect 27893 6273 27905 6276
rect 27939 6273 27951 6307
rect 28353 6307 28411 6313
rect 28353 6304 28365 6307
rect 27893 6267 27951 6273
rect 28000 6276 28365 6304
rect 28000 6236 28028 6276
rect 28353 6273 28365 6276
rect 28399 6273 28411 6307
rect 28353 6267 28411 6273
rect 28721 6307 28779 6313
rect 28721 6273 28733 6307
rect 28767 6304 28779 6307
rect 29086 6304 29092 6316
rect 28767 6276 29092 6304
rect 28767 6273 28779 6276
rect 28721 6267 28779 6273
rect 29086 6264 29092 6276
rect 29144 6264 29150 6316
rect 29178 6264 29184 6316
rect 29236 6264 29242 6316
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 32306 6304 32312 6316
rect 31803 6276 32312 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 32306 6264 32312 6276
rect 32364 6264 32370 6316
rect 32398 6264 32404 6316
rect 32456 6304 32462 6316
rect 32456 6276 33088 6304
rect 32456 6264 32462 6276
rect 27724 6208 28028 6236
rect 28077 6239 28135 6245
rect 28077 6205 28089 6239
rect 28123 6236 28135 6239
rect 28997 6239 29055 6245
rect 28997 6236 29009 6239
rect 28123 6208 29009 6236
rect 28123 6205 28135 6208
rect 28077 6199 28135 6205
rect 28997 6205 29009 6208
rect 29043 6205 29055 6239
rect 28997 6199 29055 6205
rect 29641 6239 29699 6245
rect 29641 6205 29653 6239
rect 29687 6236 29699 6239
rect 30098 6236 30104 6248
rect 29687 6208 30104 6236
rect 29687 6205 29699 6208
rect 29641 6199 29699 6205
rect 26694 6168 26700 6180
rect 24167 6140 26700 6168
rect 24167 6137 24179 6140
rect 24121 6131 24179 6137
rect 26694 6128 26700 6140
rect 26752 6168 26758 6180
rect 28092 6168 28120 6199
rect 26752 6140 28120 6168
rect 29012 6168 29040 6199
rect 30098 6196 30104 6208
rect 30156 6196 30162 6248
rect 30834 6196 30840 6248
rect 30892 6196 30898 6248
rect 31570 6196 31576 6248
rect 31628 6196 31634 6248
rect 32674 6196 32680 6248
rect 32732 6196 32738 6248
rect 33060 6236 33088 6276
rect 33134 6264 33140 6316
rect 33192 6264 33198 6316
rect 34514 6304 34520 6316
rect 33428 6276 34520 6304
rect 33428 6236 33456 6276
rect 34514 6264 34520 6276
rect 34572 6264 34578 6316
rect 33060 6208 33456 6236
rect 33505 6239 33563 6245
rect 33505 6205 33517 6239
rect 33551 6205 33563 6239
rect 33505 6199 33563 6205
rect 32398 6168 32404 6180
rect 29012 6140 32404 6168
rect 26752 6128 26758 6140
rect 32398 6128 32404 6140
rect 32456 6168 32462 6180
rect 33410 6168 33416 6180
rect 32456 6140 33416 6168
rect 32456 6128 32462 6140
rect 33410 6128 33416 6140
rect 33468 6128 33474 6180
rect 33520 6168 33548 6199
rect 34698 6196 34704 6248
rect 34756 6196 34762 6248
rect 34900 6236 34928 6344
rect 34992 6304 35020 6400
rect 35437 6307 35495 6313
rect 35437 6304 35449 6307
rect 34992 6276 35449 6304
rect 35437 6273 35449 6276
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 35618 6264 35624 6316
rect 35676 6304 35682 6316
rect 36357 6307 36415 6313
rect 36357 6304 36369 6307
rect 35676 6276 36369 6304
rect 35676 6264 35682 6276
rect 36357 6273 36369 6276
rect 36403 6273 36415 6307
rect 36357 6267 36415 6273
rect 36998 6264 37004 6316
rect 37056 6304 37062 6316
rect 37277 6307 37335 6313
rect 37277 6304 37289 6307
rect 37056 6276 37289 6304
rect 37056 6264 37062 6276
rect 37277 6273 37289 6276
rect 37323 6273 37335 6307
rect 37277 6267 37335 6273
rect 38194 6264 38200 6316
rect 38252 6264 38258 6316
rect 34900 6208 35940 6236
rect 35250 6168 35256 6180
rect 33520 6140 35256 6168
rect 35250 6128 35256 6140
rect 35308 6128 35314 6180
rect 35912 6168 35940 6208
rect 35986 6196 35992 6248
rect 36044 6236 36050 6248
rect 36173 6239 36231 6245
rect 36173 6236 36185 6239
rect 36044 6208 36185 6236
rect 36044 6196 36050 6208
rect 36173 6205 36185 6208
rect 36219 6205 36231 6239
rect 36173 6199 36231 6205
rect 36906 6196 36912 6248
rect 36964 6196 36970 6248
rect 38286 6196 38292 6248
rect 38344 6236 38350 6248
rect 38381 6239 38439 6245
rect 38381 6236 38393 6239
rect 38344 6208 38393 6236
rect 38344 6196 38350 6208
rect 38381 6205 38393 6208
rect 38427 6236 38439 6239
rect 38654 6236 38660 6248
rect 38427 6208 38660 6236
rect 38427 6205 38439 6208
rect 38381 6199 38439 6205
rect 38654 6196 38660 6208
rect 38712 6196 38718 6248
rect 35912 6140 38332 6168
rect 13446 6100 13452 6112
rect 11164 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 15102 6060 15108 6112
rect 15160 6060 15166 6112
rect 15194 6060 15200 6112
rect 15252 6060 15258 6112
rect 15286 6060 15292 6112
rect 15344 6060 15350 6112
rect 16485 6103 16543 6109
rect 16485 6069 16497 6103
rect 16531 6100 16543 6103
rect 16666 6100 16672 6112
rect 16531 6072 16672 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 16942 6060 16948 6112
rect 17000 6060 17006 6112
rect 17678 6060 17684 6112
rect 17736 6060 17742 6112
rect 19444 6100 19472 6128
rect 20533 6103 20591 6109
rect 20533 6100 20545 6103
rect 19444 6072 20545 6100
rect 20533 6069 20545 6072
rect 20579 6100 20591 6103
rect 20622 6100 20628 6112
rect 20579 6072 20628 6100
rect 20579 6069 20591 6072
rect 20533 6063 20591 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 21358 6060 21364 6112
rect 21416 6060 21422 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 23201 6103 23259 6109
rect 23201 6100 23213 6103
rect 22060 6072 23213 6100
rect 22060 6060 22066 6072
rect 23201 6069 23213 6072
rect 23247 6100 23259 6103
rect 25038 6100 25044 6112
rect 23247 6072 25044 6100
rect 23247 6069 23259 6072
rect 23201 6063 23259 6069
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 25130 6060 25136 6112
rect 25188 6060 25194 6112
rect 26142 6060 26148 6112
rect 26200 6100 26206 6112
rect 26326 6100 26332 6112
rect 26200 6072 26332 6100
rect 26200 6060 26206 6072
rect 26326 6060 26332 6072
rect 26384 6060 26390 6112
rect 26605 6103 26663 6109
rect 26605 6069 26617 6103
rect 26651 6100 26663 6103
rect 27614 6100 27620 6112
rect 26651 6072 27620 6100
rect 26651 6069 26663 6072
rect 26605 6063 26663 6069
rect 27614 6060 27620 6072
rect 27672 6060 27678 6112
rect 27706 6060 27712 6112
rect 27764 6060 27770 6112
rect 29365 6103 29423 6109
rect 29365 6069 29377 6103
rect 29411 6100 29423 6103
rect 29730 6100 29736 6112
rect 29411 6072 29736 6100
rect 29411 6069 29423 6072
rect 29365 6063 29423 6069
rect 29730 6060 29736 6072
rect 29788 6060 29794 6112
rect 30282 6060 30288 6112
rect 30340 6060 30346 6112
rect 31021 6103 31079 6109
rect 31021 6069 31033 6103
rect 31067 6100 31079 6103
rect 31202 6100 31208 6112
rect 31067 6072 31208 6100
rect 31067 6069 31079 6072
rect 31021 6063 31079 6069
rect 31202 6060 31208 6072
rect 31260 6060 31266 6112
rect 31941 6103 31999 6109
rect 31941 6069 31953 6103
rect 31987 6100 31999 6103
rect 32030 6100 32036 6112
rect 31987 6072 32036 6100
rect 31987 6069 31999 6072
rect 31941 6063 31999 6069
rect 32030 6060 32036 6072
rect 32088 6060 32094 6112
rect 32122 6060 32128 6112
rect 32180 6060 32186 6112
rect 34146 6060 34152 6112
rect 34204 6060 34210 6112
rect 34606 6060 34612 6112
rect 34664 6100 34670 6112
rect 35621 6103 35679 6109
rect 35621 6100 35633 6103
rect 34664 6072 35633 6100
rect 34664 6060 34670 6072
rect 35621 6069 35633 6072
rect 35667 6069 35679 6103
rect 35621 6063 35679 6069
rect 38010 6060 38016 6112
rect 38068 6060 38074 6112
rect 38304 6100 38332 6140
rect 38378 6100 38384 6112
rect 38304 6072 38384 6100
rect 38378 6060 38384 6072
rect 38436 6060 38442 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 4062 5896 4068 5908
rect 3651 5868 4068 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 5350 5896 5356 5908
rect 4172 5868 5356 5896
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2832 5732 3341 5760
rect 2832 5720 2838 5732
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 4062 5760 4068 5772
rect 3375 5732 4068 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 4062 5720 4068 5732
rect 4120 5760 4126 5772
rect 4172 5760 4200 5868
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5626 5856 5632 5908
rect 5684 5856 5690 5908
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 6328 5868 6377 5896
rect 6328 5856 6334 5868
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 12158 5856 12164 5908
rect 12216 5856 12222 5908
rect 12434 5896 12440 5908
rect 12268 5868 12440 5896
rect 10505 5831 10563 5837
rect 10505 5828 10517 5831
rect 10428 5800 10517 5828
rect 4120 5732 4200 5760
rect 4120 5720 4126 5732
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 7190 5760 7196 5772
rect 5224 5732 7196 5760
rect 5224 5720 5230 5732
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 9674 5760 9680 5772
rect 7484 5732 9680 5760
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 2655 5695 2713 5701
rect 2655 5661 2667 5695
rect 2701 5692 2713 5695
rect 3050 5692 3056 5704
rect 2701 5664 3056 5692
rect 2701 5661 2713 5664
rect 2655 5655 2713 5661
rect 2516 5556 2544 5655
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3510 5692 3516 5704
rect 3467 5664 3516 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 4890 5652 4896 5704
rect 4948 5701 4954 5704
rect 4948 5692 4960 5701
rect 4948 5664 4993 5692
rect 4948 5655 4960 5664
rect 4948 5652 4954 5655
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6733 5695 6791 5701
rect 6733 5692 6745 5695
rect 6052 5664 6745 5692
rect 6052 5652 6058 5664
rect 6733 5661 6745 5664
rect 6779 5692 6791 5695
rect 7484 5692 7512 5732
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 10428 5769 10456 5800
rect 10505 5797 10517 5800
rect 10551 5797 10563 5831
rect 10505 5791 10563 5797
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 12066 5828 12072 5840
rect 10928 5800 12072 5828
rect 10928 5788 10934 5800
rect 11164 5769 11192 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 11480 5732 11713 5760
rect 11480 5720 11486 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 11885 5763 11943 5769
rect 11885 5729 11897 5763
rect 11931 5760 11943 5763
rect 12176 5760 12204 5856
rect 11931 5732 12204 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 6779 5664 7512 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 2869 5627 2927 5633
rect 2869 5593 2881 5627
rect 2915 5624 2927 5627
rect 2961 5627 3019 5633
rect 2961 5624 2973 5627
rect 2915 5596 2973 5624
rect 2915 5593 2927 5596
rect 2869 5587 2927 5593
rect 2961 5593 2973 5596
rect 3007 5624 3019 5627
rect 3804 5624 3832 5652
rect 3007 5596 3832 5624
rect 3007 5593 3019 5596
rect 2961 5587 3019 5593
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 3936 5596 6224 5624
rect 3936 5584 3942 5596
rect 3234 5556 3240 5568
rect 2516 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5556 3847 5559
rect 4246 5556 4252 5568
rect 3835 5528 4252 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 5902 5516 5908 5568
rect 5960 5556 5966 5568
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 5960 5528 6009 5556
rect 5960 5516 5966 5528
rect 5997 5525 6009 5528
rect 6043 5525 6055 5559
rect 6196 5556 6224 5596
rect 7282 5584 7288 5636
rect 7340 5624 7346 5636
rect 7852 5624 7880 5655
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 10965 5695 11023 5701
rect 8680 5664 9720 5692
rect 7340 5596 7880 5624
rect 7340 5584 7346 5596
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 8680 5624 8708 5664
rect 8536 5596 8708 5624
rect 8536 5584 8542 5596
rect 9122 5584 9128 5636
rect 9180 5624 9186 5636
rect 9692 5633 9720 5664
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11330 5692 11336 5704
rect 11011 5664 11336 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11330 5652 11336 5664
rect 11388 5692 11394 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11388 5664 11989 5692
rect 11388 5652 11394 5664
rect 11977 5661 11989 5664
rect 12023 5692 12035 5695
rect 12268 5692 12296 5868
rect 12434 5856 12440 5868
rect 12492 5896 12498 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 12492 5868 12633 5896
rect 12492 5856 12498 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 12621 5859 12679 5865
rect 12986 5856 12992 5908
rect 13044 5856 13050 5908
rect 13722 5856 13728 5908
rect 13780 5856 13786 5908
rect 14461 5899 14519 5905
rect 14461 5865 14473 5899
rect 14507 5896 14519 5899
rect 14550 5896 14556 5908
rect 14507 5868 14556 5896
rect 14507 5865 14519 5868
rect 14461 5859 14519 5865
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 15838 5896 15844 5908
rect 15795 5868 15844 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17644 5868 17693 5896
rect 17644 5856 17650 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20864 5868 20913 5896
rect 20864 5856 20870 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 23474 5896 23480 5908
rect 20901 5859 20959 5865
rect 21008 5868 23480 5896
rect 12345 5831 12403 5837
rect 12345 5797 12357 5831
rect 12391 5828 12403 5831
rect 13630 5828 13636 5840
rect 12391 5800 13636 5828
rect 12391 5797 12403 5800
rect 12345 5791 12403 5797
rect 13630 5788 13636 5800
rect 13688 5788 13694 5840
rect 13740 5828 13768 5856
rect 16761 5831 16819 5837
rect 16761 5828 16773 5831
rect 13740 5800 16773 5828
rect 16761 5797 16773 5800
rect 16807 5797 16819 5831
rect 20254 5828 20260 5840
rect 16761 5791 16819 5797
rect 19628 5800 20260 5828
rect 15102 5760 15108 5772
rect 12023 5664 12296 5692
rect 12360 5732 15108 5760
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 9180 5596 9321 5624
rect 9180 5584 9186 5596
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 9677 5627 9735 5633
rect 9677 5593 9689 5627
rect 9723 5624 9735 5627
rect 9723 5596 11744 5624
rect 9723 5593 9735 5596
rect 9677 5587 9735 5593
rect 11716 5568 11744 5596
rect 12066 5584 12072 5636
rect 12124 5624 12130 5636
rect 12360 5624 12388 5732
rect 15102 5720 15108 5732
rect 15160 5760 15166 5772
rect 16301 5763 16359 5769
rect 16301 5760 16313 5763
rect 15160 5732 16313 5760
rect 15160 5720 15166 5732
rect 16301 5729 16313 5732
rect 16347 5729 16359 5763
rect 16776 5760 16804 5791
rect 16850 5760 16856 5772
rect 16776 5732 16856 5760
rect 16301 5723 16359 5729
rect 16850 5720 16856 5732
rect 16908 5760 16914 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16908 5732 17049 5760
rect 16908 5720 16914 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 19628 5704 19656 5800
rect 20254 5788 20260 5800
rect 20312 5828 20318 5840
rect 21008 5828 21036 5868
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 24394 5856 24400 5908
rect 24452 5856 24458 5908
rect 26234 5856 26240 5908
rect 26292 5896 26298 5908
rect 26329 5899 26387 5905
rect 26329 5896 26341 5899
rect 26292 5868 26341 5896
rect 26292 5856 26298 5868
rect 26329 5865 26341 5868
rect 26375 5865 26387 5899
rect 26329 5859 26387 5865
rect 30650 5856 30656 5908
rect 30708 5896 30714 5908
rect 36173 5899 36231 5905
rect 30708 5868 35572 5896
rect 30708 5856 30714 5868
rect 24946 5828 24952 5840
rect 20312 5800 21036 5828
rect 22066 5800 24952 5828
rect 20312 5788 20318 5800
rect 20073 5763 20131 5769
rect 20073 5729 20085 5763
rect 20119 5760 20131 5763
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 20119 5732 21465 5760
rect 20119 5729 20131 5732
rect 20073 5723 20131 5729
rect 21453 5729 21465 5732
rect 21499 5760 21511 5763
rect 22066 5760 22094 5800
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 33226 5788 33232 5840
rect 33284 5828 33290 5840
rect 33284 5800 35480 5828
rect 33284 5788 33290 5800
rect 24121 5763 24179 5769
rect 21499 5732 22094 5760
rect 22756 5732 24072 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 12124 5596 12388 5624
rect 12529 5627 12587 5633
rect 12124 5584 12130 5596
rect 12529 5593 12541 5627
rect 12575 5624 12587 5627
rect 12802 5624 12808 5636
rect 12575 5596 12808 5624
rect 12575 5593 12587 5596
rect 12529 5587 12587 5593
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 13464 5624 13492 5655
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15378 5692 15384 5704
rect 14783 5664 15384 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5692 15715 5695
rect 15746 5692 15752 5704
rect 15703 5664 15752 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 16206 5652 16212 5704
rect 16264 5692 16270 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 16264 5664 17233 5692
rect 16264 5652 16270 5664
rect 17221 5661 17233 5664
rect 17267 5692 17279 5695
rect 17862 5692 17868 5704
rect 17267 5664 17868 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18322 5652 18328 5704
rect 18380 5652 18386 5704
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 20640 5664 21404 5692
rect 14660 5624 14688 5652
rect 20640 5636 20668 5664
rect 13464 5596 14688 5624
rect 14921 5627 14979 5633
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 6196 5528 7665 5556
rect 5997 5519 6055 5525
rect 7653 5525 7665 5528
rect 7699 5525 7711 5559
rect 7653 5519 7711 5525
rect 8754 5516 8760 5568
rect 8812 5516 8818 5568
rect 9766 5516 9772 5568
rect 9824 5516 9830 5568
rect 10870 5516 10876 5568
rect 10928 5516 10934 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 13464 5556 13492 5596
rect 14921 5593 14933 5627
rect 14967 5624 14979 5627
rect 15470 5624 15476 5636
rect 14967 5596 15476 5624
rect 14967 5593 14979 5596
rect 14921 5587 14979 5593
rect 15470 5584 15476 5596
rect 15528 5584 15534 5636
rect 17313 5627 17371 5633
rect 17313 5593 17325 5627
rect 17359 5624 17371 5627
rect 17773 5627 17831 5633
rect 17773 5624 17785 5627
rect 17359 5596 17785 5624
rect 17359 5593 17371 5596
rect 17313 5587 17371 5593
rect 17773 5593 17785 5596
rect 17819 5593 17831 5627
rect 17773 5587 17831 5593
rect 20622 5584 20628 5636
rect 20680 5584 20686 5636
rect 20809 5627 20867 5633
rect 20809 5593 20821 5627
rect 20855 5624 20867 5627
rect 21269 5627 21327 5633
rect 21269 5624 21281 5627
rect 20855 5596 21281 5624
rect 20855 5593 20867 5596
rect 20809 5587 20867 5593
rect 21269 5593 21281 5596
rect 21315 5593 21327 5627
rect 21376 5624 21404 5664
rect 21726 5652 21732 5704
rect 21784 5692 21790 5704
rect 22756 5701 22784 5732
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 21784 5664 21833 5692
rect 21784 5652 21790 5664
rect 21821 5661 21833 5664
rect 21867 5661 21879 5695
rect 22741 5695 22799 5701
rect 22741 5692 22753 5695
rect 21821 5655 21879 5661
rect 22066 5664 22753 5692
rect 22066 5624 22094 5664
rect 22741 5661 22753 5664
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 23290 5652 23296 5704
rect 23348 5692 23354 5704
rect 23385 5695 23443 5701
rect 23385 5692 23397 5695
rect 23348 5664 23397 5692
rect 23348 5652 23354 5664
rect 23385 5661 23397 5664
rect 23431 5661 23443 5695
rect 23385 5655 23443 5661
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5661 23995 5695
rect 24044 5692 24072 5732
rect 24121 5729 24133 5763
rect 24167 5760 24179 5763
rect 26786 5760 26792 5772
rect 24167 5732 26792 5760
rect 24167 5729 24179 5732
rect 24121 5723 24179 5729
rect 26786 5720 26792 5732
rect 26844 5720 26850 5772
rect 34149 5763 34207 5769
rect 31864 5732 34100 5760
rect 24302 5692 24308 5704
rect 24044 5664 24308 5692
rect 23937 5655 23995 5661
rect 21376 5596 22094 5624
rect 22373 5627 22431 5633
rect 21269 5587 21327 5593
rect 22373 5593 22385 5627
rect 22419 5624 22431 5627
rect 23768 5624 23796 5652
rect 22419 5596 23796 5624
rect 22419 5593 22431 5596
rect 22373 5587 22431 5593
rect 11756 5528 13492 5556
rect 11756 5516 11762 5528
rect 13722 5516 13728 5568
rect 13780 5516 13786 5568
rect 15013 5559 15071 5565
rect 15013 5525 15025 5559
rect 15059 5556 15071 5559
rect 15378 5556 15384 5568
rect 15059 5528 15384 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15712 5528 16129 5556
rect 15712 5516 15718 5528
rect 16117 5525 16129 5528
rect 16163 5525 16175 5559
rect 16117 5519 16175 5525
rect 16206 5516 16212 5568
rect 16264 5556 16270 5568
rect 17126 5556 17132 5568
rect 16264 5528 17132 5556
rect 16264 5516 16270 5528
rect 17126 5516 17132 5528
rect 17184 5556 17190 5568
rect 17954 5556 17960 5568
rect 17184 5528 17960 5556
rect 17184 5516 17190 5528
rect 17954 5516 17960 5528
rect 18012 5556 18018 5568
rect 18693 5559 18751 5565
rect 18693 5556 18705 5559
rect 18012 5528 18705 5556
rect 18012 5516 18018 5528
rect 18693 5525 18705 5528
rect 18739 5525 18751 5559
rect 18693 5519 18751 5525
rect 21361 5559 21419 5565
rect 21361 5525 21373 5559
rect 21407 5556 21419 5559
rect 21450 5556 21456 5568
rect 21407 5528 21456 5556
rect 21407 5525 21419 5528
rect 21361 5519 21419 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 23753 5559 23811 5565
rect 23753 5556 23765 5559
rect 23624 5528 23765 5556
rect 23624 5516 23630 5528
rect 23753 5525 23765 5528
rect 23799 5525 23811 5559
rect 23952 5556 23980 5655
rect 24302 5652 24308 5664
rect 24360 5652 24366 5704
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 24213 5627 24271 5633
rect 24213 5593 24225 5627
rect 24259 5624 24271 5627
rect 24486 5624 24492 5636
rect 24259 5596 24492 5624
rect 24259 5593 24271 5596
rect 24213 5587 24271 5593
rect 24486 5584 24492 5596
rect 24544 5584 24550 5636
rect 24596 5624 24624 5655
rect 24762 5652 24768 5704
rect 24820 5652 24826 5704
rect 25314 5652 25320 5704
rect 25372 5652 25378 5704
rect 25685 5695 25743 5701
rect 25685 5661 25697 5695
rect 25731 5692 25743 5695
rect 25774 5692 25780 5704
rect 25731 5664 25780 5692
rect 25731 5661 25743 5664
rect 25685 5655 25743 5661
rect 25774 5652 25780 5664
rect 25832 5652 25838 5704
rect 25866 5652 25872 5704
rect 25924 5652 25930 5704
rect 27062 5652 27068 5704
rect 27120 5692 27126 5704
rect 28445 5695 28503 5701
rect 28445 5692 28457 5695
rect 27120 5664 28457 5692
rect 27120 5652 27126 5664
rect 28445 5661 28457 5664
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28626 5652 28632 5704
rect 28684 5692 28690 5704
rect 29181 5695 29239 5701
rect 29181 5692 29193 5695
rect 28684 5664 29193 5692
rect 28684 5652 28690 5664
rect 29181 5661 29193 5664
rect 29227 5661 29239 5695
rect 29181 5655 29239 5661
rect 30190 5652 30196 5704
rect 30248 5652 30254 5704
rect 31864 5692 31892 5732
rect 30300 5664 31892 5692
rect 25222 5624 25228 5636
rect 24596 5596 25228 5624
rect 25222 5584 25228 5596
rect 25280 5584 25286 5636
rect 25332 5624 25360 5652
rect 27801 5627 27859 5633
rect 27801 5624 27813 5627
rect 25332 5596 27813 5624
rect 27801 5593 27813 5596
rect 27847 5624 27859 5627
rect 29270 5624 29276 5636
rect 27847 5596 29276 5624
rect 27847 5593 27859 5596
rect 27801 5587 27859 5593
rect 29270 5584 29276 5596
rect 29328 5624 29334 5636
rect 30300 5624 30328 5664
rect 31938 5652 31944 5704
rect 31996 5652 32002 5704
rect 32033 5695 32091 5701
rect 32033 5661 32045 5695
rect 32079 5692 32091 5695
rect 32766 5692 32772 5704
rect 32079 5664 32772 5692
rect 32079 5661 32091 5664
rect 32033 5655 32091 5661
rect 32766 5652 32772 5664
rect 32824 5652 32830 5704
rect 34072 5701 34100 5732
rect 34149 5729 34161 5763
rect 34195 5760 34207 5763
rect 34238 5760 34244 5772
rect 34195 5732 34244 5760
rect 34195 5729 34207 5732
rect 34149 5723 34207 5729
rect 34238 5720 34244 5732
rect 34296 5720 34302 5772
rect 34514 5720 34520 5772
rect 34572 5760 34578 5772
rect 34572 5732 35388 5760
rect 34572 5720 34578 5732
rect 34057 5695 34115 5701
rect 34057 5661 34069 5695
rect 34103 5661 34115 5695
rect 34057 5655 34115 5661
rect 34333 5695 34391 5701
rect 34333 5661 34345 5695
rect 34379 5661 34391 5695
rect 34333 5655 34391 5661
rect 29328 5596 30328 5624
rect 31696 5627 31754 5633
rect 29328 5584 29334 5596
rect 31696 5593 31708 5627
rect 31742 5593 31754 5627
rect 31956 5624 31984 5652
rect 31956 5596 32812 5624
rect 31696 5587 31754 5593
rect 25038 5556 25044 5568
rect 23952 5528 25044 5556
rect 23753 5519 23811 5525
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 25406 5516 25412 5568
rect 25464 5516 25470 5568
rect 25498 5516 25504 5568
rect 25556 5516 25562 5568
rect 27890 5516 27896 5568
rect 27948 5516 27954 5568
rect 28534 5516 28540 5568
rect 28592 5556 28598 5568
rect 28629 5559 28687 5565
rect 28629 5556 28641 5559
rect 28592 5528 28641 5556
rect 28592 5516 28598 5528
rect 28629 5525 28641 5528
rect 28675 5525 28687 5559
rect 28629 5519 28687 5525
rect 29546 5516 29552 5568
rect 29604 5556 29610 5568
rect 29641 5559 29699 5565
rect 29641 5556 29653 5559
rect 29604 5528 29653 5556
rect 29604 5516 29610 5528
rect 29641 5525 29653 5528
rect 29687 5525 29699 5559
rect 29641 5519 29699 5525
rect 30558 5516 30564 5568
rect 30616 5516 30622 5568
rect 31726 5556 31754 5587
rect 32122 5556 32128 5568
rect 31726 5528 32128 5556
rect 32122 5516 32128 5528
rect 32180 5516 32186 5568
rect 32214 5516 32220 5568
rect 32272 5516 32278 5568
rect 32784 5565 32812 5596
rect 32858 5584 32864 5636
rect 32916 5624 32922 5636
rect 34348 5624 34376 5655
rect 34790 5652 34796 5704
rect 34848 5692 34854 5704
rect 35253 5695 35311 5701
rect 35253 5692 35265 5695
rect 34848 5664 35265 5692
rect 34848 5652 34854 5664
rect 35253 5661 35265 5664
rect 35299 5661 35311 5695
rect 35253 5655 35311 5661
rect 32916 5596 34376 5624
rect 32916 5584 32922 5596
rect 34422 5584 34428 5636
rect 34480 5624 34486 5636
rect 34701 5627 34759 5633
rect 34701 5624 34713 5627
rect 34480 5596 34713 5624
rect 34480 5584 34486 5596
rect 34701 5593 34713 5596
rect 34747 5593 34759 5627
rect 35360 5624 35388 5732
rect 35452 5692 35480 5800
rect 35544 5769 35572 5868
rect 36173 5865 36185 5899
rect 36219 5896 36231 5899
rect 36906 5896 36912 5908
rect 36219 5868 36912 5896
rect 36219 5865 36231 5868
rect 36173 5859 36231 5865
rect 36906 5856 36912 5868
rect 36964 5856 36970 5908
rect 37090 5828 37096 5840
rect 35728 5800 37096 5828
rect 35529 5763 35587 5769
rect 35529 5729 35541 5763
rect 35575 5729 35587 5763
rect 35529 5723 35587 5729
rect 35728 5692 35756 5800
rect 37090 5788 37096 5800
rect 37148 5788 37154 5840
rect 35802 5720 35808 5772
rect 35860 5720 35866 5772
rect 36170 5720 36176 5772
rect 36228 5760 36234 5772
rect 36357 5763 36415 5769
rect 36357 5760 36369 5763
rect 36228 5732 36369 5760
rect 36228 5720 36234 5732
rect 36357 5729 36369 5732
rect 36403 5760 36415 5763
rect 37734 5760 37740 5772
rect 36403 5732 37740 5760
rect 36403 5729 36415 5732
rect 36357 5723 36415 5729
rect 37734 5720 37740 5732
rect 37792 5720 37798 5772
rect 35452 5664 35756 5692
rect 35820 5692 35848 5720
rect 36541 5695 36599 5701
rect 36541 5692 36553 5695
rect 35820 5664 36553 5692
rect 36541 5661 36553 5664
rect 36587 5661 36599 5695
rect 36541 5655 36599 5661
rect 37277 5695 37335 5701
rect 37277 5661 37289 5695
rect 37323 5692 37335 5695
rect 37366 5692 37372 5704
rect 37323 5664 37372 5692
rect 37323 5661 37335 5664
rect 37277 5655 37335 5661
rect 37366 5652 37372 5664
rect 37424 5652 37430 5704
rect 38286 5652 38292 5704
rect 38344 5652 38350 5704
rect 35526 5624 35532 5636
rect 35360 5596 35532 5624
rect 34701 5587 34759 5593
rect 35526 5584 35532 5596
rect 35584 5584 35590 5636
rect 35713 5627 35771 5633
rect 35713 5593 35725 5627
rect 35759 5624 35771 5627
rect 37550 5624 37556 5636
rect 35759 5596 37556 5624
rect 35759 5593 35771 5596
rect 35713 5587 35771 5593
rect 37550 5584 37556 5596
rect 37608 5584 37614 5636
rect 32769 5559 32827 5565
rect 32769 5525 32781 5559
rect 32815 5556 32827 5559
rect 34238 5556 34244 5568
rect 32815 5528 34244 5556
rect 32815 5525 32827 5528
rect 32769 5519 32827 5525
rect 34238 5516 34244 5528
rect 34296 5516 34302 5568
rect 34514 5516 34520 5568
rect 34572 5516 34578 5568
rect 35802 5516 35808 5568
rect 35860 5556 35866 5568
rect 36078 5556 36084 5568
rect 35860 5528 36084 5556
rect 35860 5516 35866 5528
rect 36078 5516 36084 5528
rect 36136 5516 36142 5568
rect 36630 5516 36636 5568
rect 36688 5516 36694 5568
rect 36998 5516 37004 5568
rect 37056 5516 37062 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3326 5352 3332 5364
rect 2976 5324 3332 5352
rect 2976 5225 3004 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 3510 5312 3516 5364
rect 3568 5312 3574 5364
rect 4062 5312 4068 5364
rect 4120 5312 4126 5364
rect 4246 5312 4252 5364
rect 4304 5312 4310 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 4396 5324 4537 5352
rect 4396 5312 4402 5324
rect 4525 5321 4537 5324
rect 4571 5352 4583 5355
rect 4798 5352 4804 5364
rect 4571 5324 4804 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 5626 5352 5632 5364
rect 5307 5324 5632 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5626 5312 5632 5324
rect 5684 5352 5690 5364
rect 5994 5352 6000 5364
rect 5684 5324 6000 5352
rect 5684 5312 5690 5324
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6328 5324 6868 5352
rect 6328 5312 6334 5324
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3326 5225 3332 5228
rect 3152 5219 3210 5225
rect 3152 5216 3164 5219
rect 3108 5188 3164 5216
rect 3108 5176 3114 5188
rect 3152 5185 3164 5188
rect 3198 5185 3210 5219
rect 3152 5179 3210 5185
rect 3299 5219 3332 5225
rect 3299 5185 3311 5219
rect 3299 5179 3332 5185
rect 3326 5176 3332 5179
rect 3384 5176 3390 5228
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3752 5188 3801 5216
rect 3752 5176 3758 5188
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5216 4031 5219
rect 4080 5216 4108 5312
rect 4019 5188 4108 5216
rect 4264 5216 4292 5312
rect 6840 5284 6868 5324
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 7616 5324 8033 5352
rect 7616 5312 7622 5324
rect 8021 5321 8033 5324
rect 8067 5321 8079 5355
rect 8021 5315 8079 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9214 5352 9220 5364
rect 8987 5324 9220 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 10870 5352 10876 5364
rect 10551 5324 10876 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 11057 5355 11115 5361
rect 11057 5352 11069 5355
rect 11020 5324 11069 5352
rect 11020 5312 11026 5324
rect 11057 5321 11069 5324
rect 11103 5321 11115 5355
rect 11057 5315 11115 5321
rect 12345 5355 12403 5361
rect 12345 5321 12357 5355
rect 12391 5352 12403 5355
rect 12434 5352 12440 5364
rect 12391 5324 12440 5352
rect 12391 5321 12403 5324
rect 12345 5315 12403 5321
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 12805 5355 12863 5361
rect 12805 5321 12817 5355
rect 12851 5352 12863 5355
rect 13170 5352 13176 5364
rect 12851 5324 13176 5352
rect 12851 5321 12863 5324
rect 12805 5315 12863 5321
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 17954 5352 17960 5364
rect 13504 5324 17960 5352
rect 13504 5312 13510 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18230 5352 18236 5364
rect 18095 5324 18236 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 18506 5312 18512 5364
rect 18564 5312 18570 5364
rect 21818 5312 21824 5364
rect 21876 5312 21882 5364
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 25314 5352 25320 5364
rect 25004 5324 25320 5352
rect 25004 5312 25010 5324
rect 25314 5312 25320 5324
rect 25372 5312 25378 5364
rect 26237 5355 26295 5361
rect 26237 5321 26249 5355
rect 26283 5352 26295 5355
rect 26418 5352 26424 5364
rect 26283 5324 26424 5352
rect 26283 5321 26295 5324
rect 26237 5315 26295 5321
rect 26418 5312 26424 5324
rect 26476 5352 26482 5364
rect 27062 5352 27068 5364
rect 26476 5324 27068 5352
rect 26476 5312 26482 5324
rect 27062 5312 27068 5324
rect 27120 5312 27126 5364
rect 27709 5355 27767 5361
rect 27709 5321 27721 5355
rect 27755 5352 27767 5355
rect 28626 5352 28632 5364
rect 27755 5324 28632 5352
rect 27755 5321 27767 5324
rect 27709 5315 27767 5321
rect 28626 5312 28632 5324
rect 28684 5312 28690 5364
rect 29822 5312 29828 5364
rect 29880 5352 29886 5364
rect 30006 5352 30012 5364
rect 29880 5324 30012 5352
rect 29880 5312 29886 5324
rect 30006 5312 30012 5324
rect 30064 5352 30070 5364
rect 30837 5355 30895 5361
rect 30064 5324 30512 5352
rect 30064 5312 30070 5324
rect 5736 5256 6592 5284
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4264 5188 4721 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4798 5176 4804 5228
rect 4856 5176 4862 5228
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5736 5225 5764 5256
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5316 5188 5733 5216
rect 5316 5176 5322 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5902 5176 5908 5228
rect 5960 5176 5966 5228
rect 5994 5176 6000 5228
rect 6052 5176 6058 5228
rect 6564 5225 6592 5256
rect 6840 5256 12112 5284
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6840 5216 6868 5256
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6840 5188 6929 5216
rect 6549 5179 6607 5185
rect 6917 5185 6929 5188
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 2682 5108 2688 5160
rect 2740 5108 2746 5160
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 4816 5148 4844 5176
rect 6380 5148 6408 5179
rect 8662 5176 8668 5228
rect 8720 5176 8726 5228
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9876 5216 10088 5220
rect 10134 5216 10140 5228
rect 8803 5192 10140 5216
rect 8803 5188 9904 5192
rect 10060 5188 10140 5192
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11330 5216 11336 5228
rect 11011 5188 11336 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11790 5176 11796 5228
rect 11848 5176 11854 5228
rect 2915 5120 4752 5148
rect 4816 5120 6408 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 4724 5092 4752 5120
rect 7466 5108 7472 5160
rect 7524 5108 7530 5160
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5148 9275 5151
rect 9861 5151 9919 5157
rect 9263 5120 9812 5148
rect 9263 5117 9275 5120
rect 9217 5111 9275 5117
rect 2777 5083 2835 5089
rect 2777 5049 2789 5083
rect 2823 5080 2835 5083
rect 3970 5080 3976 5092
rect 2823 5052 3976 5080
rect 2823 5049 2835 5052
rect 2777 5043 2835 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 4706 5040 4712 5092
rect 4764 5040 4770 5092
rect 5629 5083 5687 5089
rect 5629 5049 5641 5083
rect 5675 5080 5687 5083
rect 5902 5080 5908 5092
rect 5675 5052 5908 5080
rect 5675 5049 5687 5052
rect 5629 5043 5687 5049
rect 5902 5040 5908 5052
rect 5960 5080 5966 5092
rect 5960 5052 7788 5080
rect 5960 5040 5966 5052
rect 7760 5024 7788 5052
rect 7926 5040 7932 5092
rect 7984 5040 7990 5092
rect 9784 5080 9812 5120
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 9950 5148 9956 5160
rect 9907 5120 9956 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10410 5108 10416 5160
rect 10468 5148 10474 5160
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 10468 5120 11161 5148
rect 10468 5108 10474 5120
rect 11149 5117 11161 5120
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 10597 5083 10655 5089
rect 10597 5080 10609 5083
rect 9784 5052 10609 5080
rect 10597 5049 10609 5052
rect 10643 5049 10655 5083
rect 12084 5080 12112 5256
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 14734 5284 14740 5296
rect 12952 5256 14740 5284
rect 12952 5244 12958 5256
rect 14734 5244 14740 5256
rect 14792 5244 14798 5296
rect 15194 5244 15200 5296
rect 15252 5284 15258 5296
rect 16485 5287 16543 5293
rect 16485 5284 16497 5287
rect 15252 5256 16497 5284
rect 15252 5244 15258 5256
rect 16485 5253 16497 5256
rect 16531 5253 16543 5287
rect 18524 5284 18552 5312
rect 21269 5287 21327 5293
rect 16485 5247 16543 5253
rect 16592 5256 18092 5284
rect 18524 5256 19104 5284
rect 12250 5216 12256 5228
rect 12176 5188 12256 5216
rect 12176 5157 12204 5188
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5185 12495 5219
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 12437 5179 12495 5185
rect 12912 5188 13645 5216
rect 12161 5151 12219 5157
rect 12161 5117 12173 5151
rect 12207 5117 12219 5151
rect 12452 5148 12480 5179
rect 12912 5148 12940 5188
rect 13633 5185 13645 5188
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 14366 5176 14372 5228
rect 14424 5176 14430 5228
rect 16592 5216 16620 5256
rect 14476 5188 16620 5216
rect 16936 5219 16994 5225
rect 12452 5120 12940 5148
rect 12161 5111 12219 5117
rect 13170 5108 13176 5160
rect 13228 5148 13234 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 13228 5120 13461 5148
rect 13228 5108 13234 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 14182 5108 14188 5160
rect 14240 5108 14246 5160
rect 12084 5052 13032 5080
rect 10597 5043 10655 5049
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 3568 4984 3617 5012
rect 3568 4972 3574 4984
rect 3605 4981 3617 4984
rect 3651 4981 3663 5015
rect 3605 4975 3663 4981
rect 3881 5015 3939 5021
rect 3881 4981 3893 5015
rect 3927 5012 3939 5015
rect 4338 5012 4344 5024
rect 3927 4984 4344 5012
rect 3927 4981 3939 4984
rect 3881 4975 3939 4981
rect 4338 4972 4344 4984
rect 4396 4972 4402 5024
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 5350 5012 5356 5024
rect 4479 4984 5356 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 6546 4972 6552 5024
rect 6604 4972 6610 5024
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 10042 5012 10048 5024
rect 9815 4984 10048 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11698 5012 11704 5024
rect 11112 4984 11704 5012
rect 11112 4972 11118 4984
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 11977 5015 12035 5021
rect 11977 4981 11989 5015
rect 12023 5012 12035 5015
rect 12434 5012 12440 5024
rect 12023 4984 12440 5012
rect 12023 4981 12035 4984
rect 11977 4975 12035 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12768 4984 12909 5012
rect 12768 4972 12774 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 13004 5012 13032 5052
rect 14476 5012 14504 5188
rect 16936 5185 16948 5219
rect 16982 5216 16994 5219
rect 17954 5216 17960 5228
rect 16982 5188 17960 5216
rect 16982 5185 16994 5188
rect 16936 5179 16994 5185
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 18064 5216 18092 5256
rect 18693 5219 18751 5225
rect 18064 5188 18644 5216
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 16632 5120 16681 5148
rect 16632 5108 16638 5120
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 17862 5108 17868 5160
rect 17920 5148 17926 5160
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 17920 5120 18521 5148
rect 17920 5108 17926 5120
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 18616 5080 18644 5188
rect 18693 5185 18705 5219
rect 18739 5216 18751 5219
rect 18966 5216 18972 5228
rect 18739 5188 18972 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19076 5225 19104 5256
rect 21269 5253 21281 5287
rect 21315 5284 21327 5287
rect 21450 5284 21456 5296
rect 21315 5256 21456 5284
rect 21315 5253 21327 5256
rect 21269 5247 21327 5253
rect 21450 5244 21456 5256
rect 21508 5284 21514 5296
rect 22278 5284 22284 5296
rect 21508 5256 22284 5284
rect 21508 5244 21514 5256
rect 22278 5244 22284 5256
rect 22336 5244 22342 5296
rect 22373 5287 22431 5293
rect 22373 5253 22385 5287
rect 22419 5284 22431 5287
rect 22462 5284 22468 5296
rect 22419 5256 22468 5284
rect 22419 5253 22431 5256
rect 22373 5247 22431 5253
rect 22462 5244 22468 5256
rect 22520 5284 22526 5296
rect 23106 5284 23112 5296
rect 22520 5256 23112 5284
rect 22520 5244 22526 5256
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 28994 5284 29000 5296
rect 24872 5256 26280 5284
rect 24872 5228 24900 5256
rect 26252 5228 26280 5256
rect 27080 5256 29000 5284
rect 19061 5219 19119 5225
rect 19061 5185 19073 5219
rect 19107 5185 19119 5219
rect 19061 5179 19119 5185
rect 22002 5176 22008 5228
rect 22060 5176 22066 5228
rect 23474 5176 23480 5228
rect 23532 5176 23538 5228
rect 24673 5219 24731 5225
rect 24673 5185 24685 5219
rect 24719 5185 24731 5219
rect 24673 5179 24731 5185
rect 19242 5108 19248 5160
rect 19300 5108 19306 5160
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 20088 5080 20116 5111
rect 20254 5108 20260 5160
rect 20312 5108 20318 5160
rect 20809 5151 20867 5157
rect 20809 5117 20821 5151
rect 20855 5148 20867 5151
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 20855 5120 21373 5148
rect 20855 5117 20867 5120
rect 20809 5111 20867 5117
rect 21361 5117 21373 5120
rect 21407 5117 21419 5151
rect 21361 5111 21419 5117
rect 21545 5151 21603 5157
rect 21545 5117 21557 5151
rect 21591 5148 21603 5151
rect 21634 5148 21640 5160
rect 21591 5120 21640 5148
rect 21591 5117 21603 5120
rect 21545 5111 21603 5117
rect 21634 5108 21640 5120
rect 21692 5108 21698 5160
rect 21726 5108 21732 5160
rect 21784 5148 21790 5160
rect 23109 5151 23167 5157
rect 23109 5148 23121 5151
rect 21784 5120 23121 5148
rect 21784 5108 21790 5120
rect 23109 5117 23121 5120
rect 23155 5148 23167 5151
rect 23842 5148 23848 5160
rect 23155 5120 23848 5148
rect 23155 5117 23167 5120
rect 23109 5111 23167 5117
rect 23842 5108 23848 5120
rect 23900 5108 23906 5160
rect 24118 5108 24124 5160
rect 24176 5148 24182 5160
rect 24213 5151 24271 5157
rect 24213 5148 24225 5151
rect 24176 5120 24225 5148
rect 24176 5108 24182 5120
rect 24213 5117 24225 5120
rect 24259 5148 24271 5151
rect 24486 5148 24492 5160
rect 24259 5120 24492 5148
rect 24259 5117 24271 5120
rect 24213 5111 24271 5117
rect 24486 5108 24492 5120
rect 24544 5108 24550 5160
rect 24688 5148 24716 5179
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 24946 5176 24952 5228
rect 25004 5176 25010 5228
rect 25130 5225 25136 5228
rect 25124 5216 25136 5225
rect 25091 5188 25136 5216
rect 25124 5179 25136 5188
rect 25130 5176 25136 5179
rect 25188 5176 25194 5228
rect 26234 5176 26240 5228
rect 26292 5176 26298 5228
rect 26510 5176 26516 5228
rect 26568 5176 26574 5228
rect 26694 5176 26700 5228
rect 26752 5176 26758 5228
rect 24964 5148 24992 5176
rect 27080 5160 27108 5256
rect 28994 5244 29000 5256
rect 29052 5284 29058 5296
rect 29178 5284 29184 5296
rect 29052 5256 29184 5284
rect 29052 5244 29058 5256
rect 29178 5244 29184 5256
rect 29236 5244 29242 5296
rect 29724 5287 29782 5293
rect 29724 5253 29736 5287
rect 29770 5284 29782 5287
rect 30282 5284 30288 5296
rect 29770 5256 30288 5284
rect 29770 5253 29782 5256
rect 29724 5247 29782 5253
rect 30282 5244 30288 5256
rect 30340 5244 30346 5296
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5216 27399 5219
rect 28537 5219 28595 5225
rect 28537 5216 28549 5219
rect 27387 5188 28549 5216
rect 27387 5185 27399 5188
rect 27341 5179 27399 5185
rect 28537 5185 28549 5188
rect 28583 5185 28595 5219
rect 29454 5216 29460 5228
rect 28537 5179 28595 5185
rect 29012 5188 29460 5216
rect 29012 5160 29040 5188
rect 29454 5176 29460 5188
rect 29512 5176 29518 5228
rect 30484 5216 30512 5324
rect 30837 5321 30849 5355
rect 30883 5352 30895 5355
rect 31570 5352 31576 5364
rect 30883 5324 31576 5352
rect 30883 5321 30895 5324
rect 30837 5315 30895 5321
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 31662 5312 31668 5364
rect 31720 5312 31726 5364
rect 32401 5355 32459 5361
rect 32401 5321 32413 5355
rect 32447 5352 32459 5355
rect 32490 5352 32496 5364
rect 32447 5324 32496 5352
rect 32447 5321 32459 5324
rect 32401 5315 32459 5321
rect 32490 5312 32496 5324
rect 32548 5312 32554 5364
rect 32858 5312 32864 5364
rect 32916 5312 32922 5364
rect 33410 5312 33416 5364
rect 33468 5352 33474 5364
rect 33468 5324 34008 5352
rect 33468 5312 33474 5324
rect 30558 5244 30564 5296
rect 30616 5284 30622 5296
rect 30616 5256 33548 5284
rect 30616 5244 30622 5256
rect 31297 5219 31355 5225
rect 31297 5216 31309 5219
rect 30484 5188 31309 5216
rect 31297 5185 31309 5188
rect 31343 5216 31355 5219
rect 31343 5188 31754 5216
rect 31343 5185 31355 5188
rect 31297 5179 31355 5185
rect 24688 5120 24992 5148
rect 27062 5108 27068 5160
rect 27120 5108 27126 5160
rect 27154 5108 27160 5160
rect 27212 5148 27218 5160
rect 27249 5151 27307 5157
rect 27249 5148 27261 5151
rect 27212 5120 27261 5148
rect 27212 5108 27218 5120
rect 27249 5117 27261 5120
rect 27295 5117 27307 5151
rect 27249 5111 27307 5117
rect 27614 5108 27620 5160
rect 27672 5148 27678 5160
rect 28353 5151 28411 5157
rect 28353 5148 28365 5151
rect 27672 5120 28365 5148
rect 27672 5108 27678 5120
rect 28353 5117 28365 5120
rect 28399 5117 28411 5151
rect 28353 5111 28411 5117
rect 28994 5108 29000 5160
rect 29052 5108 29058 5160
rect 29089 5151 29147 5157
rect 29089 5117 29101 5151
rect 29135 5117 29147 5151
rect 29089 5111 29147 5117
rect 20901 5083 20959 5089
rect 20901 5080 20913 5083
rect 18616 5052 19840 5080
rect 20088 5052 20913 5080
rect 13004 4984 14504 5012
rect 14553 5015 14611 5021
rect 12897 4975 12955 4981
rect 14553 4981 14565 5015
rect 14599 5012 14611 5015
rect 17034 5012 17040 5024
rect 14599 4984 17040 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18325 5015 18383 5021
rect 18325 5012 18337 5015
rect 18104 4984 18337 5012
rect 18104 4972 18110 4984
rect 18325 4981 18337 4984
rect 18371 4981 18383 5015
rect 18325 4975 18383 4981
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 18877 5015 18935 5021
rect 18877 5012 18889 5015
rect 18840 4984 18889 5012
rect 18840 4972 18846 4984
rect 18877 4981 18889 4984
rect 18923 4981 18935 5015
rect 18877 4975 18935 4981
rect 19429 5015 19487 5021
rect 19429 4981 19441 5015
rect 19475 5012 19487 5015
rect 19702 5012 19708 5024
rect 19475 4984 19708 5012
rect 19475 4981 19487 4984
rect 19429 4975 19487 4981
rect 19702 4972 19708 4984
rect 19760 4972 19766 5024
rect 19812 5012 19840 5052
rect 20901 5049 20913 5052
rect 20947 5049 20959 5083
rect 21652 5080 21680 5108
rect 26878 5080 26884 5092
rect 21652 5052 24900 5080
rect 20901 5043 20959 5049
rect 21266 5012 21272 5024
rect 19812 4984 21272 5012
rect 21266 4972 21272 4984
rect 21324 5012 21330 5024
rect 22462 5012 22468 5024
rect 21324 4984 22468 5012
rect 21324 4972 21330 4984
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 24486 4972 24492 5024
rect 24544 4972 24550 5024
rect 24872 5012 24900 5052
rect 25792 5052 26884 5080
rect 25792 5012 25820 5052
rect 26878 5040 26884 5052
rect 26936 5040 26942 5092
rect 27430 5040 27436 5092
rect 27488 5080 27494 5092
rect 29104 5080 29132 5111
rect 30650 5108 30656 5160
rect 30708 5148 30714 5160
rect 31021 5151 31079 5157
rect 31021 5148 31033 5151
rect 30708 5120 31033 5148
rect 30708 5108 30714 5120
rect 31021 5117 31033 5120
rect 31067 5117 31079 5151
rect 31021 5111 31079 5117
rect 31205 5151 31263 5157
rect 31205 5117 31217 5151
rect 31251 5148 31263 5151
rect 31386 5148 31392 5160
rect 31251 5120 31392 5148
rect 31251 5117 31263 5120
rect 31205 5111 31263 5117
rect 31386 5108 31392 5120
rect 31444 5108 31450 5160
rect 31726 5148 31754 5188
rect 31938 5176 31944 5228
rect 31996 5176 32002 5228
rect 32030 5176 32036 5228
rect 32088 5216 32094 5228
rect 32088 5188 32444 5216
rect 32088 5176 32094 5188
rect 31726 5120 32168 5148
rect 27488 5052 29132 5080
rect 27488 5040 27494 5052
rect 30466 5040 30472 5092
rect 30524 5080 30530 5092
rect 31757 5083 31815 5089
rect 31757 5080 31769 5083
rect 30524 5052 31769 5080
rect 30524 5040 30530 5052
rect 31757 5049 31769 5052
rect 31803 5049 31815 5083
rect 32140 5080 32168 5120
rect 32214 5108 32220 5160
rect 32272 5108 32278 5160
rect 32416 5148 32444 5188
rect 32490 5176 32496 5228
rect 32548 5176 32554 5228
rect 32582 5176 32588 5228
rect 32640 5216 32646 5228
rect 33318 5216 33324 5228
rect 32640 5188 33324 5216
rect 32640 5176 32646 5188
rect 33318 5176 33324 5188
rect 33376 5176 33382 5228
rect 33520 5225 33548 5256
rect 33505 5219 33563 5225
rect 33505 5185 33517 5219
rect 33551 5185 33563 5219
rect 33505 5179 33563 5185
rect 33870 5176 33876 5228
rect 33928 5176 33934 5228
rect 33980 5225 34008 5324
rect 34146 5312 34152 5364
rect 34204 5312 34210 5364
rect 37274 5312 37280 5364
rect 37332 5352 37338 5364
rect 37553 5355 37611 5361
rect 37553 5352 37565 5355
rect 37332 5324 37565 5352
rect 37332 5312 37338 5324
rect 37553 5321 37565 5324
rect 37599 5321 37611 5355
rect 37553 5315 37611 5321
rect 34164 5284 34192 5312
rect 34394 5287 34452 5293
rect 34394 5284 34406 5287
rect 34164 5256 34406 5284
rect 34394 5253 34406 5256
rect 34440 5253 34452 5287
rect 34394 5247 34452 5253
rect 36170 5244 36176 5296
rect 36228 5284 36234 5296
rect 36228 5256 38516 5284
rect 36228 5244 36234 5256
rect 33965 5219 34023 5225
rect 33965 5185 33977 5219
rect 34011 5185 34023 5219
rect 33965 5179 34023 5185
rect 34149 5219 34207 5225
rect 34149 5185 34161 5219
rect 34195 5216 34207 5219
rect 34238 5216 34244 5228
rect 34195 5188 34244 5216
rect 34195 5185 34207 5188
rect 34149 5179 34207 5185
rect 34238 5176 34244 5188
rect 34296 5176 34302 5228
rect 37093 5219 37151 5225
rect 37093 5185 37105 5219
rect 37139 5185 37151 5219
rect 37093 5179 37151 5185
rect 36633 5151 36691 5157
rect 32416 5120 34192 5148
rect 32858 5080 32864 5092
rect 32140 5052 32864 5080
rect 31757 5043 31815 5049
rect 32858 5040 32864 5052
rect 32916 5040 32922 5092
rect 24872 4984 25820 5012
rect 26326 4972 26332 5024
rect 26384 4972 26390 5024
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 27801 5015 27859 5021
rect 27801 5012 27813 5015
rect 26752 4984 27813 5012
rect 26752 4972 26758 4984
rect 27801 4981 27813 4984
rect 27847 4981 27859 5015
rect 27801 4975 27859 4981
rect 28902 4972 28908 5024
rect 28960 5012 28966 5024
rect 31846 5012 31852 5024
rect 28960 4984 31852 5012
rect 28960 4972 28966 4984
rect 31846 4972 31852 4984
rect 31904 4972 31910 5024
rect 32214 4972 32220 5024
rect 32272 5012 32278 5024
rect 32582 5012 32588 5024
rect 32272 4984 32588 5012
rect 32272 4972 32278 4984
rect 32582 4972 32588 4984
rect 32640 4972 32646 5024
rect 32950 4972 32956 5024
rect 33008 4972 33014 5024
rect 33042 4972 33048 5024
rect 33100 5012 33106 5024
rect 33689 5015 33747 5021
rect 33689 5012 33701 5015
rect 33100 4984 33701 5012
rect 33100 4972 33106 4984
rect 33689 4981 33701 4984
rect 33735 4981 33747 5015
rect 34164 5012 34192 5120
rect 36633 5117 36645 5151
rect 36679 5117 36691 5151
rect 37108 5148 37136 5179
rect 37274 5176 37280 5228
rect 37332 5176 37338 5228
rect 38010 5176 38016 5228
rect 38068 5176 38074 5228
rect 38488 5225 38516 5256
rect 38473 5219 38531 5225
rect 38473 5185 38485 5219
rect 38519 5185 38531 5219
rect 38473 5179 38531 5185
rect 38028 5148 38056 5176
rect 37108 5120 38056 5148
rect 38105 5151 38163 5157
rect 36633 5111 36691 5117
rect 38105 5117 38117 5151
rect 38151 5117 38163 5151
rect 38105 5111 38163 5117
rect 36446 5080 36452 5092
rect 35452 5052 36452 5080
rect 34882 5012 34888 5024
rect 34164 4984 34888 5012
rect 33689 4975 33747 4981
rect 34882 4972 34888 4984
rect 34940 5012 34946 5024
rect 35452 5012 35480 5052
rect 36446 5040 36452 5052
rect 36504 5040 36510 5092
rect 36648 5080 36676 5111
rect 37734 5080 37740 5092
rect 36648 5052 37740 5080
rect 37734 5040 37740 5052
rect 37792 5040 37798 5092
rect 37918 5040 37924 5092
rect 37976 5080 37982 5092
rect 38120 5080 38148 5111
rect 37976 5052 38148 5080
rect 37976 5040 37982 5052
rect 34940 4984 35480 5012
rect 35529 5015 35587 5021
rect 34940 4972 34946 4984
rect 35529 4981 35541 5015
rect 35575 5012 35587 5015
rect 36078 5012 36084 5024
rect 35575 4984 36084 5012
rect 35575 4981 35587 4984
rect 35529 4975 35587 4981
rect 36078 4972 36084 4984
rect 36136 4972 36142 5024
rect 37461 5015 37519 5021
rect 37461 4981 37473 5015
rect 37507 5012 37519 5015
rect 37826 5012 37832 5024
rect 37507 4984 37832 5012
rect 37507 4981 37519 4984
rect 37461 4975 37519 4981
rect 37826 4972 37832 4984
rect 37884 4972 37890 5024
rect 38286 4972 38292 5024
rect 38344 4972 38350 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 4522 4808 4528 4820
rect 3283 4780 4528 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 4522 4768 4528 4780
rect 4580 4808 4586 4820
rect 6454 4808 6460 4820
rect 4580 4780 6460 4808
rect 4580 4768 4586 4780
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 7374 4808 7380 4820
rect 7116 4780 7380 4808
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 4157 4743 4215 4749
rect 4157 4740 4169 4743
rect 3108 4712 4169 4740
rect 3108 4700 3114 4712
rect 4157 4709 4169 4712
rect 4203 4709 4215 4743
rect 4157 4703 4215 4709
rect 4985 4743 5043 4749
rect 4985 4709 4997 4743
rect 5031 4740 5043 4743
rect 7006 4740 7012 4752
rect 5031 4712 7012 4740
rect 5031 4709 5043 4712
rect 4985 4703 5043 4709
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 3605 4675 3663 4681
rect 3605 4641 3617 4675
rect 3651 4672 3663 4675
rect 4801 4675 4859 4681
rect 3651 4644 4752 4672
rect 3651 4641 3663 4644
rect 3605 4635 3663 4641
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3292 4576 3985 4604
rect 3292 4564 3298 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4356 4536 4384 4567
rect 4522 4564 4528 4616
rect 4580 4604 4586 4616
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 4580 4576 4629 4604
rect 4580 4564 4586 4576
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 4724 4604 4752 4644
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 6181 4675 6239 4681
rect 4847 4644 5488 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5460 4616 5488 4644
rect 6181 4641 6193 4675
rect 6227 4672 6239 4675
rect 6270 4672 6276 4684
rect 6227 4644 6276 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 7116 4681 7144 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 8662 4808 8668 4820
rect 8619 4780 8668 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 10008 4780 11069 4808
rect 10008 4768 10014 4780
rect 11057 4777 11069 4780
rect 11103 4808 11115 4811
rect 12158 4808 12164 4820
rect 11103 4780 12164 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 16485 4811 16543 4817
rect 16485 4808 16497 4811
rect 13504 4780 13768 4808
rect 13504 4768 13510 4780
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11296 4712 11928 4740
rect 11296 4700 11302 4712
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 9674 4672 9680 4684
rect 8352 4644 9680 4672
rect 8352 4632 8358 4644
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 9732 4644 9777 4672
rect 9732 4632 9738 4644
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11514 4672 11520 4684
rect 11204 4644 11520 4672
rect 11204 4632 11210 4644
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 11756 4644 11805 4672
rect 11756 4632 11762 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11900 4672 11928 4712
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11900 4644 12081 4672
rect 11793 4635 11851 4641
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 12158 4632 12164 4684
rect 12216 4681 12222 4684
rect 12216 4675 12244 4681
rect 12232 4641 12244 4675
rect 12216 4635 12244 4641
rect 12216 4632 12222 4635
rect 13078 4632 13084 4684
rect 13136 4672 13142 4684
rect 13740 4681 13768 4780
rect 14476 4780 16497 4808
rect 14476 4681 14504 4780
rect 16485 4777 16497 4780
rect 16531 4808 16543 4811
rect 17494 4808 17500 4820
rect 16531 4780 17500 4808
rect 16531 4777 16543 4780
rect 16485 4771 16543 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 19334 4768 19340 4820
rect 19392 4768 19398 4820
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20993 4811 21051 4817
rect 20993 4808 21005 4811
rect 20312 4780 21005 4808
rect 20312 4768 20318 4780
rect 20993 4777 21005 4780
rect 21039 4808 21051 4811
rect 21039 4780 22232 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 14734 4700 14740 4752
rect 14792 4700 14798 4752
rect 13541 4675 13599 4681
rect 13541 4672 13553 4675
rect 13136 4644 13553 4672
rect 13136 4632 13142 4644
rect 13541 4641 13553 4644
rect 13587 4641 13599 4675
rect 13541 4635 13599 4641
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4641 13783 4675
rect 13725 4635 13783 4641
rect 14461 4675 14519 4681
rect 14461 4641 14473 4675
rect 14507 4641 14519 4675
rect 14752 4672 14780 4700
rect 14752 4644 15148 4672
rect 14461 4635 14519 4641
rect 4724 4576 5212 4604
rect 4617 4567 4675 4573
rect 4706 4536 4712 4548
rect 4356 4508 4712 4536
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 4798 4496 4804 4548
rect 4856 4536 4862 4548
rect 4985 4539 5043 4545
rect 4985 4536 4997 4539
rect 4856 4508 4997 4536
rect 4856 4496 4862 4508
rect 4985 4505 4997 4508
rect 5031 4505 5043 4539
rect 4985 4499 5043 4505
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 2958 4468 2964 4480
rect 2915 4440 2964 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 4890 4468 4896 4480
rect 4479 4440 4896 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5184 4477 5212 4576
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 5316 4576 5365 4604
rect 5316 4564 5322 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5442 4564 5448 4616
rect 5500 4564 5506 4616
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 6822 4604 6828 4616
rect 6411 4576 6828 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 8312 4604 8340 4632
rect 7248 4576 8340 4604
rect 7248 4564 7254 4576
rect 9122 4564 9128 4616
rect 9180 4564 9186 4616
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 5920 4536 5948 4564
rect 5460 4508 5948 4536
rect 5460 4477 5488 4508
rect 6270 4496 6276 4548
rect 6328 4536 6334 4548
rect 6546 4536 6552 4548
rect 6328 4508 6552 4536
rect 6328 4496 6334 4508
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7438 4539 7496 4545
rect 7438 4536 7450 4539
rect 7156 4508 7450 4536
rect 7156 4496 7162 4508
rect 7438 4505 7450 4508
rect 7484 4505 7496 4539
rect 7438 4499 7496 4505
rect 7926 4496 7932 4548
rect 7984 4536 7990 4548
rect 9324 4536 9352 4567
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 9933 4607 9991 4613
rect 9933 4604 9945 4607
rect 9824 4576 9945 4604
rect 9824 4564 9830 4576
rect 9933 4573 9945 4576
rect 9979 4573 9991 4607
rect 9933 4567 9991 4573
rect 11330 4564 11336 4616
rect 11388 4564 11394 4616
rect 12342 4564 12348 4616
rect 12400 4564 12406 4616
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 13035 4576 13461 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4604 14151 4607
rect 14734 4604 14740 4616
rect 14139 4576 14740 4604
rect 14139 4573 14151 4576
rect 14093 4567 14151 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15120 4613 15148 4644
rect 17218 4632 17224 4684
rect 17276 4632 17282 4684
rect 17770 4632 17776 4684
rect 17828 4632 17834 4684
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 18322 4672 18328 4684
rect 18279 4644 18328 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18509 4675 18567 4681
rect 18509 4641 18521 4675
rect 18555 4672 18567 4675
rect 19242 4672 19248 4684
rect 18555 4644 19248 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19352 4644 19625 4672
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4604 15163 4607
rect 16574 4604 16580 4616
rect 15151 4576 16580 4604
rect 15151 4573 15163 4576
rect 15105 4567 15163 4573
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 17402 4613 17408 4616
rect 17359 4607 17408 4613
rect 17359 4573 17371 4607
rect 17405 4573 17408 4607
rect 17359 4567 17408 4573
rect 17402 4564 17408 4567
rect 17460 4564 17466 4616
rect 17494 4564 17500 4616
rect 17552 4564 17558 4616
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 10594 4536 10600 4548
rect 7984 4508 10600 4536
rect 7984 4496 7990 4508
rect 10594 4496 10600 4508
rect 10652 4496 10658 4548
rect 15378 4545 15384 4548
rect 15372 4499 15384 4545
rect 15436 4536 15442 4548
rect 15436 4508 15472 4536
rect 15378 4496 15384 4499
rect 15436 4496 15442 4508
rect 18230 4496 18236 4548
rect 18288 4536 18294 4548
rect 18432 4536 18460 4567
rect 18690 4564 18696 4616
rect 18748 4564 18754 4616
rect 19352 4604 19380 4644
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 21867 4675 21925 4681
rect 21867 4672 21879 4675
rect 19613 4635 19671 4641
rect 20824 4644 21879 4672
rect 18984 4576 19380 4604
rect 19521 4607 19579 4613
rect 18288 4508 18460 4536
rect 18288 4496 18294 4508
rect 18984 4480 19012 4576
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19536 4536 19564 4567
rect 19702 4564 19708 4616
rect 19760 4604 19766 4616
rect 19869 4607 19927 4613
rect 19869 4604 19881 4607
rect 19760 4576 19881 4604
rect 19760 4564 19766 4576
rect 19869 4573 19881 4576
rect 19915 4573 19927 4607
rect 19869 4567 19927 4573
rect 20162 4564 20168 4616
rect 20220 4604 20226 4616
rect 20824 4604 20852 4644
rect 21867 4641 21879 4644
rect 21913 4641 21925 4675
rect 21867 4635 21925 4641
rect 22005 4675 22063 4681
rect 22005 4641 22017 4675
rect 22051 4672 22063 4675
rect 22204 4672 22232 4780
rect 22278 4768 22284 4820
rect 22336 4808 22342 4820
rect 23106 4808 23112 4820
rect 22336 4780 23112 4808
rect 22336 4768 22342 4780
rect 23106 4768 23112 4780
rect 23164 4768 23170 4820
rect 24118 4808 24124 4820
rect 23492 4780 24124 4808
rect 23290 4740 23296 4752
rect 22296 4712 23296 4740
rect 22296 4681 22324 4712
rect 23290 4700 23296 4712
rect 23348 4700 23354 4752
rect 22051 4644 22232 4672
rect 22281 4675 22339 4681
rect 22051 4641 22063 4644
rect 22005 4635 22063 4641
rect 22281 4641 22293 4675
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 22741 4675 22799 4681
rect 22741 4641 22753 4675
rect 22787 4672 22799 4675
rect 23382 4672 23388 4684
rect 22787 4644 23388 4672
rect 22787 4641 22799 4644
rect 22741 4635 22799 4641
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 23492 4681 23520 4780
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24486 4768 24492 4820
rect 24544 4768 24550 4820
rect 24673 4811 24731 4817
rect 24673 4777 24685 4811
rect 24719 4808 24731 4811
rect 24762 4808 24768 4820
rect 24719 4780 24768 4808
rect 24719 4777 24731 4780
rect 24673 4771 24731 4777
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 28442 4808 28448 4820
rect 25332 4780 26648 4808
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 23658 4632 23664 4684
rect 23716 4632 23722 4684
rect 20220 4576 20852 4604
rect 20220 4564 20226 4576
rect 21726 4564 21732 4616
rect 21784 4564 21790 4616
rect 22922 4564 22928 4616
rect 22980 4564 22986 4616
rect 23201 4607 23259 4613
rect 23201 4573 23213 4607
rect 23247 4604 23259 4607
rect 24504 4604 24532 4768
rect 25332 4684 25360 4780
rect 25314 4632 25320 4684
rect 25372 4632 25378 4684
rect 26620 4672 26648 4780
rect 26712 4780 28448 4808
rect 26712 4749 26740 4780
rect 28442 4768 28448 4780
rect 28500 4768 28506 4820
rect 28902 4768 28908 4820
rect 28960 4768 28966 4820
rect 29270 4768 29276 4820
rect 29328 4768 29334 4820
rect 29641 4811 29699 4817
rect 29641 4777 29653 4811
rect 29687 4808 29699 4811
rect 30190 4808 30196 4820
rect 29687 4780 30196 4808
rect 29687 4777 29699 4780
rect 29641 4771 29699 4777
rect 30190 4768 30196 4780
rect 30248 4768 30254 4820
rect 30466 4768 30472 4820
rect 30524 4768 30530 4820
rect 31110 4768 31116 4820
rect 31168 4768 31174 4820
rect 31570 4808 31576 4820
rect 31220 4780 31576 4808
rect 26697 4743 26755 4749
rect 26697 4709 26709 4743
rect 26743 4709 26755 4743
rect 30484 4740 30512 4768
rect 26697 4703 26755 4709
rect 29288 4712 30512 4740
rect 27157 4675 27215 4681
rect 25608 4644 26188 4672
rect 26620 4644 27108 4672
rect 23247 4576 24532 4604
rect 23247 4573 23259 4576
rect 23201 4567 23259 4573
rect 25130 4564 25136 4616
rect 25188 4564 25194 4616
rect 19978 4536 19984 4548
rect 19536 4508 19984 4536
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 22940 4508 23796 4536
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 5215 4440 5457 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 5810 4428 5816 4480
rect 5868 4428 5874 4480
rect 6454 4428 6460 4480
rect 6512 4428 6518 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 10410 4468 10416 4480
rect 9539 4440 10416 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 10560 4440 13093 4468
rect 10560 4428 10566 4440
rect 13081 4437 13093 4440
rect 13127 4437 13139 4471
rect 13081 4431 13139 4437
rect 14277 4471 14335 4477
rect 14277 4437 14289 4471
rect 14323 4468 14335 4471
rect 14918 4468 14924 4480
rect 14323 4440 14924 4468
rect 14323 4437 14335 4440
rect 14277 4431 14335 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15013 4471 15071 4477
rect 15013 4437 15025 4471
rect 15059 4468 15071 4471
rect 16206 4468 16212 4480
rect 15059 4440 16212 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16577 4471 16635 4477
rect 16577 4437 16589 4471
rect 16623 4468 16635 4471
rect 18506 4468 18512 4480
rect 16623 4440 18512 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 18874 4428 18880 4480
rect 18932 4428 18938 4480
rect 18966 4428 18972 4480
rect 19024 4428 19030 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 22940 4468 22968 4508
rect 23768 4477 23796 4508
rect 23842 4496 23848 4548
rect 23900 4536 23906 4548
rect 25608 4536 25636 4644
rect 26160 4613 26188 4644
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4573 26203 4607
rect 26145 4567 26203 4573
rect 26234 4564 26240 4616
rect 26292 4613 26298 4616
rect 26292 4607 26341 4613
rect 26292 4573 26295 4607
rect 26329 4573 26341 4607
rect 26292 4567 26341 4573
rect 26292 4564 26298 4567
rect 26418 4564 26424 4616
rect 26476 4564 26482 4616
rect 27080 4604 27108 4644
rect 27157 4641 27169 4675
rect 27203 4672 27215 4675
rect 27430 4672 27436 4684
rect 27203 4644 27436 4672
rect 27203 4641 27215 4644
rect 27157 4635 27215 4641
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 27522 4632 27528 4684
rect 27580 4632 27586 4684
rect 29288 4681 29316 4712
rect 29273 4675 29331 4681
rect 29273 4641 29285 4675
rect 29319 4641 29331 4675
rect 29273 4635 29331 4641
rect 30006 4632 30012 4684
rect 30064 4672 30070 4684
rect 30101 4675 30159 4681
rect 30101 4672 30113 4675
rect 30064 4644 30113 4672
rect 30064 4632 30070 4644
rect 30101 4641 30113 4644
rect 30147 4641 30159 4675
rect 30101 4635 30159 4641
rect 30190 4632 30196 4684
rect 30248 4632 30254 4684
rect 30558 4632 30564 4684
rect 30616 4672 30622 4684
rect 31128 4681 31156 4768
rect 30653 4675 30711 4681
rect 30653 4672 30665 4675
rect 30616 4644 30665 4672
rect 30616 4632 30622 4644
rect 30653 4641 30665 4644
rect 30699 4641 30711 4675
rect 30653 4635 30711 4641
rect 31113 4675 31171 4681
rect 31113 4641 31125 4675
rect 31159 4641 31171 4675
rect 31220 4672 31248 4780
rect 31570 4768 31576 4780
rect 31628 4768 31634 4820
rect 32214 4768 32220 4820
rect 32272 4768 32278 4820
rect 32309 4811 32367 4817
rect 32309 4777 32321 4811
rect 32355 4808 32367 4811
rect 32490 4808 32496 4820
rect 32355 4780 32496 4808
rect 32355 4777 32367 4780
rect 32309 4771 32367 4777
rect 32490 4768 32496 4780
rect 32548 4768 32554 4820
rect 32674 4768 32680 4820
rect 32732 4768 32738 4820
rect 32950 4808 32956 4820
rect 32784 4780 32956 4808
rect 32232 4740 32260 4768
rect 32048 4712 32260 4740
rect 32401 4743 32459 4749
rect 31527 4675 31585 4681
rect 31527 4672 31539 4675
rect 31220 4644 31432 4672
rect 31113 4635 31171 4641
rect 27341 4607 27399 4613
rect 27080 4576 27292 4604
rect 23900 4508 25636 4536
rect 27264 4536 27292 4576
rect 27341 4573 27353 4607
rect 27387 4604 27399 4607
rect 27540 4604 27568 4632
rect 27387 4576 27568 4604
rect 27387 4573 27399 4576
rect 27341 4567 27399 4573
rect 28534 4564 28540 4616
rect 28592 4613 28598 4616
rect 28592 4604 28604 4613
rect 28813 4607 28871 4613
rect 28592 4576 28637 4604
rect 28592 4567 28604 4576
rect 28813 4573 28825 4607
rect 28859 4604 28871 4607
rect 28994 4604 29000 4616
rect 28859 4576 29000 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 28592 4564 28598 4567
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 29089 4607 29147 4613
rect 29089 4573 29101 4607
rect 29135 4604 29147 4607
rect 29822 4604 29828 4616
rect 29135 4576 29828 4604
rect 29135 4573 29147 4576
rect 29089 4567 29147 4573
rect 29822 4564 29828 4576
rect 29880 4564 29886 4616
rect 30208 4604 30236 4632
rect 29932 4576 30236 4604
rect 27264 4508 29316 4536
rect 23900 4496 23906 4508
rect 21131 4440 22968 4468
rect 23753 4471 23811 4477
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 23753 4437 23765 4471
rect 23799 4437 23811 4471
rect 23753 4431 23811 4437
rect 24118 4428 24124 4480
rect 24176 4428 24182 4480
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 25041 4471 25099 4477
rect 25041 4468 25053 4471
rect 24820 4440 25053 4468
rect 24820 4428 24826 4440
rect 25041 4437 25053 4440
rect 25087 4437 25099 4471
rect 25041 4431 25099 4437
rect 25501 4471 25559 4477
rect 25501 4437 25513 4471
rect 25547 4468 25559 4471
rect 27338 4468 27344 4480
rect 25547 4440 27344 4468
rect 25547 4437 25559 4440
rect 25501 4431 25559 4437
rect 27338 4428 27344 4440
rect 27396 4428 27402 4480
rect 27430 4428 27436 4480
rect 27488 4428 27494 4480
rect 29288 4468 29316 4508
rect 29362 4496 29368 4548
rect 29420 4496 29426 4548
rect 29454 4468 29460 4480
rect 29288 4440 29460 4468
rect 29454 4428 29460 4440
rect 29512 4468 29518 4480
rect 29932 4468 29960 4576
rect 30466 4564 30472 4616
rect 30524 4564 30530 4616
rect 31404 4613 31432 4644
rect 31521 4641 31539 4672
rect 31573 4641 31585 4675
rect 32048 4672 32076 4712
rect 32401 4709 32413 4743
rect 32447 4740 32459 4743
rect 32692 4740 32720 4768
rect 32447 4712 32720 4740
rect 32447 4709 32459 4712
rect 32401 4703 32459 4709
rect 31521 4635 31585 4641
rect 31711 4644 32076 4672
rect 31521 4616 31549 4635
rect 31389 4607 31447 4613
rect 31389 4573 31401 4607
rect 31435 4573 31447 4607
rect 31389 4567 31447 4573
rect 31478 4564 31484 4616
rect 31536 4576 31549 4616
rect 31711 4613 31739 4644
rect 32784 4613 32812 4780
rect 32950 4768 32956 4780
rect 33008 4768 33014 4820
rect 33686 4768 33692 4820
rect 33744 4768 33750 4820
rect 34517 4811 34575 4817
rect 34517 4777 34529 4811
rect 34563 4808 34575 4811
rect 34790 4808 34796 4820
rect 34563 4780 34796 4808
rect 34563 4777 34575 4780
rect 34517 4771 34575 4777
rect 34790 4768 34796 4780
rect 34848 4768 34854 4820
rect 35161 4811 35219 4817
rect 35161 4777 35173 4811
rect 35207 4808 35219 4811
rect 36630 4808 36636 4820
rect 35207 4780 36636 4808
rect 35207 4777 35219 4780
rect 35161 4771 35219 4777
rect 36630 4768 36636 4780
rect 36688 4768 36694 4820
rect 37458 4808 37464 4820
rect 37108 4780 37464 4808
rect 36357 4743 36415 4749
rect 33336 4712 35296 4740
rect 33336 4684 33364 4712
rect 32858 4632 32864 4684
rect 32916 4632 32922 4684
rect 33045 4675 33103 4681
rect 33045 4641 33057 4675
rect 33091 4672 33103 4675
rect 33226 4672 33232 4684
rect 33091 4644 33232 4672
rect 33091 4641 33103 4644
rect 33045 4635 33103 4641
rect 33226 4632 33232 4644
rect 33284 4632 33290 4684
rect 33318 4632 33324 4684
rect 33376 4632 33382 4684
rect 33502 4632 33508 4684
rect 33560 4632 33566 4684
rect 33594 4632 33600 4684
rect 33652 4632 33658 4684
rect 33870 4632 33876 4684
rect 33928 4632 33934 4684
rect 34054 4632 34060 4684
rect 34112 4632 34118 4684
rect 34330 4632 34336 4684
rect 34388 4672 34394 4684
rect 35069 4675 35127 4681
rect 35069 4672 35081 4675
rect 34388 4644 35081 4672
rect 34388 4632 34394 4644
rect 35069 4641 35081 4644
rect 35115 4672 35127 4675
rect 35158 4672 35164 4684
rect 35115 4644 35164 4672
rect 35115 4641 35127 4644
rect 35069 4635 35127 4641
rect 35158 4632 35164 4644
rect 35216 4632 35222 4684
rect 35268 4672 35296 4712
rect 36357 4709 36369 4743
rect 36403 4740 36415 4743
rect 36446 4740 36452 4752
rect 36403 4712 36452 4740
rect 36403 4709 36415 4712
rect 36357 4703 36415 4709
rect 36446 4700 36452 4712
rect 36504 4700 36510 4752
rect 35986 4681 35992 4684
rect 35805 4675 35863 4681
rect 35805 4672 35817 4675
rect 35268 4644 35817 4672
rect 35805 4641 35817 4644
rect 35851 4641 35863 4675
rect 35805 4635 35863 4641
rect 35964 4675 35992 4681
rect 35964 4641 35976 4675
rect 35964 4635 35992 4641
rect 35986 4632 35992 4635
rect 36044 4632 36050 4684
rect 37108 4681 37136 4780
rect 37458 4768 37464 4780
rect 37516 4768 37522 4820
rect 37093 4675 37151 4681
rect 37093 4641 37105 4675
rect 37139 4641 37151 4675
rect 37093 4635 37151 4641
rect 31665 4607 31739 4613
rect 31536 4564 31542 4576
rect 31665 4573 31677 4607
rect 31711 4576 31739 4607
rect 32769 4607 32827 4613
rect 31711 4573 31723 4576
rect 31665 4567 31723 4573
rect 32769 4573 32781 4607
rect 32815 4573 32827 4607
rect 32769 4567 32827 4573
rect 33410 4564 33416 4616
rect 33468 4564 33474 4616
rect 30024 4508 30696 4536
rect 30024 4477 30052 4508
rect 29512 4440 29960 4468
rect 30009 4471 30067 4477
rect 29512 4428 29518 4440
rect 30009 4437 30021 4471
rect 30055 4437 30067 4471
rect 30668 4468 30696 4508
rect 32582 4496 32588 4548
rect 32640 4536 32646 4548
rect 33520 4536 33548 4632
rect 33689 4607 33747 4613
rect 33689 4573 33701 4607
rect 33735 4604 33747 4607
rect 33962 4604 33968 4616
rect 33735 4576 33968 4604
rect 33735 4573 33747 4576
rect 33689 4567 33747 4573
rect 33962 4564 33968 4576
rect 34020 4564 34026 4616
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 34606 4604 34612 4616
rect 34195 4576 34612 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 34606 4564 34612 4576
rect 34664 4564 34670 4616
rect 34882 4564 34888 4616
rect 34940 4564 34946 4616
rect 36078 4564 36084 4616
rect 36136 4564 36142 4616
rect 36817 4607 36875 4613
rect 36817 4573 36829 4607
rect 36863 4573 36875 4607
rect 36817 4567 36875 4573
rect 37001 4607 37059 4613
rect 37001 4573 37013 4607
rect 37047 4604 37059 4607
rect 37182 4604 37188 4616
rect 37047 4576 37188 4604
rect 37047 4573 37059 4576
rect 37001 4567 37059 4573
rect 32640 4508 33272 4536
rect 33520 4508 35388 4536
rect 32640 4496 32646 4508
rect 32122 4468 32128 4480
rect 30668 4440 32128 4468
rect 30009 4431 30067 4437
rect 32122 4428 32128 4440
rect 32180 4428 32186 4480
rect 33244 4477 33272 4508
rect 33229 4471 33287 4477
rect 33229 4437 33241 4471
rect 33275 4437 33287 4471
rect 33229 4431 33287 4437
rect 34330 4428 34336 4480
rect 34388 4468 34394 4480
rect 34701 4471 34759 4477
rect 34701 4468 34713 4471
rect 34388 4440 34713 4468
rect 34388 4428 34394 4440
rect 34701 4437 34713 4440
rect 34747 4437 34759 4471
rect 35360 4468 35388 4508
rect 36832 4468 36860 4567
rect 37182 4564 37188 4576
rect 37240 4564 37246 4616
rect 36906 4496 36912 4548
rect 36964 4536 36970 4548
rect 37338 4539 37396 4545
rect 37338 4536 37350 4539
rect 36964 4508 37350 4536
rect 36964 4496 36970 4508
rect 37338 4505 37350 4508
rect 37384 4505 37396 4539
rect 37338 4499 37396 4505
rect 38473 4471 38531 4477
rect 38473 4468 38485 4471
rect 35360 4440 38485 4468
rect 34701 4431 34759 4437
rect 38473 4437 38485 4440
rect 38519 4437 38531 4471
rect 38473 4431 38531 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3786 4264 3792 4276
rect 3528 4236 3792 4264
rect 2498 4156 2504 4208
rect 2556 4196 2562 4208
rect 3528 4205 3556 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4798 4264 4804 4276
rect 4264 4236 4804 4264
rect 3053 4199 3111 4205
rect 3053 4196 3065 4199
rect 2556 4168 3065 4196
rect 2556 4156 2562 4168
rect 3053 4165 3065 4168
rect 3099 4165 3111 4199
rect 3053 4159 3111 4165
rect 3513 4199 3571 4205
rect 3513 4165 3525 4199
rect 3559 4165 3571 4199
rect 3513 4159 3571 4165
rect 2682 4088 2688 4140
rect 2740 4088 2746 4140
rect 2866 4088 2872 4140
rect 2924 4088 2930 4140
rect 3326 4088 3332 4140
rect 3384 4128 3390 4140
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3384 4100 3433 4128
rect 3384 4088 3390 4100
rect 3421 4097 3433 4100
rect 3467 4128 3479 4131
rect 3694 4128 3700 4140
rect 3467 4100 3700 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2884 4060 2912 4088
rect 4264 4069 4292 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6565 4267 6623 4273
rect 6565 4264 6577 4267
rect 5868 4236 6577 4264
rect 5868 4224 5874 4236
rect 6565 4233 6577 4236
rect 6611 4233 6623 4267
rect 6565 4227 6623 4233
rect 6822 4224 6828 4276
rect 6880 4224 6886 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 11054 4264 11060 4276
rect 7524 4236 11060 4264
rect 7524 4224 7530 4236
rect 6270 4196 6276 4208
rect 4724 4168 4936 4196
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4724 4128 4752 4168
rect 4571 4100 4752 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 4908 4128 4936 4168
rect 5184 4168 6276 4196
rect 4982 4128 4988 4140
rect 4908 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5184 4137 5212 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 6362 4156 6368 4208
rect 6420 4156 6426 4208
rect 7742 4156 7748 4208
rect 7800 4196 7806 4208
rect 9232 4205 9260 4236
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11330 4224 11336 4276
rect 11388 4264 11394 4276
rect 11609 4267 11667 4273
rect 11609 4264 11621 4267
rect 11388 4236 11621 4264
rect 11388 4224 11394 4236
rect 11609 4233 11621 4236
rect 11655 4264 11667 4267
rect 14182 4264 14188 4276
rect 11655 4236 14188 4264
rect 11655 4233 11667 4236
rect 11609 4227 11667 4233
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 16758 4264 16764 4276
rect 14976 4236 16764 4264
rect 14976 4224 14982 4236
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 18049 4267 18107 4273
rect 18049 4233 18061 4267
rect 18095 4264 18107 4267
rect 18322 4264 18328 4276
rect 18095 4236 18328 4264
rect 18095 4233 18107 4236
rect 18049 4227 18107 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 18506 4224 18512 4276
rect 18564 4224 18570 4276
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 18877 4267 18935 4273
rect 18877 4264 18889 4267
rect 18748 4236 18889 4264
rect 18748 4224 18754 4236
rect 18877 4233 18889 4236
rect 18923 4233 18935 4267
rect 19521 4267 19579 4273
rect 19521 4264 19533 4267
rect 18877 4227 18935 4233
rect 19444 4236 19533 4264
rect 9217 4199 9275 4205
rect 7800 4168 8524 4196
rect 7800 4156 7806 4168
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4128 6147 4131
rect 6454 4128 6460 4140
rect 6135 4100 6460 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7938 4131 7996 4137
rect 7938 4128 7950 4131
rect 7616 4100 7950 4128
rect 7616 4088 7622 4100
rect 7938 4097 7950 4100
rect 7984 4097 7996 4131
rect 7938 4091 7996 4097
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8294 4128 8300 4140
rect 8251 4100 8300 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8496 4137 8524 4168
rect 9217 4165 9229 4199
rect 9263 4165 9275 4199
rect 9490 4196 9496 4208
rect 9217 4159 9275 4165
rect 9324 4168 9496 4196
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 9324 4128 9352 4168
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 9640 4168 9904 4196
rect 9640 4156 9646 4168
rect 8527 4100 9352 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 9398 4088 9404 4140
rect 9456 4088 9462 4140
rect 9670 4131 9728 4137
rect 9670 4097 9682 4131
rect 9716 4128 9728 4131
rect 9766 4128 9772 4140
rect 9716 4100 9772 4128
rect 9716 4097 9728 4100
rect 9670 4091 9728 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9876 4132 9904 4168
rect 10042 4156 10048 4208
rect 10100 4196 10106 4208
rect 10198 4199 10256 4205
rect 10198 4196 10210 4199
rect 10100 4168 10210 4196
rect 10100 4156 10106 4168
rect 10198 4165 10210 4168
rect 10244 4165 10256 4199
rect 10198 4159 10256 4165
rect 12526 4156 12532 4208
rect 12584 4156 12590 4208
rect 12710 4156 12716 4208
rect 12768 4205 12774 4208
rect 12768 4196 12780 4205
rect 12768 4168 12813 4196
rect 12768 4159 12780 4168
rect 12768 4156 12774 4159
rect 14734 4156 14740 4208
rect 14792 4196 14798 4208
rect 15378 4196 15384 4208
rect 14792 4168 15384 4196
rect 14792 4156 14798 4168
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 18966 4196 18972 4208
rect 17880 4168 18972 4196
rect 9953 4132 10011 4137
rect 9876 4131 10011 4132
rect 9876 4104 9965 4131
rect 9953 4097 9965 4104
rect 9999 4097 10011 4131
rect 12158 4128 12164 4140
rect 9953 4091 10011 4097
rect 10060 4100 12164 4128
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 1820 4032 4261 4060
rect 1820 4020 1826 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 5350 4060 5356 4072
rect 4939 4032 5356 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 5184 4004 5212 4032
rect 5350 4020 5356 4032
rect 5408 4060 5414 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5408 4032 5549 4060
rect 5408 4020 5414 4032
rect 5537 4029 5549 4032
rect 5583 4060 5595 4063
rect 6178 4060 6184 4072
rect 5583 4032 6184 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 7098 4020 7104 4072
rect 7156 4020 7162 4072
rect 9490 4020 9496 4072
rect 9548 4020 9554 4072
rect 10060 4060 10088 4100
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12544 4128 12572 4156
rect 12894 4128 12900 4140
rect 12544 4100 12900 4128
rect 12894 4088 12900 4100
rect 12952 4128 12958 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12952 4100 13001 4128
rect 12952 4088 12958 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13630 4088 13636 4140
rect 13688 4088 13694 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14424 4100 14657 4128
rect 14424 4088 14430 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 15654 4088 15660 4140
rect 15712 4088 15718 4140
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16206 4088 16212 4140
rect 16264 4088 16270 4140
rect 16574 4088 16580 4140
rect 16632 4128 16638 4140
rect 16942 4137 16948 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16632 4100 16681 4128
rect 16632 4088 16638 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16936 4128 16948 4137
rect 16903 4100 16948 4128
rect 16669 4091 16727 4097
rect 16936 4091 16948 4100
rect 16942 4088 16948 4091
rect 17000 4088 17006 4140
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 17880 4128 17908 4168
rect 18966 4156 18972 4168
rect 19024 4156 19030 4208
rect 19444 4205 19472 4236
rect 19521 4233 19533 4236
rect 19567 4233 19579 4267
rect 19521 4227 19579 4233
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 20257 4267 20315 4273
rect 20257 4264 20269 4267
rect 20220 4236 20269 4264
rect 20220 4224 20226 4236
rect 20257 4233 20269 4236
rect 20303 4233 20315 4267
rect 20257 4227 20315 4233
rect 23106 4224 23112 4276
rect 23164 4264 23170 4276
rect 23661 4267 23719 4273
rect 23661 4264 23673 4267
rect 23164 4236 23673 4264
rect 23164 4224 23170 4236
rect 23661 4233 23673 4236
rect 23707 4233 23719 4267
rect 23661 4227 23719 4233
rect 24118 4224 24124 4276
rect 24176 4224 24182 4276
rect 24854 4224 24860 4276
rect 24912 4224 24918 4276
rect 26510 4224 26516 4276
rect 26568 4264 26574 4276
rect 26973 4267 27031 4273
rect 26973 4264 26985 4267
rect 26568 4236 26985 4264
rect 26568 4224 26574 4236
rect 26973 4233 26985 4236
rect 27019 4233 27031 4267
rect 26973 4227 27031 4233
rect 27338 4224 27344 4276
rect 27396 4224 27402 4276
rect 29362 4224 29368 4276
rect 29420 4264 29426 4276
rect 32030 4264 32036 4276
rect 29420 4236 32036 4264
rect 29420 4224 29426 4236
rect 32030 4224 32036 4236
rect 32088 4224 32094 4276
rect 32122 4224 32128 4276
rect 32180 4224 32186 4276
rect 32858 4224 32864 4276
rect 32916 4264 32922 4276
rect 33321 4267 33379 4273
rect 33321 4264 33333 4267
rect 32916 4236 33333 4264
rect 32916 4224 32922 4236
rect 33321 4233 33333 4236
rect 33367 4233 33379 4267
rect 33321 4227 33379 4233
rect 33410 4224 33416 4276
rect 33468 4264 33474 4276
rect 33597 4267 33655 4273
rect 33597 4264 33609 4267
rect 33468 4236 33609 4264
rect 33468 4224 33474 4236
rect 33597 4233 33609 4236
rect 33643 4233 33655 4267
rect 35894 4264 35900 4276
rect 33597 4227 33655 4233
rect 33796 4236 35900 4264
rect 19429 4199 19487 4205
rect 19429 4165 19441 4199
rect 19475 4165 19487 4199
rect 23753 4199 23811 4205
rect 19429 4159 19487 4165
rect 19628 4168 20668 4196
rect 17368 4100 17908 4128
rect 17368 4088 17374 4100
rect 18414 4088 18420 4140
rect 18472 4088 18478 4140
rect 18506 4088 18512 4140
rect 18564 4128 18570 4140
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18564 4100 19165 4128
rect 18564 4088 18570 4100
rect 19153 4097 19165 4100
rect 19199 4097 19211 4131
rect 19153 4091 19211 4097
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 19628 4128 19656 4168
rect 19300 4100 19656 4128
rect 19300 4088 19306 4100
rect 9876 4032 10088 4060
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 2958 3992 2964 4004
rect 2271 3964 2964 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 2958 3952 2964 3964
rect 3016 3992 3022 4004
rect 3016 3964 3372 3992
rect 3016 3952 3022 3964
rect 3344 3936 3372 3964
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 4985 3995 5043 4001
rect 4985 3992 4997 3995
rect 3660 3964 4752 3992
rect 3660 3952 3666 3964
rect 2590 3884 2596 3936
rect 2648 3884 2654 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4157 3887 4215 3893
rect 4614 3884 4620 3936
rect 4672 3884 4678 3936
rect 4724 3924 4752 3964
rect 4908 3964 4997 3992
rect 4908 3924 4936 3964
rect 4985 3961 4997 3964
rect 5031 3961 5043 3995
rect 4985 3955 5043 3961
rect 5166 3952 5172 4004
rect 5224 3952 5230 4004
rect 6733 3995 6791 4001
rect 6733 3961 6745 3995
rect 6779 3992 6791 3995
rect 7116 3992 7144 4020
rect 6779 3964 7144 3992
rect 6779 3961 6791 3964
rect 6733 3955 6791 3961
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 9876 4001 9904 4032
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 14461 4063 14519 4069
rect 11296 4032 11376 4060
rect 11296 4020 11302 4032
rect 9861 3995 9919 4001
rect 8352 3964 9674 3992
rect 8352 3952 8358 3964
rect 4724 3896 4936 3924
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6052 3896 6561 3924
rect 6052 3884 6058 3896
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 8812 3896 9413 3924
rect 8812 3884 8818 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9646 3924 9674 3964
rect 9861 3961 9873 3995
rect 9907 3961 9919 3995
rect 9950 3992 9956 4004
rect 9861 3955 9919 3961
rect 9948 3952 9956 3992
rect 10008 3952 10014 4004
rect 11348 4001 11376 4032
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4060 15071 4063
rect 15102 4060 15108 4072
rect 15059 4032 15108 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 11333 3995 11391 4001
rect 11333 3961 11345 3995
rect 11379 3961 11391 3995
rect 11333 3955 11391 3961
rect 13538 3952 13544 4004
rect 13596 3992 13602 4004
rect 14476 3992 14504 4023
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 15620 4032 16313 4060
rect 15620 4020 15626 4032
rect 16301 4029 16313 4032
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 18104 4032 18245 4060
rect 18104 4020 18110 4032
rect 18233 4029 18245 4032
rect 18279 4029 18291 4063
rect 18233 4023 18291 4029
rect 19337 4063 19395 4069
rect 19337 4029 19349 4063
rect 19383 4029 19395 4063
rect 19628 4060 19656 4100
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 19981 4131 20039 4137
rect 19751 4100 19932 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 19797 4063 19855 4069
rect 19797 4060 19809 4063
rect 19628 4032 19809 4060
rect 19337 4023 19395 4029
rect 19797 4029 19809 4032
rect 19843 4029 19855 4063
rect 19904 4060 19932 4100
rect 19981 4097 19993 4131
rect 20027 4128 20039 4131
rect 20530 4128 20536 4140
rect 20027 4100 20536 4128
rect 20027 4097 20039 4100
rect 19981 4091 20039 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20640 4128 20668 4168
rect 21284 4168 23244 4196
rect 21284 4128 21312 4168
rect 20640 4100 21312 4128
rect 21358 4088 21364 4140
rect 21416 4137 21422 4140
rect 21416 4128 21428 4137
rect 22088 4131 22146 4137
rect 21416 4100 21461 4128
rect 21416 4091 21428 4100
rect 22088 4097 22100 4131
rect 22134 4128 22146 4131
rect 23106 4128 23112 4140
rect 22134 4100 23112 4128
rect 22134 4097 22146 4100
rect 22088 4091 22146 4097
rect 21416 4088 21422 4091
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23216 4128 23244 4168
rect 23753 4165 23765 4199
rect 23799 4196 23811 4199
rect 24026 4196 24032 4208
rect 23799 4168 24032 4196
rect 23799 4165 23811 4168
rect 23753 4159 23811 4165
rect 24026 4156 24032 4168
rect 24084 4156 24090 4208
rect 24136 4128 24164 4224
rect 24872 4196 24900 4224
rect 24780 4168 24900 4196
rect 24305 4131 24363 4137
rect 24305 4128 24317 4131
rect 23216 4100 23980 4128
rect 24136 4100 24317 4128
rect 20254 4060 20260 4072
rect 19904 4032 20260 4060
rect 19797 4023 19855 4029
rect 13596 3964 14504 3992
rect 13596 3952 13602 3964
rect 15746 3952 15752 4004
rect 15804 3952 15810 4004
rect 19352 3992 19380 4023
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 21637 4063 21695 4069
rect 21637 4029 21649 4063
rect 21683 4060 21695 4063
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 21683 4032 21833 4060
rect 21683 4029 21695 4032
rect 21637 4023 21695 4029
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 20530 3992 20536 4004
rect 19352 3964 20536 3992
rect 20530 3952 20536 3964
rect 20588 3952 20594 4004
rect 9948 3924 9976 3952
rect 9646 3896 9976 3924
rect 9401 3887 9459 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12768 3896 13093 3924
rect 12768 3884 12774 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13081 3887 13139 3893
rect 13906 3884 13912 3936
rect 13964 3884 13970 3936
rect 14826 3884 14832 3936
rect 14884 3884 14890 3936
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 16908 3896 18981 3924
rect 16908 3884 16914 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 19334 3884 19340 3936
rect 19392 3884 19398 3936
rect 20162 3884 20168 3936
rect 20220 3884 20226 3936
rect 21836 3924 21864 4023
rect 23842 4020 23848 4072
rect 23900 4020 23906 4072
rect 23952 4060 23980 4100
rect 24305 4097 24317 4100
rect 24351 4097 24363 4131
rect 24305 4091 24363 4097
rect 24486 4088 24492 4140
rect 24544 4088 24550 4140
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24780 4128 24808 4168
rect 25130 4156 25136 4208
rect 25188 4196 25194 4208
rect 26421 4199 26479 4205
rect 26421 4196 26433 4199
rect 25188 4168 26433 4196
rect 25188 4156 25194 4168
rect 26421 4165 26433 4168
rect 26467 4196 26479 4199
rect 27154 4196 27160 4208
rect 26467 4168 27160 4196
rect 26467 4165 26479 4168
rect 26421 4159 26479 4165
rect 27154 4156 27160 4168
rect 27212 4196 27218 4208
rect 28169 4199 28227 4205
rect 28169 4196 28181 4199
rect 27212 4168 28181 4196
rect 27212 4156 27218 4168
rect 28169 4165 28181 4168
rect 28215 4165 28227 4199
rect 28169 4159 28227 4165
rect 28353 4199 28411 4205
rect 28353 4165 28365 4199
rect 28399 4196 28411 4199
rect 29178 4196 29184 4208
rect 28399 4168 29184 4196
rect 28399 4165 28411 4168
rect 28353 4159 28411 4165
rect 29178 4156 29184 4168
rect 29236 4156 29242 4208
rect 30006 4156 30012 4208
rect 30064 4196 30070 4208
rect 30064 4168 30604 4196
rect 30064 4156 30070 4168
rect 24627 4100 24808 4128
rect 24848 4131 24906 4137
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 24848 4097 24860 4131
rect 24894 4128 24906 4131
rect 25406 4128 25412 4140
rect 24894 4100 25412 4128
rect 24894 4097 24906 4100
rect 24848 4091 24906 4097
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 26513 4131 26571 4137
rect 26513 4097 26525 4131
rect 26559 4128 26571 4131
rect 27798 4128 27804 4140
rect 26559 4100 27804 4128
rect 26559 4097 26571 4100
rect 26513 4091 26571 4097
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 27982 4088 27988 4140
rect 28040 4088 28046 4140
rect 29546 4137 29552 4140
rect 29540 4128 29552 4137
rect 29507 4100 29552 4128
rect 29540 4091 29552 4100
rect 29546 4088 29552 4091
rect 29604 4088 29610 4140
rect 30576 4128 30604 4168
rect 30650 4156 30656 4208
rect 30708 4196 30714 4208
rect 31478 4196 31484 4208
rect 30708 4168 31484 4196
rect 30708 4156 30714 4168
rect 31478 4156 31484 4168
rect 31536 4156 31542 4208
rect 33796 4196 33824 4236
rect 35894 4224 35900 4236
rect 35952 4224 35958 4276
rect 37090 4224 37096 4276
rect 37148 4264 37154 4276
rect 37277 4267 37335 4273
rect 37277 4264 37289 4267
rect 37148 4236 37289 4264
rect 37148 4224 37154 4236
rect 37277 4233 37289 4236
rect 37323 4233 37335 4267
rect 37277 4227 37335 4233
rect 37458 4224 37464 4276
rect 37516 4224 37522 4276
rect 37645 4267 37703 4273
rect 37645 4233 37657 4267
rect 37691 4264 37703 4267
rect 38378 4264 38384 4276
rect 37691 4236 38384 4264
rect 37691 4233 37703 4236
rect 37645 4227 37703 4233
rect 38378 4224 38384 4236
rect 38436 4224 38442 4276
rect 34238 4196 34244 4208
rect 31956 4168 32444 4196
rect 31113 4131 31171 4137
rect 31113 4128 31125 4131
rect 30576 4100 31125 4128
rect 31113 4097 31125 4100
rect 31159 4097 31171 4131
rect 31113 4091 31171 4097
rect 31202 4088 31208 4140
rect 31260 4088 31266 4140
rect 31754 4088 31760 4140
rect 31812 4088 31818 4140
rect 31956 4137 31984 4168
rect 32416 4140 32444 4168
rect 33428 4168 33824 4196
rect 33888 4168 34244 4196
rect 31941 4131 31999 4137
rect 31941 4097 31953 4131
rect 31987 4097 31999 4131
rect 31941 4091 31999 4097
rect 32398 4088 32404 4140
rect 32456 4088 32462 4140
rect 32674 4088 32680 4140
rect 32732 4088 32738 4140
rect 33428 4137 33456 4168
rect 33888 4137 33916 4168
rect 34238 4156 34244 4168
rect 34296 4196 34302 4208
rect 37476 4196 37504 4224
rect 34296 4168 37504 4196
rect 34296 4156 34302 4168
rect 33413 4131 33471 4137
rect 33413 4097 33425 4131
rect 33459 4097 33471 4131
rect 33413 4091 33471 4097
rect 33781 4131 33839 4137
rect 33781 4097 33793 4131
rect 33827 4097 33839 4131
rect 33781 4091 33839 4097
rect 33873 4131 33931 4137
rect 33873 4097 33885 4131
rect 33919 4097 33931 4131
rect 33873 4091 33931 4097
rect 34140 4131 34198 4137
rect 34140 4097 34152 4131
rect 34186 4128 34198 4131
rect 34422 4128 34428 4140
rect 34186 4100 34428 4128
rect 34186 4097 34198 4100
rect 34140 4091 34198 4097
rect 24504 4060 24532 4088
rect 23952 4032 24532 4060
rect 26697 4063 26755 4069
rect 26697 4029 26709 4063
rect 26743 4060 26755 4063
rect 26878 4060 26884 4072
rect 26743 4032 26884 4060
rect 26743 4029 26755 4032
rect 26697 4023 26755 4029
rect 26878 4020 26884 4032
rect 26936 4020 26942 4072
rect 27430 4020 27436 4072
rect 27488 4020 27494 4072
rect 27525 4063 27583 4069
rect 27525 4029 27537 4063
rect 27571 4060 27583 4063
rect 27614 4060 27620 4072
rect 27571 4032 27620 4060
rect 27571 4029 27583 4032
rect 27525 4023 27583 4029
rect 27614 4020 27620 4032
rect 27672 4020 27678 4072
rect 27890 4020 27896 4072
rect 27948 4060 27954 4072
rect 28537 4063 28595 4069
rect 28537 4060 28549 4063
rect 27948 4032 28549 4060
rect 27948 4020 27954 4032
rect 28537 4029 28549 4032
rect 28583 4029 28595 4063
rect 28537 4023 28595 4029
rect 28994 4020 29000 4072
rect 29052 4060 29058 4072
rect 29273 4063 29331 4069
rect 29273 4060 29285 4063
rect 29052 4032 29285 4060
rect 29052 4020 29058 4032
rect 29273 4029 29285 4032
rect 29319 4029 29331 4063
rect 29273 4023 29331 4029
rect 23201 3995 23259 4001
rect 23201 3961 23213 3995
rect 23247 3992 23259 3995
rect 25961 3995 26019 4001
rect 23247 3964 23428 3992
rect 23247 3961 23259 3964
rect 23201 3955 23259 3961
rect 23400 3936 23428 3964
rect 25961 3961 25973 3995
rect 26007 3992 26019 3995
rect 26234 3992 26240 4004
rect 26007 3964 26240 3992
rect 26007 3961 26019 3964
rect 25961 3955 26019 3961
rect 26234 3952 26240 3964
rect 26292 3992 26298 4004
rect 26292 3964 27476 3992
rect 26292 3952 26298 3964
rect 27448 3936 27476 3964
rect 29086 3952 29092 4004
rect 29144 3992 29150 4004
rect 29181 3995 29239 4001
rect 29181 3992 29193 3995
rect 29144 3964 29193 3992
rect 29144 3952 29150 3964
rect 29181 3961 29193 3964
rect 29227 3961 29239 3995
rect 29181 3955 29239 3961
rect 22094 3924 22100 3936
rect 21836 3896 22100 3924
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 23290 3884 23296 3936
rect 23348 3884 23354 3936
rect 23382 3884 23388 3936
rect 23440 3884 23446 3936
rect 24118 3884 24124 3936
rect 24176 3884 24182 3936
rect 26050 3884 26056 3936
rect 26108 3884 26114 3936
rect 27430 3884 27436 3936
rect 27488 3884 27494 3936
rect 29288 3924 29316 4023
rect 31018 4020 31024 4072
rect 31076 4060 31082 4072
rect 31389 4063 31447 4069
rect 31389 4060 31401 4063
rect 31076 4032 31401 4060
rect 31076 4020 31082 4032
rect 31389 4029 31401 4032
rect 31435 4060 31447 4063
rect 31435 4032 31754 4060
rect 31435 4029 31447 4032
rect 31389 4023 31447 4029
rect 30282 3952 30288 4004
rect 30340 3992 30346 4004
rect 31573 3995 31631 4001
rect 31573 3992 31585 3995
rect 30340 3964 31585 3992
rect 30340 3952 30346 3964
rect 31573 3961 31585 3964
rect 31619 3961 31631 3995
rect 31726 3992 31754 4032
rect 32214 4020 32220 4072
rect 32272 4060 32278 4072
rect 33796 4060 33824 4091
rect 34422 4088 34428 4100
rect 34480 4088 34486 4140
rect 35360 4137 35388 4168
rect 37734 4156 37740 4208
rect 37792 4196 37798 4208
rect 38194 4196 38200 4208
rect 37792 4168 38200 4196
rect 37792 4156 37798 4168
rect 38194 4156 38200 4168
rect 38252 4156 38258 4208
rect 35618 4137 35624 4140
rect 35345 4131 35403 4137
rect 35345 4097 35357 4131
rect 35391 4097 35403 4131
rect 35612 4128 35624 4137
rect 35579 4100 35624 4128
rect 35345 4091 35403 4097
rect 35612 4091 35624 4100
rect 35618 4088 35624 4091
rect 35676 4088 35682 4140
rect 35894 4088 35900 4140
rect 35952 4128 35958 4140
rect 35952 4100 36400 4128
rect 35952 4088 35958 4100
rect 32272 4032 33824 4060
rect 36372 4060 36400 4100
rect 36814 4088 36820 4140
rect 36872 4128 36878 4140
rect 37093 4131 37151 4137
rect 37093 4128 37105 4131
rect 36872 4100 37105 4128
rect 36872 4088 36878 4100
rect 37093 4097 37105 4100
rect 37139 4097 37151 4131
rect 37093 4091 37151 4097
rect 38289 4131 38347 4137
rect 38289 4097 38301 4131
rect 38335 4128 38347 4131
rect 38562 4128 38568 4140
rect 38335 4100 38568 4128
rect 38335 4097 38347 4100
rect 38289 4091 38347 4097
rect 38562 4088 38568 4100
rect 38620 4088 38626 4140
rect 38654 4088 38660 4140
rect 38712 4088 38718 4140
rect 37737 4063 37795 4069
rect 37737 4060 37749 4063
rect 36372 4032 37749 4060
rect 32272 4020 32278 4032
rect 37737 4029 37749 4032
rect 37783 4029 37795 4063
rect 37737 4023 37795 4029
rect 37918 4020 37924 4072
rect 37976 4020 37982 4072
rect 38473 4063 38531 4069
rect 38473 4029 38485 4063
rect 38519 4060 38531 4063
rect 38672 4060 38700 4088
rect 38519 4032 38700 4060
rect 38519 4029 38531 4032
rect 38473 4023 38531 4029
rect 36725 3995 36783 4001
rect 31726 3964 33180 3992
rect 31573 3955 31631 3961
rect 29914 3924 29920 3936
rect 29288 3896 29920 3924
rect 29914 3884 29920 3896
rect 29972 3884 29978 3936
rect 30650 3884 30656 3936
rect 30708 3884 30714 3936
rect 30745 3927 30803 3933
rect 30745 3893 30757 3927
rect 30791 3924 30803 3927
rect 30834 3924 30840 3936
rect 30791 3896 30840 3924
rect 30791 3893 30803 3896
rect 30745 3887 30803 3893
rect 30834 3884 30840 3896
rect 30892 3884 30898 3936
rect 30926 3884 30932 3936
rect 30984 3924 30990 3936
rect 31938 3924 31944 3936
rect 30984 3896 31944 3924
rect 30984 3884 30990 3896
rect 31938 3884 31944 3896
rect 31996 3884 32002 3936
rect 33152 3933 33180 3964
rect 36725 3961 36737 3995
rect 36771 3992 36783 3995
rect 37182 3992 37188 4004
rect 36771 3964 37188 3992
rect 36771 3961 36783 3964
rect 36725 3955 36783 3961
rect 37182 3952 37188 3964
rect 37240 3952 37246 4004
rect 33137 3927 33195 3933
rect 33137 3893 33149 3927
rect 33183 3924 33195 3927
rect 33226 3924 33232 3936
rect 33183 3896 33232 3924
rect 33183 3893 33195 3896
rect 33137 3887 33195 3893
rect 33226 3884 33232 3896
rect 33284 3884 33290 3936
rect 35253 3927 35311 3933
rect 35253 3893 35265 3927
rect 35299 3924 35311 3927
rect 35986 3924 35992 3936
rect 35299 3896 35992 3924
rect 35299 3893 35311 3896
rect 35253 3887 35311 3893
rect 35986 3884 35992 3896
rect 36044 3884 36050 3936
rect 36262 3884 36268 3936
rect 36320 3924 36326 3936
rect 36909 3927 36967 3933
rect 36909 3924 36921 3927
rect 36320 3896 36921 3924
rect 36320 3884 36326 3896
rect 36909 3893 36921 3896
rect 36955 3893 36967 3927
rect 37200 3924 37228 3952
rect 37918 3924 37924 3936
rect 37200 3896 37924 3924
rect 36909 3887 36967 3893
rect 37918 3884 37924 3896
rect 37976 3884 37982 3936
rect 38102 3884 38108 3936
rect 38160 3884 38166 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2682 3720 2688 3732
rect 2179 3692 2688 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 2866 3680 2872 3732
rect 2924 3680 2930 3732
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 2406 3612 2412 3664
rect 2464 3652 2470 3664
rect 3436 3652 3464 3683
rect 3602 3680 3608 3732
rect 3660 3680 3666 3732
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4154 3720 4160 3732
rect 3752 3692 4160 3720
rect 3752 3680 3758 3692
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4304 3692 5488 3720
rect 4304 3680 4310 3692
rect 5460 3664 5488 3692
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 9125 3723 9183 3729
rect 6052 3692 7604 3720
rect 6052 3680 6058 3692
rect 2464 3624 5028 3652
rect 2464 3612 2470 3624
rect 5000 3596 5028 3624
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 5500 3624 5948 3652
rect 5500 3612 5506 3624
rect 3053 3587 3111 3593
rect 3053 3553 3065 3587
rect 3099 3584 3111 3587
rect 3694 3584 3700 3596
rect 3099 3556 3700 3584
rect 3099 3553 3111 3556
rect 3053 3547 3111 3553
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3584 3847 3587
rect 3835 3556 4200 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 1854 3476 1860 3528
rect 1912 3476 1918 3528
rect 1946 3476 1952 3528
rect 2004 3476 2010 3528
rect 2222 3476 2228 3528
rect 2280 3476 2286 3528
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2866 3516 2872 3528
rect 2731 3488 2872 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3878 3476 3884 3528
rect 3936 3476 3942 3528
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 4028 3488 4077 3516
rect 4028 3476 4034 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4172 3516 4200 3556
rect 4356 3556 4660 3584
rect 4246 3516 4252 3528
rect 4172 3488 4252 3516
rect 4065 3479 4123 3485
rect 4080 3448 4108 3479
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4356 3525 4384 3556
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4632 3516 4660 3556
rect 4982 3544 4988 3596
rect 5040 3544 5046 3596
rect 5442 3516 5448 3528
rect 4632 3488 5448 3516
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 5920 3525 5948 3624
rect 7374 3612 7380 3664
rect 7432 3612 7438 3664
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 7190 3584 7196 3596
rect 6043 3556 7196 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3510 5963 3519
rect 5951 3485 6040 3510
rect 5905 3482 6040 3485
rect 5905 3479 5963 3482
rect 2332 3420 4108 3448
rect 2332 3392 2360 3420
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4709 3451 4767 3457
rect 4709 3448 4721 3451
rect 4212 3420 4721 3448
rect 4212 3408 4218 3420
rect 4709 3417 4721 3420
rect 4755 3417 4767 3451
rect 4709 3411 4767 3417
rect 5166 3408 5172 3460
rect 5224 3408 5230 3460
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 6012 3448 6040 3482
rect 6270 3476 6276 3528
rect 6328 3476 6334 3528
rect 6086 3448 6092 3460
rect 5316 3420 5948 3448
rect 6012 3420 6092 3448
rect 5316 3408 5322 3420
rect 1670 3340 1676 3392
rect 1728 3340 1734 3392
rect 2314 3340 2320 3392
rect 2372 3340 2378 3392
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 3326 3380 3332 3392
rect 2648 3352 3332 3380
rect 2648 3340 2654 3352
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 3421 3383 3479 3389
rect 3421 3349 3433 3383
rect 3467 3380 3479 3383
rect 3510 3380 3516 3392
rect 3467 3352 3516 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3510 3340 3516 3352
rect 3568 3380 3574 3392
rect 5368 3389 5396 3420
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 3568 3352 5089 3380
rect 3568 3340 3574 3352
rect 5077 3349 5089 3352
rect 5123 3349 5135 3383
rect 5077 3343 5135 3349
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 5534 3340 5540 3392
rect 5592 3340 5598 3392
rect 5920 3380 5948 3420
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 7466 3380 7472 3392
rect 5920 3352 7472 3380
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7576 3380 7604 3692
rect 9125 3689 9137 3723
rect 9171 3720 9183 3723
rect 9398 3720 9404 3732
rect 9171 3692 9404 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 14369 3723 14427 3729
rect 14369 3720 14381 3723
rect 12216 3692 14381 3720
rect 12216 3680 12222 3692
rect 14369 3689 14381 3692
rect 14415 3689 14427 3723
rect 16850 3720 16856 3732
rect 14369 3683 14427 3689
rect 14844 3692 16856 3720
rect 8297 3655 8355 3661
rect 8297 3621 8309 3655
rect 8343 3652 8355 3655
rect 9950 3652 9956 3664
rect 8343 3624 9956 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 10045 3655 10103 3661
rect 10045 3621 10057 3655
rect 10091 3652 10103 3655
rect 10134 3652 10140 3664
rect 10091 3624 10140 3652
rect 10091 3621 10103 3624
rect 10045 3615 10103 3621
rect 10134 3612 10140 3624
rect 10192 3612 10198 3664
rect 11057 3655 11115 3661
rect 11057 3621 11069 3655
rect 11103 3652 11115 3655
rect 11146 3652 11152 3664
rect 11103 3624 11152 3652
rect 11103 3621 11115 3624
rect 11057 3615 11115 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 12618 3612 12624 3664
rect 12676 3612 12682 3664
rect 13906 3612 13912 3664
rect 13964 3612 13970 3664
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8478 3584 8484 3596
rect 8435 3556 8484 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8294 3516 8300 3528
rect 8159 3488 8300 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8036 3448 8064 3479
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8404 3448 8432 3547
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 10502 3584 10508 3596
rect 8588 3556 10508 3584
rect 8588 3525 8616 3556
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12526 3584 12532 3596
rect 12483 3556 12532 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12894 3544 12900 3596
rect 12952 3544 12958 3596
rect 13924 3584 13952 3612
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 13372 3556 13952 3584
rect 14200 3556 14749 3584
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3518 8999 3519
rect 8987 3490 9076 3518
rect 8987 3485 8999 3490
rect 8941 3479 8999 3485
rect 9048 3448 9076 3490
rect 9214 3476 9220 3528
rect 9272 3476 9278 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9456 3488 9781 3516
rect 9456 3476 9462 3488
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10284 3488 10609 3516
rect 10284 3476 10290 3488
rect 10597 3485 10609 3488
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10778 3476 10784 3528
rect 10836 3476 10842 3528
rect 12181 3519 12239 3525
rect 12181 3485 12193 3519
rect 12227 3516 12239 3519
rect 12710 3516 12716 3528
rect 12227 3488 12716 3516
rect 12227 3485 12239 3488
rect 12181 3479 12239 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3516 12863 3519
rect 13372 3516 13400 3556
rect 12851 3488 13400 3516
rect 13449 3519 13507 3525
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14200 3516 14228 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 13771 3488 14228 3516
rect 14369 3519 14427 3525
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14369 3485 14381 3519
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14844 3516 14872 3692
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17954 3680 17960 3732
rect 18012 3680 18018 3732
rect 19242 3680 19248 3732
rect 19300 3680 19306 3732
rect 20717 3723 20775 3729
rect 20717 3689 20729 3723
rect 20763 3720 20775 3723
rect 22002 3720 22008 3732
rect 20763 3692 22008 3720
rect 20763 3689 20775 3692
rect 20717 3683 20775 3689
rect 22002 3680 22008 3692
rect 22060 3680 22066 3732
rect 22189 3723 22247 3729
rect 22189 3689 22201 3723
rect 22235 3720 22247 3723
rect 22922 3720 22928 3732
rect 22235 3692 22928 3720
rect 22235 3689 22247 3692
rect 22189 3683 22247 3689
rect 22922 3680 22928 3692
rect 22980 3720 22986 3732
rect 22980 3692 23796 3720
rect 22980 3680 22986 3692
rect 17865 3655 17923 3661
rect 17865 3621 17877 3655
rect 17911 3652 17923 3655
rect 17911 3624 18552 3652
rect 17911 3621 17923 3624
rect 17865 3615 17923 3621
rect 17218 3544 17224 3596
rect 17276 3544 17282 3596
rect 17405 3587 17463 3593
rect 17405 3553 17417 3587
rect 17451 3584 17463 3587
rect 17678 3584 17684 3596
rect 17451 3556 17684 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 18524 3593 18552 3624
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3553 18567 3587
rect 18509 3547 18567 3553
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3584 18751 3587
rect 19260 3584 19288 3680
rect 23017 3655 23075 3661
rect 23017 3621 23029 3655
rect 23063 3652 23075 3655
rect 23768 3652 23796 3692
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 24397 3723 24455 3729
rect 24397 3720 24409 3723
rect 24084 3692 24409 3720
rect 24084 3680 24090 3692
rect 24397 3689 24409 3692
rect 24443 3689 24455 3723
rect 24397 3683 24455 3689
rect 24762 3680 24768 3732
rect 24820 3680 24826 3732
rect 25038 3680 25044 3732
rect 25096 3720 25102 3732
rect 25133 3723 25191 3729
rect 25133 3720 25145 3723
rect 25096 3692 25145 3720
rect 25096 3680 25102 3692
rect 25133 3689 25145 3692
rect 25179 3689 25191 3723
rect 26881 3723 26939 3729
rect 26881 3720 26893 3723
rect 25133 3683 25191 3689
rect 25424 3692 26893 3720
rect 24780 3652 24808 3680
rect 25424 3652 25452 3692
rect 26881 3689 26893 3692
rect 26927 3689 26939 3723
rect 26881 3683 26939 3689
rect 27522 3680 27528 3732
rect 27580 3680 27586 3732
rect 29178 3680 29184 3732
rect 29236 3680 29242 3732
rect 29638 3680 29644 3732
rect 29696 3680 29702 3732
rect 30006 3680 30012 3732
rect 30064 3720 30070 3732
rect 30926 3720 30932 3732
rect 30064 3692 30932 3720
rect 30064 3680 30070 3692
rect 30926 3680 30932 3692
rect 30984 3680 30990 3732
rect 31389 3723 31447 3729
rect 31389 3689 31401 3723
rect 31435 3720 31447 3723
rect 31570 3720 31576 3732
rect 31435 3692 31576 3720
rect 31435 3689 31447 3692
rect 31389 3683 31447 3689
rect 31570 3680 31576 3692
rect 31628 3680 31634 3732
rect 32030 3680 32036 3732
rect 32088 3720 32094 3732
rect 32861 3723 32919 3729
rect 32861 3720 32873 3723
rect 32088 3692 32873 3720
rect 32088 3680 32094 3692
rect 32861 3689 32873 3692
rect 32907 3689 32919 3723
rect 32861 3683 32919 3689
rect 33042 3680 33048 3732
rect 33100 3680 33106 3732
rect 34698 3680 34704 3732
rect 34756 3680 34762 3732
rect 35342 3680 35348 3732
rect 35400 3720 35406 3732
rect 37274 3720 37280 3732
rect 35400 3692 37280 3720
rect 35400 3680 35406 3692
rect 37274 3680 37280 3692
rect 37332 3680 37338 3732
rect 37737 3723 37795 3729
rect 37737 3689 37749 3723
rect 37783 3689 37795 3723
rect 37737 3683 37795 3689
rect 23063 3624 23704 3652
rect 23768 3624 24532 3652
rect 24780 3624 25452 3652
rect 26789 3655 26847 3661
rect 23063 3621 23075 3624
rect 23017 3615 23075 3621
rect 18739 3556 19288 3584
rect 18739 3553 18751 3556
rect 18693 3547 18751 3553
rect 22370 3544 22376 3596
rect 22428 3544 22434 3596
rect 23676 3593 23704 3624
rect 23661 3587 23719 3593
rect 23661 3553 23673 3587
rect 23707 3553 23719 3587
rect 23661 3547 23719 3553
rect 23768 3556 24440 3584
rect 14507 3488 14872 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 10870 3448 10876 3460
rect 8036 3420 8432 3448
rect 8496 3420 8892 3448
rect 9048 3420 10876 3448
rect 8496 3380 8524 3420
rect 7576 3352 8524 3380
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 8864 3380 8892 3420
rect 10870 3408 10876 3420
rect 10928 3408 10934 3460
rect 10980 3420 12434 3448
rect 10318 3380 10324 3392
rect 8864 3352 10324 3380
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10980 3389 11008 3420
rect 10965 3383 11023 3389
rect 10965 3349 10977 3383
rect 11011 3349 11023 3383
rect 12406 3380 12434 3420
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 13464 3448 13492 3479
rect 13998 3448 14004 3460
rect 12676 3420 13492 3448
rect 13924 3420 14004 3448
rect 12676 3408 12682 3420
rect 13814 3380 13820 3392
rect 12406 3352 13820 3380
rect 10965 3343 11023 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 13924 3389 13952 3420
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 14384 3448 14412 3479
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 14976 3488 15301 3516
rect 14976 3476 14982 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 15289 3479 15347 3485
rect 16592 3488 17049 3516
rect 16592 3460 16620 3488
rect 17037 3485 17049 3488
rect 17083 3516 17095 3519
rect 17310 3516 17316 3528
rect 17083 3488 17316 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 17862 3516 17868 3528
rect 17543 3488 17868 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 18966 3516 18972 3528
rect 18923 3488 18972 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 14550 3448 14556 3460
rect 14384 3420 14556 3448
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 14642 3408 14648 3460
rect 14700 3408 14706 3460
rect 16574 3408 16580 3460
rect 16632 3408 16638 3460
rect 16666 3408 16672 3460
rect 16724 3448 16730 3460
rect 16770 3451 16828 3457
rect 16770 3448 16782 3451
rect 16724 3420 16782 3448
rect 16724 3408 16730 3420
rect 16770 3417 16782 3420
rect 16816 3417 16828 3451
rect 16770 3411 16828 3417
rect 17402 3408 17408 3460
rect 17460 3408 17466 3460
rect 17954 3408 17960 3460
rect 18012 3448 18018 3460
rect 19260 3448 19288 3479
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 22094 3516 22100 3528
rect 20855 3488 22100 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 23014 3516 23020 3528
rect 22603 3488 23020 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 23768 3516 23796 3556
rect 23164 3488 23796 3516
rect 24029 3519 24087 3525
rect 23164 3476 23170 3488
rect 24029 3485 24041 3519
rect 24075 3485 24087 3519
rect 24029 3479 24087 3485
rect 24213 3519 24271 3525
rect 24213 3485 24225 3519
rect 24259 3485 24271 3519
rect 24213 3479 24271 3485
rect 18012 3420 19288 3448
rect 21076 3451 21134 3457
rect 18012 3408 18018 3420
rect 21076 3417 21088 3451
rect 21122 3448 21134 3451
rect 21122 3420 22140 3448
rect 21122 3417 21134 3420
rect 21076 3411 21134 3417
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3349 13967 3383
rect 13909 3343 13967 3349
rect 14182 3340 14188 3392
rect 14240 3340 14246 3392
rect 15102 3340 15108 3392
rect 15160 3380 15166 3392
rect 15657 3383 15715 3389
rect 15657 3380 15669 3383
rect 15160 3352 15669 3380
rect 15160 3340 15166 3352
rect 15657 3349 15669 3352
rect 15703 3380 15715 3383
rect 17420 3380 17448 3408
rect 22112 3392 22140 3420
rect 22738 3408 22744 3460
rect 22796 3448 22802 3460
rect 24044 3448 24072 3479
rect 22796 3420 24072 3448
rect 22796 3408 22802 3420
rect 15703 3352 17448 3380
rect 15703 3349 15715 3352
rect 15657 3343 15715 3349
rect 19058 3340 19064 3392
rect 19116 3340 19122 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 19484 3352 19901 3380
rect 19484 3340 19490 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 19889 3343 19947 3349
rect 22094 3340 22100 3392
rect 22152 3340 22158 3392
rect 22646 3340 22652 3392
rect 22704 3340 22710 3392
rect 23109 3383 23167 3389
rect 23109 3349 23121 3383
rect 23155 3380 23167 3383
rect 23198 3380 23204 3392
rect 23155 3352 23204 3380
rect 23155 3349 23167 3352
rect 23109 3343 23167 3349
rect 23198 3340 23204 3352
rect 23256 3340 23262 3392
rect 23474 3340 23480 3392
rect 23532 3380 23538 3392
rect 23845 3383 23903 3389
rect 23845 3380 23857 3383
rect 23532 3352 23857 3380
rect 23532 3340 23538 3352
rect 23845 3349 23857 3352
rect 23891 3349 23903 3383
rect 24228 3380 24256 3479
rect 24412 3448 24440 3556
rect 24504 3516 24532 3624
rect 26789 3621 26801 3655
rect 26835 3652 26847 3655
rect 27540 3652 27568 3680
rect 26835 3624 27568 3652
rect 26835 3621 26847 3624
rect 26789 3615 26847 3621
rect 31938 3612 31944 3664
rect 31996 3652 32002 3664
rect 33060 3652 33088 3680
rect 35434 3652 35440 3664
rect 31996 3624 33088 3652
rect 33152 3624 35440 3652
rect 31996 3612 32002 3624
rect 24854 3544 24860 3596
rect 24912 3584 24918 3596
rect 25409 3587 25467 3593
rect 25409 3584 25421 3587
rect 24912 3556 25421 3584
rect 24912 3544 24918 3556
rect 25409 3553 25421 3556
rect 25455 3553 25467 3587
rect 25409 3547 25467 3553
rect 27430 3544 27436 3596
rect 27488 3544 27494 3596
rect 28997 3587 29055 3593
rect 28997 3553 29009 3587
rect 29043 3584 29055 3587
rect 29043 3556 29868 3584
rect 29043 3553 29055 3556
rect 28997 3547 29055 3553
rect 24949 3519 25007 3525
rect 24949 3516 24961 3519
rect 24504 3488 24961 3516
rect 24949 3485 24961 3488
rect 24995 3485 25007 3519
rect 24949 3479 25007 3485
rect 25317 3519 25375 3525
rect 25317 3485 25329 3519
rect 25363 3485 25375 3519
rect 25317 3479 25375 3485
rect 25332 3448 25360 3479
rect 25958 3476 25964 3528
rect 26016 3516 26022 3528
rect 27617 3519 27675 3525
rect 27617 3516 27629 3519
rect 26016 3488 27629 3516
rect 26016 3476 26022 3488
rect 27617 3485 27629 3488
rect 27663 3485 27675 3519
rect 27617 3479 27675 3485
rect 28353 3519 28411 3525
rect 28353 3485 28365 3519
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 24412 3420 25360 3448
rect 25676 3451 25734 3457
rect 25676 3417 25688 3451
rect 25722 3448 25734 3451
rect 26694 3448 26700 3460
rect 25722 3420 26700 3448
rect 25722 3417 25734 3420
rect 25676 3411 25734 3417
rect 26694 3408 26700 3420
rect 26752 3408 26758 3460
rect 26970 3408 26976 3460
rect 27028 3448 27034 3460
rect 28368 3448 28396 3479
rect 29362 3476 29368 3528
rect 29420 3476 29426 3528
rect 29840 3525 29868 3556
rect 31662 3544 31668 3596
rect 31720 3584 31726 3596
rect 32677 3587 32735 3593
rect 32677 3584 32689 3587
rect 31720 3556 32689 3584
rect 31720 3544 31726 3556
rect 32677 3553 32689 3556
rect 32723 3553 32735 3587
rect 32677 3547 32735 3553
rect 32950 3544 32956 3596
rect 33008 3584 33014 3596
rect 33152 3584 33180 3624
rect 35434 3612 35440 3624
rect 35492 3612 35498 3664
rect 35802 3652 35808 3664
rect 35636 3624 35808 3652
rect 33008 3556 33180 3584
rect 33008 3544 33014 3556
rect 33226 3544 33232 3596
rect 33284 3584 33290 3596
rect 35253 3587 35311 3593
rect 35253 3584 35265 3587
rect 33284 3556 35265 3584
rect 33284 3544 33290 3556
rect 35253 3553 35265 3556
rect 35299 3553 35311 3587
rect 35253 3547 35311 3553
rect 35526 3544 35532 3596
rect 35584 3544 35590 3596
rect 29825 3519 29883 3525
rect 29825 3485 29837 3519
rect 29871 3485 29883 3519
rect 29825 3479 29883 3485
rect 29914 3476 29920 3528
rect 29972 3516 29978 3528
rect 31297 3519 31355 3525
rect 31297 3516 31309 3519
rect 29972 3488 31309 3516
rect 29972 3476 29978 3488
rect 31297 3485 31309 3488
rect 31343 3485 31355 3519
rect 31297 3479 31355 3485
rect 31386 3476 31392 3528
rect 31444 3516 31450 3528
rect 31941 3519 31999 3525
rect 31941 3516 31953 3519
rect 31444 3488 31953 3516
rect 31444 3476 31450 3488
rect 31941 3485 31953 3488
rect 31987 3485 31999 3519
rect 31941 3479 31999 3485
rect 32030 3476 32036 3528
rect 32088 3516 32094 3528
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 32088 3488 33057 3516
rect 32088 3476 32094 3488
rect 33045 3485 33057 3488
rect 33091 3485 33103 3519
rect 33045 3479 33103 3485
rect 34422 3476 34428 3528
rect 34480 3476 34486 3528
rect 35069 3519 35127 3525
rect 35069 3485 35081 3519
rect 35115 3516 35127 3519
rect 35636 3516 35664 3624
rect 35802 3612 35808 3624
rect 35860 3612 35866 3664
rect 36354 3612 36360 3664
rect 36412 3652 36418 3664
rect 37752 3652 37780 3683
rect 38102 3680 38108 3732
rect 38160 3680 38166 3732
rect 36412 3624 37780 3652
rect 36412 3612 36418 3624
rect 35894 3544 35900 3596
rect 35952 3544 35958 3596
rect 38120 3584 38148 3680
rect 37476 3556 38148 3584
rect 38197 3587 38255 3593
rect 35115 3488 35664 3516
rect 35115 3485 35127 3488
rect 35069 3479 35127 3485
rect 35710 3476 35716 3528
rect 35768 3476 35774 3528
rect 37476 3525 37504 3556
rect 38197 3553 38209 3587
rect 38243 3584 38255 3587
rect 38286 3584 38292 3596
rect 38243 3556 38292 3584
rect 38243 3553 38255 3556
rect 38197 3547 38255 3553
rect 38286 3544 38292 3556
rect 38344 3544 38350 3596
rect 37461 3519 37519 3525
rect 37461 3485 37473 3519
rect 37507 3485 37519 3519
rect 37461 3479 37519 3485
rect 37737 3519 37795 3525
rect 37737 3485 37749 3519
rect 37783 3485 37795 3519
rect 37737 3479 37795 3485
rect 30466 3448 30472 3460
rect 27028 3420 28396 3448
rect 29932 3420 30472 3448
rect 27028 3408 27034 3420
rect 24486 3380 24492 3392
rect 24228 3352 24492 3380
rect 23845 3343 23903 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 28258 3340 28264 3392
rect 28316 3340 28322 3392
rect 29932 3389 29960 3420
rect 30466 3408 30472 3420
rect 30524 3448 30530 3460
rect 30650 3448 30656 3460
rect 30524 3420 30656 3448
rect 30524 3408 30530 3420
rect 30650 3408 30656 3420
rect 30708 3408 30714 3460
rect 31052 3451 31110 3457
rect 31052 3417 31064 3451
rect 31098 3448 31110 3451
rect 32125 3451 32183 3457
rect 32125 3448 32137 3451
rect 31098 3420 32137 3448
rect 31098 3417 31110 3420
rect 31052 3411 31110 3417
rect 32125 3417 32137 3420
rect 32171 3417 32183 3451
rect 32125 3411 32183 3417
rect 33594 3408 33600 3460
rect 33652 3408 33658 3460
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 36265 3451 36323 3457
rect 36265 3448 36277 3451
rect 36044 3420 36277 3448
rect 36044 3408 36050 3420
rect 36265 3417 36277 3420
rect 36311 3417 36323 3451
rect 36265 3411 36323 3417
rect 36538 3408 36544 3460
rect 36596 3448 36602 3460
rect 37752 3448 37780 3479
rect 37826 3476 37832 3528
rect 37884 3516 37890 3528
rect 38105 3519 38163 3525
rect 38105 3516 38117 3519
rect 37884 3488 38117 3516
rect 37884 3476 37890 3488
rect 38105 3485 38117 3488
rect 38151 3485 38163 3519
rect 38105 3479 38163 3485
rect 36596 3420 37780 3448
rect 36596 3408 36602 3420
rect 29917 3383 29975 3389
rect 29917 3349 29929 3383
rect 29963 3349 29975 3383
rect 29917 3343 29975 3349
rect 30098 3340 30104 3392
rect 30156 3380 30162 3392
rect 34146 3380 34152 3392
rect 30156 3352 34152 3380
rect 30156 3340 30162 3352
rect 34146 3340 34152 3352
rect 34204 3340 34210 3392
rect 35158 3340 35164 3392
rect 35216 3340 35222 3392
rect 36354 3340 36360 3392
rect 36412 3380 36418 3392
rect 37553 3383 37611 3389
rect 37553 3380 37565 3383
rect 36412 3352 37565 3380
rect 36412 3340 36418 3352
rect 37553 3349 37565 3352
rect 37599 3349 37611 3383
rect 37553 3343 37611 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 1762 3136 1768 3188
rect 1820 3136 1826 3188
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 2409 3179 2467 3185
rect 2409 3176 2421 3179
rect 1912 3148 2421 3176
rect 1912 3136 1918 3148
rect 2409 3145 2421 3148
rect 2455 3145 2467 3179
rect 4246 3176 4252 3188
rect 2409 3139 2467 3145
rect 3528 3148 4252 3176
rect 2314 3068 2320 3120
rect 2372 3068 2378 3120
rect 2774 3068 2780 3120
rect 2832 3068 2838 3120
rect 1026 3000 1032 3052
rect 1084 3040 1090 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 1084 3012 1501 3040
rect 1084 3000 1090 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 1489 3003 1547 3009
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2056 2972 2084 3003
rect 2590 3000 2596 3052
rect 2648 3000 2654 3052
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 2792 3040 2820 3068
rect 2731 3012 2820 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 3142 3000 3148 3052
rect 3200 3000 3206 3052
rect 3418 3000 3424 3052
rect 3476 3000 3482 3052
rect 2958 2972 2964 2984
rect 2056 2944 2964 2972
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3050 2932 3056 2984
rect 3108 2932 3114 2984
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2972 3295 2975
rect 3528 2972 3556 3148
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5537 3179 5595 3185
rect 5537 3176 5549 3179
rect 4856 3148 5549 3176
rect 4856 3136 4862 3148
rect 5537 3145 5549 3148
rect 5583 3145 5595 3179
rect 5537 3139 5595 3145
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6328 3148 6377 3176
rect 6328 3136 6334 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3176 7159 3179
rect 7558 3176 7564 3188
rect 7147 3148 7564 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 8812 3148 11008 3176
rect 8812 3136 8818 3148
rect 3605 3111 3663 3117
rect 3605 3077 3617 3111
rect 3651 3108 3663 3111
rect 6638 3108 6644 3120
rect 3651 3080 6644 3108
rect 3651 3077 3663 3080
rect 3605 3071 3663 3077
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 9214 3108 9220 3120
rect 7208 3080 9220 3108
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 4890 3000 4896 3052
rect 4948 3000 4954 3052
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 7208 3040 7236 3080
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 10778 3068 10784 3120
rect 10836 3068 10842 3120
rect 5307 3012 7236 3040
rect 7285 3043 7343 3049
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 3283 2944 3556 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3660 2944 3893 2972
rect 3660 2932 3666 2944
rect 3881 2941 3893 2944
rect 3927 2941 3939 2975
rect 3881 2935 3939 2941
rect 2498 2864 2504 2916
rect 2556 2864 2562 2916
rect 2682 2864 2688 2916
rect 2740 2864 2746 2916
rect 2777 2907 2835 2913
rect 2777 2873 2789 2907
rect 2823 2904 2835 2907
rect 4080 2904 4108 3000
rect 5350 2932 5356 2984
rect 5408 2932 5414 2984
rect 6178 2932 6184 2984
rect 6236 2932 6242 2984
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 2823 2876 4108 2904
rect 5368 2904 5396 2932
rect 6932 2904 6960 2935
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7300 2972 7328 3003
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7742 3040 7748 3052
rect 7607 3012 7748 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7834 3000 7840 3052
rect 7892 3000 7898 3052
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3040 8079 3043
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 8067 3012 8125 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 10410 3040 10416 3052
rect 9723 3012 10416 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 7064 2944 7328 2972
rect 7653 2975 7711 2981
rect 7064 2932 7070 2944
rect 7653 2941 7665 2975
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 5368 2876 6960 2904
rect 7668 2904 7696 2935
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 8260 2944 8585 2972
rect 8260 2932 8266 2944
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 9048 2904 9076 3000
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9640 2944 10057 2972
rect 9640 2932 9646 2944
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 7668 2876 9076 2904
rect 2823 2873 2835 2876
rect 2777 2867 2835 2873
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2700 2836 2728 2864
rect 2271 2808 2728 2836
rect 3145 2839 3203 2845
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 3145 2805 3157 2839
rect 3191 2836 3203 2839
rect 3786 2836 3792 2848
rect 3191 2808 3792 2836
rect 3191 2805 3203 2808
rect 3145 2799 3203 2805
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5994 2836 6000 2848
rect 5491 2808 6000 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6086 2796 6092 2848
rect 6144 2836 6150 2848
rect 7668 2836 7696 2876
rect 6144 2808 7696 2836
rect 10796 2836 10824 3068
rect 10980 2972 11008 3148
rect 11238 3136 11244 3188
rect 11296 3136 11302 3188
rect 11701 3179 11759 3185
rect 11701 3145 11713 3179
rect 11747 3176 11759 3179
rect 14182 3176 14188 3188
rect 11747 3148 14188 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 14550 3136 14556 3188
rect 14608 3176 14614 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 14608 3148 17141 3176
rect 14608 3136 14614 3148
rect 17129 3145 17141 3148
rect 17175 3145 17187 3179
rect 17129 3139 17187 3145
rect 18782 3136 18788 3188
rect 18840 3136 18846 3188
rect 19058 3136 19064 3188
rect 19116 3136 19122 3188
rect 19429 3179 19487 3185
rect 19429 3145 19441 3179
rect 19475 3176 19487 3179
rect 19978 3176 19984 3188
rect 19475 3148 19984 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 20530 3136 20536 3188
rect 20588 3176 20594 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 20588 3148 21833 3176
rect 20588 3136 20594 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 22094 3136 22100 3188
rect 22152 3136 22158 3188
rect 23566 3136 23572 3188
rect 23624 3176 23630 3188
rect 23624 3148 24532 3176
rect 23624 3136 23630 3148
rect 16574 3108 16580 3120
rect 13280 3080 16580 3108
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3040 11115 3043
rect 11422 3040 11428 3052
rect 11103 3012 11428 3040
rect 11103 3009 11115 3012
rect 11057 3003 11115 3009
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 11514 3000 11520 3052
rect 11572 3000 11578 3052
rect 13280 3049 13308 3080
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 16669 3111 16727 3117
rect 16669 3077 16681 3111
rect 16715 3108 16727 3111
rect 16758 3108 16764 3120
rect 16715 3080 16764 3108
rect 16715 3077 16727 3080
rect 16669 3071 16727 3077
rect 16758 3068 16764 3080
rect 16816 3068 16822 3120
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 11808 2972 11836 3003
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 14458 3040 14464 3052
rect 14016 3012 14464 3040
rect 10980 2944 11836 2972
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 12032 2944 12265 2972
rect 12032 2932 12038 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 11422 2864 11428 2916
rect 11480 2904 11486 2916
rect 12894 2904 12900 2916
rect 11480 2876 12900 2904
rect 11480 2864 11486 2876
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 14016 2904 14044 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3040 15347 3043
rect 15470 3040 15476 3052
rect 15335 3012 15476 3040
rect 15335 3009 15347 3012
rect 15289 3003 15347 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17034 3040 17040 3052
rect 16991 3012 17040 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 18800 3040 18828 3136
rect 18739 3012 18828 3040
rect 19076 3040 19104 3136
rect 22370 3068 22376 3120
rect 22428 3108 22434 3120
rect 22428 3080 24440 3108
rect 22428 3068 22434 3080
rect 19521 3043 19579 3049
rect 19521 3040 19533 3043
rect 19076 3012 19533 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 19521 3009 19533 3012
rect 19567 3009 19579 3043
rect 19521 3003 19579 3009
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20254 3040 20260 3052
rect 20036 3012 20260 3040
rect 20036 3000 20042 3012
rect 20254 3000 20260 3012
rect 20312 3000 20318 3052
rect 20898 3000 20904 3052
rect 20956 3040 20962 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 20956 3012 22017 3040
rect 20956 3000 20962 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3040 22707 3043
rect 23290 3040 23296 3052
rect 22695 3012 23296 3040
rect 22695 3009 22707 3012
rect 22649 3003 22707 3009
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 24118 3000 24124 3052
rect 24176 3000 24182 3052
rect 14090 2932 14096 2984
rect 14148 2932 14154 2984
rect 14182 2932 14188 2984
rect 14240 2932 14246 2984
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15068 2944 15577 2972
rect 15068 2932 15074 2944
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2941 16819 2975
rect 16761 2935 16819 2941
rect 13740 2876 14044 2904
rect 14200 2904 14228 2932
rect 16776 2904 16804 2935
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 17276 2944 17509 2972
rect 17276 2932 17282 2944
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 18874 2932 18880 2984
rect 18932 2932 18938 2984
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 14200 2876 16804 2904
rect 13170 2836 13176 2848
rect 10796 2808 13176 2836
rect 6144 2796 6150 2808
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13449 2839 13507 2845
rect 13449 2805 13461 2839
rect 13495 2836 13507 2839
rect 13740 2836 13768 2876
rect 13495 2808 13768 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 13872 2808 16681 2836
rect 13872 2796 13878 2808
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 16669 2799 16727 2805
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 20088 2836 20116 2935
rect 21082 2932 21088 2984
rect 21140 2932 21146 2984
rect 22738 2932 22744 2984
rect 22796 2972 22802 2984
rect 24412 2981 24440 3080
rect 24504 3040 24532 3148
rect 24946 3136 24952 3188
rect 25004 3136 25010 3188
rect 26602 3136 26608 3188
rect 26660 3136 26666 3188
rect 26786 3136 26792 3188
rect 26844 3176 26850 3188
rect 26973 3179 27031 3185
rect 26973 3176 26985 3179
rect 26844 3148 26985 3176
rect 26844 3136 26850 3148
rect 26973 3145 26985 3148
rect 27019 3145 27031 3179
rect 26973 3139 27031 3145
rect 27706 3136 27712 3188
rect 27764 3136 27770 3188
rect 28258 3136 28264 3188
rect 28316 3136 28322 3188
rect 30190 3136 30196 3188
rect 30248 3136 30254 3188
rect 30834 3136 30840 3188
rect 30892 3176 30898 3188
rect 34514 3176 34520 3188
rect 30892 3148 34520 3176
rect 30892 3136 30898 3148
rect 34514 3136 34520 3148
rect 34572 3136 34578 3188
rect 35158 3136 35164 3188
rect 35216 3176 35222 3188
rect 36449 3179 36507 3185
rect 36449 3176 36461 3179
rect 35216 3148 36461 3176
rect 35216 3136 35222 3148
rect 36449 3145 36461 3148
rect 36495 3145 36507 3179
rect 36449 3139 36507 3145
rect 36814 3136 36820 3188
rect 36872 3136 36878 3188
rect 36998 3136 37004 3188
rect 37056 3176 37062 3188
rect 37056 3148 38240 3176
rect 37056 3136 37062 3148
rect 25314 3068 25320 3120
rect 25372 3108 25378 3120
rect 25372 3080 27200 3108
rect 25372 3068 25378 3080
rect 24504 3012 25360 3040
rect 23017 2975 23075 2981
rect 23017 2972 23029 2975
rect 22796 2944 23029 2972
rect 22796 2932 22802 2944
rect 23017 2941 23029 2944
rect 23063 2941 23075 2975
rect 23017 2935 23075 2941
rect 24397 2975 24455 2981
rect 24397 2941 24409 2975
rect 24443 2941 24455 2975
rect 24397 2935 24455 2941
rect 24946 2932 24952 2984
rect 25004 2972 25010 2984
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 25004 2944 25237 2972
rect 25004 2932 25010 2944
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 25332 2972 25360 3012
rect 26326 3000 26332 3052
rect 26384 3000 26390 3052
rect 27172 3049 27200 3080
rect 26789 3043 26847 3049
rect 26789 3009 26801 3043
rect 26835 3009 26847 3043
rect 26789 3003 26847 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 27433 3043 27491 3049
rect 27433 3009 27445 3043
rect 27479 3040 27491 3043
rect 27724 3040 27752 3136
rect 28276 3108 28304 3136
rect 28276 3080 30420 3108
rect 27479 3012 27752 3040
rect 30101 3043 30159 3049
rect 27479 3009 27491 3012
rect 27433 3003 27491 3009
rect 30101 3009 30113 3043
rect 30147 3040 30159 3043
rect 30282 3040 30288 3052
rect 30147 3012 30288 3040
rect 30147 3009 30159 3012
rect 30101 3003 30159 3009
rect 26418 2972 26424 2984
rect 25332 2944 26424 2972
rect 25225 2935 25283 2941
rect 26418 2932 26424 2944
rect 26476 2932 26482 2984
rect 21637 2907 21695 2913
rect 21637 2873 21649 2907
rect 21683 2904 21695 2907
rect 26804 2904 26832 3003
rect 30282 3000 30288 3012
rect 30340 3000 30346 3052
rect 30392 3049 30420 3080
rect 30650 3068 30656 3120
rect 30708 3108 30714 3120
rect 31386 3108 31392 3120
rect 30708 3080 31392 3108
rect 30708 3068 30714 3080
rect 31386 3068 31392 3080
rect 31444 3068 31450 3120
rect 31938 3108 31944 3120
rect 31772 3080 31944 3108
rect 31772 3049 31800 3080
rect 31938 3068 31944 3080
rect 31996 3068 32002 3120
rect 32306 3068 32312 3120
rect 32364 3108 32370 3120
rect 35802 3108 35808 3120
rect 32364 3080 35808 3108
rect 32364 3068 32370 3080
rect 35802 3068 35808 3080
rect 35860 3068 35866 3120
rect 36832 3108 36860 3136
rect 36004 3080 36860 3108
rect 37277 3111 37335 3117
rect 30377 3043 30435 3049
rect 30377 3009 30389 3043
rect 30423 3009 30435 3043
rect 30377 3003 30435 3009
rect 31757 3043 31815 3049
rect 31757 3009 31769 3043
rect 31803 3009 31815 3043
rect 31757 3003 31815 3009
rect 31846 3000 31852 3052
rect 31904 3040 31910 3052
rect 32585 3043 32643 3049
rect 32585 3040 32597 3043
rect 31904 3012 32597 3040
rect 31904 3000 31910 3012
rect 32585 3009 32597 3012
rect 32631 3009 32643 3043
rect 34054 3040 34060 3052
rect 32585 3003 32643 3009
rect 32876 3012 34060 3040
rect 27338 2932 27344 2984
rect 27396 2972 27402 2984
rect 27709 2975 27767 2981
rect 27709 2972 27721 2975
rect 27396 2944 27721 2972
rect 27396 2932 27402 2944
rect 27709 2941 27721 2944
rect 27755 2941 27767 2975
rect 27709 2935 27767 2941
rect 28258 2932 28264 2984
rect 28316 2972 28322 2984
rect 28905 2975 28963 2981
rect 28905 2972 28917 2975
rect 28316 2944 28917 2972
rect 28316 2932 28322 2944
rect 28905 2941 28917 2944
rect 28951 2941 28963 2975
rect 28905 2935 28963 2941
rect 30466 2932 30472 2984
rect 30524 2972 30530 2984
rect 30745 2975 30803 2981
rect 30745 2972 30757 2975
rect 30524 2944 30757 2972
rect 30524 2932 30530 2944
rect 30745 2941 30757 2944
rect 30791 2941 30803 2975
rect 30745 2935 30803 2941
rect 31202 2932 31208 2984
rect 31260 2972 31266 2984
rect 32493 2975 32551 2981
rect 31260 2944 32168 2972
rect 31260 2932 31266 2944
rect 21683 2876 26832 2904
rect 21683 2873 21695 2876
rect 21637 2867 21695 2873
rect 26878 2864 26884 2916
rect 26936 2904 26942 2916
rect 29178 2904 29184 2916
rect 26936 2876 29184 2904
rect 26936 2864 26942 2876
rect 29178 2864 29184 2876
rect 29236 2864 29242 2916
rect 29288 2876 31754 2904
rect 19392 2808 20116 2836
rect 19392 2796 19398 2808
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 24026 2836 24032 2848
rect 22060 2808 24032 2836
rect 22060 2796 22066 2808
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 24302 2796 24308 2848
rect 24360 2836 24366 2848
rect 26510 2836 26516 2848
rect 24360 2808 26516 2836
rect 24360 2796 24366 2808
rect 26510 2796 26516 2808
rect 26568 2796 26574 2848
rect 28626 2796 28632 2848
rect 28684 2836 28690 2848
rect 29288 2836 29316 2876
rect 28684 2808 29316 2836
rect 31726 2836 31754 2876
rect 32030 2836 32036 2848
rect 31726 2808 32036 2836
rect 28684 2796 28690 2808
rect 32030 2796 32036 2808
rect 32088 2796 32094 2848
rect 32140 2836 32168 2944
rect 32493 2941 32505 2975
rect 32539 2972 32551 2975
rect 32876 2972 32904 3012
rect 34054 3000 34060 3012
rect 34112 3000 34118 3052
rect 34149 3043 34207 3049
rect 34149 3009 34161 3043
rect 34195 3040 34207 3043
rect 34330 3040 34336 3052
rect 34195 3012 34336 3040
rect 34195 3009 34207 3012
rect 34149 3003 34207 3009
rect 34330 3000 34336 3012
rect 34388 3000 34394 3052
rect 34885 3043 34943 3049
rect 34885 3009 34897 3043
rect 34931 3040 34943 3043
rect 36004 3040 36032 3080
rect 37277 3077 37289 3111
rect 37323 3108 37335 3111
rect 37550 3108 37556 3120
rect 37323 3080 37556 3108
rect 37323 3077 37335 3080
rect 37277 3071 37335 3077
rect 37550 3068 37556 3080
rect 37608 3068 37614 3120
rect 38212 3049 38240 3148
rect 34931 3012 36032 3040
rect 36357 3043 36415 3049
rect 34931 3009 34943 3012
rect 34885 3003 34943 3009
rect 36357 3009 36369 3043
rect 36403 3040 36415 3043
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 36403 3012 38025 3040
rect 36403 3009 36415 3012
rect 36357 3003 36415 3009
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 38197 3043 38255 3049
rect 38197 3009 38209 3043
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 38381 3043 38439 3049
rect 38381 3009 38393 3043
rect 38427 3040 38439 3043
rect 38654 3040 38660 3052
rect 38427 3012 38660 3040
rect 38427 3009 38439 3012
rect 38381 3003 38439 3009
rect 38654 3000 38660 3012
rect 38712 3000 38718 3052
rect 32539 2944 32904 2972
rect 32539 2941 32551 2944
rect 32493 2935 32551 2941
rect 32950 2932 32956 2984
rect 33008 2932 33014 2984
rect 34241 2975 34299 2981
rect 34241 2941 34253 2975
rect 34287 2941 34299 2975
rect 34241 2935 34299 2941
rect 32214 2864 32220 2916
rect 32272 2864 32278 2916
rect 34256 2904 34284 2935
rect 34790 2932 34796 2984
rect 34848 2972 34854 2984
rect 35161 2975 35219 2981
rect 35161 2972 35173 2975
rect 34848 2944 35173 2972
rect 34848 2932 34854 2944
rect 35161 2941 35173 2944
rect 35207 2941 35219 2975
rect 35161 2935 35219 2941
rect 36078 2932 36084 2984
rect 36136 2972 36142 2984
rect 37001 2975 37059 2981
rect 37001 2972 37013 2975
rect 36136 2944 37013 2972
rect 36136 2932 36142 2944
rect 37001 2941 37013 2944
rect 37047 2941 37059 2975
rect 37001 2935 37059 2941
rect 37918 2932 37924 2984
rect 37976 2932 37982 2984
rect 32324 2876 34284 2904
rect 34348 2876 37872 2904
rect 32324 2836 32352 2876
rect 32140 2808 32352 2836
rect 32582 2796 32588 2848
rect 32640 2796 32646 2848
rect 33410 2796 33416 2848
rect 33468 2836 33474 2848
rect 34348 2836 34376 2876
rect 37844 2848 37872 2876
rect 33468 2808 34376 2836
rect 33468 2796 33474 2808
rect 36078 2796 36084 2848
rect 36136 2836 36142 2848
rect 36630 2836 36636 2848
rect 36136 2808 36636 2836
rect 36136 2796 36142 2808
rect 36630 2796 36636 2808
rect 36688 2796 36694 2848
rect 37826 2796 37832 2848
rect 37884 2796 37890 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2866 2592 2872 2644
rect 2924 2592 2930 2644
rect 2958 2592 2964 2644
rect 3016 2592 3022 2644
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3200 2604 3801 2632
rect 3200 2592 3206 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 8444 2604 8769 2632
rect 8444 2592 8450 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 9490 2632 9496 2644
rect 9171 2604 9496 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 12802 2632 12808 2644
rect 11747 2604 12808 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13078 2592 13084 2644
rect 13136 2592 13142 2644
rect 14366 2592 14372 2644
rect 14424 2592 14430 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 16945 2635 17003 2641
rect 16945 2632 16957 2635
rect 16632 2604 16957 2632
rect 16632 2592 16638 2604
rect 16945 2601 16957 2604
rect 16991 2601 17003 2635
rect 16945 2595 17003 2601
rect 18506 2592 18512 2644
rect 18564 2592 18570 2644
rect 19150 2592 19156 2644
rect 19208 2632 19214 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 19208 2604 19257 2632
rect 19208 2592 19214 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19245 2595 19303 2601
rect 20165 2635 20223 2641
rect 20165 2601 20177 2635
rect 20211 2632 20223 2635
rect 20438 2632 20444 2644
rect 20211 2604 20444 2632
rect 20211 2601 20223 2604
rect 20165 2595 20223 2601
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 22646 2592 22652 2644
rect 22704 2632 22710 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 22704 2604 23305 2632
rect 22704 2592 22710 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 23293 2595 23351 2601
rect 24210 2592 24216 2644
rect 24268 2592 24274 2644
rect 25222 2592 25228 2644
rect 25280 2632 25286 2644
rect 25869 2635 25927 2641
rect 25869 2632 25881 2635
rect 25280 2604 25881 2632
rect 25280 2592 25286 2604
rect 25869 2601 25881 2604
rect 25915 2601 25927 2635
rect 25869 2595 25927 2601
rect 26602 2592 26608 2644
rect 26660 2592 26666 2644
rect 29089 2635 29147 2641
rect 29089 2601 29101 2635
rect 29135 2632 29147 2635
rect 29362 2632 29368 2644
rect 29135 2604 29368 2632
rect 29135 2601 29147 2604
rect 29089 2595 29147 2601
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 29822 2592 29828 2644
rect 29880 2592 29886 2644
rect 30374 2592 30380 2644
rect 30432 2632 30438 2644
rect 31021 2635 31079 2641
rect 31021 2632 31033 2635
rect 30432 2604 31033 2632
rect 30432 2592 30438 2604
rect 31021 2601 31033 2604
rect 31067 2601 31079 2635
rect 31021 2595 31079 2601
rect 33134 2592 33140 2644
rect 33192 2632 33198 2644
rect 33597 2635 33655 2641
rect 33597 2632 33609 2635
rect 33192 2604 33609 2632
rect 33192 2592 33198 2604
rect 33597 2601 33609 2604
rect 33643 2601 33655 2635
rect 33597 2595 33655 2601
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 34333 2635 34391 2641
rect 34333 2632 34345 2635
rect 33744 2604 34345 2632
rect 33744 2592 33750 2604
rect 34333 2601 34345 2604
rect 34379 2601 34391 2635
rect 34333 2595 34391 2601
rect 35526 2592 35532 2644
rect 35584 2592 35590 2644
rect 36078 2592 36084 2644
rect 36136 2632 36142 2644
rect 36173 2635 36231 2641
rect 36173 2632 36185 2635
rect 36136 2604 36185 2632
rect 36136 2592 36142 2604
rect 36173 2601 36185 2604
rect 36219 2601 36231 2635
rect 36173 2595 36231 2601
rect 36906 2592 36912 2644
rect 36964 2592 36970 2644
rect 37277 2635 37335 2641
rect 37277 2601 37289 2635
rect 37323 2632 37335 2635
rect 37642 2632 37648 2644
rect 37323 2604 37648 2632
rect 37323 2601 37335 2604
rect 37277 2595 37335 2601
rect 37642 2592 37648 2604
rect 37700 2592 37706 2644
rect 38010 2592 38016 2644
rect 38068 2592 38074 2644
rect 2884 2564 2912 2592
rect 4065 2567 4123 2573
rect 4065 2564 4077 2567
rect 2884 2536 4077 2564
rect 4065 2533 4077 2536
rect 4111 2533 4123 2567
rect 4065 2527 4123 2533
rect 6549 2567 6607 2573
rect 6549 2533 6561 2567
rect 6595 2564 6607 2567
rect 12066 2564 12072 2576
rect 6595 2536 8294 2564
rect 6595 2533 6607 2536
rect 6549 2527 6607 2533
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1452 2468 1961 2496
rect 1452 2456 1458 2468
rect 1949 2465 1961 2468
rect 1995 2465 2007 2499
rect 5626 2496 5632 2508
rect 1949 2459 2007 2465
rect 3988 2468 5632 2496
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3988 2437 4016 2468
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6880 2468 7113 2496
rect 6880 2456 6886 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3292 2400 3525 2428
rect 3292 2388 3298 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5592 2400 6009 2428
rect 5592 2388 5598 2400
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 7650 2388 7656 2440
rect 7708 2428 7714 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7708 2400 8125 2428
rect 7708 2388 7714 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 5074 2320 5080 2372
rect 5132 2320 5138 2372
rect 8266 2360 8294 2536
rect 8956 2536 12072 2564
rect 8956 2437 8984 2536
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 13096 2564 13124 2592
rect 12483 2536 13124 2564
rect 16853 2567 16911 2573
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 18524 2564 18552 2592
rect 16899 2536 18552 2564
rect 19797 2567 19855 2573
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 19797 2533 19809 2567
rect 19843 2564 19855 2567
rect 23934 2564 23940 2576
rect 19843 2536 23940 2564
rect 19843 2533 19855 2536
rect 19797 2527 19855 2533
rect 23934 2524 23940 2536
rect 23992 2524 23998 2576
rect 29840 2564 29868 2592
rect 31757 2567 31815 2573
rect 31757 2564 31769 2567
rect 29840 2536 31769 2564
rect 31757 2533 31769 2536
rect 31803 2533 31815 2567
rect 35544 2564 35572 2592
rect 31757 2527 31815 2533
rect 33980 2536 35572 2564
rect 9766 2496 9772 2508
rect 9048 2468 9772 2496
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9048 2360 9076 2468
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10594 2456 10600 2508
rect 10652 2456 10658 2508
rect 12986 2456 12992 2508
rect 13044 2456 13050 2508
rect 17310 2496 17316 2508
rect 14108 2468 17316 2496
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 8266 2332 9076 2360
rect 9324 2292 9352 2391
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12342 2428 12348 2440
rect 12115 2400 12348 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 9861 2363 9919 2369
rect 9861 2329 9873 2363
rect 9907 2360 9919 2363
rect 11532 2360 11560 2391
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 14108 2437 14136 2468
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 18322 2456 18328 2508
rect 18380 2456 18386 2508
rect 19242 2456 19248 2508
rect 19300 2456 19306 2508
rect 20714 2456 20720 2508
rect 20772 2456 20778 2508
rect 23382 2456 23388 2508
rect 23440 2496 23446 2508
rect 23845 2499 23903 2505
rect 23845 2496 23857 2499
rect 23440 2468 23857 2496
rect 23440 2456 23446 2468
rect 23845 2465 23857 2468
rect 23891 2465 23903 2499
rect 23845 2459 23903 2465
rect 26142 2456 26148 2508
rect 26200 2496 26206 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26200 2468 27629 2496
rect 26200 2456 26206 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 29362 2456 29368 2508
rect 29420 2496 29426 2508
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 29420 2468 30021 2496
rect 29420 2456 29426 2468
rect 30009 2465 30021 2468
rect 30055 2465 30067 2499
rect 30009 2459 30067 2465
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 9907 2332 11560 2360
rect 15028 2360 15056 2391
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 15746 2360 15752 2372
rect 15028 2332 15752 2360
rect 9907 2329 9919 2332
rect 9861 2323 9919 2329
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 16114 2320 16120 2372
rect 16172 2320 16178 2372
rect 16684 2360 16712 2391
rect 16850 2388 16856 2440
rect 16908 2428 16914 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 16908 2400 17509 2428
rect 16908 2388 16914 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 18874 2388 18880 2440
rect 18932 2388 18938 2440
rect 18690 2360 18696 2372
rect 16684 2332 18696 2360
rect 18690 2320 18696 2332
rect 18748 2320 18754 2372
rect 11146 2292 11152 2304
rect 9324 2264 11152 2292
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 19260 2292 19288 2456
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23474 2428 23480 2440
rect 23247 2400 23480 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 24026 2388 24032 2440
rect 24084 2388 24090 2440
rect 25498 2388 25504 2440
rect 25556 2428 25562 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25556 2400 25605 2428
rect 25556 2388 25562 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26418 2388 26424 2440
rect 26476 2388 26482 2440
rect 26510 2388 26516 2440
rect 26568 2428 26574 2440
rect 26789 2431 26847 2437
rect 26789 2428 26801 2431
rect 26568 2400 26801 2428
rect 26568 2388 26574 2400
rect 26789 2397 26801 2400
rect 26835 2397 26847 2431
rect 26789 2391 26847 2397
rect 26973 2431 27031 2437
rect 26973 2397 26985 2431
rect 27019 2428 27031 2431
rect 27246 2428 27252 2440
rect 27019 2400 27252 2428
rect 27019 2397 27031 2400
rect 26973 2391 27031 2397
rect 27246 2388 27252 2400
rect 27304 2388 27310 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 27632 2400 28457 2428
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 22097 2363 22155 2369
rect 22097 2360 22109 2363
rect 21968 2332 22109 2360
rect 21968 2320 21974 2332
rect 22097 2329 22109 2332
rect 22143 2329 22155 2363
rect 22097 2323 22155 2329
rect 24118 2320 24124 2372
rect 24176 2360 24182 2372
rect 24581 2363 24639 2369
rect 24581 2360 24593 2363
rect 24176 2332 24593 2360
rect 24176 2320 24182 2332
rect 24581 2329 24593 2332
rect 24627 2329 24639 2363
rect 24581 2323 24639 2329
rect 24762 2320 24768 2372
rect 24820 2360 24826 2372
rect 27632 2360 27660 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 29178 2388 29184 2440
rect 29236 2388 29242 2440
rect 29730 2388 29736 2440
rect 29788 2388 29794 2440
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2397 31631 2431
rect 31573 2391 31631 2397
rect 24820 2332 27660 2360
rect 24820 2320 24826 2332
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 31588 2360 31616 2391
rect 31938 2388 31944 2440
rect 31996 2388 32002 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 33980 2428 34008 2536
rect 34054 2456 34060 2508
rect 34112 2496 34118 2508
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 34112 2468 35173 2496
rect 34112 2456 34118 2468
rect 35161 2465 35173 2468
rect 35207 2465 35219 2499
rect 35161 2459 35219 2465
rect 35802 2456 35808 2508
rect 35860 2496 35866 2508
rect 36725 2499 36783 2505
rect 36725 2496 36737 2499
rect 35860 2468 36737 2496
rect 35860 2456 35866 2468
rect 36725 2465 36737 2468
rect 36771 2465 36783 2499
rect 36725 2459 36783 2465
rect 37826 2456 37832 2508
rect 37884 2456 37890 2508
rect 38470 2496 38476 2508
rect 38212 2468 38476 2496
rect 33551 2400 34008 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 34146 2388 34152 2440
rect 34204 2388 34210 2440
rect 34514 2388 34520 2440
rect 34572 2388 34578 2440
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 38212 2437 38240 2468
rect 38470 2456 38476 2468
rect 38528 2456 38534 2508
rect 38654 2456 38660 2508
rect 38712 2456 38718 2508
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34664 2400 34713 2428
rect 34664 2388 34670 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 37093 2431 37151 2437
rect 37093 2428 37105 2431
rect 34701 2391 34759 2397
rect 35866 2400 37105 2428
rect 29052 2332 31616 2360
rect 29052 2320 29058 2332
rect 31662 2320 31668 2372
rect 31720 2360 31726 2372
rect 32309 2363 32367 2369
rect 32309 2360 32321 2363
rect 31720 2332 32321 2360
rect 31720 2320 31726 2332
rect 32309 2329 32321 2332
rect 32355 2329 32367 2363
rect 32309 2323 32367 2329
rect 34422 2320 34428 2372
rect 34480 2360 34486 2372
rect 35866 2360 35894 2400
rect 37093 2397 37105 2400
rect 37139 2397 37151 2431
rect 37093 2391 37151 2397
rect 38197 2431 38255 2437
rect 38197 2397 38209 2431
rect 38243 2397 38255 2431
rect 38197 2391 38255 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2428 38439 2431
rect 38672 2428 38700 2456
rect 38427 2400 38700 2428
rect 38427 2397 38439 2400
rect 38381 2391 38439 2397
rect 34480 2332 35894 2360
rect 34480 2320 34486 2332
rect 14323 2264 19288 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 29270 2252 29276 2304
rect 29328 2292 29334 2304
rect 29365 2295 29423 2301
rect 29365 2292 29377 2295
rect 29328 2264 29377 2292
rect 29328 2252 29334 2264
rect 29365 2261 29377 2264
rect 29411 2261 29423 2295
rect 29365 2255 29423 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 6362 2048 6368 2100
rect 6420 2088 6426 2100
rect 9858 2088 9864 2100
rect 6420 2060 9864 2088
rect 6420 2048 6426 2060
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 33594 1708 33600 1760
rect 33652 1748 33658 1760
rect 39298 1748 39304 1760
rect 33652 1720 39304 1748
rect 33652 1708 33658 1720
rect 39298 1708 39304 1720
rect 39356 1708 39362 1760
rect 11514 1504 11520 1556
rect 11572 1544 11578 1556
rect 16482 1544 16488 1556
rect 11572 1516 16488 1544
rect 11572 1504 11578 1516
rect 16482 1504 16488 1516
rect 16540 1504 16546 1556
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 37372 32376 37424 32428
rect 14096 32351 14148 32360
rect 14096 32317 14105 32351
rect 14105 32317 14139 32351
rect 14139 32317 14148 32351
rect 14096 32308 14148 32317
rect 15016 32308 15068 32360
rect 24584 32351 24636 32360
rect 24584 32317 24593 32351
rect 24593 32317 24627 32351
rect 24627 32317 24636 32351
rect 24584 32308 24636 32317
rect 23940 32240 23992 32292
rect 28448 32308 28500 32360
rect 28816 32351 28868 32360
rect 28816 32317 28825 32351
rect 28825 32317 28859 32351
rect 28859 32317 28868 32351
rect 28816 32308 28868 32317
rect 36636 32308 36688 32360
rect 10048 32172 10100 32224
rect 13452 32215 13504 32224
rect 13452 32181 13461 32215
rect 13461 32181 13495 32215
rect 13495 32181 13504 32215
rect 13452 32172 13504 32181
rect 14280 32215 14332 32224
rect 14280 32181 14289 32215
rect 14289 32181 14323 32215
rect 14323 32181 14332 32215
rect 14280 32172 14332 32181
rect 24032 32215 24084 32224
rect 24032 32181 24041 32215
rect 24041 32181 24075 32215
rect 24075 32181 24084 32215
rect 24032 32172 24084 32181
rect 25412 32215 25464 32224
rect 25412 32181 25421 32215
rect 25421 32181 25455 32215
rect 25455 32181 25464 32215
rect 25412 32172 25464 32181
rect 26608 32172 26660 32224
rect 27068 32172 27120 32224
rect 27528 32215 27580 32224
rect 27528 32181 27537 32215
rect 27537 32181 27571 32215
rect 27571 32181 27580 32215
rect 27528 32172 27580 32181
rect 28264 32215 28316 32224
rect 28264 32181 28273 32215
rect 28273 32181 28307 32215
rect 28307 32181 28316 32215
rect 28264 32172 28316 32181
rect 36360 32215 36412 32224
rect 36360 32181 36369 32215
rect 36369 32181 36403 32215
rect 36403 32181 36412 32215
rect 36360 32172 36412 32181
rect 37740 32172 37792 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 14096 32011 14148 32020
rect 14096 31977 14105 32011
rect 14105 31977 14139 32011
rect 14139 31977 14148 32011
rect 14096 31968 14148 31977
rect 14280 31968 14332 32020
rect 23940 32011 23992 32020
rect 23940 31977 23949 32011
rect 23949 31977 23983 32011
rect 23983 31977 23992 32011
rect 23940 31968 23992 31977
rect 24032 31968 24084 32020
rect 28264 31968 28316 32020
rect 28448 32011 28500 32020
rect 28448 31977 28457 32011
rect 28457 31977 28491 32011
rect 28491 31977 28500 32011
rect 28448 31968 28500 31977
rect 10048 31900 10100 31952
rect 10416 31764 10468 31816
rect 11244 31807 11296 31816
rect 11244 31773 11253 31807
rect 11253 31773 11287 31807
rect 11287 31773 11296 31807
rect 11244 31764 11296 31773
rect 13912 31807 13964 31816
rect 13912 31773 13921 31807
rect 13921 31773 13955 31807
rect 13955 31773 13964 31807
rect 13912 31764 13964 31773
rect 15568 31807 15620 31816
rect 15568 31773 15577 31807
rect 15577 31773 15611 31807
rect 15611 31773 15620 31807
rect 15568 31764 15620 31773
rect 19064 31807 19116 31816
rect 19064 31773 19073 31807
rect 19073 31773 19107 31807
rect 19107 31773 19116 31807
rect 19064 31764 19116 31773
rect 19248 31764 19300 31816
rect 24768 31832 24820 31884
rect 26608 31832 26660 31884
rect 27068 31832 27120 31884
rect 14740 31696 14792 31748
rect 23940 31696 23992 31748
rect 25228 31764 25280 31816
rect 26332 31764 26384 31816
rect 34704 31832 34756 31884
rect 29184 31807 29236 31816
rect 29184 31773 29193 31807
rect 29193 31773 29227 31807
rect 29227 31773 29236 31807
rect 29184 31764 29236 31773
rect 31760 31764 31812 31816
rect 32036 31764 32088 31816
rect 35440 31764 35492 31816
rect 36452 31764 36504 31816
rect 36728 31807 36780 31816
rect 36728 31773 36737 31807
rect 36737 31773 36771 31807
rect 36771 31773 36780 31807
rect 36728 31764 36780 31773
rect 36912 31764 36964 31816
rect 37464 31807 37516 31816
rect 37464 31773 37473 31807
rect 37473 31773 37507 31807
rect 37507 31773 37516 31807
rect 37464 31764 37516 31773
rect 38108 31807 38160 31816
rect 38108 31773 38117 31807
rect 38117 31773 38151 31807
rect 38151 31773 38160 31807
rect 38108 31764 38160 31773
rect 29276 31696 29328 31748
rect 9680 31671 9732 31680
rect 9680 31637 9689 31671
rect 9689 31637 9723 31671
rect 9723 31637 9732 31671
rect 9680 31628 9732 31637
rect 10600 31671 10652 31680
rect 10600 31637 10609 31671
rect 10609 31637 10643 31671
rect 10643 31637 10652 31671
rect 10600 31628 10652 31637
rect 13268 31671 13320 31680
rect 13268 31637 13277 31671
rect 13277 31637 13311 31671
rect 13311 31637 13320 31671
rect 13268 31628 13320 31637
rect 13636 31628 13688 31680
rect 14648 31628 14700 31680
rect 18512 31628 18564 31680
rect 19340 31628 19392 31680
rect 20352 31671 20404 31680
rect 20352 31637 20361 31671
rect 20361 31637 20395 31671
rect 20395 31637 20404 31671
rect 20352 31628 20404 31637
rect 23664 31628 23716 31680
rect 24400 31671 24452 31680
rect 24400 31637 24409 31671
rect 24409 31637 24443 31671
rect 24443 31637 24452 31671
rect 24400 31628 24452 31637
rect 25136 31671 25188 31680
rect 25136 31637 25145 31671
rect 25145 31637 25179 31671
rect 25179 31637 25188 31671
rect 25136 31628 25188 31637
rect 28448 31628 28500 31680
rect 28540 31671 28592 31680
rect 28540 31637 28549 31671
rect 28549 31637 28583 31671
rect 28583 31637 28592 31671
rect 28540 31628 28592 31637
rect 29736 31671 29788 31680
rect 29736 31637 29745 31671
rect 29745 31637 29779 31671
rect 29779 31637 29788 31671
rect 29736 31628 29788 31637
rect 35348 31628 35400 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 9680 31424 9732 31476
rect 13268 31424 13320 31476
rect 16120 31424 16172 31476
rect 14740 31356 14792 31408
rect 11060 31288 11112 31340
rect 14096 31331 14148 31340
rect 14096 31297 14130 31331
rect 14130 31297 14148 31331
rect 14096 31288 14148 31297
rect 18512 31331 18564 31340
rect 18512 31297 18546 31331
rect 18546 31297 18564 31331
rect 18512 31288 18564 31297
rect 10048 31263 10100 31272
rect 10048 31229 10057 31263
rect 10057 31229 10091 31263
rect 10091 31229 10100 31263
rect 10048 31220 10100 31229
rect 10876 31263 10928 31272
rect 10876 31229 10885 31263
rect 10885 31229 10919 31263
rect 10919 31229 10928 31263
rect 10876 31220 10928 31229
rect 11520 31263 11572 31272
rect 11520 31229 11529 31263
rect 11529 31229 11563 31263
rect 11563 31229 11572 31263
rect 11520 31220 11572 31229
rect 13636 31263 13688 31272
rect 13636 31229 13645 31263
rect 13645 31229 13679 31263
rect 13679 31229 13688 31263
rect 13636 31220 13688 31229
rect 13728 31220 13780 31272
rect 15844 31263 15896 31272
rect 15844 31229 15853 31263
rect 15853 31229 15887 31263
rect 15887 31229 15896 31263
rect 15844 31220 15896 31229
rect 18236 31263 18288 31272
rect 18236 31229 18245 31263
rect 18245 31229 18279 31263
rect 18279 31229 18288 31263
rect 18236 31220 18288 31229
rect 19340 31424 19392 31476
rect 20352 31424 20404 31476
rect 23848 31424 23900 31476
rect 25136 31356 25188 31408
rect 22284 31288 22336 31340
rect 24768 31288 24820 31340
rect 28080 31424 28132 31476
rect 28816 31424 28868 31476
rect 29184 31467 29236 31476
rect 29184 31433 29193 31467
rect 29193 31433 29227 31467
rect 29227 31433 29236 31467
rect 29184 31424 29236 31433
rect 29276 31467 29328 31476
rect 29276 31433 29285 31467
rect 29285 31433 29319 31467
rect 29319 31433 29328 31467
rect 29276 31424 29328 31433
rect 19984 31263 20036 31272
rect 19984 31229 19993 31263
rect 19993 31229 20027 31263
rect 20027 31229 20036 31263
rect 19984 31220 20036 31229
rect 8760 31127 8812 31136
rect 8760 31093 8769 31127
rect 8769 31093 8803 31127
rect 8803 31093 8812 31127
rect 8760 31084 8812 31093
rect 10324 31127 10376 31136
rect 10324 31093 10333 31127
rect 10333 31093 10367 31127
rect 10367 31093 10376 31127
rect 10324 31084 10376 31093
rect 11336 31127 11388 31136
rect 11336 31093 11345 31127
rect 11345 31093 11379 31127
rect 11379 31093 11388 31127
rect 11336 31084 11388 31093
rect 12164 31127 12216 31136
rect 12164 31093 12173 31127
rect 12173 31093 12207 31127
rect 12207 31093 12216 31127
rect 12164 31084 12216 31093
rect 12900 31127 12952 31136
rect 12900 31093 12909 31127
rect 12909 31093 12943 31127
rect 12943 31093 12952 31127
rect 12900 31084 12952 31093
rect 15292 31127 15344 31136
rect 15292 31093 15301 31127
rect 15301 31093 15335 31127
rect 15335 31093 15344 31127
rect 15292 31084 15344 31093
rect 19156 31084 19208 31136
rect 19616 31127 19668 31136
rect 19616 31093 19625 31127
rect 19625 31093 19659 31127
rect 19659 31093 19668 31127
rect 19616 31084 19668 31093
rect 20536 31127 20588 31136
rect 20536 31093 20545 31127
rect 20545 31093 20579 31127
rect 20579 31093 20588 31127
rect 20536 31084 20588 31093
rect 21916 31084 21968 31136
rect 24676 31220 24728 31272
rect 26148 31288 26200 31340
rect 27528 31356 27580 31408
rect 33324 31356 33376 31408
rect 36360 31356 36412 31408
rect 28448 31288 28500 31340
rect 29460 31288 29512 31340
rect 24860 31152 24912 31204
rect 24952 31084 25004 31136
rect 25872 31127 25924 31136
rect 25872 31093 25881 31127
rect 25881 31093 25915 31127
rect 25915 31093 25924 31127
rect 25872 31084 25924 31093
rect 28632 31220 28684 31272
rect 29920 31220 29972 31272
rect 29736 31084 29788 31136
rect 31116 31084 31168 31136
rect 34152 31263 34204 31272
rect 34152 31229 34161 31263
rect 34161 31229 34195 31263
rect 34195 31229 34204 31263
rect 34152 31220 34204 31229
rect 33784 31152 33836 31204
rect 32312 31084 32364 31136
rect 34336 31127 34388 31136
rect 34336 31093 34345 31127
rect 34345 31093 34379 31127
rect 34379 31093 34388 31127
rect 34336 31084 34388 31093
rect 36820 31220 36872 31272
rect 35808 31084 35860 31136
rect 36176 31084 36228 31136
rect 36544 31127 36596 31136
rect 36544 31093 36553 31127
rect 36553 31093 36587 31127
rect 36587 31093 36596 31127
rect 36544 31084 36596 31093
rect 37924 31127 37976 31136
rect 37924 31093 37933 31127
rect 37933 31093 37967 31127
rect 37967 31093 37976 31127
rect 37924 31084 37976 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 10876 30880 10928 30932
rect 11520 30880 11572 30932
rect 15016 30880 15068 30932
rect 15568 30923 15620 30932
rect 15568 30889 15577 30923
rect 15577 30889 15611 30923
rect 15611 30889 15620 30923
rect 15568 30880 15620 30889
rect 19248 30923 19300 30932
rect 19248 30889 19257 30923
rect 19257 30889 19291 30923
rect 19291 30889 19300 30923
rect 19248 30880 19300 30889
rect 23756 30880 23808 30932
rect 23940 30880 23992 30932
rect 24584 30880 24636 30932
rect 15752 30812 15804 30864
rect 11336 30787 11388 30796
rect 11336 30753 11345 30787
rect 11345 30753 11379 30787
rect 11379 30753 11388 30787
rect 11336 30744 11388 30753
rect 9312 30719 9364 30728
rect 9312 30685 9321 30719
rect 9321 30685 9355 30719
rect 9355 30685 9364 30719
rect 9312 30676 9364 30685
rect 10600 30676 10652 30728
rect 11428 30676 11480 30728
rect 10140 30540 10192 30592
rect 11060 30540 11112 30592
rect 11704 30540 11756 30592
rect 13728 30744 13780 30796
rect 12624 30676 12676 30728
rect 14648 30676 14700 30728
rect 13452 30608 13504 30660
rect 14740 30608 14792 30660
rect 16120 30787 16172 30796
rect 16120 30753 16129 30787
rect 16129 30753 16163 30787
rect 16163 30753 16172 30787
rect 16120 30744 16172 30753
rect 19616 30744 19668 30796
rect 21916 30787 21968 30796
rect 21916 30753 21925 30787
rect 21925 30753 21959 30787
rect 21959 30753 21968 30787
rect 21916 30744 21968 30753
rect 26608 30880 26660 30932
rect 27988 30880 28040 30932
rect 28632 30880 28684 30932
rect 29000 30880 29052 30932
rect 29920 30880 29972 30932
rect 17224 30676 17276 30728
rect 18236 30676 18288 30728
rect 17960 30651 18012 30660
rect 17960 30617 17994 30651
rect 17994 30617 18012 30651
rect 17960 30608 18012 30617
rect 20536 30676 20588 30728
rect 22468 30676 22520 30728
rect 29460 30744 29512 30796
rect 24400 30676 24452 30728
rect 24952 30676 25004 30728
rect 26148 30676 26200 30728
rect 28540 30676 28592 30728
rect 33140 30880 33192 30932
rect 36452 30880 36504 30932
rect 37924 30880 37976 30932
rect 33968 30744 34020 30796
rect 16120 30540 16172 30592
rect 16580 30540 16632 30592
rect 23572 30608 23624 30660
rect 25412 30608 25464 30660
rect 26332 30608 26384 30660
rect 31024 30676 31076 30728
rect 32312 30676 32364 30728
rect 35808 30676 35860 30728
rect 30472 30608 30524 30660
rect 31300 30608 31352 30660
rect 33232 30608 33284 30660
rect 35348 30608 35400 30660
rect 36912 30608 36964 30660
rect 19340 30540 19392 30592
rect 19432 30540 19484 30592
rect 20720 30583 20772 30592
rect 20720 30549 20729 30583
rect 20729 30549 20763 30583
rect 20763 30549 20772 30583
rect 20720 30540 20772 30549
rect 23664 30583 23716 30592
rect 23664 30549 23673 30583
rect 23673 30549 23707 30583
rect 23707 30549 23716 30583
rect 23664 30540 23716 30549
rect 24124 30583 24176 30592
rect 24124 30549 24133 30583
rect 24133 30549 24167 30583
rect 24167 30549 24176 30583
rect 24124 30540 24176 30549
rect 29368 30540 29420 30592
rect 29552 30583 29604 30592
rect 29552 30549 29561 30583
rect 29561 30549 29595 30583
rect 29595 30549 29604 30583
rect 29552 30540 29604 30549
rect 33048 30540 33100 30592
rect 33876 30583 33928 30592
rect 33876 30549 33885 30583
rect 33885 30549 33919 30583
rect 33919 30549 33928 30583
rect 33876 30540 33928 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 8760 30268 8812 30320
rect 11428 30336 11480 30388
rect 12164 30336 12216 30388
rect 13912 30336 13964 30388
rect 14924 30336 14976 30388
rect 16120 30336 16172 30388
rect 12900 30311 12952 30320
rect 12900 30277 12934 30311
rect 12934 30277 12952 30311
rect 12900 30268 12952 30277
rect 10416 30243 10468 30252
rect 10416 30209 10425 30243
rect 10425 30209 10459 30243
rect 10459 30209 10468 30243
rect 10416 30200 10468 30209
rect 11152 30243 11204 30252
rect 11152 30209 11161 30243
rect 11161 30209 11195 30243
rect 11195 30209 11204 30243
rect 11152 30200 11204 30209
rect 11520 30200 11572 30252
rect 11612 30200 11664 30252
rect 12624 30243 12676 30252
rect 12624 30209 12633 30243
rect 12633 30209 12667 30243
rect 12667 30209 12676 30243
rect 12624 30200 12676 30209
rect 14924 30243 14976 30252
rect 14924 30209 14942 30243
rect 14942 30209 14976 30243
rect 14924 30200 14976 30209
rect 15016 30243 15068 30252
rect 15016 30209 15025 30243
rect 15025 30209 15059 30243
rect 15059 30209 15068 30243
rect 15016 30200 15068 30209
rect 15752 30243 15804 30252
rect 15752 30209 15761 30243
rect 15761 30209 15795 30243
rect 15795 30209 15804 30243
rect 15752 30200 15804 30209
rect 15844 30200 15896 30252
rect 17224 30200 17276 30252
rect 17408 30243 17460 30252
rect 17408 30209 17442 30243
rect 17442 30209 17460 30243
rect 17408 30200 17460 30209
rect 19248 30336 19300 30388
rect 19340 30336 19392 30388
rect 19800 30243 19852 30252
rect 19800 30209 19809 30243
rect 19809 30209 19843 30243
rect 19843 30209 19852 30243
rect 19800 30200 19852 30209
rect 22284 30336 22336 30388
rect 24584 30336 24636 30388
rect 24952 30336 25004 30388
rect 30472 30379 30524 30388
rect 30472 30345 30481 30379
rect 30481 30345 30515 30379
rect 30515 30345 30524 30379
rect 30472 30336 30524 30345
rect 31024 30336 31076 30388
rect 32312 30336 32364 30388
rect 33324 30336 33376 30388
rect 33600 30336 33652 30388
rect 34428 30336 34480 30388
rect 36912 30336 36964 30388
rect 23756 30243 23808 30252
rect 23756 30209 23774 30243
rect 23774 30209 23808 30243
rect 23756 30200 23808 30209
rect 23848 30243 23900 30252
rect 23848 30209 23857 30243
rect 23857 30209 23891 30243
rect 23891 30209 23900 30243
rect 23848 30200 23900 30209
rect 24860 30200 24912 30252
rect 26424 30200 26476 30252
rect 27804 30243 27856 30252
rect 27804 30209 27813 30243
rect 27813 30209 27847 30243
rect 27847 30209 27856 30243
rect 27804 30200 27856 30209
rect 27988 30243 28040 30252
rect 27988 30209 28006 30243
rect 28006 30209 28040 30243
rect 27988 30200 28040 30209
rect 28080 30243 28132 30252
rect 28080 30209 28089 30243
rect 28089 30209 28123 30243
rect 28123 30209 28132 30243
rect 28080 30200 28132 30209
rect 28816 30243 28868 30252
rect 28816 30209 28825 30243
rect 28825 30209 28859 30243
rect 28859 30209 28868 30243
rect 28816 30200 28868 30209
rect 7840 30132 7892 30184
rect 10140 30175 10192 30184
rect 10140 30141 10149 30175
rect 10149 30141 10183 30175
rect 10183 30141 10192 30175
rect 10140 30132 10192 30141
rect 10600 30132 10652 30184
rect 11244 30132 11296 30184
rect 9496 30039 9548 30048
rect 9496 30005 9505 30039
rect 9505 30005 9539 30039
rect 9539 30005 9548 30039
rect 9496 29996 9548 30005
rect 10784 30064 10836 30116
rect 10416 29996 10468 30048
rect 14556 30132 14608 30184
rect 19156 30132 19208 30184
rect 19340 30132 19392 30184
rect 19616 30175 19668 30184
rect 19616 30141 19650 30175
rect 19650 30141 19668 30175
rect 19616 30132 19668 30141
rect 22744 30175 22796 30184
rect 22744 30141 22753 30175
rect 22753 30141 22787 30175
rect 22787 30141 22796 30175
rect 22744 30132 22796 30141
rect 15200 30064 15252 30116
rect 12900 29996 12952 30048
rect 16028 29996 16080 30048
rect 21088 30064 21140 30116
rect 19616 29996 19668 30048
rect 19708 29996 19760 30048
rect 23848 29996 23900 30048
rect 29000 30175 29052 30184
rect 29000 30141 29009 30175
rect 29009 30141 29043 30175
rect 29043 30141 29052 30175
rect 29000 30132 29052 30141
rect 29552 30200 29604 30252
rect 34704 30268 34756 30320
rect 30656 30200 30708 30252
rect 32956 30243 33008 30252
rect 32956 30209 32974 30243
rect 32974 30209 33008 30243
rect 32956 30200 33008 30209
rect 33048 30243 33100 30252
rect 33048 30209 33057 30243
rect 33057 30209 33091 30243
rect 33091 30209 33100 30243
rect 33048 30200 33100 30209
rect 33784 30243 33836 30252
rect 33784 30209 33793 30243
rect 33793 30209 33827 30243
rect 33827 30209 33836 30243
rect 33784 30200 33836 30209
rect 33968 30243 34020 30252
rect 33968 30209 33977 30243
rect 33977 30209 34011 30243
rect 34011 30209 34020 30243
rect 33968 30200 34020 30209
rect 36176 30243 36228 30252
rect 36176 30209 36185 30243
rect 36185 30209 36219 30243
rect 36219 30209 36228 30243
rect 36176 30200 36228 30209
rect 37740 30311 37792 30320
rect 37740 30277 37749 30311
rect 37749 30277 37783 30311
rect 37783 30277 37792 30311
rect 37740 30268 37792 30277
rect 37464 30200 37516 30252
rect 37648 30243 37700 30252
rect 37648 30209 37657 30243
rect 37657 30209 37691 30243
rect 37691 30209 37700 30243
rect 37648 30200 37700 30209
rect 32772 30175 32824 30184
rect 32772 30141 32781 30175
rect 32781 30141 32815 30175
rect 32815 30141 32824 30175
rect 32772 30132 32824 30141
rect 26240 30064 26292 30116
rect 33324 30107 33376 30116
rect 33324 30073 33333 30107
rect 33333 30073 33367 30107
rect 33367 30073 33376 30107
rect 33324 30064 33376 30073
rect 34612 30175 34664 30184
rect 34612 30141 34621 30175
rect 34621 30141 34655 30175
rect 34655 30141 34664 30175
rect 34612 30132 34664 30141
rect 34704 30175 34756 30184
rect 34704 30141 34713 30175
rect 34713 30141 34747 30175
rect 34747 30141 34756 30175
rect 34704 30132 34756 30141
rect 36360 30132 36412 30184
rect 37832 30175 37884 30184
rect 37832 30141 37841 30175
rect 37841 30141 37875 30175
rect 37875 30141 37884 30175
rect 37832 30132 37884 30141
rect 34796 30064 34848 30116
rect 35440 30064 35492 30116
rect 24584 29996 24636 30048
rect 27988 29996 28040 30048
rect 29092 30039 29144 30048
rect 29092 30005 29101 30039
rect 29101 30005 29135 30039
rect 29135 30005 29144 30039
rect 29092 29996 29144 30005
rect 32036 29996 32088 30048
rect 33416 29996 33468 30048
rect 35716 29996 35768 30048
rect 35900 29996 35952 30048
rect 37372 30064 37424 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 9496 29792 9548 29844
rect 11152 29792 11204 29844
rect 14556 29792 14608 29844
rect 16580 29792 16632 29844
rect 17408 29792 17460 29844
rect 19064 29792 19116 29844
rect 22744 29835 22796 29844
rect 22744 29801 22753 29835
rect 22753 29801 22787 29835
rect 22787 29801 22796 29835
rect 22744 29792 22796 29801
rect 23572 29835 23624 29844
rect 23572 29801 23581 29835
rect 23581 29801 23615 29835
rect 23615 29801 23624 29835
rect 23572 29792 23624 29801
rect 25228 29792 25280 29844
rect 28816 29792 28868 29844
rect 29092 29792 29144 29844
rect 30656 29835 30708 29844
rect 30656 29801 30665 29835
rect 30665 29801 30699 29835
rect 30699 29801 30708 29835
rect 30656 29792 30708 29801
rect 32036 29792 32088 29844
rect 32956 29792 33008 29844
rect 33232 29792 33284 29844
rect 34152 29792 34204 29844
rect 11244 29724 11296 29776
rect 6000 29631 6052 29640
rect 6000 29597 6009 29631
rect 6009 29597 6043 29631
rect 6043 29597 6052 29631
rect 6000 29588 6052 29597
rect 6368 29588 6420 29640
rect 8760 29588 8812 29640
rect 9312 29588 9364 29640
rect 10324 29588 10376 29640
rect 11796 29656 11848 29708
rect 12900 29699 12952 29708
rect 12900 29665 12909 29699
rect 12909 29665 12943 29699
rect 12943 29665 12952 29699
rect 12900 29656 12952 29665
rect 13360 29656 13412 29708
rect 15292 29656 15344 29708
rect 13728 29588 13780 29640
rect 18144 29631 18196 29640
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 18880 29699 18932 29708
rect 18880 29665 18889 29699
rect 18889 29665 18923 29699
rect 18923 29665 18932 29699
rect 18880 29656 18932 29665
rect 27068 29724 27120 29776
rect 20720 29656 20772 29708
rect 23940 29656 23992 29708
rect 24124 29699 24176 29708
rect 24124 29665 24133 29699
rect 24133 29665 24167 29699
rect 24167 29665 24176 29699
rect 24124 29656 24176 29665
rect 24676 29656 24728 29708
rect 24768 29656 24820 29708
rect 26148 29656 26200 29708
rect 26976 29656 27028 29708
rect 19616 29588 19668 29640
rect 25872 29588 25924 29640
rect 16856 29520 16908 29572
rect 18880 29520 18932 29572
rect 19800 29520 19852 29572
rect 20076 29520 20128 29572
rect 23664 29520 23716 29572
rect 31760 29631 31812 29640
rect 31760 29597 31769 29631
rect 31769 29597 31803 29631
rect 31803 29597 31812 29631
rect 31760 29588 31812 29597
rect 32772 29699 32824 29708
rect 32772 29665 32781 29699
rect 32781 29665 32815 29699
rect 32815 29665 32824 29699
rect 32772 29656 32824 29665
rect 33140 29699 33192 29708
rect 33140 29665 33149 29699
rect 33149 29665 33183 29699
rect 33183 29665 33192 29699
rect 33140 29656 33192 29665
rect 37464 29792 37516 29844
rect 37280 29656 37332 29708
rect 34336 29588 34388 29640
rect 34428 29631 34480 29640
rect 34428 29597 34437 29631
rect 34437 29597 34471 29631
rect 34471 29597 34480 29631
rect 34428 29588 34480 29597
rect 35808 29631 35860 29640
rect 35808 29597 35817 29631
rect 35817 29597 35851 29631
rect 35851 29597 35860 29631
rect 35808 29588 35860 29597
rect 36636 29588 36688 29640
rect 38108 29588 38160 29640
rect 5356 29495 5408 29504
rect 5356 29461 5365 29495
rect 5365 29461 5399 29495
rect 5399 29461 5408 29495
rect 5356 29452 5408 29461
rect 6184 29495 6236 29504
rect 6184 29461 6193 29495
rect 6193 29461 6227 29495
rect 6227 29461 6236 29495
rect 6184 29452 6236 29461
rect 8208 29452 8260 29504
rect 9864 29452 9916 29504
rect 10784 29452 10836 29504
rect 11060 29495 11112 29504
rect 11060 29461 11069 29495
rect 11069 29461 11103 29495
rect 11103 29461 11112 29495
rect 11060 29452 11112 29461
rect 11152 29452 11204 29504
rect 11336 29452 11388 29504
rect 11612 29452 11664 29504
rect 14740 29495 14792 29504
rect 14740 29461 14749 29495
rect 14749 29461 14783 29495
rect 14783 29461 14792 29495
rect 14740 29452 14792 29461
rect 15108 29495 15160 29504
rect 15108 29461 15117 29495
rect 15117 29461 15151 29495
rect 15151 29461 15160 29495
rect 15108 29452 15160 29461
rect 18328 29495 18380 29504
rect 18328 29461 18337 29495
rect 18337 29461 18371 29495
rect 18371 29461 18380 29495
rect 18328 29452 18380 29461
rect 19340 29452 19392 29504
rect 19984 29452 20036 29504
rect 24124 29452 24176 29504
rect 24768 29452 24820 29504
rect 24952 29452 25004 29504
rect 26240 29452 26292 29504
rect 26424 29495 26476 29504
rect 26424 29461 26433 29495
rect 26433 29461 26467 29495
rect 26467 29461 26476 29495
rect 26424 29452 26476 29461
rect 32220 29495 32272 29504
rect 32220 29461 32229 29495
rect 32229 29461 32263 29495
rect 32263 29461 32272 29495
rect 32220 29452 32272 29461
rect 32588 29495 32640 29504
rect 32588 29461 32597 29495
rect 32597 29461 32631 29495
rect 32631 29461 32640 29495
rect 32588 29452 32640 29461
rect 32680 29495 32732 29504
rect 32680 29461 32689 29495
rect 32689 29461 32723 29495
rect 32723 29461 32732 29495
rect 32680 29452 32732 29461
rect 32956 29520 33008 29572
rect 34704 29520 34756 29572
rect 34612 29452 34664 29504
rect 36452 29452 36504 29504
rect 37648 29452 37700 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 6184 29248 6236 29300
rect 10600 29248 10652 29300
rect 11796 29248 11848 29300
rect 5080 29180 5132 29232
rect 5816 29155 5868 29164
rect 5816 29121 5825 29155
rect 5825 29121 5859 29155
rect 5859 29121 5868 29155
rect 5816 29112 5868 29121
rect 12624 29248 12676 29300
rect 14096 29248 14148 29300
rect 17960 29248 18012 29300
rect 18144 29248 18196 29300
rect 18328 29248 18380 29300
rect 19340 29248 19392 29300
rect 19432 29248 19484 29300
rect 31300 29291 31352 29300
rect 31300 29257 31309 29291
rect 31309 29257 31343 29291
rect 31343 29257 31352 29291
rect 31300 29248 31352 29257
rect 32220 29248 32272 29300
rect 32680 29248 32732 29300
rect 33876 29248 33928 29300
rect 34428 29248 34480 29300
rect 34520 29248 34572 29300
rect 13728 29180 13780 29232
rect 11060 29112 11112 29164
rect 15200 29112 15252 29164
rect 6460 29044 6512 29096
rect 8760 29087 8812 29096
rect 8760 29053 8769 29087
rect 8769 29053 8803 29087
rect 8803 29053 8812 29087
rect 8760 29044 8812 29053
rect 15108 29044 15160 29096
rect 32588 29112 32640 29164
rect 32956 29112 33008 29164
rect 33048 29112 33100 29164
rect 32220 29087 32272 29096
rect 7932 28976 7984 29028
rect 4620 28951 4672 28960
rect 4620 28917 4629 28951
rect 4629 28917 4663 28951
rect 4663 28917 4672 28951
rect 4620 28908 4672 28917
rect 4712 28951 4764 28960
rect 4712 28917 4721 28951
rect 4721 28917 4755 28951
rect 4755 28917 4764 28951
rect 4712 28908 4764 28917
rect 8024 28908 8076 28960
rect 32220 29053 32229 29087
rect 32229 29053 32263 29087
rect 32263 29053 32272 29087
rect 32220 29044 32272 29053
rect 33140 29044 33192 29096
rect 23940 28976 23992 29028
rect 24584 28976 24636 29028
rect 27804 28976 27856 29028
rect 28540 28976 28592 29028
rect 30748 29019 30800 29028
rect 30748 28985 30757 29019
rect 30757 28985 30791 29019
rect 30791 28985 30800 29019
rect 30748 28976 30800 28985
rect 13820 28908 13872 28960
rect 31116 29019 31168 29028
rect 31116 28985 31125 29019
rect 31125 28985 31159 29019
rect 31159 28985 31168 29019
rect 31116 28976 31168 28985
rect 32772 28976 32824 29028
rect 34796 29180 34848 29232
rect 36728 29248 36780 29300
rect 36820 29291 36872 29300
rect 36820 29257 36829 29291
rect 36829 29257 36863 29291
rect 36863 29257 36872 29291
rect 36820 29248 36872 29257
rect 35900 29180 35952 29232
rect 36084 29112 36136 29164
rect 36452 29155 36504 29164
rect 36452 29121 36461 29155
rect 36461 29121 36495 29155
rect 36495 29121 36504 29155
rect 36452 29112 36504 29121
rect 35900 29019 35952 29028
rect 35900 28985 35909 29019
rect 35909 28985 35943 29019
rect 35943 28985 35952 29019
rect 37648 29044 37700 29096
rect 35900 28976 35952 28985
rect 36268 28976 36320 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 10784 28704 10836 28756
rect 15016 28704 15068 28756
rect 3792 28543 3844 28552
rect 3792 28509 3801 28543
rect 3801 28509 3835 28543
rect 3835 28509 3844 28543
rect 3792 28500 3844 28509
rect 4712 28500 4764 28552
rect 6184 28500 6236 28552
rect 5448 28432 5500 28484
rect 7196 28543 7248 28552
rect 7196 28509 7205 28543
rect 7205 28509 7239 28543
rect 7239 28509 7248 28543
rect 7196 28500 7248 28509
rect 9772 28543 9824 28552
rect 9772 28509 9781 28543
rect 9781 28509 9815 28543
rect 9815 28509 9824 28543
rect 9772 28500 9824 28509
rect 9956 28500 10008 28552
rect 14464 28543 14516 28552
rect 14464 28509 14473 28543
rect 14473 28509 14507 28543
rect 14507 28509 14516 28543
rect 14464 28500 14516 28509
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 19432 28500 19484 28552
rect 23572 28500 23624 28552
rect 23664 28500 23716 28552
rect 25044 28543 25096 28552
rect 25044 28509 25053 28543
rect 25053 28509 25087 28543
rect 25087 28509 25096 28543
rect 25044 28500 25096 28509
rect 27344 28543 27396 28552
rect 27344 28509 27353 28543
rect 27353 28509 27387 28543
rect 27387 28509 27396 28543
rect 27344 28500 27396 28509
rect 27436 28500 27488 28552
rect 28356 28500 28408 28552
rect 33140 28500 33192 28552
rect 34244 28543 34296 28552
rect 34244 28509 34253 28543
rect 34253 28509 34287 28543
rect 34287 28509 34296 28543
rect 34244 28500 34296 28509
rect 37924 28543 37976 28552
rect 37924 28509 37933 28543
rect 37933 28509 37967 28543
rect 37967 28509 37976 28543
rect 37924 28500 37976 28509
rect 13820 28432 13872 28484
rect 14648 28432 14700 28484
rect 4620 28364 4672 28416
rect 4712 28407 4764 28416
rect 4712 28373 4721 28407
rect 4721 28373 4755 28407
rect 4755 28373 4764 28407
rect 4712 28364 4764 28373
rect 5540 28364 5592 28416
rect 6368 28407 6420 28416
rect 6368 28373 6377 28407
rect 6377 28373 6411 28407
rect 6411 28373 6420 28407
rect 6368 28364 6420 28373
rect 7104 28407 7156 28416
rect 7104 28373 7113 28407
rect 7113 28373 7147 28407
rect 7147 28373 7156 28407
rect 7104 28364 7156 28373
rect 7656 28364 7708 28416
rect 10416 28364 10468 28416
rect 10508 28407 10560 28416
rect 10508 28373 10517 28407
rect 10517 28373 10551 28407
rect 10551 28373 10560 28407
rect 10508 28364 10560 28373
rect 15016 28364 15068 28416
rect 15292 28364 15344 28416
rect 18512 28364 18564 28416
rect 18972 28407 19024 28416
rect 18972 28373 18981 28407
rect 18981 28373 19015 28407
rect 19015 28373 19024 28407
rect 18972 28364 19024 28373
rect 19340 28407 19392 28416
rect 19340 28373 19349 28407
rect 19349 28373 19383 28407
rect 19383 28373 19392 28407
rect 19340 28364 19392 28373
rect 22836 28407 22888 28416
rect 22836 28373 22845 28407
rect 22845 28373 22879 28407
rect 22879 28373 22888 28407
rect 22836 28364 22888 28373
rect 23756 28407 23808 28416
rect 23756 28373 23765 28407
rect 23765 28373 23799 28407
rect 23799 28373 23808 28407
rect 23756 28364 23808 28373
rect 26792 28407 26844 28416
rect 26792 28373 26801 28407
rect 26801 28373 26835 28407
rect 26835 28373 26844 28407
rect 26792 28364 26844 28373
rect 27528 28407 27580 28416
rect 27528 28373 27537 28407
rect 27537 28373 27571 28407
rect 27571 28373 27580 28407
rect 27528 28364 27580 28373
rect 28264 28407 28316 28416
rect 28264 28373 28273 28407
rect 28273 28373 28307 28407
rect 28307 28373 28316 28407
rect 28264 28364 28316 28373
rect 28632 28364 28684 28416
rect 31024 28407 31076 28416
rect 31024 28373 31033 28407
rect 31033 28373 31067 28407
rect 31067 28373 31076 28407
rect 31024 28364 31076 28373
rect 32404 28407 32456 28416
rect 32404 28373 32413 28407
rect 32413 28373 32447 28407
rect 32447 28373 32456 28407
rect 32404 28364 32456 28373
rect 32956 28407 33008 28416
rect 32956 28373 32965 28407
rect 32965 28373 32999 28407
rect 32999 28373 33008 28407
rect 32956 28364 33008 28373
rect 33692 28407 33744 28416
rect 33692 28373 33701 28407
rect 33701 28373 33735 28407
rect 33735 28373 33744 28407
rect 33692 28364 33744 28373
rect 36636 28364 36688 28416
rect 36912 28364 36964 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 5356 28160 5408 28212
rect 6000 28160 6052 28212
rect 7196 28160 7248 28212
rect 7656 28160 7708 28212
rect 8208 28160 8260 28212
rect 9772 28203 9824 28212
rect 9772 28169 9781 28203
rect 9781 28169 9815 28203
rect 9815 28169 9824 28203
rect 9772 28160 9824 28169
rect 10508 28160 10560 28212
rect 14464 28203 14516 28212
rect 14464 28169 14473 28203
rect 14473 28169 14507 28203
rect 14507 28169 14516 28203
rect 14464 28160 14516 28169
rect 15200 28160 15252 28212
rect 3700 28024 3752 28076
rect 5724 28092 5776 28144
rect 2780 27956 2832 28008
rect 3608 27999 3660 28008
rect 3608 27965 3617 27999
rect 3617 27965 3651 27999
rect 3651 27965 3660 27999
rect 3608 27956 3660 27965
rect 4528 27956 4580 28008
rect 6920 28024 6972 28076
rect 11336 28024 11388 28076
rect 14740 28092 14792 28144
rect 18236 28160 18288 28212
rect 19340 28160 19392 28212
rect 22744 28160 22796 28212
rect 19340 28067 19392 28076
rect 19340 28033 19349 28067
rect 19349 28033 19383 28067
rect 19383 28033 19392 28067
rect 19340 28024 19392 28033
rect 23664 28092 23716 28144
rect 27528 28160 27580 28212
rect 27988 28160 28040 28212
rect 32956 28160 33008 28212
rect 36268 28203 36320 28212
rect 36268 28169 36277 28203
rect 36277 28169 36311 28203
rect 36311 28169 36320 28203
rect 36268 28160 36320 28169
rect 37740 28092 37792 28144
rect 26976 28067 27028 28076
rect 26976 28033 26985 28067
rect 26985 28033 27019 28067
rect 27019 28033 27028 28067
rect 26976 28024 27028 28033
rect 28080 28024 28132 28076
rect 6184 27999 6236 28008
rect 6184 27965 6193 27999
rect 6193 27965 6227 27999
rect 6227 27965 6236 27999
rect 6184 27956 6236 27965
rect 8024 27956 8076 28008
rect 9680 27999 9732 28008
rect 9680 27965 9689 27999
rect 9689 27965 9723 27999
rect 9723 27965 9732 27999
rect 9680 27956 9732 27965
rect 10692 27956 10744 28008
rect 11060 27956 11112 28008
rect 11520 27999 11572 28008
rect 11520 27965 11529 27999
rect 11529 27965 11563 27999
rect 11563 27965 11572 27999
rect 11520 27956 11572 27965
rect 13820 27956 13872 28008
rect 14004 27956 14056 28008
rect 2964 27863 3016 27872
rect 2964 27829 2973 27863
rect 2973 27829 3007 27863
rect 3007 27829 3016 27863
rect 2964 27820 3016 27829
rect 3056 27863 3108 27872
rect 3056 27829 3065 27863
rect 3065 27829 3099 27863
rect 3099 27829 3108 27863
rect 3056 27820 3108 27829
rect 5448 27820 5500 27872
rect 9036 27863 9088 27872
rect 9036 27829 9045 27863
rect 9045 27829 9079 27863
rect 9079 27829 9088 27863
rect 9036 27820 9088 27829
rect 10600 27863 10652 27872
rect 10600 27829 10609 27863
rect 10609 27829 10643 27863
rect 10643 27829 10652 27863
rect 10600 27820 10652 27829
rect 12164 27863 12216 27872
rect 12164 27829 12173 27863
rect 12173 27829 12207 27863
rect 12207 27829 12216 27863
rect 12164 27820 12216 27829
rect 12532 27820 12584 27872
rect 12992 27863 13044 27872
rect 12992 27829 13001 27863
rect 13001 27829 13035 27863
rect 13035 27829 13044 27863
rect 12992 27820 13044 27829
rect 13544 27820 13596 27872
rect 14280 27820 14332 27872
rect 15016 27999 15068 28008
rect 15016 27965 15025 27999
rect 15025 27965 15059 27999
rect 15059 27965 15068 27999
rect 15016 27956 15068 27965
rect 15568 27956 15620 28008
rect 18144 27956 18196 28008
rect 18972 27956 19024 28008
rect 14924 27820 14976 27872
rect 20720 27863 20772 27872
rect 20720 27829 20729 27863
rect 20729 27829 20763 27863
rect 20763 27829 20772 27863
rect 20720 27820 20772 27829
rect 22376 27863 22428 27872
rect 22376 27829 22385 27863
rect 22385 27829 22419 27863
rect 22419 27829 22428 27863
rect 22376 27820 22428 27829
rect 23480 27820 23532 27872
rect 24492 27999 24544 28008
rect 24492 27965 24501 27999
rect 24501 27965 24535 27999
rect 24535 27965 24544 27999
rect 24492 27956 24544 27965
rect 26148 27956 26200 28008
rect 28632 27999 28684 28008
rect 28632 27965 28641 27999
rect 28641 27965 28675 27999
rect 28675 27965 28684 27999
rect 28632 27956 28684 27965
rect 29000 28024 29052 28076
rect 29184 28024 29236 28076
rect 32588 28024 32640 28076
rect 36084 28024 36136 28076
rect 24676 27888 24728 27940
rect 28356 27931 28408 27940
rect 28356 27897 28365 27931
rect 28365 27897 28399 27931
rect 28399 27897 28408 27931
rect 28356 27888 28408 27897
rect 28724 27888 28776 27940
rect 33232 27956 33284 28008
rect 33784 27999 33836 28008
rect 33784 27965 33793 27999
rect 33793 27965 33827 27999
rect 33827 27965 33836 27999
rect 33784 27956 33836 27965
rect 34520 27999 34572 28008
rect 34520 27965 34529 27999
rect 34529 27965 34563 27999
rect 34563 27965 34572 27999
rect 34520 27956 34572 27965
rect 35348 27956 35400 28008
rect 35900 27956 35952 28008
rect 24032 27820 24084 27872
rect 25320 27863 25372 27872
rect 25320 27829 25329 27863
rect 25329 27829 25363 27863
rect 25363 27829 25372 27863
rect 25320 27820 25372 27829
rect 26056 27863 26108 27872
rect 26056 27829 26065 27863
rect 26065 27829 26099 27863
rect 26099 27829 26108 27863
rect 26056 27820 26108 27829
rect 27712 27820 27764 27872
rect 29276 27863 29328 27872
rect 29276 27829 29285 27863
rect 29285 27829 29319 27863
rect 29319 27829 29328 27863
rect 29276 27820 29328 27829
rect 31392 27820 31444 27872
rect 32956 27863 33008 27872
rect 32956 27829 32965 27863
rect 32965 27829 32999 27863
rect 32999 27829 33008 27863
rect 32956 27820 33008 27829
rect 34336 27863 34388 27872
rect 34336 27829 34345 27863
rect 34345 27829 34379 27863
rect 34379 27829 34388 27863
rect 34336 27820 34388 27829
rect 35808 27863 35860 27872
rect 35808 27829 35817 27863
rect 35817 27829 35851 27863
rect 35851 27829 35860 27863
rect 35808 27820 35860 27829
rect 37372 27820 37424 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2780 27659 2832 27668
rect 2780 27625 2789 27659
rect 2789 27625 2823 27659
rect 2823 27625 2832 27659
rect 2780 27616 2832 27625
rect 4988 27548 5040 27600
rect 5264 27480 5316 27532
rect 5448 27480 5500 27532
rect 5908 27480 5960 27532
rect 6552 27480 6604 27532
rect 6920 27616 6972 27668
rect 9956 27616 10008 27668
rect 10876 27616 10928 27668
rect 12624 27616 12676 27668
rect 14740 27616 14792 27668
rect 18052 27616 18104 27668
rect 19432 27616 19484 27668
rect 23112 27616 23164 27668
rect 24032 27616 24084 27668
rect 24492 27616 24544 27668
rect 27344 27616 27396 27668
rect 29000 27659 29052 27668
rect 29000 27625 29009 27659
rect 29009 27625 29043 27659
rect 29043 27625 29052 27659
rect 29000 27616 29052 27625
rect 5080 27412 5132 27464
rect 5540 27412 5592 27464
rect 6092 27455 6144 27464
rect 6092 27421 6101 27455
rect 6101 27421 6135 27455
rect 6135 27421 6144 27455
rect 6092 27412 6144 27421
rect 6368 27455 6420 27464
rect 6368 27421 6377 27455
rect 6377 27421 6411 27455
rect 6411 27421 6420 27455
rect 6368 27412 6420 27421
rect 8392 27455 8444 27464
rect 8392 27421 8401 27455
rect 8401 27421 8435 27455
rect 8435 27421 8444 27455
rect 8392 27412 8444 27421
rect 10416 27455 10468 27464
rect 10416 27421 10434 27455
rect 10434 27421 10468 27455
rect 10416 27412 10468 27421
rect 9220 27387 9272 27396
rect 9220 27353 9229 27387
rect 9229 27353 9263 27387
rect 9263 27353 9272 27387
rect 11244 27523 11296 27532
rect 11244 27489 11253 27523
rect 11253 27489 11287 27523
rect 11287 27489 11296 27523
rect 11244 27480 11296 27489
rect 12256 27455 12308 27464
rect 12256 27421 12265 27455
rect 12265 27421 12299 27455
rect 12299 27421 12308 27455
rect 12256 27412 12308 27421
rect 12532 27412 12584 27464
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 16028 27523 16080 27532
rect 16028 27489 16037 27523
rect 16037 27489 16071 27523
rect 16071 27489 16080 27523
rect 16028 27480 16080 27489
rect 25688 27548 25740 27600
rect 9220 27344 9272 27353
rect 14004 27344 14056 27396
rect 15384 27344 15436 27396
rect 20720 27412 20772 27464
rect 21364 27455 21416 27464
rect 21364 27421 21373 27455
rect 21373 27421 21407 27455
rect 21407 27421 21416 27455
rect 21364 27412 21416 27421
rect 23756 27480 23808 27532
rect 23848 27480 23900 27532
rect 22100 27412 22152 27464
rect 22836 27412 22888 27464
rect 23296 27412 23348 27464
rect 25412 27412 25464 27464
rect 21272 27344 21324 27396
rect 2044 27276 2096 27328
rect 3700 27276 3752 27328
rect 7012 27319 7064 27328
rect 7012 27285 7021 27319
rect 7021 27285 7055 27319
rect 7055 27285 7064 27319
rect 7012 27276 7064 27285
rect 7656 27276 7708 27328
rect 9404 27276 9456 27328
rect 10416 27276 10468 27328
rect 10784 27319 10836 27328
rect 10784 27285 10793 27319
rect 10793 27285 10827 27319
rect 10827 27285 10836 27319
rect 10784 27276 10836 27285
rect 11152 27319 11204 27328
rect 11152 27285 11161 27319
rect 11161 27285 11195 27319
rect 11195 27285 11204 27319
rect 11152 27276 11204 27285
rect 11612 27319 11664 27328
rect 11612 27285 11621 27319
rect 11621 27285 11655 27319
rect 11655 27285 11664 27319
rect 11612 27276 11664 27285
rect 12716 27276 12768 27328
rect 12808 27276 12860 27328
rect 13912 27276 13964 27328
rect 15476 27276 15528 27328
rect 15844 27276 15896 27328
rect 15936 27319 15988 27328
rect 15936 27285 15945 27319
rect 15945 27285 15979 27319
rect 15979 27285 15988 27319
rect 15936 27276 15988 27285
rect 17684 27276 17736 27328
rect 18972 27276 19024 27328
rect 19340 27276 19392 27328
rect 21916 27319 21968 27328
rect 21916 27285 21925 27319
rect 21925 27285 21959 27319
rect 21959 27285 21968 27319
rect 21916 27276 21968 27285
rect 22284 27276 22336 27328
rect 23388 27319 23440 27328
rect 23388 27285 23397 27319
rect 23397 27285 23431 27319
rect 23431 27285 23440 27319
rect 23388 27276 23440 27285
rect 23756 27319 23808 27328
rect 23756 27285 23765 27319
rect 23765 27285 23799 27319
rect 23799 27285 23808 27319
rect 23756 27276 23808 27285
rect 24400 27319 24452 27328
rect 24400 27285 24409 27319
rect 24409 27285 24443 27319
rect 24443 27285 24452 27319
rect 24400 27276 24452 27285
rect 24768 27319 24820 27328
rect 24768 27285 24777 27319
rect 24777 27285 24811 27319
rect 24811 27285 24820 27319
rect 24768 27276 24820 27285
rect 24952 27276 25004 27328
rect 26976 27480 27028 27532
rect 27712 27480 27764 27532
rect 27804 27523 27856 27532
rect 27804 27489 27813 27523
rect 27813 27489 27847 27523
rect 27847 27489 27856 27523
rect 27804 27480 27856 27489
rect 28908 27548 28960 27600
rect 29184 27548 29236 27600
rect 28540 27480 28592 27532
rect 29000 27480 29052 27532
rect 31576 27616 31628 27668
rect 27068 27412 27120 27464
rect 28080 27455 28132 27464
rect 28080 27421 28089 27455
rect 28089 27421 28123 27455
rect 28123 27421 28132 27455
rect 28080 27412 28132 27421
rect 29184 27412 29236 27464
rect 30564 27412 30616 27464
rect 26056 27344 26108 27396
rect 28632 27276 28684 27328
rect 29552 27319 29604 27328
rect 29552 27285 29561 27319
rect 29561 27285 29595 27319
rect 29595 27285 29604 27319
rect 29552 27276 29604 27285
rect 30656 27276 30708 27328
rect 32404 27412 32456 27464
rect 33324 27548 33376 27600
rect 33692 27480 33744 27532
rect 35900 27616 35952 27668
rect 34244 27480 34296 27532
rect 34796 27412 34848 27464
rect 36636 27455 36688 27464
rect 36636 27421 36645 27455
rect 36645 27421 36679 27455
rect 36679 27421 36688 27455
rect 36636 27412 36688 27421
rect 36912 27344 36964 27396
rect 38016 27344 38068 27396
rect 32128 27276 32180 27328
rect 32588 27276 32640 27328
rect 34152 27276 34204 27328
rect 34520 27276 34572 27328
rect 36636 27276 36688 27328
rect 37096 27276 37148 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 3608 27072 3660 27124
rect 4620 27072 4672 27124
rect 6460 27072 6512 27124
rect 9404 27115 9456 27124
rect 9404 27081 9413 27115
rect 9413 27081 9447 27115
rect 9447 27081 9456 27115
rect 9404 27072 9456 27081
rect 2964 27004 3016 27056
rect 5356 27004 5408 27056
rect 6184 27047 6236 27056
rect 6184 27013 6193 27047
rect 6193 27013 6227 27047
rect 6227 27013 6236 27047
rect 6184 27004 6236 27013
rect 2044 26775 2096 26784
rect 2044 26741 2053 26775
rect 2053 26741 2087 26775
rect 2087 26741 2096 26775
rect 2044 26732 2096 26741
rect 2320 26732 2372 26784
rect 3700 26936 3752 26988
rect 6092 26936 6144 26988
rect 7656 26936 7708 26988
rect 9036 27004 9088 27056
rect 7840 26936 7892 26988
rect 8024 26979 8076 26988
rect 8024 26945 8033 26979
rect 8033 26945 8067 26979
rect 8067 26945 8076 26979
rect 8024 26936 8076 26945
rect 9956 27072 10008 27124
rect 10416 27072 10468 27124
rect 10968 27072 11020 27124
rect 11152 27072 11204 27124
rect 11612 27072 11664 27124
rect 12164 27072 12216 27124
rect 12256 27115 12308 27124
rect 12256 27081 12265 27115
rect 12265 27081 12299 27115
rect 12299 27081 12308 27115
rect 12256 27072 12308 27081
rect 12624 27072 12676 27124
rect 12716 27072 12768 27124
rect 13820 27115 13872 27124
rect 13820 27081 13829 27115
rect 13829 27081 13863 27115
rect 13863 27081 13872 27115
rect 13820 27072 13872 27081
rect 14832 27072 14884 27124
rect 15384 27072 15436 27124
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 10508 26979 10560 26988
rect 10508 26945 10542 26979
rect 10542 26945 10560 26979
rect 10508 26936 10560 26945
rect 3608 26868 3660 26920
rect 4712 26868 4764 26920
rect 9588 26868 9640 26920
rect 9864 26868 9916 26920
rect 11244 26868 11296 26920
rect 15936 27072 15988 27124
rect 16580 27072 16632 27124
rect 18052 27072 18104 27124
rect 18236 27072 18288 27124
rect 11704 26911 11756 26920
rect 11704 26877 11713 26911
rect 11713 26877 11747 26911
rect 11747 26877 11756 26911
rect 11704 26868 11756 26877
rect 10232 26800 10284 26852
rect 13912 26911 13964 26920
rect 13912 26877 13921 26911
rect 13921 26877 13955 26911
rect 13955 26877 13964 26911
rect 13912 26868 13964 26877
rect 10692 26732 10744 26784
rect 11796 26732 11848 26784
rect 14832 26979 14884 26988
rect 14832 26945 14841 26979
rect 14841 26945 14875 26979
rect 14875 26945 14884 26979
rect 14832 26936 14884 26945
rect 14924 26979 14976 26988
rect 14924 26945 14958 26979
rect 14958 26945 14976 26979
rect 14924 26936 14976 26945
rect 14188 26868 14240 26920
rect 18512 26936 18564 26988
rect 19432 27072 19484 27124
rect 21088 27115 21140 27124
rect 21088 27081 21097 27115
rect 21097 27081 21131 27115
rect 21131 27081 21140 27115
rect 21088 27072 21140 27081
rect 21364 27072 21416 27124
rect 22284 27115 22336 27124
rect 22284 27081 22293 27115
rect 22293 27081 22327 27115
rect 22327 27081 22336 27115
rect 22284 27072 22336 27081
rect 16396 26911 16448 26920
rect 16396 26877 16405 26911
rect 16405 26877 16439 26911
rect 16439 26877 16448 26911
rect 16396 26868 16448 26877
rect 14096 26800 14148 26852
rect 14648 26800 14700 26852
rect 18880 26800 18932 26852
rect 16120 26732 16172 26784
rect 17684 26732 17736 26784
rect 19708 26911 19760 26920
rect 19708 26877 19742 26911
rect 19742 26877 19760 26911
rect 19708 26868 19760 26877
rect 20076 26868 20128 26920
rect 21272 26911 21324 26920
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 19340 26843 19392 26852
rect 19340 26809 19349 26843
rect 19349 26809 19383 26843
rect 19383 26809 19392 26843
rect 19340 26800 19392 26809
rect 20628 26775 20680 26784
rect 20628 26741 20637 26775
rect 20637 26741 20671 26775
rect 20671 26741 20680 26775
rect 20628 26732 20680 26741
rect 24768 27072 24820 27124
rect 25320 27072 25372 27124
rect 26148 27072 26200 27124
rect 26792 27072 26844 27124
rect 28080 27072 28132 27124
rect 28724 27115 28776 27124
rect 28724 27081 28733 27115
rect 28733 27081 28767 27115
rect 28767 27081 28776 27115
rect 28724 27072 28776 27081
rect 29184 27115 29236 27124
rect 29184 27081 29193 27115
rect 29193 27081 29227 27115
rect 29227 27081 29236 27115
rect 29184 27072 29236 27081
rect 29552 27072 29604 27124
rect 30656 27072 30708 27124
rect 33232 27072 33284 27124
rect 34336 27072 34388 27124
rect 37924 27072 37976 27124
rect 22744 26936 22796 26988
rect 24584 26936 24636 26988
rect 26056 26936 26108 26988
rect 22376 26911 22428 26920
rect 22376 26877 22385 26911
rect 22385 26877 22419 26911
rect 22419 26877 22428 26911
rect 22376 26868 22428 26877
rect 22652 26911 22704 26920
rect 22652 26877 22661 26911
rect 22661 26877 22695 26911
rect 22695 26877 22704 26911
rect 22652 26868 22704 26877
rect 23296 26911 23348 26920
rect 23296 26877 23305 26911
rect 23305 26877 23339 26911
rect 23339 26877 23348 26911
rect 23296 26868 23348 26877
rect 23664 26911 23716 26920
rect 23664 26877 23698 26911
rect 23698 26877 23716 26911
rect 23664 26868 23716 26877
rect 24032 26868 24084 26920
rect 24676 26911 24728 26920
rect 24676 26877 24685 26911
rect 24685 26877 24719 26911
rect 24719 26877 24728 26911
rect 24676 26868 24728 26877
rect 24952 26868 25004 26920
rect 26976 26979 27028 26988
rect 26976 26945 26985 26979
rect 26985 26945 27019 26979
rect 27019 26945 27028 26979
rect 26976 26936 27028 26945
rect 35808 27004 35860 27056
rect 37740 27047 37792 27056
rect 37740 27013 37749 27047
rect 37749 27013 37783 27047
rect 37783 27013 37792 27047
rect 37740 27004 37792 27013
rect 29092 26936 29144 26988
rect 29460 26936 29512 26988
rect 29644 26979 29696 26988
rect 29644 26945 29653 26979
rect 29653 26945 29687 26979
rect 29687 26945 29696 26979
rect 29644 26936 29696 26945
rect 32772 26979 32824 26988
rect 32772 26945 32781 26979
rect 32781 26945 32815 26979
rect 32815 26945 32824 26979
rect 32772 26936 32824 26945
rect 26516 26868 26568 26920
rect 28908 26868 28960 26920
rect 23388 26800 23440 26852
rect 23848 26732 23900 26784
rect 25044 26800 25096 26852
rect 27712 26732 27764 26784
rect 30288 26911 30340 26920
rect 30288 26877 30297 26911
rect 30297 26877 30331 26911
rect 30331 26877 30340 26911
rect 30288 26868 30340 26877
rect 31576 26868 31628 26920
rect 33048 26979 33100 26988
rect 33048 26945 33057 26979
rect 33057 26945 33091 26979
rect 33091 26945 33100 26979
rect 33048 26936 33100 26945
rect 34244 26936 34296 26988
rect 36084 26936 36136 26988
rect 37924 26936 37976 26988
rect 33232 26868 33284 26920
rect 33784 26911 33836 26920
rect 33784 26877 33793 26911
rect 33793 26877 33827 26911
rect 33827 26877 33836 26911
rect 33784 26868 33836 26877
rect 34704 26911 34756 26920
rect 34704 26877 34713 26911
rect 34713 26877 34747 26911
rect 34747 26877 34756 26911
rect 34704 26868 34756 26877
rect 34796 26868 34848 26920
rect 36268 26868 36320 26920
rect 33600 26800 33652 26852
rect 34244 26800 34296 26852
rect 30012 26775 30064 26784
rect 30012 26741 30021 26775
rect 30021 26741 30055 26775
rect 30055 26741 30064 26775
rect 30012 26732 30064 26741
rect 30564 26732 30616 26784
rect 33232 26732 33284 26784
rect 34520 26732 34572 26784
rect 36544 26732 36596 26784
rect 37280 26732 37332 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2044 26528 2096 26580
rect 3792 26435 3844 26444
rect 3792 26401 3801 26435
rect 3801 26401 3835 26435
rect 3835 26401 3844 26435
rect 3792 26392 3844 26401
rect 5908 26528 5960 26580
rect 8392 26528 8444 26580
rect 9588 26528 9640 26580
rect 11520 26528 11572 26580
rect 12808 26528 12860 26580
rect 13084 26528 13136 26580
rect 14096 26571 14148 26580
rect 14096 26537 14105 26571
rect 14105 26537 14139 26571
rect 14139 26537 14148 26571
rect 14096 26528 14148 26537
rect 15568 26528 15620 26580
rect 17500 26528 17552 26580
rect 19340 26528 19392 26580
rect 9864 26460 9916 26512
rect 5540 26392 5592 26444
rect 6368 26392 6420 26444
rect 11336 26460 11388 26512
rect 2320 26324 2372 26376
rect 3056 26324 3108 26376
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 4712 26367 4764 26376
rect 4712 26333 4721 26367
rect 4721 26333 4755 26367
rect 4755 26333 4764 26367
rect 4712 26324 4764 26333
rect 7104 26324 7156 26376
rect 9496 26324 9548 26376
rect 11428 26392 11480 26444
rect 12532 26460 12584 26512
rect 10876 26367 10928 26376
rect 10876 26333 10885 26367
rect 10885 26333 10919 26367
rect 10919 26333 10928 26367
rect 10876 26324 10928 26333
rect 12992 26392 13044 26444
rect 15476 26435 15528 26444
rect 15476 26401 15485 26435
rect 15485 26401 15519 26435
rect 15519 26401 15528 26435
rect 15476 26392 15528 26401
rect 3700 26188 3752 26240
rect 5816 26256 5868 26308
rect 8760 26256 8812 26308
rect 10232 26256 10284 26308
rect 11244 26256 11296 26308
rect 5632 26231 5684 26240
rect 5632 26197 5641 26231
rect 5641 26197 5675 26231
rect 5675 26197 5684 26231
rect 5632 26188 5684 26197
rect 7656 26188 7708 26240
rect 10968 26231 11020 26240
rect 10968 26197 10977 26231
rect 10977 26197 11011 26231
rect 11011 26197 11020 26231
rect 10968 26188 11020 26197
rect 11152 26188 11204 26240
rect 11796 26256 11848 26308
rect 14740 26324 14792 26376
rect 11612 26188 11664 26240
rect 14648 26256 14700 26308
rect 16120 26367 16172 26376
rect 16120 26333 16129 26367
rect 16129 26333 16163 26367
rect 16163 26333 16172 26367
rect 16120 26324 16172 26333
rect 17500 26324 17552 26376
rect 19432 26392 19484 26444
rect 22100 26528 22152 26580
rect 23204 26528 23256 26580
rect 23480 26528 23532 26580
rect 23572 26528 23624 26580
rect 23848 26528 23900 26580
rect 26516 26571 26568 26580
rect 26516 26537 26525 26571
rect 26525 26537 26559 26571
rect 26559 26537 26568 26571
rect 26516 26528 26568 26537
rect 29644 26528 29696 26580
rect 30288 26528 30340 26580
rect 23388 26392 23440 26444
rect 24216 26392 24268 26444
rect 27068 26503 27120 26512
rect 27068 26469 27077 26503
rect 27077 26469 27111 26503
rect 27111 26469 27120 26503
rect 27068 26460 27120 26469
rect 18236 26324 18288 26376
rect 21272 26367 21324 26376
rect 21272 26333 21281 26367
rect 21281 26333 21315 26367
rect 21315 26333 21324 26367
rect 21272 26324 21324 26333
rect 21916 26324 21968 26376
rect 13084 26231 13136 26240
rect 13084 26197 13093 26231
rect 13093 26197 13127 26231
rect 13127 26197 13136 26231
rect 13084 26188 13136 26197
rect 14004 26188 14056 26240
rect 14556 26188 14608 26240
rect 15292 26256 15344 26308
rect 17960 26299 18012 26308
rect 17960 26265 17994 26299
rect 17994 26265 18012 26299
rect 17960 26256 18012 26265
rect 18880 26256 18932 26308
rect 15568 26231 15620 26240
rect 15568 26197 15577 26231
rect 15577 26197 15611 26231
rect 15611 26197 15620 26231
rect 15568 26188 15620 26197
rect 20260 26188 20312 26240
rect 23664 26324 23716 26376
rect 30564 26392 30616 26444
rect 28724 26324 28776 26376
rect 25412 26256 25464 26308
rect 26240 26256 26292 26308
rect 27804 26256 27856 26308
rect 30012 26324 30064 26376
rect 31392 26367 31444 26376
rect 31392 26333 31426 26367
rect 31426 26333 31444 26367
rect 31392 26324 31444 26333
rect 33784 26528 33836 26580
rect 35348 26528 35400 26580
rect 34796 26392 34848 26444
rect 33140 26324 33192 26376
rect 34704 26324 34756 26376
rect 35532 26435 35584 26444
rect 35532 26401 35541 26435
rect 35541 26401 35575 26435
rect 35575 26401 35584 26435
rect 35532 26392 35584 26401
rect 36084 26392 36136 26444
rect 36452 26435 36504 26444
rect 36452 26401 36461 26435
rect 36461 26401 36495 26435
rect 36495 26401 36504 26435
rect 36452 26392 36504 26401
rect 37280 26460 37332 26512
rect 37004 26435 37056 26444
rect 37004 26401 37013 26435
rect 37013 26401 37047 26435
rect 37047 26401 37056 26435
rect 37004 26392 37056 26401
rect 37096 26392 37148 26444
rect 37648 26435 37700 26444
rect 37648 26401 37657 26435
rect 37657 26401 37691 26435
rect 37691 26401 37700 26435
rect 37648 26392 37700 26401
rect 38200 26392 38252 26444
rect 24952 26188 25004 26240
rect 33968 26256 34020 26308
rect 35348 26299 35400 26308
rect 35348 26265 35357 26299
rect 35357 26265 35391 26299
rect 35391 26265 35400 26299
rect 35348 26256 35400 26265
rect 36728 26367 36780 26376
rect 36728 26333 36737 26367
rect 36737 26333 36771 26367
rect 36771 26333 36780 26367
rect 36728 26324 36780 26333
rect 37832 26324 37884 26376
rect 37924 26324 37976 26376
rect 33600 26188 33652 26240
rect 35900 26256 35952 26308
rect 37188 26188 37240 26240
rect 37740 26231 37792 26240
rect 37740 26197 37749 26231
rect 37749 26197 37783 26231
rect 37783 26197 37792 26231
rect 37740 26188 37792 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5632 25984 5684 26036
rect 7012 25984 7064 26036
rect 2320 25916 2372 25968
rect 3976 25916 4028 25968
rect 2044 25848 2096 25900
rect 4712 25848 4764 25900
rect 5356 25848 5408 25900
rect 8116 25984 8168 26036
rect 9220 25984 9272 26036
rect 9680 25984 9732 26036
rect 10600 25984 10652 26036
rect 11152 25984 11204 26036
rect 11704 25984 11756 26036
rect 13084 25984 13136 26036
rect 15568 25984 15620 26036
rect 17960 25984 18012 26036
rect 21272 25984 21324 26036
rect 25688 25984 25740 26036
rect 11244 25959 11296 25968
rect 11244 25925 11253 25959
rect 11253 25925 11287 25959
rect 11287 25925 11296 25959
rect 11244 25916 11296 25925
rect 13544 25916 13596 25968
rect 23112 25916 23164 25968
rect 7840 25848 7892 25900
rect 10048 25848 10100 25900
rect 9772 25780 9824 25832
rect 10692 25848 10744 25900
rect 14556 25848 14608 25900
rect 15292 25848 15344 25900
rect 11152 25780 11204 25832
rect 11612 25780 11664 25832
rect 4804 25712 4856 25764
rect 10508 25712 10560 25764
rect 14280 25780 14332 25832
rect 14740 25823 14792 25832
rect 14740 25789 14749 25823
rect 14749 25789 14783 25823
rect 14783 25789 14792 25823
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 18972 25848 19024 25900
rect 14740 25780 14792 25789
rect 16396 25780 16448 25832
rect 18144 25780 18196 25832
rect 20260 25848 20312 25900
rect 14924 25712 14976 25764
rect 4896 25687 4948 25696
rect 4896 25653 4905 25687
rect 4905 25653 4939 25687
rect 4939 25653 4948 25687
rect 4896 25644 4948 25653
rect 6092 25687 6144 25696
rect 6092 25653 6101 25687
rect 6101 25653 6135 25687
rect 6135 25653 6144 25687
rect 6092 25644 6144 25653
rect 6736 25644 6788 25696
rect 17132 25644 17184 25696
rect 23204 25823 23256 25832
rect 23204 25789 23213 25823
rect 23213 25789 23247 25823
rect 23247 25789 23256 25823
rect 23204 25780 23256 25789
rect 18972 25712 19024 25764
rect 20260 25712 20312 25764
rect 27436 25984 27488 26036
rect 28264 25984 28316 26036
rect 28448 26027 28500 26036
rect 28448 25993 28457 26027
rect 28457 25993 28491 26027
rect 28491 25993 28500 26027
rect 28448 25984 28500 25993
rect 28908 25984 28960 26036
rect 31576 26027 31628 26036
rect 31576 25993 31585 26027
rect 31585 25993 31619 26027
rect 31619 25993 31628 26027
rect 31576 25984 31628 25993
rect 32128 26027 32180 26036
rect 32128 25993 32137 26027
rect 32137 25993 32171 26027
rect 32171 25993 32180 26027
rect 32128 25984 32180 25993
rect 32956 25984 33008 26036
rect 33232 25984 33284 26036
rect 33600 25984 33652 26036
rect 33968 26027 34020 26036
rect 33968 25993 33977 26027
rect 33977 25993 34011 26027
rect 34011 25993 34020 26027
rect 33968 25984 34020 25993
rect 35348 25984 35400 26036
rect 38200 26027 38252 26036
rect 38200 25993 38209 26027
rect 38209 25993 38243 26027
rect 38243 25993 38252 26027
rect 38200 25984 38252 25993
rect 28632 25916 28684 25968
rect 29092 25848 29144 25900
rect 32588 25959 32640 25968
rect 32588 25925 32597 25959
rect 32597 25925 32631 25959
rect 32631 25925 32640 25959
rect 32588 25916 32640 25925
rect 35440 25959 35492 25968
rect 35440 25925 35449 25959
rect 35449 25925 35483 25959
rect 35483 25925 35492 25959
rect 35440 25916 35492 25925
rect 32864 25848 32916 25900
rect 27620 25780 27672 25832
rect 34520 25891 34572 25900
rect 34520 25857 34529 25891
rect 34529 25857 34563 25891
rect 34563 25857 34572 25891
rect 34520 25848 34572 25857
rect 34796 25848 34848 25900
rect 37372 25916 37424 25968
rect 36820 25848 36872 25900
rect 37004 25848 37056 25900
rect 37832 25891 37884 25900
rect 37832 25857 37841 25891
rect 37841 25857 37875 25891
rect 37875 25857 37884 25891
rect 37832 25848 37884 25857
rect 33416 25780 33468 25832
rect 37648 25780 37700 25832
rect 35532 25712 35584 25764
rect 22560 25644 22612 25696
rect 24768 25687 24820 25696
rect 24768 25653 24777 25687
rect 24777 25653 24811 25687
rect 24811 25653 24820 25687
rect 24768 25644 24820 25653
rect 24860 25644 24912 25696
rect 26424 25644 26476 25696
rect 31944 25687 31996 25696
rect 31944 25653 31953 25687
rect 31953 25653 31987 25687
rect 31987 25653 31996 25687
rect 31944 25644 31996 25653
rect 33692 25687 33744 25696
rect 33692 25653 33701 25687
rect 33701 25653 33735 25687
rect 33735 25653 33744 25687
rect 33692 25644 33744 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2044 25483 2096 25492
rect 2044 25449 2053 25483
rect 2053 25449 2087 25483
rect 2087 25449 2096 25483
rect 2044 25440 2096 25449
rect 3976 25415 4028 25424
rect 3976 25381 3985 25415
rect 3985 25381 4019 25415
rect 4019 25381 4028 25415
rect 3976 25372 4028 25381
rect 3884 25304 3936 25356
rect 4896 25440 4948 25492
rect 5540 25440 5592 25492
rect 7656 25440 7708 25492
rect 10048 25483 10100 25492
rect 10048 25449 10057 25483
rect 10057 25449 10091 25483
rect 10091 25449 10100 25483
rect 10048 25440 10100 25449
rect 5080 25372 5132 25424
rect 14188 25440 14240 25492
rect 14464 25483 14516 25492
rect 14464 25449 14473 25483
rect 14473 25449 14507 25483
rect 14507 25449 14516 25483
rect 14464 25440 14516 25449
rect 14740 25440 14792 25492
rect 15016 25440 15068 25492
rect 18696 25440 18748 25492
rect 23756 25440 23808 25492
rect 24216 25483 24268 25492
rect 24216 25449 24225 25483
rect 24225 25449 24259 25483
rect 24259 25449 24268 25483
rect 24216 25440 24268 25449
rect 25228 25440 25280 25492
rect 28448 25440 28500 25492
rect 32864 25483 32916 25492
rect 32864 25449 32873 25483
rect 32873 25449 32907 25483
rect 32907 25449 32916 25483
rect 32864 25440 32916 25449
rect 18972 25415 19024 25424
rect 18972 25381 18981 25415
rect 18981 25381 19015 25415
rect 19015 25381 19024 25415
rect 18972 25372 19024 25381
rect 4804 25304 4856 25356
rect 10968 25304 11020 25356
rect 11244 25304 11296 25356
rect 19432 25304 19484 25356
rect 22652 25304 22704 25356
rect 23940 25304 23992 25356
rect 29644 25304 29696 25356
rect 30748 25304 30800 25356
rect 7012 25279 7064 25288
rect 7012 25245 7021 25279
rect 7021 25245 7055 25279
rect 7055 25245 7064 25279
rect 7012 25236 7064 25245
rect 8392 25279 8444 25288
rect 8392 25245 8401 25279
rect 8401 25245 8435 25279
rect 8435 25245 8444 25279
rect 8392 25236 8444 25245
rect 13268 25279 13320 25288
rect 13268 25245 13277 25279
rect 13277 25245 13311 25279
rect 13311 25245 13320 25279
rect 13268 25236 13320 25245
rect 16764 25236 16816 25288
rect 18052 25279 18104 25288
rect 18052 25245 18061 25279
rect 18061 25245 18095 25279
rect 18095 25245 18104 25279
rect 18052 25236 18104 25245
rect 26424 25279 26476 25288
rect 26424 25245 26433 25279
rect 26433 25245 26467 25279
rect 26467 25245 26476 25279
rect 26424 25236 26476 25245
rect 29276 25236 29328 25288
rect 30196 25279 30248 25288
rect 30196 25245 30205 25279
rect 30205 25245 30239 25279
rect 30239 25245 30248 25279
rect 30196 25236 30248 25245
rect 35440 25483 35492 25492
rect 35440 25449 35449 25483
rect 35449 25449 35483 25483
rect 35483 25449 35492 25483
rect 35440 25440 35492 25449
rect 37188 25440 37240 25492
rect 38016 25483 38068 25492
rect 38016 25449 38025 25483
rect 38025 25449 38059 25483
rect 38059 25449 38068 25483
rect 38016 25440 38068 25449
rect 37096 25372 37148 25424
rect 37740 25304 37792 25356
rect 35900 25236 35952 25288
rect 11152 25168 11204 25220
rect 35716 25168 35768 25220
rect 3700 25100 3752 25152
rect 4896 25100 4948 25152
rect 7564 25143 7616 25152
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 7564 25100 7616 25109
rect 7748 25143 7800 25152
rect 7748 25109 7757 25143
rect 7757 25109 7791 25143
rect 7791 25109 7800 25143
rect 7748 25100 7800 25109
rect 11428 25100 11480 25152
rect 12716 25143 12768 25152
rect 12716 25109 12725 25143
rect 12725 25109 12759 25143
rect 12759 25109 12768 25143
rect 12716 25100 12768 25109
rect 16396 25143 16448 25152
rect 16396 25109 16405 25143
rect 16405 25109 16439 25143
rect 16439 25109 16448 25143
rect 16396 25100 16448 25109
rect 18696 25100 18748 25152
rect 25688 25100 25740 25152
rect 29552 25143 29604 25152
rect 29552 25109 29561 25143
rect 29561 25109 29595 25143
rect 29595 25109 29604 25143
rect 29552 25100 29604 25109
rect 38292 25100 38344 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4712 24896 4764 24948
rect 5080 24896 5132 24948
rect 5264 24896 5316 24948
rect 7012 24939 7064 24948
rect 7012 24905 7021 24939
rect 7021 24905 7055 24939
rect 7055 24905 7064 24939
rect 7012 24896 7064 24905
rect 12716 24896 12768 24948
rect 31116 24896 31168 24948
rect 3976 24803 4028 24812
rect 3976 24769 3985 24803
rect 3985 24769 4019 24803
rect 4019 24769 4028 24803
rect 3976 24760 4028 24769
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 7012 24692 7064 24744
rect 8852 24735 8904 24744
rect 8852 24701 8861 24735
rect 8861 24701 8895 24735
rect 8895 24701 8904 24735
rect 8852 24692 8904 24701
rect 26240 24828 26292 24880
rect 10140 24760 10192 24812
rect 7196 24624 7248 24676
rect 11060 24692 11112 24744
rect 13636 24760 13688 24812
rect 12992 24735 13044 24744
rect 12992 24701 13001 24735
rect 13001 24701 13035 24735
rect 13035 24701 13044 24735
rect 12992 24692 13044 24701
rect 13912 24692 13964 24744
rect 16120 24735 16172 24744
rect 16120 24701 16129 24735
rect 16129 24701 16163 24735
rect 16163 24701 16172 24735
rect 16120 24692 16172 24701
rect 16856 24692 16908 24744
rect 18236 24760 18288 24812
rect 22468 24760 22520 24812
rect 18880 24735 18932 24744
rect 18880 24701 18889 24735
rect 18889 24701 18923 24735
rect 18923 24701 18932 24735
rect 18880 24692 18932 24701
rect 23756 24692 23808 24744
rect 18052 24624 18104 24676
rect 24124 24624 24176 24676
rect 3884 24556 3936 24608
rect 8208 24599 8260 24608
rect 8208 24565 8217 24599
rect 8217 24565 8251 24599
rect 8251 24565 8260 24599
rect 8208 24556 8260 24565
rect 9588 24599 9640 24608
rect 9588 24565 9597 24599
rect 9597 24565 9631 24599
rect 9631 24565 9640 24599
rect 9588 24556 9640 24565
rect 10876 24556 10928 24608
rect 12072 24599 12124 24608
rect 12072 24565 12081 24599
rect 12081 24565 12115 24599
rect 12115 24565 12124 24599
rect 12072 24556 12124 24565
rect 13452 24556 13504 24608
rect 14280 24599 14332 24608
rect 14280 24565 14289 24599
rect 14289 24565 14323 24599
rect 14323 24565 14332 24599
rect 14280 24556 14332 24565
rect 15384 24556 15436 24608
rect 23848 24599 23900 24608
rect 23848 24565 23857 24599
rect 23857 24565 23891 24599
rect 23891 24565 23900 24599
rect 23848 24556 23900 24565
rect 25228 24735 25280 24744
rect 25228 24701 25237 24735
rect 25237 24701 25271 24735
rect 25271 24701 25280 24735
rect 25228 24692 25280 24701
rect 25780 24692 25832 24744
rect 26148 24735 26200 24744
rect 26148 24701 26157 24735
rect 26157 24701 26191 24735
rect 26191 24701 26200 24735
rect 26148 24692 26200 24701
rect 29368 24760 29420 24812
rect 29276 24735 29328 24744
rect 29276 24701 29285 24735
rect 29285 24701 29319 24735
rect 29319 24701 29328 24735
rect 29276 24692 29328 24701
rect 29828 24692 29880 24744
rect 34704 24692 34756 24744
rect 35900 24735 35952 24744
rect 35900 24701 35909 24735
rect 35909 24701 35943 24735
rect 35943 24701 35952 24735
rect 35900 24692 35952 24701
rect 37004 24735 37056 24744
rect 37004 24701 37013 24735
rect 37013 24701 37047 24735
rect 37047 24701 37056 24735
rect 37004 24692 37056 24701
rect 37096 24692 37148 24744
rect 29736 24624 29788 24676
rect 26332 24556 26384 24608
rect 26516 24556 26568 24608
rect 28356 24599 28408 24608
rect 28356 24565 28365 24599
rect 28365 24565 28399 24599
rect 28399 24565 28408 24599
rect 28356 24556 28408 24565
rect 28724 24556 28776 24608
rect 29920 24599 29972 24608
rect 29920 24565 29929 24599
rect 29929 24565 29963 24599
rect 29963 24565 29972 24599
rect 29920 24556 29972 24565
rect 30748 24599 30800 24608
rect 30748 24565 30757 24599
rect 30757 24565 30791 24599
rect 30791 24565 30800 24599
rect 30748 24556 30800 24565
rect 34336 24556 34388 24608
rect 35348 24599 35400 24608
rect 35348 24565 35357 24599
rect 35357 24565 35391 24599
rect 35391 24565 35400 24599
rect 35348 24556 35400 24565
rect 36360 24599 36412 24608
rect 36360 24565 36369 24599
rect 36369 24565 36403 24599
rect 36403 24565 36412 24599
rect 36360 24556 36412 24565
rect 36912 24556 36964 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 5080 24352 5132 24404
rect 7380 24352 7432 24404
rect 13912 24352 13964 24404
rect 16120 24352 16172 24404
rect 17316 24352 17368 24404
rect 24032 24352 24084 24404
rect 25044 24352 25096 24404
rect 26148 24352 26200 24404
rect 26424 24352 26476 24404
rect 27620 24395 27672 24404
rect 27620 24361 27629 24395
rect 27629 24361 27663 24395
rect 27663 24361 27672 24395
rect 27620 24352 27672 24361
rect 12072 24284 12124 24336
rect 16212 24284 16264 24336
rect 29828 24352 29880 24404
rect 30196 24352 30248 24404
rect 31116 24395 31168 24404
rect 31116 24361 31125 24395
rect 31125 24361 31159 24395
rect 31159 24361 31168 24395
rect 31116 24352 31168 24361
rect 34612 24352 34664 24404
rect 37740 24395 37792 24404
rect 37740 24361 37749 24395
rect 37749 24361 37783 24395
rect 37783 24361 37792 24395
rect 37740 24352 37792 24361
rect 32588 24284 32640 24336
rect 33324 24284 33376 24336
rect 3424 24191 3476 24200
rect 3424 24157 3433 24191
rect 3433 24157 3467 24191
rect 3467 24157 3476 24191
rect 3424 24148 3476 24157
rect 4620 24148 4672 24200
rect 6368 24191 6420 24200
rect 6368 24157 6377 24191
rect 6377 24157 6411 24191
rect 6411 24157 6420 24191
rect 6368 24148 6420 24157
rect 7104 24148 7156 24200
rect 9036 24191 9088 24200
rect 9036 24157 9045 24191
rect 9045 24157 9079 24191
rect 9079 24157 9088 24191
rect 9036 24148 9088 24157
rect 10876 24148 10928 24200
rect 13544 24148 13596 24200
rect 14556 24148 14608 24200
rect 14648 24191 14700 24200
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 16396 24148 16448 24200
rect 18512 24216 18564 24268
rect 25964 24259 26016 24268
rect 25964 24225 25973 24259
rect 25973 24225 26007 24259
rect 26007 24225 26016 24259
rect 25964 24216 26016 24225
rect 6828 24080 6880 24132
rect 2872 24055 2924 24064
rect 2872 24021 2881 24055
rect 2881 24021 2915 24055
rect 2915 24021 2924 24055
rect 2872 24012 2924 24021
rect 3792 24055 3844 24064
rect 3792 24021 3801 24055
rect 3801 24021 3835 24055
rect 3835 24021 3844 24055
rect 3792 24012 3844 24021
rect 5264 24012 5316 24064
rect 8668 24012 8720 24064
rect 9312 24012 9364 24064
rect 11612 24012 11664 24064
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 17960 24191 18012 24200
rect 17960 24157 17969 24191
rect 17969 24157 18003 24191
rect 18003 24157 18012 24191
rect 17960 24148 18012 24157
rect 18604 24191 18656 24200
rect 18604 24157 18613 24191
rect 18613 24157 18647 24191
rect 18647 24157 18656 24191
rect 18604 24148 18656 24157
rect 24768 24148 24820 24200
rect 29644 24259 29696 24268
rect 29644 24225 29653 24259
rect 29653 24225 29687 24259
rect 29687 24225 29696 24259
rect 29644 24216 29696 24225
rect 29736 24216 29788 24268
rect 29920 24216 29972 24268
rect 35624 24216 35676 24268
rect 26516 24148 26568 24200
rect 16764 24080 16816 24132
rect 13360 24012 13412 24064
rect 13728 24012 13780 24064
rect 15568 24012 15620 24064
rect 17040 24012 17092 24064
rect 25688 24080 25740 24132
rect 29552 24148 29604 24200
rect 30748 24148 30800 24200
rect 30932 24191 30984 24200
rect 30932 24157 30941 24191
rect 30941 24157 30975 24191
rect 30975 24157 30984 24191
rect 30932 24148 30984 24157
rect 17868 24012 17920 24064
rect 25228 24012 25280 24064
rect 26240 24055 26292 24064
rect 26240 24021 26249 24055
rect 26249 24021 26283 24055
rect 26283 24021 26292 24055
rect 26240 24012 26292 24021
rect 26332 24012 26384 24064
rect 27344 24055 27396 24064
rect 27344 24021 27353 24055
rect 27353 24021 27387 24055
rect 27387 24021 27396 24055
rect 27344 24012 27396 24021
rect 30288 24080 30340 24132
rect 33784 24148 33836 24200
rect 35716 24148 35768 24200
rect 36176 24191 36228 24200
rect 36176 24157 36185 24191
rect 36185 24157 36219 24191
rect 36219 24157 36228 24191
rect 36176 24148 36228 24157
rect 36912 24148 36964 24200
rect 29276 24012 29328 24064
rect 30196 24012 30248 24064
rect 30380 24055 30432 24064
rect 30380 24021 30389 24055
rect 30389 24021 30423 24055
rect 30423 24021 30432 24055
rect 30380 24012 30432 24021
rect 31852 24055 31904 24064
rect 31852 24021 31861 24055
rect 31861 24021 31895 24055
rect 31895 24021 31904 24055
rect 31852 24012 31904 24021
rect 35716 24012 35768 24064
rect 36636 24012 36688 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3424 23808 3476 23860
rect 4988 23808 5040 23860
rect 5172 23808 5224 23860
rect 5724 23808 5776 23860
rect 4712 23672 4764 23724
rect 3056 23647 3108 23656
rect 3056 23613 3065 23647
rect 3065 23613 3099 23647
rect 3099 23613 3108 23647
rect 3056 23604 3108 23613
rect 3884 23647 3936 23656
rect 3884 23613 3893 23647
rect 3893 23613 3927 23647
rect 3927 23613 3936 23647
rect 3884 23604 3936 23613
rect 3976 23604 4028 23656
rect 4804 23647 4856 23656
rect 4804 23613 4813 23647
rect 4813 23613 4847 23647
rect 4847 23613 4856 23647
rect 4804 23604 4856 23613
rect 5264 23604 5316 23656
rect 7748 23808 7800 23860
rect 8208 23808 8260 23860
rect 8576 23851 8628 23860
rect 8576 23817 8585 23851
rect 8585 23817 8619 23851
rect 8619 23817 8628 23851
rect 8576 23808 8628 23817
rect 9036 23808 9088 23860
rect 9588 23808 9640 23860
rect 10324 23740 10376 23792
rect 12532 23740 12584 23792
rect 13820 23808 13872 23860
rect 14280 23808 14332 23860
rect 14648 23808 14700 23860
rect 16764 23808 16816 23860
rect 13452 23740 13504 23792
rect 14556 23740 14608 23792
rect 6276 23604 6328 23656
rect 5356 23536 5408 23588
rect 7012 23672 7064 23724
rect 12716 23672 12768 23724
rect 13636 23672 13688 23724
rect 14188 23672 14240 23724
rect 16304 23740 16356 23792
rect 15384 23715 15436 23724
rect 15384 23681 15418 23715
rect 15418 23681 15436 23715
rect 15384 23672 15436 23681
rect 18052 23808 18104 23860
rect 18512 23808 18564 23860
rect 18696 23808 18748 23860
rect 18880 23808 18932 23860
rect 22192 23808 22244 23860
rect 22468 23808 22520 23860
rect 23848 23808 23900 23860
rect 25044 23808 25096 23860
rect 26332 23808 26384 23860
rect 17868 23715 17920 23724
rect 17868 23681 17902 23715
rect 17902 23681 17920 23715
rect 17868 23672 17920 23681
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 27344 23851 27396 23860
rect 27344 23817 27353 23851
rect 27353 23817 27387 23851
rect 27387 23817 27396 23851
rect 27344 23808 27396 23817
rect 28356 23808 28408 23860
rect 29736 23808 29788 23860
rect 28172 23740 28224 23792
rect 25228 23672 25280 23724
rect 25780 23715 25832 23724
rect 25780 23681 25789 23715
rect 25789 23681 25823 23715
rect 25823 23681 25832 23715
rect 25780 23672 25832 23681
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 30932 23808 30984 23860
rect 37004 23808 37056 23860
rect 29368 23715 29420 23724
rect 29368 23681 29386 23715
rect 29386 23681 29420 23715
rect 29368 23672 29420 23681
rect 30288 23672 30340 23724
rect 34336 23715 34388 23724
rect 34336 23681 34370 23715
rect 34370 23681 34388 23715
rect 34336 23672 34388 23681
rect 35624 23672 35676 23724
rect 7104 23604 7156 23656
rect 2504 23511 2556 23520
rect 2504 23477 2513 23511
rect 2513 23477 2547 23511
rect 2547 23477 2556 23511
rect 2504 23468 2556 23477
rect 4068 23511 4120 23520
rect 4068 23477 4077 23511
rect 4077 23477 4111 23511
rect 4111 23477 4120 23511
rect 4068 23468 4120 23477
rect 5448 23511 5500 23520
rect 5448 23477 5457 23511
rect 5457 23477 5491 23511
rect 5491 23477 5500 23511
rect 5448 23468 5500 23477
rect 7104 23511 7156 23520
rect 7104 23477 7113 23511
rect 7113 23477 7147 23511
rect 7147 23477 7156 23511
rect 7104 23468 7156 23477
rect 8392 23604 8444 23656
rect 10232 23604 10284 23656
rect 13728 23647 13780 23656
rect 13728 23613 13737 23647
rect 13737 23613 13771 23647
rect 13771 23613 13780 23647
rect 13728 23604 13780 23613
rect 13820 23604 13872 23656
rect 17040 23647 17092 23656
rect 17040 23613 17049 23647
rect 17049 23613 17083 23647
rect 17083 23613 17092 23647
rect 17040 23604 17092 23613
rect 14556 23536 14608 23588
rect 17500 23579 17552 23588
rect 17500 23545 17509 23579
rect 17509 23545 17543 23579
rect 17543 23545 17552 23579
rect 17500 23536 17552 23545
rect 7840 23468 7892 23520
rect 13728 23468 13780 23520
rect 15384 23468 15436 23520
rect 16212 23468 16264 23520
rect 18236 23604 18288 23656
rect 18696 23604 18748 23656
rect 23388 23647 23440 23656
rect 23388 23613 23397 23647
rect 23397 23613 23431 23647
rect 23431 23613 23440 23647
rect 23388 23604 23440 23613
rect 25872 23647 25924 23656
rect 25872 23613 25906 23647
rect 25906 23613 25924 23647
rect 25872 23604 25924 23613
rect 27712 23604 27764 23656
rect 29000 23604 29052 23656
rect 29828 23604 29880 23656
rect 30104 23604 30156 23656
rect 19340 23468 19392 23520
rect 19616 23511 19668 23520
rect 19616 23477 19625 23511
rect 19625 23477 19659 23511
rect 19659 23477 19668 23511
rect 19616 23468 19668 23477
rect 22468 23511 22520 23520
rect 22468 23477 22477 23511
rect 22477 23477 22511 23511
rect 22511 23477 22520 23511
rect 22468 23468 22520 23477
rect 23756 23468 23808 23520
rect 24952 23468 25004 23520
rect 25136 23468 25188 23520
rect 25412 23468 25464 23520
rect 27620 23536 27672 23588
rect 28724 23536 28776 23588
rect 30472 23604 30524 23656
rect 31116 23604 31168 23656
rect 33876 23647 33928 23656
rect 33876 23613 33885 23647
rect 33885 23613 33919 23647
rect 33919 23613 33928 23647
rect 33876 23604 33928 23613
rect 36544 23604 36596 23656
rect 26976 23511 27028 23520
rect 26976 23477 26985 23511
rect 26985 23477 27019 23511
rect 27019 23477 27028 23511
rect 26976 23468 27028 23477
rect 27988 23468 28040 23520
rect 28540 23511 28592 23520
rect 28540 23477 28549 23511
rect 28549 23477 28583 23511
rect 28583 23477 28592 23511
rect 28540 23468 28592 23477
rect 33324 23511 33376 23520
rect 33324 23477 33333 23511
rect 33333 23477 33367 23511
rect 33367 23477 33376 23511
rect 33324 23468 33376 23477
rect 35900 23468 35952 23520
rect 36452 23468 36504 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4620 23307 4672 23316
rect 4620 23273 4629 23307
rect 4629 23273 4663 23307
rect 4663 23273 4672 23307
rect 4620 23264 4672 23273
rect 4712 23264 4764 23316
rect 6828 23307 6880 23316
rect 6828 23273 6837 23307
rect 6837 23273 6871 23307
rect 6871 23273 6880 23307
rect 6828 23264 6880 23273
rect 4252 23196 4304 23248
rect 4344 23196 4396 23248
rect 2044 23060 2096 23112
rect 3792 23060 3844 23112
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 4436 22992 4488 23044
rect 4804 22992 4856 23044
rect 5172 23171 5224 23180
rect 5172 23137 5181 23171
rect 5181 23137 5215 23171
rect 5215 23137 5224 23171
rect 5172 23128 5224 23137
rect 6920 23128 6972 23180
rect 7656 23264 7708 23316
rect 7380 23128 7432 23180
rect 5448 23060 5500 23112
rect 8392 23196 8444 23248
rect 8852 23264 8904 23316
rect 9588 23264 9640 23316
rect 12716 23264 12768 23316
rect 7665 23103 7717 23112
rect 7665 23069 7711 23103
rect 7711 23069 7717 23103
rect 8576 23171 8628 23180
rect 8576 23137 8585 23171
rect 8585 23137 8619 23171
rect 8619 23137 8628 23171
rect 8576 23128 8628 23137
rect 8668 23128 8720 23180
rect 9588 23171 9640 23180
rect 9588 23137 9597 23171
rect 9597 23137 9631 23171
rect 9631 23137 9640 23171
rect 9588 23128 9640 23137
rect 13268 23264 13320 23316
rect 15200 23264 15252 23316
rect 13360 23196 13412 23248
rect 15384 23196 15436 23248
rect 13728 23171 13780 23180
rect 13728 23137 13737 23171
rect 13737 23137 13771 23171
rect 13771 23137 13780 23171
rect 13728 23128 13780 23137
rect 7665 23060 7717 23069
rect 5356 22992 5408 23044
rect 9312 23103 9364 23112
rect 9312 23069 9321 23103
rect 9321 23069 9355 23103
rect 9355 23069 9364 23103
rect 9312 23060 9364 23069
rect 10232 23060 10284 23112
rect 12716 23103 12768 23112
rect 12716 23069 12725 23103
rect 12725 23069 12759 23103
rect 12759 23069 12768 23103
rect 12716 23060 12768 23069
rect 12900 23103 12952 23112
rect 12900 23069 12918 23103
rect 12918 23069 12952 23103
rect 12900 23060 12952 23069
rect 13912 23103 13964 23112
rect 13912 23069 13921 23103
rect 13921 23069 13955 23103
rect 13955 23069 13964 23103
rect 13912 23060 13964 23069
rect 15568 23264 15620 23316
rect 16304 23264 16356 23316
rect 17960 23264 18012 23316
rect 18604 23264 18656 23316
rect 18696 23239 18748 23248
rect 18696 23205 18705 23239
rect 18705 23205 18739 23239
rect 18739 23205 18748 23239
rect 18696 23196 18748 23205
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 22468 23128 22520 23180
rect 22744 23128 22796 23180
rect 25412 23264 25464 23316
rect 25688 23128 25740 23180
rect 26608 23264 26660 23316
rect 27712 23307 27764 23316
rect 27712 23273 27721 23307
rect 27721 23273 27755 23307
rect 27755 23273 27764 23307
rect 27712 23264 27764 23273
rect 29368 23264 29420 23316
rect 30288 23264 30340 23316
rect 32588 23307 32640 23316
rect 32588 23273 32597 23307
rect 32597 23273 32631 23307
rect 32631 23273 32640 23307
rect 32588 23264 32640 23273
rect 34704 23307 34756 23316
rect 34704 23273 34713 23307
rect 34713 23273 34747 23307
rect 34747 23273 34756 23307
rect 34704 23264 34756 23273
rect 34796 23264 34848 23316
rect 36452 23264 36504 23316
rect 31116 23196 31168 23248
rect 35992 23196 36044 23248
rect 26240 23128 26292 23180
rect 26976 23128 27028 23180
rect 32588 23128 32640 23180
rect 34612 23128 34664 23180
rect 35900 23128 35952 23180
rect 37004 23264 37056 23316
rect 37004 23171 37056 23180
rect 37004 23137 37013 23171
rect 37013 23137 37047 23171
rect 37047 23137 37056 23171
rect 37004 23128 37056 23137
rect 37740 23128 37792 23180
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 19616 23060 19668 23112
rect 21272 23103 21324 23112
rect 21272 23069 21281 23103
rect 21281 23069 21315 23103
rect 21315 23069 21324 23103
rect 21272 23060 21324 23069
rect 22100 23060 22152 23112
rect 23388 23060 23440 23112
rect 27896 23103 27948 23112
rect 27896 23069 27905 23103
rect 27905 23069 27939 23103
rect 27939 23069 27948 23103
rect 27896 23060 27948 23069
rect 27988 23060 28040 23112
rect 32312 23060 32364 23112
rect 32772 23060 32824 23112
rect 35348 23060 35400 23112
rect 36452 23103 36504 23112
rect 36452 23069 36461 23103
rect 36461 23069 36495 23103
rect 36495 23069 36504 23103
rect 36452 23060 36504 23069
rect 37464 23103 37516 23112
rect 37464 23069 37473 23103
rect 37473 23069 37507 23103
rect 37507 23069 37516 23103
rect 37464 23060 37516 23069
rect 10692 22992 10744 23044
rect 23296 22992 23348 23044
rect 26056 22992 26108 23044
rect 26332 22992 26384 23044
rect 31852 22992 31904 23044
rect 33600 22992 33652 23044
rect 4528 22967 4580 22976
rect 4528 22933 4537 22967
rect 4537 22933 4571 22967
rect 4571 22933 4580 22967
rect 4528 22924 4580 22933
rect 6920 22967 6972 22976
rect 6920 22933 6929 22967
rect 6929 22933 6963 22967
rect 6963 22933 6972 22967
rect 6920 22924 6972 22933
rect 7012 22924 7064 22976
rect 9864 22924 9916 22976
rect 13176 22924 13228 22976
rect 14096 22967 14148 22976
rect 14096 22933 14105 22967
rect 14105 22933 14139 22967
rect 14139 22933 14148 22967
rect 14096 22924 14148 22933
rect 17960 22967 18012 22976
rect 17960 22933 17969 22967
rect 17969 22933 18003 22967
rect 18003 22933 18012 22967
rect 17960 22924 18012 22933
rect 18512 22924 18564 22976
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 21916 22967 21968 22976
rect 21916 22933 21925 22967
rect 21925 22933 21959 22967
rect 21959 22933 21968 22967
rect 21916 22924 21968 22933
rect 22376 22967 22428 22976
rect 22376 22933 22385 22967
rect 22385 22933 22419 22967
rect 22419 22933 22428 22967
rect 22376 22924 22428 22933
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 23940 22924 23992 22976
rect 25780 22967 25832 22976
rect 25780 22933 25789 22967
rect 25789 22933 25823 22967
rect 25823 22933 25832 22967
rect 25780 22924 25832 22933
rect 26240 22967 26292 22976
rect 26240 22933 26249 22967
rect 26249 22933 26283 22967
rect 26283 22933 26292 22967
rect 26240 22924 26292 22933
rect 26608 22967 26660 22976
rect 26608 22933 26617 22967
rect 26617 22933 26651 22967
rect 26651 22933 26660 22967
rect 26608 22924 26660 22933
rect 32588 22924 32640 22976
rect 33048 22924 33100 22976
rect 33968 22967 34020 22976
rect 33968 22933 33977 22967
rect 33977 22933 34011 22967
rect 34011 22933 34020 22967
rect 33968 22924 34020 22933
rect 35532 22924 35584 22976
rect 36912 22924 36964 22976
rect 37188 22924 37240 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4528 22720 4580 22772
rect 2504 22652 2556 22704
rect 2044 22584 2096 22636
rect 4344 22627 4396 22636
rect 4344 22593 4353 22627
rect 4353 22593 4387 22627
rect 4387 22593 4396 22627
rect 4344 22584 4396 22593
rect 4436 22627 4488 22636
rect 6368 22720 6420 22772
rect 6920 22720 6972 22772
rect 9864 22763 9916 22772
rect 9864 22729 9873 22763
rect 9873 22729 9907 22763
rect 9907 22729 9916 22763
rect 9864 22720 9916 22729
rect 10324 22720 10376 22772
rect 10692 22763 10744 22772
rect 10692 22729 10701 22763
rect 10701 22729 10735 22763
rect 10735 22729 10744 22763
rect 10692 22720 10744 22729
rect 12992 22763 13044 22772
rect 12992 22729 13001 22763
rect 13001 22729 13035 22763
rect 13035 22729 13044 22763
rect 12992 22720 13044 22729
rect 14096 22720 14148 22772
rect 17868 22720 17920 22772
rect 18236 22720 18288 22772
rect 21272 22720 21324 22772
rect 21364 22720 21416 22772
rect 21916 22720 21968 22772
rect 22468 22720 22520 22772
rect 25228 22720 25280 22772
rect 26056 22763 26108 22772
rect 26056 22729 26065 22763
rect 26065 22729 26099 22763
rect 26099 22729 26108 22763
rect 26056 22720 26108 22729
rect 26332 22720 26384 22772
rect 26608 22720 26660 22772
rect 27620 22720 27672 22772
rect 28540 22720 28592 22772
rect 30104 22720 30156 22772
rect 33784 22763 33836 22772
rect 33784 22729 33793 22763
rect 33793 22729 33827 22763
rect 33827 22729 33836 22763
rect 33784 22720 33836 22729
rect 7564 22652 7616 22704
rect 4436 22593 4470 22627
rect 4470 22593 4488 22627
rect 4436 22584 4488 22593
rect 8576 22652 8628 22704
rect 11612 22652 11664 22704
rect 11796 22695 11848 22704
rect 11796 22661 11830 22695
rect 11830 22661 11848 22695
rect 11796 22652 11848 22661
rect 12440 22652 12492 22704
rect 13636 22652 13688 22704
rect 3976 22516 4028 22568
rect 3884 22448 3936 22500
rect 7840 22584 7892 22636
rect 8668 22584 8720 22636
rect 10232 22584 10284 22636
rect 12532 22584 12584 22636
rect 13360 22584 13412 22636
rect 8116 22516 8168 22568
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 11336 22559 11388 22568
rect 11336 22525 11345 22559
rect 11345 22525 11379 22559
rect 11379 22525 11388 22559
rect 11336 22516 11388 22525
rect 13268 22516 13320 22568
rect 16304 22584 16356 22636
rect 17684 22584 17736 22636
rect 22376 22652 22428 22704
rect 6184 22448 6236 22500
rect 4620 22380 4672 22432
rect 5356 22423 5408 22432
rect 5356 22389 5365 22423
rect 5365 22389 5399 22423
rect 5399 22389 5408 22423
rect 5356 22380 5408 22389
rect 8760 22448 8812 22500
rect 8024 22423 8076 22432
rect 8024 22389 8033 22423
rect 8033 22389 8067 22423
rect 8067 22389 8076 22423
rect 8024 22380 8076 22389
rect 8300 22380 8352 22432
rect 9588 22380 9640 22432
rect 21364 22559 21416 22568
rect 21364 22525 21373 22559
rect 21373 22525 21407 22559
rect 21407 22525 21416 22559
rect 21364 22516 21416 22525
rect 18144 22423 18196 22432
rect 18144 22389 18153 22423
rect 18153 22389 18187 22423
rect 18187 22389 18196 22423
rect 18144 22380 18196 22389
rect 20168 22423 20220 22432
rect 20168 22389 20177 22423
rect 20177 22389 20211 22423
rect 20211 22389 20220 22423
rect 20168 22380 20220 22389
rect 22560 22516 22612 22568
rect 23388 22584 23440 22636
rect 27896 22652 27948 22704
rect 28908 22652 28960 22704
rect 28632 22584 28684 22636
rect 30380 22652 30432 22704
rect 35348 22720 35400 22772
rect 35624 22720 35676 22772
rect 36544 22720 36596 22772
rect 36636 22763 36688 22772
rect 36636 22729 36645 22763
rect 36645 22729 36679 22763
rect 36679 22729 36688 22763
rect 36636 22720 36688 22729
rect 37096 22763 37148 22772
rect 37096 22729 37105 22763
rect 37105 22729 37139 22763
rect 37139 22729 37148 22763
rect 37096 22720 37148 22729
rect 29000 22516 29052 22568
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 32588 22627 32640 22636
rect 32588 22593 32622 22627
rect 32622 22593 32640 22627
rect 32588 22584 32640 22593
rect 35532 22652 35584 22704
rect 36452 22652 36504 22704
rect 35992 22584 36044 22636
rect 36912 22652 36964 22704
rect 37556 22652 37608 22704
rect 23480 22448 23532 22500
rect 24216 22448 24268 22500
rect 35440 22559 35492 22568
rect 35440 22525 35449 22559
rect 35449 22525 35483 22559
rect 35483 22525 35492 22559
rect 35440 22516 35492 22525
rect 36360 22516 36412 22568
rect 36728 22516 36780 22568
rect 37280 22516 37332 22568
rect 37648 22627 37700 22636
rect 37648 22593 37657 22627
rect 37657 22593 37691 22627
rect 37691 22593 37700 22627
rect 37648 22584 37700 22593
rect 37740 22516 37792 22568
rect 35716 22448 35768 22500
rect 22192 22380 22244 22432
rect 22836 22380 22888 22432
rect 28540 22423 28592 22432
rect 28540 22389 28549 22423
rect 28549 22389 28583 22423
rect 28583 22389 28592 22423
rect 28540 22380 28592 22389
rect 30380 22423 30432 22432
rect 30380 22389 30389 22423
rect 30389 22389 30423 22423
rect 30423 22389 30432 22423
rect 30380 22380 30432 22389
rect 33876 22380 33928 22432
rect 34520 22380 34572 22432
rect 35440 22380 35492 22432
rect 35624 22380 35676 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3976 22176 4028 22228
rect 5632 22219 5684 22228
rect 3884 22108 3936 22160
rect 5632 22185 5641 22219
rect 5641 22185 5675 22219
rect 5675 22185 5684 22219
rect 5632 22176 5684 22185
rect 5908 22176 5960 22228
rect 6920 22176 6972 22228
rect 11336 22176 11388 22228
rect 16856 22176 16908 22228
rect 17684 22219 17736 22228
rect 17684 22185 17693 22219
rect 17693 22185 17727 22219
rect 17727 22185 17736 22219
rect 17684 22176 17736 22185
rect 18052 22176 18104 22228
rect 5172 22083 5224 22092
rect 5172 22049 5181 22083
rect 5181 22049 5215 22083
rect 5215 22049 5224 22083
rect 5172 22040 5224 22049
rect 7840 22040 7892 22092
rect 7932 22040 7984 22092
rect 8484 22083 8536 22092
rect 8484 22049 8493 22083
rect 8493 22049 8527 22083
rect 8527 22049 8536 22083
rect 8484 22040 8536 22049
rect 10876 22040 10928 22092
rect 12900 22040 12952 22092
rect 18144 22040 18196 22092
rect 21824 22176 21876 22228
rect 25688 22219 25740 22228
rect 25688 22185 25697 22219
rect 25697 22185 25731 22219
rect 25731 22185 25740 22219
rect 25688 22176 25740 22185
rect 26240 22176 26292 22228
rect 22560 22108 22612 22160
rect 23020 22108 23072 22160
rect 2044 21972 2096 22024
rect 7104 21972 7156 22024
rect 2872 21904 2924 21956
rect 4068 21904 4120 21956
rect 5356 21904 5408 21956
rect 5448 21904 5500 21956
rect 5908 21904 5960 21956
rect 6276 21904 6328 21956
rect 9956 21904 10008 21956
rect 6184 21836 6236 21888
rect 8300 21836 8352 21888
rect 10324 21836 10376 21888
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 19984 22015 20036 22024
rect 19984 21981 20018 22015
rect 20018 21981 20036 22015
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 12440 21836 12492 21888
rect 17224 21879 17276 21888
rect 17224 21845 17233 21879
rect 17233 21845 17267 21879
rect 17267 21845 17276 21879
rect 17224 21836 17276 21845
rect 19984 21972 20036 21981
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 22744 22040 22796 22092
rect 22100 22015 22152 22024
rect 22100 21981 22109 22015
rect 22109 21981 22143 22015
rect 22143 21981 22152 22015
rect 22100 21972 22152 21981
rect 18788 21836 18840 21888
rect 21180 21879 21232 21888
rect 21180 21845 21189 21879
rect 21189 21845 21223 21879
rect 21223 21845 21232 21879
rect 21180 21836 21232 21845
rect 23296 22040 23348 22092
rect 24032 22108 24084 22160
rect 24124 22040 24176 22092
rect 25780 22040 25832 22092
rect 26148 22040 26200 22092
rect 28816 22176 28868 22228
rect 29368 22176 29420 22228
rect 34796 22176 34848 22228
rect 35440 22219 35492 22228
rect 35440 22185 35449 22219
rect 35449 22185 35483 22219
rect 35483 22185 35492 22219
rect 35440 22176 35492 22185
rect 37464 22176 37516 22228
rect 37648 22176 37700 22228
rect 28448 22108 28500 22160
rect 30380 22108 30432 22160
rect 33876 22151 33928 22160
rect 33876 22117 33885 22151
rect 33885 22117 33919 22151
rect 33919 22117 33928 22151
rect 33876 22108 33928 22117
rect 23204 21904 23256 21956
rect 25688 21904 25740 21956
rect 28448 21904 28500 21956
rect 32220 22040 32272 22092
rect 34428 22040 34480 22092
rect 36268 22108 36320 22160
rect 35992 22040 36044 22092
rect 33048 21972 33100 22024
rect 31944 21904 31996 21956
rect 35256 21972 35308 22024
rect 35348 21972 35400 22024
rect 36360 22015 36412 22024
rect 36360 21981 36369 22015
rect 36369 21981 36403 22015
rect 36403 21981 36412 22015
rect 36360 21972 36412 21981
rect 37188 21972 37240 22024
rect 22100 21836 22152 21888
rect 23020 21836 23072 21888
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 23572 21879 23624 21888
rect 23572 21845 23581 21879
rect 23581 21845 23615 21879
rect 23615 21845 23624 21879
rect 23572 21836 23624 21845
rect 24124 21836 24176 21888
rect 28816 21836 28868 21888
rect 29368 21836 29420 21888
rect 32404 21879 32456 21888
rect 32404 21845 32413 21879
rect 32413 21845 32447 21879
rect 32447 21845 32456 21879
rect 32404 21836 32456 21845
rect 34980 21879 35032 21888
rect 34980 21845 34989 21879
rect 34989 21845 35023 21879
rect 35023 21845 35032 21879
rect 34980 21836 35032 21845
rect 35900 21947 35952 21956
rect 35900 21913 35909 21947
rect 35909 21913 35943 21947
rect 35943 21913 35952 21947
rect 35900 21904 35952 21913
rect 36452 21904 36504 21956
rect 36176 21836 36228 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3056 21632 3108 21684
rect 5172 21632 5224 21684
rect 7932 21675 7984 21684
rect 7932 21641 7941 21675
rect 7941 21641 7975 21675
rect 7975 21641 7984 21675
rect 7932 21632 7984 21641
rect 8576 21632 8628 21684
rect 13728 21632 13780 21684
rect 21180 21632 21232 21684
rect 22376 21632 22428 21684
rect 22560 21675 22612 21684
rect 22560 21641 22569 21675
rect 22569 21641 22603 21675
rect 22603 21641 22612 21675
rect 22560 21632 22612 21641
rect 23388 21632 23440 21684
rect 24032 21632 24084 21684
rect 24308 21632 24360 21684
rect 32772 21675 32824 21684
rect 32772 21641 32781 21675
rect 32781 21641 32815 21675
rect 32815 21641 32824 21675
rect 32772 21632 32824 21641
rect 33324 21632 33376 21684
rect 33600 21632 33652 21684
rect 5908 21564 5960 21616
rect 11704 21564 11756 21616
rect 3424 21471 3476 21480
rect 3424 21437 3433 21471
rect 3433 21437 3467 21471
rect 3467 21437 3476 21471
rect 3424 21428 3476 21437
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 12440 21496 12492 21548
rect 12624 21496 12676 21548
rect 20720 21564 20772 21616
rect 22468 21564 22520 21616
rect 37556 21675 37608 21684
rect 37556 21641 37565 21675
rect 37565 21641 37599 21675
rect 37599 21641 37608 21675
rect 37556 21632 37608 21641
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17960 21496 18012 21548
rect 19984 21496 20036 21548
rect 10600 21471 10652 21480
rect 10600 21437 10609 21471
rect 10609 21437 10643 21471
rect 10643 21437 10652 21471
rect 10600 21428 10652 21437
rect 12348 21471 12400 21480
rect 12348 21437 12357 21471
rect 12357 21437 12391 21471
rect 12391 21437 12400 21471
rect 12348 21428 12400 21437
rect 15844 21471 15896 21480
rect 15844 21437 15853 21471
rect 15853 21437 15887 21471
rect 15887 21437 15896 21471
rect 15844 21428 15896 21437
rect 12440 21360 12492 21412
rect 6092 21292 6144 21344
rect 8300 21292 8352 21344
rect 9956 21335 10008 21344
rect 9956 21301 9965 21335
rect 9965 21301 9999 21335
rect 9999 21301 10008 21335
rect 9956 21292 10008 21301
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 11428 21292 11480 21344
rect 17224 21360 17276 21412
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 18236 21428 18288 21480
rect 19156 21471 19208 21480
rect 19156 21437 19165 21471
rect 19165 21437 19199 21471
rect 19199 21437 19208 21471
rect 19156 21428 19208 21437
rect 18328 21360 18380 21412
rect 12716 21292 12768 21344
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 19892 21292 19944 21344
rect 20904 21292 20956 21344
rect 30196 21496 30248 21548
rect 31944 21496 31996 21548
rect 24860 21292 24912 21344
rect 27988 21292 28040 21344
rect 29276 21292 29328 21344
rect 30472 21428 30524 21480
rect 33784 21539 33836 21548
rect 33784 21505 33793 21539
rect 33793 21505 33827 21539
rect 33827 21505 33836 21539
rect 33784 21496 33836 21505
rect 34796 21539 34848 21548
rect 34796 21505 34805 21539
rect 34805 21505 34839 21539
rect 34839 21505 34848 21539
rect 34796 21496 34848 21505
rect 35440 21496 35492 21548
rect 34152 21428 34204 21480
rect 33416 21360 33468 21412
rect 30932 21292 30984 21344
rect 33876 21292 33928 21344
rect 34612 21471 34664 21480
rect 34612 21437 34646 21471
rect 34646 21437 34664 21471
rect 34612 21428 34664 21437
rect 34980 21428 35032 21480
rect 35256 21360 35308 21412
rect 37464 21471 37516 21480
rect 37464 21437 37473 21471
rect 37473 21437 37507 21471
rect 37507 21437 37516 21471
rect 37464 21428 37516 21437
rect 38016 21335 38068 21344
rect 38016 21301 38025 21335
rect 38025 21301 38059 21335
rect 38059 21301 38068 21335
rect 38016 21292 38068 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3424 21088 3476 21140
rect 10600 21088 10652 21140
rect 11060 21088 11112 21140
rect 11704 21131 11756 21140
rect 11704 21097 11713 21131
rect 11713 21097 11747 21131
rect 11747 21097 11756 21131
rect 11704 21088 11756 21097
rect 16764 21088 16816 21140
rect 17132 21088 17184 21140
rect 17868 21088 17920 21140
rect 18328 21088 18380 21140
rect 23020 21088 23072 21140
rect 3608 21063 3660 21072
rect 3608 21029 3617 21063
rect 3617 21029 3651 21063
rect 3651 21029 3660 21063
rect 3608 21020 3660 21029
rect 4896 21020 4948 21072
rect 4620 20952 4672 21004
rect 4528 20748 4580 20800
rect 5264 20952 5316 21004
rect 6644 20927 6696 20936
rect 6644 20893 6653 20927
rect 6653 20893 6687 20927
rect 6687 20893 6696 20927
rect 6644 20884 6696 20893
rect 7748 20884 7800 20936
rect 6460 20816 6512 20868
rect 8392 20816 8444 20868
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 13176 20952 13228 21004
rect 13728 20995 13780 21004
rect 13728 20961 13737 20995
rect 13737 20961 13771 20995
rect 13771 20961 13780 20995
rect 13728 20952 13780 20961
rect 19432 21020 19484 21072
rect 23204 21063 23256 21072
rect 23204 21029 23213 21063
rect 23213 21029 23247 21063
rect 23247 21029 23256 21063
rect 23204 21020 23256 21029
rect 12440 20884 12492 20936
rect 7196 20791 7248 20800
rect 7196 20757 7205 20791
rect 7205 20757 7239 20791
rect 7239 20757 7248 20791
rect 7196 20748 7248 20757
rect 8300 20748 8352 20800
rect 11060 20816 11112 20868
rect 12624 20816 12676 20868
rect 12808 20859 12860 20868
rect 12808 20825 12826 20859
rect 12826 20825 12860 20859
rect 12808 20816 12860 20825
rect 13452 20884 13504 20936
rect 13820 20884 13872 20936
rect 18788 20952 18840 21004
rect 19340 20952 19392 21004
rect 19892 20995 19944 21004
rect 19892 20961 19901 20995
rect 19901 20961 19935 20995
rect 19935 20961 19944 20995
rect 19892 20952 19944 20961
rect 20260 20952 20312 21004
rect 23572 21088 23624 21140
rect 29368 21131 29420 21140
rect 29368 21097 29377 21131
rect 29377 21097 29411 21131
rect 29411 21097 29420 21131
rect 29368 21088 29420 21097
rect 31300 21088 31352 21140
rect 32404 21088 32456 21140
rect 34152 21131 34204 21140
rect 34152 21097 34161 21131
rect 34161 21097 34195 21131
rect 34195 21097 34204 21131
rect 34152 21088 34204 21097
rect 34612 21088 34664 21140
rect 35808 21088 35860 21140
rect 36360 21088 36412 21140
rect 36728 21131 36780 21140
rect 36728 21097 36737 21131
rect 36737 21097 36771 21131
rect 36771 21097 36780 21131
rect 36728 21088 36780 21097
rect 37280 21088 37332 21140
rect 37464 21063 37516 21072
rect 37464 21029 37473 21063
rect 37473 21029 37507 21063
rect 37507 21029 37516 21063
rect 37464 21020 37516 21029
rect 16212 20816 16264 20868
rect 18604 20884 18656 20936
rect 20904 20884 20956 20936
rect 21548 20884 21600 20936
rect 22560 20884 22612 20936
rect 27252 20927 27304 20936
rect 27252 20893 27261 20927
rect 27261 20893 27295 20927
rect 27295 20893 27304 20927
rect 27252 20884 27304 20893
rect 27344 20884 27396 20936
rect 27436 20884 27488 20936
rect 21916 20816 21968 20868
rect 22836 20816 22888 20868
rect 24952 20816 25004 20868
rect 31208 20859 31260 20868
rect 31208 20825 31226 20859
rect 31226 20825 31260 20859
rect 31208 20816 31260 20825
rect 31392 20884 31444 20936
rect 34428 20927 34480 20936
rect 34428 20893 34437 20927
rect 34437 20893 34471 20927
rect 34471 20893 34480 20927
rect 34428 20884 34480 20893
rect 34704 20859 34756 20868
rect 9680 20748 9732 20800
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 13176 20791 13228 20800
rect 13176 20757 13185 20791
rect 13185 20757 13219 20791
rect 13219 20757 13228 20791
rect 13176 20748 13228 20757
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 16120 20791 16172 20800
rect 16120 20757 16129 20791
rect 16129 20757 16163 20791
rect 16163 20757 16172 20791
rect 16120 20748 16172 20757
rect 16488 20748 16540 20800
rect 18052 20748 18104 20800
rect 18236 20748 18288 20800
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 19340 20748 19392 20800
rect 26516 20791 26568 20800
rect 26516 20757 26525 20791
rect 26525 20757 26559 20791
rect 26559 20757 26568 20791
rect 26516 20748 26568 20757
rect 27896 20791 27948 20800
rect 27896 20757 27905 20791
rect 27905 20757 27939 20791
rect 27939 20757 27948 20791
rect 27896 20748 27948 20757
rect 27988 20748 28040 20800
rect 31024 20748 31076 20800
rect 34704 20825 34713 20859
rect 34713 20825 34747 20859
rect 34747 20825 34756 20859
rect 34704 20816 34756 20825
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 10416 20544 10468 20596
rect 11060 20544 11112 20596
rect 11612 20544 11664 20596
rect 12900 20544 12952 20596
rect 13544 20544 13596 20596
rect 15844 20544 15896 20596
rect 18144 20544 18196 20596
rect 18236 20544 18288 20596
rect 5264 20476 5316 20528
rect 7196 20476 7248 20528
rect 9956 20476 10008 20528
rect 5080 20408 5132 20460
rect 7472 20408 7524 20460
rect 8392 20408 8444 20460
rect 11428 20408 11480 20460
rect 11704 20408 11756 20460
rect 16120 20476 16172 20528
rect 16488 20476 16540 20528
rect 19156 20544 19208 20596
rect 19340 20544 19392 20596
rect 19984 20544 20036 20596
rect 21916 20587 21968 20596
rect 21916 20553 21925 20587
rect 21925 20553 21959 20587
rect 21959 20553 21968 20587
rect 21916 20544 21968 20553
rect 26516 20544 26568 20596
rect 30472 20544 30524 20596
rect 12256 20408 12308 20460
rect 12900 20451 12952 20460
rect 12900 20417 12934 20451
rect 12934 20417 12952 20451
rect 12900 20408 12952 20417
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 14188 20451 14240 20460
rect 14188 20417 14197 20451
rect 14197 20417 14231 20451
rect 14231 20417 14240 20451
rect 14188 20408 14240 20417
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 3884 20340 3936 20392
rect 4528 20340 4580 20392
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 6368 20340 6420 20392
rect 2504 20204 2556 20256
rect 4896 20247 4948 20256
rect 4896 20213 4905 20247
rect 4905 20213 4939 20247
rect 4939 20213 4948 20247
rect 4896 20204 4948 20213
rect 5540 20247 5592 20256
rect 5540 20213 5549 20247
rect 5549 20213 5583 20247
rect 5583 20213 5592 20247
rect 9680 20340 9732 20392
rect 12440 20340 12492 20392
rect 12532 20383 12584 20392
rect 12532 20349 12541 20383
rect 12541 20349 12575 20383
rect 12575 20349 12584 20383
rect 12532 20340 12584 20349
rect 9864 20272 9916 20324
rect 5540 20204 5592 20213
rect 7748 20204 7800 20256
rect 11980 20204 12032 20256
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 14280 20340 14332 20392
rect 13820 20204 13872 20256
rect 14556 20247 14608 20256
rect 14556 20213 14565 20247
rect 14565 20213 14599 20247
rect 14599 20213 14608 20247
rect 14556 20204 14608 20213
rect 15844 20204 15896 20256
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 18144 20451 18196 20460
rect 18144 20417 18178 20451
rect 18178 20417 18196 20451
rect 18144 20408 18196 20417
rect 18328 20451 18380 20460
rect 18328 20417 18337 20451
rect 18337 20417 18371 20451
rect 18371 20417 18380 20451
rect 18328 20408 18380 20417
rect 27712 20476 27764 20528
rect 30932 20519 30984 20528
rect 30932 20485 30972 20519
rect 30972 20485 30984 20519
rect 31208 20544 31260 20596
rect 33416 20544 33468 20596
rect 33968 20544 34020 20596
rect 34704 20544 34756 20596
rect 30932 20476 30984 20485
rect 35992 20476 36044 20528
rect 23112 20408 23164 20460
rect 27528 20408 27580 20460
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 27988 20408 28040 20417
rect 31116 20408 31168 20460
rect 33416 20408 33468 20460
rect 34612 20451 34664 20460
rect 34612 20417 34621 20451
rect 34621 20417 34655 20451
rect 34655 20417 34664 20451
rect 34612 20408 34664 20417
rect 18972 20340 19024 20392
rect 23296 20383 23348 20392
rect 23296 20349 23305 20383
rect 23305 20349 23339 20383
rect 23339 20349 23348 20383
rect 23296 20340 23348 20349
rect 23940 20383 23992 20392
rect 23940 20349 23949 20383
rect 23949 20349 23983 20383
rect 23983 20349 23992 20383
rect 23940 20340 23992 20349
rect 25780 20383 25832 20392
rect 25780 20349 25789 20383
rect 25789 20349 25823 20383
rect 25823 20349 25832 20383
rect 25780 20340 25832 20349
rect 27436 20340 27488 20392
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 22928 20272 22980 20324
rect 18052 20204 18104 20256
rect 18144 20204 18196 20256
rect 18328 20204 18380 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23388 20247 23440 20256
rect 23388 20213 23397 20247
rect 23397 20213 23431 20247
rect 23431 20213 23440 20247
rect 23388 20204 23440 20213
rect 25228 20204 25280 20256
rect 25688 20204 25740 20256
rect 25872 20247 25924 20256
rect 25872 20213 25881 20247
rect 25881 20213 25915 20247
rect 25915 20213 25924 20247
rect 25872 20204 25924 20213
rect 26976 20247 27028 20256
rect 26976 20213 26985 20247
rect 26985 20213 27019 20247
rect 27019 20213 27028 20247
rect 26976 20204 27028 20213
rect 28908 20204 28960 20256
rect 31392 20340 31444 20392
rect 31760 20340 31812 20392
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4252 20000 4304 20052
rect 4620 20000 4672 20052
rect 6644 20000 6696 20052
rect 8852 20000 8904 20052
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 11980 20043 12032 20052
rect 11980 20009 11989 20043
rect 11989 20009 12023 20043
rect 12023 20009 12032 20043
rect 11980 20000 12032 20009
rect 17960 20000 18012 20052
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 2044 19864 2096 19916
rect 4896 19864 4948 19916
rect 2504 19839 2556 19848
rect 2504 19805 2538 19839
rect 2538 19805 2556 19839
rect 2504 19796 2556 19805
rect 4620 19796 4672 19848
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 4712 19660 4764 19712
rect 5080 19660 5132 19712
rect 5356 19703 5408 19712
rect 5356 19669 5365 19703
rect 5365 19669 5399 19703
rect 5399 19669 5408 19703
rect 5356 19660 5408 19669
rect 6092 19864 6144 19916
rect 6368 19864 6420 19916
rect 9680 19864 9732 19916
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 10692 19796 10744 19848
rect 12624 19796 12676 19848
rect 14280 19796 14332 19848
rect 14556 19796 14608 19848
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19432 19864 19484 19916
rect 23204 20000 23256 20052
rect 23296 20000 23348 20052
rect 23940 20000 23992 20052
rect 22928 19864 22980 19916
rect 23112 19864 23164 19916
rect 23480 19864 23532 19916
rect 25872 20000 25924 20052
rect 27068 20000 27120 20052
rect 27252 20000 27304 20052
rect 27620 20000 27672 20052
rect 30380 20000 30432 20052
rect 31852 20000 31904 20052
rect 30656 19932 30708 19984
rect 31116 19932 31168 19984
rect 31300 19932 31352 19984
rect 26700 19864 26752 19916
rect 27896 19864 27948 19916
rect 29368 19864 29420 19916
rect 30472 19907 30524 19916
rect 30472 19873 30481 19907
rect 30481 19873 30515 19907
rect 30515 19873 30524 19907
rect 30472 19864 30524 19873
rect 15844 19796 15896 19848
rect 6276 19728 6328 19780
rect 16488 19728 16540 19780
rect 6460 19703 6512 19712
rect 6460 19669 6469 19703
rect 6469 19669 6503 19703
rect 6503 19669 6512 19703
rect 6460 19660 6512 19669
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 8576 19660 8628 19712
rect 10232 19660 10284 19712
rect 12440 19660 12492 19712
rect 12900 19660 12952 19712
rect 14004 19660 14056 19712
rect 18788 19796 18840 19848
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 22560 19796 22612 19848
rect 23296 19796 23348 19848
rect 25136 19796 25188 19848
rect 28080 19796 28132 19848
rect 30380 19839 30432 19848
rect 30380 19805 30398 19839
rect 30398 19805 30432 19839
rect 30380 19796 30432 19805
rect 31024 19796 31076 19848
rect 31300 19796 31352 19848
rect 18052 19660 18104 19712
rect 20812 19660 20864 19712
rect 21364 19660 21416 19712
rect 21732 19703 21784 19712
rect 21732 19669 21741 19703
rect 21741 19669 21775 19703
rect 21775 19669 21784 19703
rect 21732 19660 21784 19669
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 23204 19660 23256 19712
rect 25504 19660 25556 19712
rect 26976 19728 27028 19780
rect 28540 19728 28592 19780
rect 32036 19839 32088 19848
rect 32036 19805 32045 19839
rect 32045 19805 32079 19839
rect 32079 19805 32088 19839
rect 32036 19796 32088 19805
rect 34888 19796 34940 19848
rect 35348 19839 35400 19848
rect 35348 19805 35357 19839
rect 35357 19805 35391 19839
rect 35391 19805 35400 19839
rect 35348 19796 35400 19805
rect 36452 19796 36504 19848
rect 36820 19839 36872 19848
rect 36820 19805 36829 19839
rect 36829 19805 36863 19839
rect 36863 19805 36872 19839
rect 36820 19796 36872 19805
rect 38476 19839 38528 19848
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 38476 19796 38528 19805
rect 25964 19660 26016 19712
rect 27528 19660 27580 19712
rect 29920 19660 29972 19712
rect 30380 19660 30432 19712
rect 32220 19703 32272 19712
rect 32220 19669 32229 19703
rect 32229 19669 32263 19703
rect 32263 19669 32272 19703
rect 32220 19660 32272 19669
rect 32956 19703 33008 19712
rect 32956 19669 32965 19703
rect 32965 19669 32999 19703
rect 32999 19669 33008 19703
rect 32956 19660 33008 19669
rect 33784 19660 33836 19712
rect 34704 19703 34756 19712
rect 34704 19669 34713 19703
rect 34713 19669 34747 19703
rect 34747 19669 34756 19703
rect 34704 19660 34756 19669
rect 35440 19703 35492 19712
rect 35440 19669 35449 19703
rect 35449 19669 35483 19703
rect 35483 19669 35492 19703
rect 35440 19660 35492 19669
rect 36176 19703 36228 19712
rect 36176 19669 36185 19703
rect 36185 19669 36219 19703
rect 36219 19669 36228 19703
rect 36176 19660 36228 19669
rect 37832 19703 37884 19712
rect 37832 19669 37841 19703
rect 37841 19669 37875 19703
rect 37875 19669 37884 19703
rect 37832 19660 37884 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2044 19456 2096 19508
rect 2964 19320 3016 19372
rect 3424 19252 3476 19304
rect 5172 19456 5224 19508
rect 5356 19456 5408 19508
rect 9496 19456 9548 19508
rect 12256 19456 12308 19508
rect 5080 19388 5132 19440
rect 6276 19388 6328 19440
rect 6920 19388 6972 19440
rect 4252 19363 4304 19372
rect 4252 19329 4261 19363
rect 4261 19329 4295 19363
rect 4295 19329 4304 19363
rect 4252 19320 4304 19329
rect 5632 19320 5684 19372
rect 7748 19363 7800 19372
rect 4068 19184 4120 19236
rect 5172 19159 5224 19168
rect 5172 19125 5181 19159
rect 5181 19125 5215 19159
rect 5215 19125 5224 19159
rect 5172 19116 5224 19125
rect 5540 19116 5592 19168
rect 5632 19116 5684 19168
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 7748 19329 7766 19363
rect 7766 19329 7800 19363
rect 7748 19320 7800 19329
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 8668 19320 8720 19372
rect 8852 19320 8904 19372
rect 7104 19116 7156 19168
rect 7564 19295 7616 19304
rect 7564 19261 7573 19295
rect 7573 19261 7607 19295
rect 7607 19261 7616 19295
rect 7564 19252 7616 19261
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9496 19295 9548 19304
rect 9496 19261 9505 19295
rect 9505 19261 9539 19295
rect 9539 19261 9548 19295
rect 9496 19252 9548 19261
rect 12716 19499 12768 19508
rect 12716 19465 12725 19499
rect 12725 19465 12759 19499
rect 12759 19465 12768 19499
rect 12716 19456 12768 19465
rect 13084 19456 13136 19508
rect 14188 19456 14240 19508
rect 18696 19499 18748 19508
rect 18696 19465 18705 19499
rect 18705 19465 18739 19499
rect 18739 19465 18748 19499
rect 18696 19456 18748 19465
rect 21272 19456 21324 19508
rect 22192 19456 22244 19508
rect 14372 19431 14424 19440
rect 14372 19397 14381 19431
rect 14381 19397 14415 19431
rect 14415 19397 14424 19431
rect 14372 19388 14424 19397
rect 15660 19388 15712 19440
rect 11888 19252 11940 19304
rect 8300 19184 8352 19236
rect 11520 19184 11572 19236
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12900 19320 12952 19372
rect 12256 19252 12308 19304
rect 13820 19252 13872 19304
rect 14464 19252 14516 19304
rect 17408 19295 17460 19304
rect 17408 19261 17417 19295
rect 17417 19261 17451 19295
rect 17451 19261 17460 19295
rect 17408 19252 17460 19261
rect 17592 19295 17644 19304
rect 17592 19261 17601 19295
rect 17601 19261 17635 19295
rect 17635 19261 17644 19295
rect 17592 19252 17644 19261
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 18236 19320 18288 19372
rect 18880 19320 18932 19372
rect 21364 19363 21416 19372
rect 21364 19329 21373 19363
rect 21373 19329 21407 19363
rect 21407 19329 21416 19363
rect 21364 19320 21416 19329
rect 21548 19320 21600 19372
rect 22652 19388 22704 19440
rect 25228 19456 25280 19508
rect 25964 19456 26016 19508
rect 26424 19456 26476 19508
rect 26700 19499 26752 19508
rect 26700 19465 26709 19499
rect 26709 19465 26743 19499
rect 26743 19465 26752 19499
rect 26700 19456 26752 19465
rect 28080 19456 28132 19508
rect 28908 19456 28960 19508
rect 25136 19320 25188 19372
rect 27068 19320 27120 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 27896 19363 27948 19372
rect 27896 19329 27905 19363
rect 27905 19329 27939 19363
rect 27939 19329 27948 19363
rect 27896 19320 27948 19329
rect 21732 19252 21784 19304
rect 23296 19252 23348 19304
rect 12256 19159 12308 19168
rect 12256 19125 12265 19159
rect 12265 19125 12299 19159
rect 12299 19125 12308 19159
rect 12256 19116 12308 19125
rect 15844 19116 15896 19168
rect 16028 19116 16080 19168
rect 16948 19159 17000 19168
rect 16948 19125 16957 19159
rect 16957 19125 16991 19159
rect 16991 19125 17000 19159
rect 16948 19116 17000 19125
rect 22560 19116 22612 19168
rect 22836 19116 22888 19168
rect 24584 19295 24636 19304
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 24584 19252 24636 19261
rect 26884 19252 26936 19304
rect 28172 19295 28224 19304
rect 28172 19261 28181 19295
rect 28181 19261 28215 19295
rect 28215 19261 28224 19295
rect 29368 19456 29420 19508
rect 30380 19456 30432 19508
rect 32220 19456 32272 19508
rect 34704 19456 34756 19508
rect 34888 19499 34940 19508
rect 34888 19465 34897 19499
rect 34897 19465 34931 19499
rect 34931 19465 34940 19499
rect 34888 19456 34940 19465
rect 35440 19456 35492 19508
rect 36176 19456 36228 19508
rect 31024 19388 31076 19440
rect 28172 19252 28224 19261
rect 25412 19116 25464 19168
rect 28908 19184 28960 19236
rect 30932 19320 30984 19372
rect 30748 19252 30800 19304
rect 32036 19388 32088 19440
rect 31852 19363 31904 19372
rect 31852 19329 31861 19363
rect 31861 19329 31895 19363
rect 31895 19329 31904 19363
rect 31852 19320 31904 19329
rect 34704 19320 34756 19372
rect 36544 19388 36596 19440
rect 30012 19116 30064 19168
rect 31300 19159 31352 19168
rect 31300 19125 31309 19159
rect 31309 19125 31343 19159
rect 31343 19125 31352 19159
rect 31300 19116 31352 19125
rect 33324 19159 33376 19168
rect 33324 19125 33333 19159
rect 33333 19125 33367 19159
rect 33367 19125 33376 19159
rect 33324 19116 33376 19125
rect 33416 19116 33468 19168
rect 34612 19116 34664 19168
rect 35992 19252 36044 19304
rect 35348 19116 35400 19168
rect 35900 19116 35952 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4620 18955 4672 18964
rect 4620 18921 4629 18955
rect 4629 18921 4663 18955
rect 4663 18921 4672 18955
rect 4620 18912 4672 18921
rect 5172 18912 5224 18964
rect 3424 18844 3476 18896
rect 2044 18776 2096 18828
rect 4620 18776 4672 18828
rect 3792 18708 3844 18760
rect 4712 18708 4764 18760
rect 6920 18912 6972 18964
rect 7932 18912 7984 18964
rect 8576 18912 8628 18964
rect 6092 18776 6144 18828
rect 6368 18708 6420 18760
rect 8576 18708 8628 18760
rect 10048 18912 10100 18964
rect 12716 18912 12768 18964
rect 12808 18955 12860 18964
rect 12808 18921 12817 18955
rect 12817 18921 12851 18955
rect 12851 18921 12860 18955
rect 12808 18912 12860 18921
rect 16488 18955 16540 18964
rect 16488 18921 16497 18955
rect 16497 18921 16531 18955
rect 16531 18921 16540 18955
rect 16488 18912 16540 18921
rect 17408 18912 17460 18964
rect 22376 18912 22428 18964
rect 23296 18912 23348 18964
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 24308 18912 24360 18964
rect 24584 18912 24636 18964
rect 8852 18776 8904 18828
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 5080 18572 5132 18624
rect 5724 18572 5776 18624
rect 6184 18615 6236 18624
rect 6184 18581 6193 18615
rect 6193 18581 6227 18615
rect 6227 18581 6236 18615
rect 6184 18572 6236 18581
rect 6828 18572 6880 18624
rect 9220 18572 9272 18624
rect 9496 18572 9548 18624
rect 12256 18819 12308 18828
rect 12256 18785 12265 18819
rect 12265 18785 12299 18819
rect 12299 18785 12308 18819
rect 12256 18776 12308 18785
rect 16948 18776 17000 18828
rect 17960 18819 18012 18828
rect 17960 18785 17969 18819
rect 17969 18785 18003 18819
rect 18003 18785 18012 18819
rect 17960 18776 18012 18785
rect 21548 18776 21600 18828
rect 22836 18844 22888 18896
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 22928 18708 22980 18760
rect 20720 18640 20772 18692
rect 23296 18751 23348 18760
rect 23296 18717 23305 18751
rect 23305 18717 23339 18751
rect 23339 18717 23348 18751
rect 23296 18708 23348 18717
rect 24032 18683 24084 18692
rect 24032 18649 24041 18683
rect 24041 18649 24075 18683
rect 24075 18649 24084 18683
rect 25412 18912 25464 18964
rect 27344 18912 27396 18964
rect 27896 18912 27948 18964
rect 28816 18912 28868 18964
rect 30656 18912 30708 18964
rect 31760 18912 31812 18964
rect 35348 18912 35400 18964
rect 35440 18912 35492 18964
rect 35808 18912 35860 18964
rect 28724 18844 28776 18896
rect 36820 18844 36872 18896
rect 25136 18776 25188 18828
rect 28080 18819 28132 18828
rect 28080 18785 28089 18819
rect 28089 18785 28123 18819
rect 28123 18785 28132 18819
rect 28080 18776 28132 18785
rect 28816 18776 28868 18828
rect 30840 18776 30892 18828
rect 31760 18776 31812 18828
rect 25504 18751 25556 18760
rect 25504 18717 25538 18751
rect 25538 18717 25556 18751
rect 25504 18708 25556 18717
rect 28264 18708 28316 18760
rect 32956 18708 33008 18760
rect 33232 18708 33284 18760
rect 35624 18776 35676 18828
rect 35900 18776 35952 18828
rect 36728 18776 36780 18828
rect 38476 18955 38528 18964
rect 38476 18921 38485 18955
rect 38485 18921 38519 18955
rect 38519 18921 38528 18955
rect 38476 18912 38528 18921
rect 24032 18640 24084 18649
rect 10508 18572 10560 18624
rect 17592 18572 17644 18624
rect 20076 18572 20128 18624
rect 22652 18572 22704 18624
rect 22744 18572 22796 18624
rect 25596 18572 25648 18624
rect 27160 18572 27212 18624
rect 27436 18572 27488 18624
rect 27528 18572 27580 18624
rect 29552 18615 29604 18624
rect 29552 18581 29561 18615
rect 29561 18581 29595 18615
rect 29595 18581 29604 18615
rect 29552 18572 29604 18581
rect 31300 18640 31352 18692
rect 33324 18640 33376 18692
rect 30196 18572 30248 18624
rect 30932 18572 30984 18624
rect 33048 18615 33100 18624
rect 33048 18581 33057 18615
rect 33057 18581 33091 18615
rect 33091 18581 33100 18615
rect 36084 18751 36136 18760
rect 36084 18717 36093 18751
rect 36093 18717 36127 18751
rect 36127 18717 36136 18751
rect 36084 18708 36136 18717
rect 37372 18683 37424 18692
rect 37372 18649 37406 18683
rect 37406 18649 37424 18683
rect 37372 18640 37424 18649
rect 33048 18572 33100 18581
rect 34612 18572 34664 18624
rect 37648 18572 37700 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2044 18232 2096 18284
rect 3332 18232 3384 18284
rect 4160 18368 4212 18420
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 7564 18368 7616 18420
rect 7840 18368 7892 18420
rect 10048 18368 10100 18420
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 12348 18368 12400 18420
rect 4068 18300 4120 18352
rect 20904 18300 20956 18352
rect 6368 18275 6420 18284
rect 6368 18241 6377 18275
rect 6377 18241 6411 18275
rect 6411 18241 6420 18275
rect 6368 18232 6420 18241
rect 6644 18275 6696 18284
rect 6644 18241 6678 18275
rect 6678 18241 6696 18275
rect 6644 18232 6696 18241
rect 20076 18232 20128 18284
rect 20812 18232 20864 18284
rect 22100 18300 22152 18352
rect 23664 18368 23716 18420
rect 25780 18411 25832 18420
rect 25780 18377 25789 18411
rect 25789 18377 25823 18411
rect 25823 18377 25832 18411
rect 25780 18368 25832 18377
rect 27528 18368 27580 18420
rect 28264 18368 28316 18420
rect 28540 18368 28592 18420
rect 29552 18368 29604 18420
rect 29920 18411 29972 18420
rect 29920 18377 29929 18411
rect 29929 18377 29963 18411
rect 29963 18377 29972 18411
rect 29920 18368 29972 18377
rect 30012 18411 30064 18420
rect 30012 18377 30021 18411
rect 30021 18377 30055 18411
rect 30055 18377 30064 18411
rect 30012 18368 30064 18377
rect 35440 18368 35492 18420
rect 36820 18368 36872 18420
rect 37832 18368 37884 18420
rect 22836 18300 22888 18352
rect 23388 18300 23440 18352
rect 24032 18300 24084 18352
rect 26332 18300 26384 18352
rect 23296 18232 23348 18284
rect 4252 18164 4304 18216
rect 11336 18207 11388 18216
rect 11336 18173 11345 18207
rect 11345 18173 11379 18207
rect 11379 18173 11388 18207
rect 11336 18164 11388 18173
rect 4712 18096 4764 18148
rect 12256 18164 12308 18216
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 15660 18207 15712 18216
rect 15660 18173 15669 18207
rect 15669 18173 15703 18207
rect 15703 18173 15712 18207
rect 15660 18164 15712 18173
rect 16488 18207 16540 18216
rect 16488 18173 16497 18207
rect 16497 18173 16531 18207
rect 16531 18173 16540 18207
rect 16488 18164 16540 18173
rect 17776 18207 17828 18216
rect 17776 18173 17785 18207
rect 17785 18173 17819 18207
rect 17819 18173 17828 18207
rect 17776 18164 17828 18173
rect 23204 18207 23256 18216
rect 23204 18173 23213 18207
rect 23213 18173 23247 18207
rect 23247 18173 23256 18207
rect 23204 18164 23256 18173
rect 6092 18071 6144 18080
rect 6092 18037 6101 18071
rect 6101 18037 6135 18071
rect 6135 18037 6144 18071
rect 6092 18028 6144 18037
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 10232 18028 10284 18080
rect 14740 18096 14792 18148
rect 10692 18071 10744 18080
rect 10692 18037 10701 18071
rect 10701 18037 10735 18071
rect 10735 18037 10744 18071
rect 10692 18028 10744 18037
rect 12348 18071 12400 18080
rect 12348 18037 12357 18071
rect 12357 18037 12391 18071
rect 12391 18037 12400 18071
rect 12348 18028 12400 18037
rect 15016 18028 15068 18080
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 17224 18071 17276 18080
rect 17224 18037 17233 18071
rect 17233 18037 17267 18071
rect 17267 18037 17276 18071
rect 17224 18028 17276 18037
rect 17868 18028 17920 18080
rect 24584 18275 24636 18284
rect 24584 18241 24593 18275
rect 24593 18241 24627 18275
rect 24627 18241 24636 18275
rect 24584 18232 24636 18241
rect 33232 18300 33284 18352
rect 33784 18275 33836 18284
rect 33784 18241 33818 18275
rect 33818 18241 33836 18275
rect 33784 18232 33836 18241
rect 35624 18300 35676 18352
rect 36176 18300 36228 18352
rect 36544 18300 36596 18352
rect 25596 18164 25648 18216
rect 26516 18164 26568 18216
rect 27436 18164 27488 18216
rect 29000 18164 29052 18216
rect 29736 18207 29788 18216
rect 29736 18173 29745 18207
rect 29745 18173 29779 18207
rect 29779 18173 29788 18207
rect 29736 18164 29788 18173
rect 37556 18164 37608 18216
rect 37832 18207 37884 18216
rect 37832 18173 37841 18207
rect 37841 18173 37875 18207
rect 37875 18173 37884 18207
rect 37832 18164 37884 18173
rect 27712 18096 27764 18148
rect 28724 18071 28776 18080
rect 28724 18037 28733 18071
rect 28733 18037 28767 18071
rect 28767 18037 28776 18071
rect 28724 18028 28776 18037
rect 30380 18071 30432 18080
rect 30380 18037 30389 18071
rect 30389 18037 30423 18071
rect 30423 18037 30432 18071
rect 30380 18028 30432 18037
rect 30748 18071 30800 18080
rect 30748 18037 30757 18071
rect 30757 18037 30791 18071
rect 30791 18037 30800 18071
rect 30748 18028 30800 18037
rect 36084 18028 36136 18080
rect 36452 18028 36504 18080
rect 36728 18071 36780 18080
rect 36728 18037 36737 18071
rect 36737 18037 36771 18071
rect 36771 18037 36780 18071
rect 36728 18028 36780 18037
rect 37280 18071 37332 18080
rect 37280 18037 37289 18071
rect 37289 18037 37323 18071
rect 37323 18037 37332 18071
rect 37280 18028 37332 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2964 17867 3016 17876
rect 2964 17833 2973 17867
rect 2973 17833 3007 17867
rect 3007 17833 3016 17867
rect 2964 17824 3016 17833
rect 3332 17824 3384 17876
rect 6644 17824 6696 17876
rect 15660 17824 15712 17876
rect 17776 17824 17828 17876
rect 20904 17867 20956 17876
rect 20904 17833 20913 17867
rect 20913 17833 20947 17867
rect 20947 17833 20956 17867
rect 20904 17824 20956 17833
rect 6828 17756 6880 17808
rect 3792 17688 3844 17740
rect 4712 17688 4764 17740
rect 6184 17688 6236 17740
rect 7840 17731 7892 17740
rect 7840 17697 7849 17731
rect 7849 17697 7883 17731
rect 7883 17697 7892 17731
rect 7840 17688 7892 17697
rect 10692 17731 10744 17740
rect 10692 17697 10701 17731
rect 10701 17697 10735 17731
rect 10735 17697 10744 17731
rect 10692 17688 10744 17697
rect 10048 17620 10100 17672
rect 12348 17620 12400 17672
rect 12716 17731 12768 17740
rect 12716 17697 12725 17731
rect 12725 17697 12759 17731
rect 12759 17697 12768 17731
rect 12716 17688 12768 17697
rect 14740 17688 14792 17740
rect 4620 17552 4672 17604
rect 18144 17756 18196 17808
rect 16028 17620 16080 17672
rect 4160 17484 4212 17536
rect 5172 17484 5224 17536
rect 5264 17484 5316 17536
rect 10048 17484 10100 17536
rect 17500 17552 17552 17604
rect 18604 17552 18656 17604
rect 11060 17527 11112 17536
rect 11060 17493 11069 17527
rect 11069 17493 11103 17527
rect 11103 17493 11112 17527
rect 11060 17484 11112 17493
rect 12440 17484 12492 17536
rect 12900 17527 12952 17536
rect 12900 17493 12909 17527
rect 12909 17493 12943 17527
rect 12943 17493 12952 17527
rect 12900 17484 12952 17493
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 14740 17484 14792 17536
rect 15476 17527 15528 17536
rect 15476 17493 15485 17527
rect 15485 17493 15519 17527
rect 15519 17493 15528 17527
rect 15476 17484 15528 17493
rect 16580 17484 16632 17536
rect 24952 17824 25004 17876
rect 26332 17867 26384 17876
rect 26332 17833 26341 17867
rect 26341 17833 26375 17867
rect 26375 17833 26384 17867
rect 26332 17824 26384 17833
rect 26792 17824 26844 17876
rect 22468 17688 22520 17740
rect 23664 17688 23716 17740
rect 24308 17688 24360 17740
rect 26884 17731 26936 17740
rect 26884 17697 26893 17731
rect 26893 17697 26927 17731
rect 26927 17697 26936 17731
rect 26884 17688 26936 17697
rect 28172 17688 28224 17740
rect 37372 17867 37424 17876
rect 37372 17833 37381 17867
rect 37381 17833 37415 17867
rect 37415 17833 37424 17867
rect 37372 17824 37424 17833
rect 37832 17756 37884 17808
rect 19432 17552 19484 17604
rect 21364 17552 21416 17604
rect 18972 17484 19024 17536
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 22652 17595 22704 17604
rect 22652 17561 22661 17595
rect 22661 17561 22695 17595
rect 22695 17561 22704 17595
rect 22652 17552 22704 17561
rect 24492 17552 24544 17604
rect 25688 17620 25740 17672
rect 27712 17663 27764 17672
rect 27712 17629 27721 17663
rect 27721 17629 27755 17663
rect 27755 17629 27764 17663
rect 27712 17620 27764 17629
rect 28264 17620 28316 17672
rect 28632 17620 28684 17672
rect 35256 17688 35308 17740
rect 35348 17731 35400 17740
rect 35348 17697 35357 17731
rect 35357 17697 35391 17731
rect 35391 17697 35400 17731
rect 35348 17688 35400 17697
rect 36544 17688 36596 17740
rect 37280 17688 37332 17740
rect 36176 17620 36228 17672
rect 36452 17620 36504 17672
rect 36912 17663 36964 17672
rect 36912 17629 36921 17663
rect 36921 17629 36955 17663
rect 36955 17629 36964 17663
rect 36912 17620 36964 17629
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 22008 17484 22060 17536
rect 22744 17484 22796 17536
rect 34980 17552 35032 17604
rect 36084 17552 36136 17604
rect 29000 17484 29052 17536
rect 29184 17484 29236 17536
rect 29736 17527 29788 17536
rect 29736 17493 29745 17527
rect 29745 17493 29779 17527
rect 29779 17493 29788 17527
rect 29736 17484 29788 17493
rect 33324 17527 33376 17536
rect 33324 17493 33333 17527
rect 33333 17493 33367 17527
rect 33367 17493 33376 17527
rect 33324 17484 33376 17493
rect 33784 17527 33836 17536
rect 33784 17493 33793 17527
rect 33793 17493 33827 17527
rect 33827 17493 33836 17527
rect 33784 17484 33836 17493
rect 33876 17527 33928 17536
rect 33876 17493 33885 17527
rect 33885 17493 33919 17527
rect 33919 17493 33928 17527
rect 33876 17484 33928 17493
rect 34704 17484 34756 17536
rect 36268 17527 36320 17536
rect 36268 17493 36277 17527
rect 36277 17493 36311 17527
rect 36311 17493 36320 17527
rect 36268 17484 36320 17493
rect 37556 17484 37608 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4988 17280 5040 17332
rect 4620 17255 4672 17264
rect 4620 17221 4629 17255
rect 4629 17221 4663 17255
rect 4663 17221 4672 17255
rect 26792 17280 26844 17332
rect 29000 17280 29052 17332
rect 29092 17280 29144 17332
rect 33876 17280 33928 17332
rect 36084 17280 36136 17332
rect 36912 17280 36964 17332
rect 37648 17323 37700 17332
rect 37648 17289 37657 17323
rect 37657 17289 37691 17323
rect 37691 17289 37700 17323
rect 37648 17280 37700 17289
rect 4620 17212 4672 17221
rect 7840 17212 7892 17264
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 10048 17144 10100 17196
rect 3424 17119 3476 17128
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 4712 17076 4764 17128
rect 7012 17076 7064 17128
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 8392 17076 8444 17128
rect 2780 16983 2832 16992
rect 2780 16949 2789 16983
rect 2789 16949 2823 16983
rect 2823 16949 2832 16983
rect 2780 16940 2832 16949
rect 3148 16940 3200 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 6920 16983 6972 16992
rect 6920 16949 6929 16983
rect 6929 16949 6963 16983
rect 6963 16949 6972 16983
rect 6920 16940 6972 16949
rect 7656 16983 7708 16992
rect 7656 16949 7665 16983
rect 7665 16949 7699 16983
rect 7699 16949 7708 16983
rect 7656 16940 7708 16949
rect 8484 17008 8536 17060
rect 8668 17051 8720 17060
rect 8668 17017 8677 17051
rect 8677 17017 8711 17051
rect 8711 17017 8720 17051
rect 8668 17008 8720 17017
rect 9864 17008 9916 17060
rect 13268 17212 13320 17264
rect 15476 17212 15528 17264
rect 18604 17255 18656 17264
rect 18604 17221 18613 17255
rect 18613 17221 18647 17255
rect 18647 17221 18656 17255
rect 18604 17212 18656 17221
rect 20720 17212 20772 17264
rect 21456 17212 21508 17264
rect 21916 17212 21968 17264
rect 33048 17212 33100 17264
rect 15200 17144 15252 17196
rect 15384 17187 15436 17196
rect 15384 17153 15418 17187
rect 15418 17153 15436 17187
rect 15384 17144 15436 17153
rect 17307 17187 17359 17196
rect 17307 17153 17315 17187
rect 17315 17153 17349 17187
rect 17349 17153 17359 17187
rect 17307 17144 17359 17153
rect 18144 17144 18196 17196
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 22376 17187 22428 17196
rect 22376 17153 22385 17187
rect 22385 17153 22419 17187
rect 22419 17153 22428 17187
rect 22376 17144 22428 17153
rect 29920 17144 29972 17196
rect 35256 17212 35308 17264
rect 36084 17187 36136 17196
rect 36084 17153 36118 17187
rect 36118 17153 36136 17187
rect 36084 17144 36136 17153
rect 11060 17076 11112 17128
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 10968 17008 11020 17060
rect 9312 16940 9364 16992
rect 9956 16940 10008 16992
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 12624 17076 12676 17128
rect 13084 17076 13136 17128
rect 13268 17008 13320 17060
rect 11336 16940 11388 16949
rect 13360 16983 13412 16992
rect 13360 16949 13369 16983
rect 13369 16949 13403 16983
rect 13403 16949 13412 16983
rect 13360 16940 13412 16949
rect 15108 17119 15160 17128
rect 15108 17085 15117 17119
rect 15117 17085 15151 17119
rect 15151 17085 15160 17119
rect 15108 17076 15160 17085
rect 16212 17076 16264 17128
rect 16488 17051 16540 17060
rect 16488 17017 16497 17051
rect 16497 17017 16531 17051
rect 16531 17017 16540 17051
rect 16488 17008 16540 17017
rect 16304 16940 16356 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 23388 17076 23440 17128
rect 23848 17119 23900 17128
rect 23848 17085 23857 17119
rect 23857 17085 23891 17119
rect 23891 17085 23900 17119
rect 23848 17076 23900 17085
rect 26516 17076 26568 17128
rect 27436 17076 27488 17128
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 27896 17076 27948 17128
rect 33140 17076 33192 17128
rect 35440 17076 35492 17128
rect 35624 17076 35676 17128
rect 36452 17076 36504 17128
rect 38108 17076 38160 17128
rect 17868 17051 17920 17060
rect 17868 17017 17877 17051
rect 17877 17017 17911 17051
rect 17911 17017 17920 17051
rect 17868 17008 17920 17017
rect 24584 17008 24636 17060
rect 22560 16983 22612 16992
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 23296 16983 23348 16992
rect 23296 16949 23305 16983
rect 23305 16949 23339 16983
rect 23339 16949 23348 16983
rect 23296 16940 23348 16949
rect 24308 16983 24360 16992
rect 24308 16949 24317 16983
rect 24317 16949 24351 16983
rect 24351 16949 24360 16983
rect 24308 16940 24360 16949
rect 25504 16940 25556 16992
rect 26240 16940 26292 16992
rect 26792 16940 26844 16992
rect 27068 16940 27120 16992
rect 30932 16940 30984 16992
rect 36728 16940 36780 16992
rect 38200 16940 38252 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3148 16736 3200 16788
rect 3424 16736 3476 16788
rect 7012 16779 7064 16788
rect 7012 16745 7021 16779
rect 7021 16745 7055 16779
rect 7055 16745 7064 16779
rect 7012 16736 7064 16745
rect 7564 16736 7616 16788
rect 9956 16736 10008 16788
rect 12440 16736 12492 16788
rect 2964 16643 3016 16652
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 4528 16600 4580 16652
rect 7104 16600 7156 16652
rect 8668 16600 8720 16652
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 3884 16532 3936 16584
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 6184 16532 6236 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 10508 16532 10560 16584
rect 12900 16779 12952 16788
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 15108 16736 15160 16788
rect 15200 16736 15252 16788
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 16304 16736 16356 16788
rect 17316 16736 17368 16788
rect 18328 16736 18380 16788
rect 20168 16736 20220 16788
rect 23848 16736 23900 16788
rect 16028 16600 16080 16652
rect 22560 16600 22612 16652
rect 24952 16736 25004 16788
rect 11704 16532 11756 16584
rect 13636 16532 13688 16584
rect 15108 16575 15160 16584
rect 15108 16541 15142 16575
rect 15142 16541 15160 16575
rect 15108 16532 15160 16541
rect 17224 16532 17276 16584
rect 17500 16532 17552 16584
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 2412 16464 2464 16516
rect 2596 16396 2648 16448
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 4804 16464 4856 16516
rect 5448 16396 5500 16448
rect 7748 16396 7800 16448
rect 13268 16464 13320 16516
rect 12716 16396 12768 16448
rect 17592 16464 17644 16516
rect 25044 16532 25096 16584
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 21272 16507 21324 16516
rect 21272 16473 21281 16507
rect 21281 16473 21315 16507
rect 21315 16473 21324 16507
rect 21272 16464 21324 16473
rect 23572 16396 23624 16448
rect 26056 16600 26108 16652
rect 26424 16736 26476 16788
rect 26240 16668 26292 16720
rect 27988 16668 28040 16720
rect 29552 16668 29604 16720
rect 27068 16600 27120 16652
rect 27436 16643 27488 16652
rect 27436 16609 27445 16643
rect 27445 16609 27479 16643
rect 27479 16609 27488 16643
rect 27436 16600 27488 16609
rect 28264 16643 28316 16652
rect 28264 16609 28273 16643
rect 28273 16609 28307 16643
rect 28307 16609 28316 16643
rect 28264 16600 28316 16609
rect 28540 16600 28592 16652
rect 33140 16643 33192 16652
rect 26332 16464 26384 16516
rect 30380 16532 30432 16584
rect 33140 16609 33149 16643
rect 33149 16609 33183 16643
rect 33183 16609 33192 16643
rect 33140 16600 33192 16609
rect 36176 16600 36228 16652
rect 32588 16575 32640 16584
rect 32588 16541 32597 16575
rect 32597 16541 32631 16575
rect 32631 16541 32640 16575
rect 32588 16532 32640 16541
rect 35440 16532 35492 16584
rect 37740 16532 37792 16584
rect 38384 16575 38436 16584
rect 38384 16541 38393 16575
rect 38393 16541 38427 16575
rect 38427 16541 38436 16575
rect 38384 16532 38436 16541
rect 33876 16464 33928 16516
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 27620 16396 27672 16448
rect 27988 16396 28040 16448
rect 28080 16439 28132 16448
rect 28080 16405 28089 16439
rect 28089 16405 28123 16439
rect 28123 16405 28132 16439
rect 28080 16396 28132 16405
rect 29092 16396 29144 16448
rect 31852 16439 31904 16448
rect 31852 16405 31861 16439
rect 31861 16405 31895 16439
rect 31895 16405 31904 16439
rect 31852 16396 31904 16405
rect 35624 16464 35676 16516
rect 36084 16464 36136 16516
rect 35348 16396 35400 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3792 16192 3844 16244
rect 4988 16192 5040 16244
rect 5540 16192 5592 16244
rect 2780 16124 2832 16176
rect 4528 16124 4580 16176
rect 5264 16124 5316 16176
rect 6920 16124 6972 16176
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 4620 16056 4672 16108
rect 5356 16056 5408 16108
rect 5448 15988 5500 16040
rect 6000 15920 6052 15972
rect 6184 15988 6236 16040
rect 6368 15920 6420 15972
rect 3056 15852 3108 15904
rect 4712 15852 4764 15904
rect 7748 16192 7800 16244
rect 8392 16192 8444 16244
rect 8484 16192 8536 16244
rect 9864 16192 9916 16244
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 9220 15988 9272 16040
rect 12256 16192 12308 16244
rect 15844 16192 15896 16244
rect 16580 16192 16632 16244
rect 18696 16192 18748 16244
rect 18880 16192 18932 16244
rect 16948 16124 17000 16176
rect 18420 16124 18472 16176
rect 23296 16192 23348 16244
rect 11060 16056 11112 16108
rect 12532 16056 12584 16108
rect 18144 16099 18196 16108
rect 18144 16065 18153 16099
rect 18153 16065 18187 16099
rect 18187 16065 18196 16099
rect 18144 16056 18196 16065
rect 23204 16056 23256 16108
rect 26240 16124 26292 16176
rect 29552 16192 29604 16244
rect 34704 16235 34756 16244
rect 34704 16201 34713 16235
rect 34713 16201 34747 16235
rect 34747 16201 34756 16235
rect 34704 16192 34756 16201
rect 35992 16235 36044 16244
rect 35992 16201 36001 16235
rect 36001 16201 36035 16235
rect 36035 16201 36044 16235
rect 35992 16192 36044 16201
rect 36084 16235 36136 16244
rect 36084 16201 36093 16235
rect 36093 16201 36127 16235
rect 36127 16201 36136 16235
rect 36084 16192 36136 16201
rect 37188 16192 37240 16244
rect 38384 16192 38436 16244
rect 8208 15920 8260 15972
rect 16212 15988 16264 16040
rect 16764 16031 16816 16040
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 26148 16056 26200 16108
rect 28632 16167 28684 16176
rect 28632 16133 28641 16167
rect 28641 16133 28675 16167
rect 28675 16133 28684 16167
rect 28632 16124 28684 16133
rect 31852 16124 31904 16176
rect 27712 16056 27764 16108
rect 35348 16099 35400 16108
rect 35348 16065 35357 16099
rect 35357 16065 35391 16099
rect 35391 16065 35400 16099
rect 35348 16056 35400 16065
rect 36268 16056 36320 16108
rect 24952 15988 25004 16040
rect 29736 15988 29788 16040
rect 30380 15988 30432 16040
rect 32404 15988 32456 16040
rect 31576 15920 31628 15972
rect 34796 16031 34848 16040
rect 34796 15997 34805 16031
rect 34805 15997 34839 16031
rect 34839 15997 34848 16031
rect 34796 15988 34848 15997
rect 35716 15988 35768 16040
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 37372 16031 37424 16040
rect 37372 15997 37381 16031
rect 37381 15997 37415 16031
rect 37415 15997 37424 16031
rect 37372 15988 37424 15997
rect 37556 16031 37608 16040
rect 37556 15997 37565 16031
rect 37565 15997 37599 16031
rect 37599 15997 37608 16031
rect 37556 15988 37608 15997
rect 38384 15988 38436 16040
rect 8852 15852 8904 15904
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 23296 15852 23348 15904
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 28448 15852 28500 15904
rect 32864 15895 32916 15904
rect 32864 15861 32873 15895
rect 32873 15861 32907 15895
rect 32907 15861 32916 15895
rect 32864 15852 32916 15861
rect 32956 15852 33008 15904
rect 33600 15895 33652 15904
rect 33600 15861 33609 15895
rect 33609 15861 33643 15895
rect 33643 15861 33652 15895
rect 33600 15852 33652 15861
rect 34336 15895 34388 15904
rect 34336 15861 34345 15895
rect 34345 15861 34379 15895
rect 34379 15861 34388 15895
rect 34336 15852 34388 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 4804 15648 4856 15700
rect 9772 15648 9824 15700
rect 15384 15648 15436 15700
rect 15752 15648 15804 15700
rect 3608 15580 3660 15632
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 7840 15580 7892 15632
rect 2320 15444 2372 15496
rect 2780 15444 2832 15496
rect 2596 15376 2648 15428
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 2412 15308 2464 15360
rect 3332 15308 3384 15360
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 4160 15308 4212 15360
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 6460 15351 6512 15360
rect 6460 15317 6469 15351
rect 6469 15317 6503 15351
rect 6503 15317 6512 15351
rect 6460 15308 6512 15317
rect 6920 15512 6972 15564
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 8208 15512 8260 15564
rect 8484 15512 8536 15564
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 13820 15512 13872 15564
rect 11244 15444 11296 15453
rect 12532 15444 12584 15496
rect 12900 15444 12952 15496
rect 13544 15444 13596 15496
rect 17040 15648 17092 15700
rect 17500 15580 17552 15632
rect 16672 15512 16724 15564
rect 16948 15555 17000 15564
rect 16948 15521 16957 15555
rect 16957 15521 16991 15555
rect 16991 15521 17000 15555
rect 16948 15512 17000 15521
rect 17040 15555 17092 15564
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 7104 15308 7156 15360
rect 9312 15376 9364 15428
rect 9956 15419 10008 15428
rect 9956 15385 9965 15419
rect 9965 15385 9999 15419
rect 9999 15385 10008 15419
rect 9956 15376 10008 15385
rect 12808 15376 12860 15428
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 9680 15308 9732 15360
rect 11612 15308 11664 15360
rect 13912 15308 13964 15360
rect 15476 15419 15528 15428
rect 15476 15385 15485 15419
rect 15485 15385 15519 15419
rect 15519 15385 15528 15419
rect 18420 15512 18472 15564
rect 22836 15512 22888 15564
rect 23388 15512 23440 15564
rect 23572 15555 23624 15564
rect 23572 15521 23581 15555
rect 23581 15521 23615 15555
rect 23615 15521 23624 15555
rect 23572 15512 23624 15521
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 23204 15444 23256 15496
rect 24308 15444 24360 15496
rect 15476 15376 15528 15385
rect 20076 15376 20128 15428
rect 21916 15419 21968 15428
rect 21916 15385 21950 15419
rect 21950 15385 21968 15419
rect 21916 15376 21968 15385
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 17316 15351 17368 15360
rect 17316 15317 17325 15351
rect 17325 15317 17359 15351
rect 17359 15317 17368 15351
rect 17316 15308 17368 15317
rect 17408 15308 17460 15360
rect 18420 15351 18472 15360
rect 18420 15317 18429 15351
rect 18429 15317 18463 15351
rect 18463 15317 18472 15351
rect 18420 15308 18472 15317
rect 19340 15308 19392 15360
rect 20444 15308 20496 15360
rect 23112 15351 23164 15360
rect 23112 15317 23121 15351
rect 23121 15317 23155 15351
rect 23155 15317 23164 15351
rect 23112 15308 23164 15317
rect 23848 15308 23900 15360
rect 23940 15308 23992 15360
rect 25688 15555 25740 15564
rect 25688 15521 25697 15555
rect 25697 15521 25731 15555
rect 25731 15521 25740 15555
rect 25688 15512 25740 15521
rect 26240 15648 26292 15700
rect 27804 15648 27856 15700
rect 28540 15648 28592 15700
rect 29092 15648 29144 15700
rect 30104 15648 30156 15700
rect 27896 15580 27948 15632
rect 26792 15444 26844 15496
rect 31852 15580 31904 15632
rect 30288 15555 30340 15564
rect 30288 15521 30297 15555
rect 30297 15521 30331 15555
rect 30331 15521 30340 15555
rect 30288 15512 30340 15521
rect 30932 15512 30984 15564
rect 31392 15555 31444 15564
rect 31392 15521 31401 15555
rect 31401 15521 31435 15555
rect 31435 15521 31444 15555
rect 31392 15512 31444 15521
rect 31576 15512 31628 15564
rect 33876 15691 33928 15700
rect 33876 15657 33885 15691
rect 33885 15657 33919 15691
rect 33919 15657 33928 15691
rect 33876 15648 33928 15657
rect 34336 15648 34388 15700
rect 34796 15648 34848 15700
rect 35624 15648 35676 15700
rect 35716 15691 35768 15700
rect 35716 15657 35725 15691
rect 35725 15657 35759 15691
rect 35759 15657 35768 15691
rect 35716 15648 35768 15657
rect 36360 15691 36412 15700
rect 36360 15657 36369 15691
rect 36369 15657 36403 15691
rect 36403 15657 36412 15691
rect 36360 15648 36412 15657
rect 37648 15648 37700 15700
rect 33140 15580 33192 15632
rect 29736 15444 29788 15496
rect 31208 15444 31260 15496
rect 32312 15487 32364 15496
rect 32312 15453 32321 15487
rect 32321 15453 32355 15487
rect 32355 15453 32364 15487
rect 32312 15444 32364 15453
rect 28816 15376 28868 15428
rect 30564 15376 30616 15428
rect 32680 15512 32732 15564
rect 33324 15512 33376 15564
rect 37740 15512 37792 15564
rect 36452 15419 36504 15428
rect 36452 15385 36461 15419
rect 36461 15385 36495 15419
rect 36495 15385 36504 15419
rect 36452 15376 36504 15385
rect 25228 15308 25280 15360
rect 29920 15308 29972 15360
rect 30104 15351 30156 15360
rect 30104 15317 30113 15351
rect 30113 15317 30147 15351
rect 30147 15317 30156 15351
rect 30104 15308 30156 15317
rect 32128 15308 32180 15360
rect 32496 15308 32548 15360
rect 33232 15308 33284 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1584 15036 1636 15088
rect 2412 15079 2464 15088
rect 2412 15045 2421 15079
rect 2421 15045 2455 15079
rect 2455 15045 2464 15079
rect 2412 15036 2464 15045
rect 3056 15079 3108 15088
rect 3056 15045 3068 15079
rect 3068 15045 3108 15079
rect 3056 15036 3108 15045
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 4436 15104 4488 15156
rect 4896 15036 4948 15088
rect 5632 15104 5684 15156
rect 6460 15104 6512 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 7840 15104 7892 15156
rect 8208 15104 8260 15156
rect 8392 15104 8444 15156
rect 10968 15147 11020 15156
rect 10968 15113 10977 15147
rect 10977 15113 11011 15147
rect 11011 15113 11020 15147
rect 10968 15104 11020 15113
rect 2872 14968 2924 15020
rect 4436 15011 4488 15020
rect 4436 14977 4445 15011
rect 4445 14977 4479 15011
rect 4479 14977 4488 15011
rect 4436 14968 4488 14977
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 7656 15036 7708 15088
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 4252 14764 4304 14816
rect 4804 14764 4856 14816
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 9312 14968 9364 15020
rect 6092 14900 6144 14909
rect 6184 14832 6236 14884
rect 8484 14943 8536 14952
rect 8484 14909 8493 14943
rect 8493 14909 8527 14943
rect 8527 14909 8536 14943
rect 8484 14900 8536 14909
rect 8576 14900 8628 14952
rect 11336 14900 11388 14952
rect 12440 15036 12492 15088
rect 12900 15147 12952 15156
rect 12900 15113 12909 15147
rect 12909 15113 12943 15147
rect 12943 15113 12952 15147
rect 12900 15104 12952 15113
rect 13360 15104 13412 15156
rect 11612 14968 11664 15020
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 15476 15104 15528 15156
rect 16856 15104 16908 15156
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 17960 15104 18012 15156
rect 19524 15104 19576 15156
rect 20076 15104 20128 15156
rect 21916 15104 21968 15156
rect 16488 14968 16540 15020
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 17868 14900 17920 14952
rect 18512 14900 18564 14952
rect 18604 14943 18656 14952
rect 18604 14909 18613 14943
rect 18613 14909 18647 14943
rect 18647 14909 18656 14943
rect 18604 14900 18656 14909
rect 8208 14764 8260 14816
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 12992 14832 13044 14884
rect 17408 14832 17460 14884
rect 12256 14764 12308 14816
rect 13084 14764 13136 14816
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 16672 14764 16724 14816
rect 17040 14764 17092 14816
rect 19248 14943 19300 14952
rect 19248 14909 19257 14943
rect 19257 14909 19291 14943
rect 19291 14909 19300 14943
rect 19248 14900 19300 14909
rect 20444 15011 20496 15020
rect 20444 14977 20473 15011
rect 20473 14977 20496 15011
rect 20444 14968 20496 14977
rect 20720 15011 20772 15020
rect 20720 14977 20729 15011
rect 20729 14977 20763 15011
rect 20763 14977 20772 15011
rect 20720 14968 20772 14977
rect 21640 14968 21692 15020
rect 23112 15104 23164 15156
rect 23756 15104 23808 15156
rect 26056 15036 26108 15088
rect 23756 15011 23808 15020
rect 23756 14977 23765 15011
rect 23765 14977 23799 15011
rect 23799 14977 23808 15011
rect 23756 14968 23808 14977
rect 22284 14900 22336 14952
rect 22744 14943 22796 14952
rect 22744 14909 22753 14943
rect 22753 14909 22787 14943
rect 22787 14909 22796 14943
rect 22744 14900 22796 14909
rect 23296 14900 23348 14952
rect 23664 14900 23716 14952
rect 19708 14764 19760 14816
rect 22652 14832 22704 14884
rect 23756 14764 23808 14816
rect 24768 14968 24820 15020
rect 25228 14900 25280 14952
rect 26056 14943 26108 14952
rect 26056 14909 26065 14943
rect 26065 14909 26099 14943
rect 26099 14909 26108 14943
rect 26056 14900 26108 14909
rect 26700 15104 26752 15156
rect 30288 15104 30340 15156
rect 31484 15104 31536 15156
rect 32404 15104 32456 15156
rect 32864 15104 32916 15156
rect 33600 15104 33652 15156
rect 34244 15104 34296 15156
rect 34428 15147 34480 15156
rect 34428 15113 34437 15147
rect 34437 15113 34471 15147
rect 34471 15113 34480 15147
rect 34428 15104 34480 15113
rect 37372 15104 37424 15156
rect 38292 15147 38344 15156
rect 38292 15113 38301 15147
rect 38301 15113 38335 15147
rect 38335 15113 38344 15147
rect 38292 15104 38344 15113
rect 38568 15104 38620 15156
rect 29552 15036 29604 15088
rect 27804 15011 27856 15020
rect 27804 14977 27822 15011
rect 27822 14977 27856 15011
rect 27804 14968 27856 14977
rect 27068 14900 27120 14952
rect 28448 14900 28500 14952
rect 32404 14968 32456 15020
rect 33876 15011 33928 15020
rect 33876 14977 33885 15011
rect 33885 14977 33919 15011
rect 33919 14977 33928 15011
rect 33876 14968 33928 14977
rect 28632 14943 28684 14952
rect 28632 14909 28641 14943
rect 28641 14909 28675 14943
rect 28675 14909 28684 14943
rect 28632 14900 28684 14909
rect 28816 14943 28868 14952
rect 28816 14909 28825 14943
rect 28825 14909 28859 14943
rect 28859 14909 28868 14943
rect 28816 14900 28868 14909
rect 27160 14832 27212 14884
rect 24400 14807 24452 14816
rect 24400 14773 24409 14807
rect 24409 14773 24443 14807
rect 24443 14773 24452 14807
rect 24400 14764 24452 14773
rect 24676 14764 24728 14816
rect 27620 14764 27672 14816
rect 31576 14832 31628 14884
rect 34796 14900 34848 14952
rect 35900 14943 35952 14952
rect 35900 14909 35909 14943
rect 35909 14909 35943 14943
rect 35943 14909 35952 14943
rect 35900 14900 35952 14909
rect 36544 14943 36596 14952
rect 36544 14909 36553 14943
rect 36553 14909 36587 14943
rect 36587 14909 36596 14943
rect 36544 14900 36596 14909
rect 37924 14943 37976 14952
rect 37924 14909 37933 14943
rect 37933 14909 37967 14943
rect 37967 14909 37976 14943
rect 37924 14900 37976 14909
rect 32772 14832 32824 14884
rect 30656 14764 30708 14816
rect 31024 14764 31076 14816
rect 32588 14764 32640 14816
rect 34520 14807 34572 14816
rect 34520 14773 34529 14807
rect 34529 14773 34563 14807
rect 34563 14773 34572 14807
rect 34520 14764 34572 14773
rect 35348 14764 35400 14816
rect 37188 14764 37240 14816
rect 37280 14807 37332 14816
rect 37280 14773 37289 14807
rect 37289 14773 37323 14807
rect 37323 14773 37332 14807
rect 37280 14764 37332 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1952 14560 2004 14612
rect 3608 14603 3660 14612
rect 3608 14569 3617 14603
rect 3617 14569 3651 14603
rect 3651 14569 3660 14603
rect 3608 14560 3660 14569
rect 4620 14560 4672 14612
rect 7380 14560 7432 14612
rect 8484 14560 8536 14612
rect 9036 14560 9088 14612
rect 2780 14356 2832 14408
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 10140 14356 10192 14408
rect 11336 14560 11388 14612
rect 13360 14560 13412 14612
rect 15292 14560 15344 14612
rect 12256 14424 12308 14476
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 12992 14467 13044 14476
rect 12992 14433 13001 14467
rect 13001 14433 13035 14467
rect 13035 14433 13044 14467
rect 12992 14424 13044 14433
rect 14096 14424 14148 14476
rect 15568 14424 15620 14476
rect 18144 14560 18196 14612
rect 19248 14560 19300 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 20076 14560 20128 14612
rect 12624 14356 12676 14408
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 13544 14356 13596 14408
rect 7012 14288 7064 14340
rect 8576 14288 8628 14340
rect 9128 14331 9180 14340
rect 9128 14297 9137 14331
rect 9137 14297 9171 14331
rect 9171 14297 9180 14331
rect 9128 14288 9180 14297
rect 11428 14288 11480 14340
rect 16304 14356 16356 14408
rect 17408 14356 17460 14408
rect 17592 14356 17644 14408
rect 20720 14492 20772 14544
rect 23756 14560 23808 14612
rect 24308 14560 24360 14612
rect 19524 14467 19576 14476
rect 19524 14433 19533 14467
rect 19533 14433 19567 14467
rect 19567 14433 19576 14467
rect 19524 14424 19576 14433
rect 19708 14424 19760 14476
rect 23848 14424 23900 14476
rect 25688 14424 25740 14476
rect 26240 14424 26292 14476
rect 8208 14220 8260 14272
rect 11244 14220 11296 14272
rect 12716 14220 12768 14272
rect 12808 14220 12860 14272
rect 14188 14288 14240 14340
rect 16488 14331 16540 14340
rect 16488 14297 16522 14331
rect 16522 14297 16540 14331
rect 16488 14288 16540 14297
rect 18788 14331 18840 14340
rect 18788 14297 18806 14331
rect 18806 14297 18840 14331
rect 18788 14288 18840 14297
rect 23296 14288 23348 14340
rect 24032 14288 24084 14340
rect 14096 14263 14148 14272
rect 14096 14229 14105 14263
rect 14105 14229 14139 14263
rect 14139 14229 14148 14263
rect 14096 14220 14148 14229
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 18512 14220 18564 14272
rect 20168 14220 20220 14272
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 22744 14220 22796 14272
rect 27528 14356 27580 14408
rect 28080 14560 28132 14612
rect 28632 14492 28684 14544
rect 27988 14424 28040 14476
rect 30748 14560 30800 14612
rect 31208 14560 31260 14612
rect 32312 14560 32364 14612
rect 33232 14603 33284 14612
rect 33232 14569 33241 14603
rect 33241 14569 33275 14603
rect 33275 14569 33284 14603
rect 33232 14560 33284 14569
rect 34796 14603 34848 14612
rect 34796 14569 34805 14603
rect 34805 14569 34839 14603
rect 34839 14569 34848 14603
rect 34796 14560 34848 14569
rect 35348 14560 35400 14612
rect 36544 14560 36596 14612
rect 37280 14560 37332 14612
rect 37372 14560 37424 14612
rect 33140 14467 33192 14476
rect 33140 14433 33149 14467
rect 33149 14433 33183 14467
rect 33183 14433 33192 14467
rect 33140 14424 33192 14433
rect 31024 14399 31076 14408
rect 24768 14288 24820 14340
rect 24216 14220 24268 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 26332 14263 26384 14272
rect 26332 14229 26341 14263
rect 26341 14229 26375 14263
rect 26375 14229 26384 14263
rect 26332 14220 26384 14229
rect 31024 14365 31033 14399
rect 31033 14365 31067 14399
rect 31067 14365 31076 14399
rect 31024 14356 31076 14365
rect 30104 14288 30156 14340
rect 36176 14356 36228 14408
rect 26976 14220 27028 14272
rect 29736 14220 29788 14272
rect 31484 14220 31536 14272
rect 33784 14220 33836 14272
rect 38292 14492 38344 14544
rect 37832 14356 37884 14408
rect 37648 14288 37700 14340
rect 37372 14220 37424 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 14016 1728 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6644 14016 6696 14068
rect 9404 14016 9456 14068
rect 1584 13948 1636 14000
rect 7012 13991 7064 14000
rect 7012 13957 7021 13991
rect 7021 13957 7055 13991
rect 7055 13957 7064 13991
rect 7012 13948 7064 13957
rect 8300 13948 8352 14000
rect 11980 14016 12032 14068
rect 12532 14016 12584 14068
rect 14096 14016 14148 14068
rect 16672 14016 16724 14068
rect 17868 14016 17920 14068
rect 18144 14016 18196 14068
rect 18788 14016 18840 14068
rect 20076 14016 20128 14068
rect 20168 14016 20220 14068
rect 23940 14016 23992 14068
rect 24032 14059 24084 14068
rect 24032 14025 24041 14059
rect 24041 14025 24075 14059
rect 24075 14025 24084 14059
rect 24032 14016 24084 14025
rect 24676 14016 24728 14068
rect 24952 14059 25004 14068
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 25228 14016 25280 14068
rect 25964 14059 26016 14068
rect 25964 14025 25973 14059
rect 25973 14025 26007 14059
rect 26007 14025 26016 14059
rect 25964 14016 26016 14025
rect 26700 14016 26752 14068
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 3424 13880 3476 13932
rect 3976 13923 4028 13932
rect 3976 13889 3985 13923
rect 3985 13889 4019 13923
rect 4019 13889 4028 13923
rect 3976 13880 4028 13889
rect 2964 13812 3016 13864
rect 4620 13744 4672 13796
rect 5080 13744 5132 13796
rect 5632 13676 5684 13728
rect 6092 13676 6144 13728
rect 7932 13812 7984 13864
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 9496 13812 9548 13864
rect 7840 13744 7892 13796
rect 10416 13880 10468 13932
rect 9220 13676 9272 13728
rect 9404 13719 9456 13728
rect 9404 13685 9413 13719
rect 9413 13685 9447 13719
rect 9447 13685 9456 13719
rect 9404 13676 9456 13685
rect 11796 13880 11848 13932
rect 12808 13880 12860 13932
rect 12532 13812 12584 13864
rect 14280 13948 14332 14000
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 16304 13812 16356 13864
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 19340 13880 19392 13932
rect 22192 13948 22244 14000
rect 23664 13948 23716 14000
rect 24216 13948 24268 14000
rect 18420 13812 18472 13864
rect 20720 13812 20772 13864
rect 21732 13812 21784 13864
rect 23572 13923 23624 13932
rect 23572 13889 23581 13923
rect 23581 13889 23615 13923
rect 23615 13889 23624 13923
rect 23572 13880 23624 13889
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 26976 14059 27028 14068
rect 26976 14025 26985 14059
rect 26985 14025 27019 14059
rect 27019 14025 27028 14059
rect 26976 14016 27028 14025
rect 27712 14059 27764 14068
rect 27712 14025 27721 14059
rect 27721 14025 27755 14059
rect 27755 14025 27764 14059
rect 27712 14016 27764 14025
rect 29552 14059 29604 14068
rect 29552 14025 29561 14059
rect 29561 14025 29595 14059
rect 29595 14025 29604 14059
rect 29552 14016 29604 14025
rect 30104 14016 30156 14068
rect 30564 14059 30616 14068
rect 30564 14025 30573 14059
rect 30573 14025 30607 14059
rect 30607 14025 30616 14059
rect 30564 14016 30616 14025
rect 32772 14016 32824 14068
rect 35900 14016 35952 14068
rect 36544 14016 36596 14068
rect 27436 13948 27488 14000
rect 30288 13948 30340 14000
rect 29920 13880 29972 13932
rect 31208 13923 31260 13932
rect 31208 13889 31217 13923
rect 31217 13889 31251 13923
rect 31251 13889 31260 13923
rect 31208 13880 31260 13889
rect 34520 13880 34572 13932
rect 10416 13744 10468 13796
rect 10968 13744 11020 13796
rect 23480 13744 23532 13796
rect 23848 13744 23900 13796
rect 25688 13812 25740 13864
rect 35992 13880 36044 13932
rect 37188 14016 37240 14068
rect 37648 14059 37700 14068
rect 37648 14025 37657 14059
rect 37657 14025 37691 14059
rect 37691 14025 37700 14059
rect 37648 14016 37700 14025
rect 37924 14016 37976 14068
rect 37648 13880 37700 13932
rect 24308 13744 24360 13796
rect 24584 13744 24636 13796
rect 27436 13812 27488 13864
rect 27528 13855 27580 13864
rect 27528 13821 27537 13855
rect 27537 13821 27571 13855
rect 27571 13821 27580 13855
rect 27528 13812 27580 13821
rect 34796 13812 34848 13864
rect 26516 13744 26568 13796
rect 10508 13676 10560 13728
rect 10600 13719 10652 13728
rect 10600 13685 10609 13719
rect 10609 13685 10643 13719
rect 10643 13685 10652 13719
rect 10600 13676 10652 13685
rect 13636 13719 13688 13728
rect 13636 13685 13645 13719
rect 13645 13685 13679 13719
rect 13679 13685 13688 13719
rect 13636 13676 13688 13685
rect 30472 13676 30524 13728
rect 30932 13676 30984 13728
rect 36360 13812 36412 13864
rect 37004 13744 37056 13796
rect 37740 13744 37792 13796
rect 37464 13676 37516 13728
rect 38752 13676 38804 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2872 13472 2924 13524
rect 10508 13515 10560 13524
rect 10508 13481 10517 13515
rect 10517 13481 10551 13515
rect 10551 13481 10560 13515
rect 10508 13472 10560 13481
rect 12624 13472 12676 13524
rect 13452 13472 13504 13524
rect 14464 13472 14516 13524
rect 16488 13472 16540 13524
rect 3608 13379 3660 13388
rect 3608 13345 3617 13379
rect 3617 13345 3651 13379
rect 3651 13345 3660 13379
rect 3608 13336 3660 13345
rect 6552 13336 6604 13388
rect 10232 13336 10284 13388
rect 8760 13311 8812 13320
rect 8760 13277 8769 13311
rect 8769 13277 8803 13311
rect 8803 13277 8812 13311
rect 8760 13268 8812 13277
rect 6920 13200 6972 13252
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 11336 13200 11388 13252
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 13636 13268 13688 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 23296 13472 23348 13524
rect 23848 13472 23900 13524
rect 26056 13472 26108 13524
rect 26332 13472 26384 13524
rect 26608 13515 26660 13524
rect 26608 13481 26617 13515
rect 26617 13481 26651 13515
rect 26651 13481 26660 13515
rect 26608 13472 26660 13481
rect 27068 13515 27120 13524
rect 27068 13481 27077 13515
rect 27077 13481 27111 13515
rect 27111 13481 27120 13515
rect 27068 13472 27120 13481
rect 28356 13472 28408 13524
rect 36176 13472 36228 13524
rect 28724 13404 28776 13456
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 18512 13379 18564 13388
rect 18512 13345 18521 13379
rect 18521 13345 18555 13379
rect 18555 13345 18564 13379
rect 18512 13336 18564 13345
rect 22284 13336 22336 13388
rect 25780 13336 25832 13388
rect 28172 13336 28224 13388
rect 34796 13336 34848 13388
rect 37740 13472 37792 13524
rect 37924 13472 37976 13524
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 22100 13268 22152 13320
rect 23204 13268 23256 13320
rect 27712 13268 27764 13320
rect 30656 13311 30708 13320
rect 30656 13277 30665 13311
rect 30665 13277 30699 13311
rect 30699 13277 30708 13311
rect 30656 13268 30708 13277
rect 31944 13311 31996 13320
rect 31944 13277 31953 13311
rect 31953 13277 31987 13311
rect 31987 13277 31996 13311
rect 31944 13268 31996 13277
rect 32036 13268 32088 13320
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22100 13132 22152 13141
rect 25044 13200 25096 13252
rect 26516 13132 26568 13184
rect 26792 13132 26844 13184
rect 27344 13175 27396 13184
rect 27344 13141 27353 13175
rect 27353 13141 27387 13175
rect 27387 13141 27396 13175
rect 27344 13132 27396 13141
rect 27528 13132 27580 13184
rect 28632 13200 28684 13252
rect 29736 13200 29788 13252
rect 30564 13200 30616 13252
rect 34336 13200 34388 13252
rect 37280 13200 37332 13252
rect 29276 13132 29328 13184
rect 31208 13175 31260 13184
rect 31208 13141 31217 13175
rect 31217 13141 31251 13175
rect 31251 13141 31260 13175
rect 31208 13132 31260 13141
rect 31300 13175 31352 13184
rect 31300 13141 31309 13175
rect 31309 13141 31343 13175
rect 31343 13141 31352 13175
rect 31300 13132 31352 13141
rect 33784 13132 33836 13184
rect 37004 13132 37056 13184
rect 37464 13132 37516 13184
rect 37740 13132 37792 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 11336 12971 11388 12980
rect 11336 12937 11345 12971
rect 11345 12937 11379 12971
rect 11379 12937 11388 12971
rect 11336 12928 11388 12937
rect 1952 12792 2004 12844
rect 3148 12792 3200 12844
rect 3240 12792 3292 12844
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 6368 12792 6420 12844
rect 8300 12792 8352 12844
rect 9220 12860 9272 12912
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 9864 12792 9916 12844
rect 10600 12792 10652 12844
rect 12532 12903 12584 12912
rect 12532 12869 12541 12903
rect 12541 12869 12575 12903
rect 12575 12869 12584 12903
rect 12532 12860 12584 12869
rect 12716 12860 12768 12912
rect 13728 12860 13780 12912
rect 15660 12860 15712 12912
rect 17684 12928 17736 12980
rect 23572 12928 23624 12980
rect 27344 12928 27396 12980
rect 18236 12860 18288 12912
rect 18328 12860 18380 12912
rect 22100 12903 22152 12912
rect 22100 12869 22134 12903
rect 22134 12869 22152 12903
rect 22100 12860 22152 12869
rect 23020 12860 23072 12912
rect 2872 12724 2924 12776
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 10140 12724 10192 12776
rect 12440 12724 12492 12776
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 19340 12792 19392 12844
rect 21916 12792 21968 12844
rect 23204 12792 23256 12844
rect 24124 12835 24176 12844
rect 24124 12801 24133 12835
rect 24133 12801 24167 12835
rect 24167 12801 24176 12835
rect 24124 12792 24176 12801
rect 24768 12792 24820 12844
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 11796 12699 11848 12708
rect 11796 12665 11805 12699
rect 11805 12665 11839 12699
rect 11839 12665 11848 12699
rect 16764 12724 16816 12776
rect 20904 12767 20956 12776
rect 20904 12733 20913 12767
rect 20913 12733 20947 12767
rect 20947 12733 20956 12767
rect 20904 12724 20956 12733
rect 11796 12656 11848 12665
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 7656 12588 7708 12640
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 15844 12588 15896 12640
rect 16856 12588 16908 12640
rect 21548 12631 21600 12640
rect 21548 12597 21557 12631
rect 21557 12597 21591 12631
rect 21591 12597 21600 12631
rect 21548 12588 21600 12597
rect 22560 12588 22612 12640
rect 28448 12860 28500 12912
rect 30472 12860 30524 12912
rect 30656 12971 30708 12980
rect 30656 12937 30665 12971
rect 30665 12937 30699 12971
rect 30699 12937 30708 12971
rect 30656 12928 30708 12937
rect 31300 12928 31352 12980
rect 32128 12928 32180 12980
rect 36360 12928 36412 12980
rect 37280 12971 37332 12980
rect 37280 12937 37289 12971
rect 37289 12937 37323 12971
rect 37323 12937 37332 12971
rect 37280 12928 37332 12937
rect 38292 12971 38344 12980
rect 38292 12937 38301 12971
rect 38301 12937 38335 12971
rect 38335 12937 38344 12971
rect 38292 12928 38344 12937
rect 33692 12860 33744 12912
rect 34520 12903 34572 12912
rect 34520 12869 34529 12903
rect 34529 12869 34563 12903
rect 34563 12869 34572 12903
rect 34520 12860 34572 12869
rect 37556 12860 37608 12912
rect 38108 12860 38160 12912
rect 31024 12835 31076 12844
rect 31024 12801 31033 12835
rect 31033 12801 31067 12835
rect 31067 12801 31076 12835
rect 31024 12792 31076 12801
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 34796 12792 34848 12844
rect 37372 12792 37424 12844
rect 27436 12724 27488 12776
rect 27528 12767 27580 12776
rect 27528 12733 27537 12767
rect 27537 12733 27571 12767
rect 27571 12733 27580 12767
rect 27528 12724 27580 12733
rect 28356 12767 28408 12776
rect 28356 12733 28365 12767
rect 28365 12733 28399 12767
rect 28399 12733 28408 12767
rect 28356 12724 28408 12733
rect 28816 12724 28868 12776
rect 30472 12767 30524 12776
rect 30472 12733 30481 12767
rect 30481 12733 30515 12767
rect 30515 12733 30524 12767
rect 30472 12724 30524 12733
rect 30564 12724 30616 12776
rect 32128 12724 32180 12776
rect 33140 12724 33192 12776
rect 36728 12767 36780 12776
rect 36728 12733 36737 12767
rect 36737 12733 36771 12767
rect 36771 12733 36780 12767
rect 36728 12724 36780 12733
rect 32772 12656 32824 12708
rect 22836 12588 22888 12640
rect 24952 12588 25004 12640
rect 26332 12588 26384 12640
rect 26700 12588 26752 12640
rect 28540 12631 28592 12640
rect 28540 12597 28549 12631
rect 28549 12597 28583 12631
rect 28583 12597 28592 12631
rect 28540 12588 28592 12597
rect 29920 12631 29972 12640
rect 29920 12597 29929 12631
rect 29929 12597 29963 12631
rect 29963 12597 29972 12631
rect 29920 12588 29972 12597
rect 34244 12656 34296 12708
rect 32956 12631 33008 12640
rect 32956 12597 32965 12631
rect 32965 12597 32999 12631
rect 32999 12597 33008 12631
rect 32956 12588 33008 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2872 12427 2924 12436
rect 2872 12393 2881 12427
rect 2881 12393 2915 12427
rect 2915 12393 2924 12427
rect 2872 12384 2924 12393
rect 2504 12316 2556 12368
rect 3976 12384 4028 12436
rect 4620 12384 4672 12436
rect 5908 12384 5960 12436
rect 8300 12384 8352 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 12440 12384 12492 12436
rect 15752 12384 15804 12436
rect 18236 12427 18288 12436
rect 18236 12393 18245 12427
rect 18245 12393 18279 12427
rect 18279 12393 18288 12427
rect 18236 12384 18288 12393
rect 3516 12316 3568 12368
rect 4804 12316 4856 12368
rect 18604 12316 18656 12368
rect 6184 12248 6236 12300
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 12164 12248 12216 12300
rect 13912 12248 13964 12300
rect 14740 12248 14792 12300
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 3608 12223 3660 12232
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 4804 12180 4856 12232
rect 7656 12223 7708 12232
rect 7656 12189 7690 12223
rect 7690 12189 7708 12223
rect 2412 12044 2464 12096
rect 4988 12112 5040 12164
rect 7656 12180 7708 12189
rect 8392 12180 8444 12232
rect 9588 12180 9640 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 13452 12180 13504 12232
rect 8484 12112 8536 12164
rect 9220 12112 9272 12164
rect 12164 12112 12216 12164
rect 16672 12248 16724 12300
rect 20720 12248 20772 12300
rect 22560 12248 22612 12300
rect 22652 12291 22704 12300
rect 22652 12257 22661 12291
rect 22661 12257 22695 12291
rect 22695 12257 22704 12291
rect 22652 12248 22704 12257
rect 28356 12427 28408 12436
rect 28356 12393 28365 12427
rect 28365 12393 28399 12427
rect 28399 12393 28408 12427
rect 28356 12384 28408 12393
rect 28448 12427 28500 12436
rect 28448 12393 28457 12427
rect 28457 12393 28491 12427
rect 28491 12393 28500 12427
rect 28448 12384 28500 12393
rect 32496 12384 32548 12436
rect 32772 12384 32824 12436
rect 28816 12316 28868 12368
rect 30932 12316 30984 12368
rect 24216 12248 24268 12300
rect 24768 12248 24820 12300
rect 25228 12248 25280 12300
rect 25504 12248 25556 12300
rect 16856 12180 16908 12232
rect 21640 12223 21692 12232
rect 21640 12189 21658 12223
rect 21658 12189 21692 12223
rect 21640 12180 21692 12189
rect 21824 12180 21876 12232
rect 8208 12044 8260 12096
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13820 12044 13872 12096
rect 14004 12044 14056 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 15292 12044 15344 12096
rect 15384 12044 15436 12096
rect 17500 12044 17552 12096
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 22928 12223 22980 12232
rect 22928 12189 22937 12223
rect 22937 12189 22971 12223
rect 22971 12189 22980 12223
rect 22928 12180 22980 12189
rect 24400 12180 24452 12232
rect 27712 12291 27764 12300
rect 27712 12257 27721 12291
rect 27721 12257 27755 12291
rect 27755 12257 27764 12291
rect 27712 12248 27764 12257
rect 28540 12248 28592 12300
rect 26240 12180 26292 12232
rect 31852 12248 31904 12300
rect 32036 12248 32088 12300
rect 32956 12291 33008 12300
rect 32956 12257 32965 12291
rect 32965 12257 32999 12291
rect 32999 12257 33008 12291
rect 32956 12248 33008 12257
rect 33140 12248 33192 12300
rect 26700 12112 26752 12164
rect 27068 12112 27120 12164
rect 28448 12112 28500 12164
rect 30104 12223 30156 12232
rect 30104 12189 30113 12223
rect 30113 12189 30147 12223
rect 30147 12189 30156 12223
rect 30104 12180 30156 12189
rect 31668 12223 31720 12232
rect 31668 12189 31677 12223
rect 31677 12189 31711 12223
rect 31711 12189 31720 12223
rect 31668 12180 31720 12189
rect 36728 12384 36780 12436
rect 37464 12427 37516 12436
rect 37464 12393 37473 12427
rect 37473 12393 37507 12427
rect 37507 12393 37516 12427
rect 37464 12384 37516 12393
rect 37832 12427 37884 12436
rect 37832 12393 37841 12427
rect 37841 12393 37875 12427
rect 37875 12393 37884 12427
rect 37832 12384 37884 12393
rect 36452 12291 36504 12300
rect 36452 12257 36461 12291
rect 36461 12257 36495 12291
rect 36495 12257 36504 12291
rect 36452 12248 36504 12257
rect 37924 12248 37976 12300
rect 33784 12180 33836 12232
rect 38016 12112 38068 12164
rect 22836 12044 22888 12096
rect 23204 12044 23256 12096
rect 24400 12087 24452 12096
rect 24400 12053 24409 12087
rect 24409 12053 24443 12087
rect 24443 12053 24452 12087
rect 24400 12044 24452 12053
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 24860 12087 24912 12096
rect 24860 12053 24869 12087
rect 24869 12053 24903 12087
rect 24903 12053 24912 12087
rect 24860 12044 24912 12053
rect 25780 12044 25832 12096
rect 27436 12044 27488 12096
rect 27988 12087 28040 12096
rect 27988 12053 27997 12087
rect 27997 12053 28031 12087
rect 28031 12053 28040 12087
rect 27988 12044 28040 12053
rect 29092 12044 29144 12096
rect 30564 12087 30616 12096
rect 30564 12053 30573 12087
rect 30573 12053 30607 12087
rect 30607 12053 30616 12087
rect 30564 12044 30616 12053
rect 31116 12044 31168 12096
rect 31668 12044 31720 12096
rect 31944 12044 31996 12096
rect 32404 12044 32456 12096
rect 32496 12044 32548 12096
rect 33232 12044 33284 12096
rect 34520 12087 34572 12096
rect 34520 12053 34529 12087
rect 34529 12053 34563 12087
rect 34563 12053 34572 12087
rect 34520 12044 34572 12053
rect 36084 12044 36136 12096
rect 37188 12087 37240 12096
rect 37188 12053 37197 12087
rect 37197 12053 37231 12087
rect 37231 12053 37240 12087
rect 37188 12044 37240 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2320 11840 2372 11892
rect 3608 11840 3660 11892
rect 1768 11815 1820 11824
rect 1768 11781 1777 11815
rect 1777 11781 1811 11815
rect 1811 11781 1820 11815
rect 1768 11772 1820 11781
rect 1860 11772 1912 11824
rect 3056 11772 3108 11824
rect 5264 11840 5316 11892
rect 6460 11840 6512 11892
rect 6736 11840 6788 11892
rect 7288 11840 7340 11892
rect 8116 11840 8168 11892
rect 9680 11840 9732 11892
rect 5172 11772 5224 11824
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 8392 11772 8444 11824
rect 2320 11568 2372 11620
rect 2504 11500 2556 11552
rect 4804 11636 4856 11688
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8024 11704 8076 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10968 11840 11020 11892
rect 2780 11500 2832 11552
rect 6736 11636 6788 11688
rect 6644 11568 6696 11620
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 8760 11636 8812 11688
rect 9220 11679 9272 11688
rect 9220 11645 9254 11679
rect 9254 11645 9272 11679
rect 9220 11636 9272 11645
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 9588 11636 9640 11688
rect 8576 11568 8628 11620
rect 10324 11568 10376 11620
rect 5172 11500 5224 11552
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 7932 11500 7984 11552
rect 9128 11500 9180 11552
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 14096 11840 14148 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 17132 11840 17184 11892
rect 17408 11840 17460 11892
rect 17500 11840 17552 11892
rect 13728 11772 13780 11824
rect 16212 11815 16264 11824
rect 16212 11781 16252 11815
rect 16252 11781 16264 11815
rect 16212 11772 16264 11781
rect 11980 11704 12032 11756
rect 13176 11704 13228 11756
rect 15384 11704 15436 11756
rect 16672 11704 16724 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 18052 11636 18104 11688
rect 18420 11679 18472 11688
rect 13912 11500 13964 11552
rect 14096 11500 14148 11552
rect 15292 11500 15344 11552
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 17592 11500 17644 11552
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 18604 11840 18656 11892
rect 20444 11840 20496 11892
rect 20904 11883 20956 11892
rect 20904 11849 20913 11883
rect 20913 11849 20947 11883
rect 20947 11849 20956 11883
rect 20904 11840 20956 11849
rect 22284 11840 22336 11892
rect 23204 11840 23256 11892
rect 27712 11840 27764 11892
rect 27988 11840 28040 11892
rect 30104 11840 30156 11892
rect 33140 11840 33192 11892
rect 38292 11883 38344 11892
rect 22376 11772 22428 11824
rect 22652 11772 22704 11824
rect 23572 11772 23624 11824
rect 24768 11772 24820 11824
rect 27068 11772 27120 11824
rect 29920 11772 29972 11824
rect 32036 11772 32088 11824
rect 38292 11849 38301 11883
rect 38301 11849 38335 11883
rect 38335 11849 38344 11883
rect 38292 11840 38344 11849
rect 37740 11772 37792 11824
rect 23388 11747 23440 11756
rect 23388 11713 23397 11747
rect 23397 11713 23431 11747
rect 23431 11713 23440 11747
rect 23388 11704 23440 11713
rect 24952 11747 25004 11756
rect 24952 11713 24961 11747
rect 24961 11713 24995 11747
rect 24995 11713 25004 11747
rect 24952 11704 25004 11713
rect 26148 11704 26200 11756
rect 19248 11679 19300 11688
rect 19248 11645 19257 11679
rect 19257 11645 19291 11679
rect 19291 11645 19300 11679
rect 19248 11636 19300 11645
rect 21732 11636 21784 11688
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 23296 11636 23348 11688
rect 23848 11636 23900 11688
rect 24584 11636 24636 11688
rect 27804 11747 27856 11756
rect 27804 11713 27822 11747
rect 27822 11713 27856 11747
rect 27804 11704 27856 11713
rect 28448 11704 28500 11756
rect 28816 11747 28868 11756
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 29276 11747 29328 11756
rect 29276 11713 29285 11747
rect 29285 11713 29319 11747
rect 29319 11713 29328 11747
rect 29276 11704 29328 11713
rect 33232 11747 33284 11756
rect 33232 11713 33250 11747
rect 33250 11713 33284 11747
rect 33232 11704 33284 11713
rect 33508 11747 33560 11756
rect 33508 11713 33517 11747
rect 33517 11713 33551 11747
rect 33551 11713 33560 11747
rect 33508 11704 33560 11713
rect 18696 11543 18748 11552
rect 18696 11509 18705 11543
rect 18705 11509 18739 11543
rect 18739 11509 18748 11543
rect 18696 11500 18748 11509
rect 22928 11500 22980 11552
rect 23204 11543 23256 11552
rect 23204 11509 23213 11543
rect 23213 11509 23247 11543
rect 23247 11509 23256 11543
rect 23204 11500 23256 11509
rect 23480 11500 23532 11552
rect 27896 11679 27948 11688
rect 27896 11645 27905 11679
rect 27905 11645 27939 11679
rect 27939 11645 27948 11679
rect 27896 11636 27948 11645
rect 28724 11636 28776 11688
rect 29000 11679 29052 11688
rect 29000 11645 29009 11679
rect 29009 11645 29043 11679
rect 29043 11645 29052 11679
rect 29000 11636 29052 11645
rect 29828 11636 29880 11688
rect 28080 11568 28132 11620
rect 29736 11568 29788 11620
rect 34704 11679 34756 11688
rect 34704 11645 34713 11679
rect 34713 11645 34747 11679
rect 34747 11645 34756 11679
rect 34704 11636 34756 11645
rect 34796 11636 34848 11688
rect 35532 11679 35584 11688
rect 35532 11645 35541 11679
rect 35541 11645 35575 11679
rect 35575 11645 35584 11679
rect 35532 11636 35584 11645
rect 37188 11636 37240 11688
rect 37464 11636 37516 11688
rect 25596 11500 25648 11552
rect 28264 11500 28316 11552
rect 31852 11500 31904 11552
rect 35348 11500 35400 11552
rect 37372 11568 37424 11620
rect 37924 11636 37976 11688
rect 37096 11500 37148 11552
rect 37832 11500 37884 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1860 11296 1912 11348
rect 4896 11296 4948 11348
rect 6368 11296 6420 11348
rect 6552 11296 6604 11348
rect 6736 11296 6788 11348
rect 8300 11296 8352 11348
rect 8392 11296 8444 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 9220 11296 9272 11348
rect 9404 11296 9456 11348
rect 5264 11228 5316 11280
rect 5540 11228 5592 11280
rect 8944 11271 8996 11280
rect 8944 11237 8953 11271
rect 8953 11237 8987 11271
rect 8987 11237 8996 11271
rect 8944 11228 8996 11237
rect 11980 11296 12032 11348
rect 12992 11296 13044 11348
rect 14096 11228 14148 11280
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 2780 11092 2832 11144
rect 2596 11024 2648 11076
rect 3332 11024 3384 11076
rect 7196 11092 7248 11144
rect 14004 11160 14056 11212
rect 14924 11296 14976 11348
rect 15108 11296 15160 11348
rect 16580 11296 16632 11348
rect 17132 11296 17184 11348
rect 21180 11296 21232 11348
rect 21732 11339 21784 11348
rect 21732 11305 21741 11339
rect 21741 11305 21775 11339
rect 21775 11305 21784 11339
rect 21732 11296 21784 11305
rect 22560 11296 22612 11348
rect 24860 11296 24912 11348
rect 28816 11296 28868 11348
rect 29000 11296 29052 11348
rect 31116 11296 31168 11348
rect 31300 11296 31352 11348
rect 32772 11296 32824 11348
rect 33508 11296 33560 11348
rect 34704 11339 34756 11348
rect 34704 11305 34713 11339
rect 34713 11305 34747 11339
rect 34747 11305 34756 11339
rect 34704 11296 34756 11305
rect 37648 11296 37700 11348
rect 38292 11296 38344 11348
rect 16212 11228 16264 11280
rect 16672 11160 16724 11212
rect 22284 11228 22336 11280
rect 27804 11228 27856 11280
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 25596 11160 25648 11212
rect 29828 11160 29880 11212
rect 34244 11228 34296 11280
rect 35716 11228 35768 11280
rect 33968 11160 34020 11212
rect 34520 11160 34572 11212
rect 36820 11160 36872 11212
rect 37096 11228 37148 11280
rect 37004 11160 37056 11212
rect 37372 11203 37424 11212
rect 37372 11169 37381 11203
rect 37381 11169 37415 11203
rect 37415 11169 37424 11203
rect 37372 11160 37424 11169
rect 14280 11092 14332 11144
rect 17500 11092 17552 11144
rect 1676 10956 1728 11008
rect 3424 10956 3476 11008
rect 3608 10999 3660 11008
rect 3608 10965 3617 10999
rect 3617 10965 3651 10999
rect 3651 10965 3660 10999
rect 3608 10956 3660 10965
rect 4804 10956 4856 11008
rect 10048 11067 10100 11076
rect 10048 11033 10066 11067
rect 10066 11033 10100 11067
rect 10048 11024 10100 11033
rect 11520 11024 11572 11076
rect 13452 11024 13504 11076
rect 13820 11024 13872 11076
rect 15384 11024 15436 11076
rect 15844 11024 15896 11076
rect 18880 11067 18932 11076
rect 18880 11033 18889 11067
rect 18889 11033 18923 11067
rect 18923 11033 18932 11067
rect 18880 11024 18932 11033
rect 19248 11024 19300 11076
rect 22008 11092 22060 11144
rect 23020 11135 23072 11144
rect 23020 11101 23038 11135
rect 23038 11101 23072 11135
rect 23020 11092 23072 11101
rect 23204 11092 23256 11144
rect 25504 11092 25556 11144
rect 26056 11092 26108 11144
rect 26240 11135 26292 11144
rect 26240 11101 26274 11135
rect 26274 11101 26292 11135
rect 26240 11092 26292 11101
rect 29092 11092 29144 11144
rect 31208 11135 31260 11144
rect 31208 11101 31226 11135
rect 31226 11101 31260 11135
rect 31208 11092 31260 11101
rect 31944 11092 31996 11144
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 14096 10956 14148 11008
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 18604 10999 18656 11008
rect 18604 10965 18613 10999
rect 18613 10965 18647 10999
rect 18647 10965 18656 10999
rect 18604 10956 18656 10965
rect 23388 10956 23440 11008
rect 23940 11067 23992 11076
rect 23940 11033 23949 11067
rect 23949 11033 23983 11067
rect 23983 11033 23992 11067
rect 23940 11024 23992 11033
rect 25228 11024 25280 11076
rect 28080 11024 28132 11076
rect 32404 11092 32456 11144
rect 36360 11092 36412 11144
rect 36452 11135 36504 11144
rect 36452 11101 36461 11135
rect 36461 11101 36495 11135
rect 36495 11101 36504 11135
rect 36452 11092 36504 11101
rect 37464 11092 37516 11144
rect 37924 11092 37976 11144
rect 26792 10956 26844 11008
rect 32956 11024 33008 11076
rect 33048 10999 33100 11008
rect 33048 10965 33057 10999
rect 33057 10965 33091 10999
rect 33091 10965 33100 10999
rect 33048 10956 33100 10965
rect 36084 10956 36136 11008
rect 38660 11024 38712 11076
rect 37924 10999 37976 11008
rect 37924 10965 37933 10999
rect 37933 10965 37967 10999
rect 37967 10965 37976 10999
rect 37924 10956 37976 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 2320 10752 2372 10804
rect 3240 10752 3292 10804
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 4712 10752 4764 10804
rect 1952 10727 2004 10736
rect 1952 10693 1961 10727
rect 1961 10693 1995 10727
rect 1995 10693 2004 10727
rect 1952 10684 2004 10693
rect 3424 10727 3476 10736
rect 3424 10693 3433 10727
rect 3433 10693 3467 10727
rect 3467 10693 3476 10727
rect 5080 10752 5132 10804
rect 5264 10752 5316 10804
rect 5356 10795 5408 10804
rect 5356 10761 5365 10795
rect 5365 10761 5399 10795
rect 5399 10761 5408 10795
rect 5356 10752 5408 10761
rect 6828 10752 6880 10804
rect 6920 10752 6972 10804
rect 7932 10752 7984 10804
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 9036 10752 9088 10804
rect 10048 10752 10100 10804
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 13084 10752 13136 10804
rect 3424 10684 3476 10693
rect 3148 10616 3200 10668
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2228 10548 2280 10557
rect 2412 10591 2464 10600
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 2872 10480 2924 10532
rect 3700 10616 3752 10668
rect 4804 10659 4856 10668
rect 4804 10625 4813 10659
rect 4813 10625 4847 10659
rect 4847 10625 4856 10659
rect 4804 10616 4856 10625
rect 4712 10480 4764 10532
rect 8760 10616 8812 10668
rect 5172 10548 5224 10600
rect 8944 10616 8996 10668
rect 10140 10616 10192 10668
rect 12440 10616 12492 10668
rect 15108 10616 15160 10668
rect 17592 10752 17644 10804
rect 18420 10795 18472 10804
rect 18420 10761 18429 10795
rect 18429 10761 18463 10795
rect 18463 10761 18472 10795
rect 18420 10752 18472 10761
rect 22192 10795 22244 10804
rect 22192 10761 22201 10795
rect 22201 10761 22235 10795
rect 22235 10761 22244 10795
rect 22192 10752 22244 10761
rect 22652 10752 22704 10804
rect 23480 10752 23532 10804
rect 23848 10752 23900 10804
rect 24216 10795 24268 10804
rect 24216 10761 24225 10795
rect 24225 10761 24259 10795
rect 24259 10761 24268 10795
rect 24216 10752 24268 10761
rect 26148 10795 26200 10804
rect 26148 10761 26157 10795
rect 26157 10761 26191 10795
rect 26191 10761 26200 10795
rect 26148 10752 26200 10761
rect 27620 10752 27672 10804
rect 28264 10795 28316 10804
rect 28264 10761 28273 10795
rect 28273 10761 28307 10795
rect 28307 10761 28316 10795
rect 28264 10752 28316 10761
rect 29276 10795 29328 10804
rect 29276 10761 29285 10795
rect 29285 10761 29319 10795
rect 29319 10761 29328 10795
rect 29276 10752 29328 10761
rect 30196 10752 30248 10804
rect 30472 10795 30524 10804
rect 30472 10761 30481 10795
rect 30481 10761 30515 10795
rect 30515 10761 30524 10795
rect 30472 10752 30524 10761
rect 31024 10752 31076 10804
rect 33048 10752 33100 10804
rect 33968 10752 34020 10804
rect 22376 10684 22428 10736
rect 23388 10684 23440 10736
rect 16672 10616 16724 10668
rect 18696 10616 18748 10668
rect 32312 10684 32364 10736
rect 32956 10727 33008 10736
rect 32956 10693 32965 10727
rect 32965 10693 32999 10727
rect 32999 10693 33008 10727
rect 32956 10684 33008 10693
rect 24400 10616 24452 10668
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 9864 10548 9916 10600
rect 10508 10548 10560 10600
rect 4804 10412 4856 10464
rect 9588 10480 9640 10532
rect 12716 10548 12768 10600
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 13176 10591 13228 10600
rect 13176 10557 13185 10591
rect 13185 10557 13219 10591
rect 13219 10557 13228 10591
rect 13176 10548 13228 10557
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14096 10548 14148 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 31852 10659 31904 10668
rect 31852 10625 31861 10659
rect 31861 10625 31895 10659
rect 31895 10625 31904 10659
rect 31852 10616 31904 10625
rect 14188 10548 14240 10557
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 15568 10591 15620 10600
rect 15568 10557 15577 10591
rect 15577 10557 15611 10591
rect 15611 10557 15620 10591
rect 15568 10548 15620 10557
rect 23020 10548 23072 10600
rect 12808 10480 12860 10532
rect 16028 10480 16080 10532
rect 6000 10412 6052 10464
rect 6828 10412 6880 10464
rect 8576 10412 8628 10464
rect 9036 10412 9088 10464
rect 14924 10455 14976 10464
rect 14924 10421 14933 10455
rect 14933 10421 14967 10455
rect 14967 10421 14976 10455
rect 14924 10412 14976 10421
rect 24676 10455 24728 10464
rect 24676 10421 24685 10455
rect 24685 10421 24719 10455
rect 24719 10421 24728 10455
rect 24676 10412 24728 10421
rect 25044 10412 25096 10464
rect 28264 10548 28316 10600
rect 28356 10591 28408 10600
rect 28356 10557 28365 10591
rect 28365 10557 28399 10591
rect 28399 10557 28408 10591
rect 28356 10548 28408 10557
rect 30472 10480 30524 10532
rect 27804 10455 27856 10464
rect 27804 10421 27813 10455
rect 27813 10421 27847 10455
rect 27847 10421 27856 10455
rect 27804 10412 27856 10421
rect 29368 10412 29420 10464
rect 30288 10412 30340 10464
rect 34520 10616 34572 10668
rect 32220 10591 32272 10600
rect 32220 10557 32229 10591
rect 32229 10557 32263 10591
rect 32263 10557 32272 10591
rect 32220 10548 32272 10557
rect 32404 10591 32456 10600
rect 32404 10557 32413 10591
rect 32413 10557 32447 10591
rect 32447 10557 32456 10591
rect 32404 10548 32456 10557
rect 35348 10727 35400 10736
rect 35348 10693 35366 10727
rect 35366 10693 35400 10727
rect 36084 10795 36136 10804
rect 36084 10761 36093 10795
rect 36093 10761 36127 10795
rect 36127 10761 36136 10795
rect 36084 10752 36136 10761
rect 37004 10752 37056 10804
rect 37556 10795 37608 10804
rect 37556 10761 37565 10795
rect 37565 10761 37599 10795
rect 37599 10761 37608 10795
rect 37556 10752 37608 10761
rect 37648 10795 37700 10804
rect 37648 10761 37657 10795
rect 37657 10761 37691 10795
rect 37691 10761 37700 10795
rect 37648 10752 37700 10761
rect 35348 10684 35400 10693
rect 37188 10684 37240 10736
rect 35532 10616 35584 10668
rect 33048 10480 33100 10532
rect 36176 10591 36228 10600
rect 36176 10557 36185 10591
rect 36185 10557 36219 10591
rect 36219 10557 36228 10591
rect 36176 10548 36228 10557
rect 36268 10591 36320 10600
rect 36268 10557 36277 10591
rect 36277 10557 36311 10591
rect 36311 10557 36320 10591
rect 36268 10548 36320 10557
rect 37280 10548 37332 10600
rect 37648 10548 37700 10600
rect 31024 10412 31076 10464
rect 31392 10412 31444 10464
rect 35900 10412 35952 10464
rect 38476 10480 38528 10532
rect 38292 10455 38344 10464
rect 38292 10421 38301 10455
rect 38301 10421 38335 10455
rect 38335 10421 38344 10455
rect 38292 10412 38344 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3608 10140 3660 10192
rect 3424 10004 3476 10056
rect 5264 10208 5316 10260
rect 10232 10208 10284 10260
rect 4712 10140 4764 10192
rect 5080 10183 5132 10192
rect 5080 10149 5089 10183
rect 5089 10149 5123 10183
rect 5123 10149 5132 10183
rect 5080 10140 5132 10149
rect 5540 10140 5592 10192
rect 7656 10140 7708 10192
rect 7840 10183 7892 10192
rect 7840 10149 7849 10183
rect 7849 10149 7883 10183
rect 7883 10149 7892 10183
rect 7840 10140 7892 10149
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 13176 10208 13228 10260
rect 14188 10208 14240 10260
rect 14924 10208 14976 10260
rect 15844 10251 15896 10260
rect 15844 10217 15853 10251
rect 15853 10217 15887 10251
rect 15887 10217 15896 10251
rect 15844 10208 15896 10217
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 18144 10208 18196 10260
rect 27068 10251 27120 10260
rect 27068 10217 27077 10251
rect 27077 10217 27111 10251
rect 27111 10217 27120 10251
rect 27068 10208 27120 10217
rect 27344 10208 27396 10260
rect 30932 10208 30984 10260
rect 31300 10251 31352 10260
rect 31300 10217 31309 10251
rect 31309 10217 31343 10251
rect 31343 10217 31352 10251
rect 31300 10208 31352 10217
rect 31668 10208 31720 10260
rect 36268 10208 36320 10260
rect 37464 10208 37516 10260
rect 37924 10208 37976 10260
rect 4804 10072 4856 10124
rect 8668 10072 8720 10124
rect 12900 10072 12952 10124
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 8852 10004 8904 10056
rect 16672 10115 16724 10124
rect 16672 10081 16681 10115
rect 16681 10081 16715 10115
rect 16715 10081 16724 10115
rect 16672 10072 16724 10081
rect 27528 10140 27580 10192
rect 28356 10140 28408 10192
rect 29184 10140 29236 10192
rect 31852 10140 31904 10192
rect 32128 10140 32180 10192
rect 27712 10115 27764 10124
rect 27712 10081 27721 10115
rect 27721 10081 27755 10115
rect 27755 10081 27764 10115
rect 27712 10072 27764 10081
rect 29828 10072 29880 10124
rect 34336 10140 34388 10192
rect 33048 10115 33100 10124
rect 33048 10081 33057 10115
rect 33057 10081 33091 10115
rect 33091 10081 33100 10115
rect 33048 10072 33100 10081
rect 33784 10115 33836 10124
rect 33784 10081 33793 10115
rect 33793 10081 33827 10115
rect 33827 10081 33836 10115
rect 33784 10072 33836 10081
rect 37372 10072 37424 10124
rect 14280 10004 14332 10056
rect 15108 10004 15160 10056
rect 30932 10004 30984 10056
rect 31576 10047 31628 10056
rect 31576 10013 31585 10047
rect 31585 10013 31619 10047
rect 31619 10013 31628 10047
rect 31576 10004 31628 10013
rect 1768 9936 1820 9988
rect 3700 9936 3752 9988
rect 3056 9868 3108 9920
rect 4712 9868 4764 9920
rect 8484 9868 8536 9920
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12808 9936 12860 9988
rect 17684 9936 17736 9988
rect 32220 10004 32272 10056
rect 34520 10004 34572 10056
rect 12072 9868 12124 9877
rect 15568 9868 15620 9920
rect 16856 9868 16908 9920
rect 23020 9911 23072 9920
rect 23020 9877 23029 9911
rect 23029 9877 23063 9911
rect 23063 9877 23072 9911
rect 23020 9868 23072 9877
rect 26792 9868 26844 9920
rect 30748 9911 30800 9920
rect 30748 9877 30757 9911
rect 30757 9877 30791 9911
rect 30791 9877 30800 9911
rect 30748 9868 30800 9877
rect 32036 9868 32088 9920
rect 32128 9868 32180 9920
rect 35348 9936 35400 9988
rect 36820 10004 36872 10056
rect 37280 9936 37332 9988
rect 36452 9868 36504 9920
rect 36820 9868 36872 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2412 9664 2464 9716
rect 3056 9707 3108 9716
rect 3056 9673 3065 9707
rect 3065 9673 3099 9707
rect 3099 9673 3108 9707
rect 3056 9664 3108 9673
rect 3608 9664 3660 9716
rect 5172 9664 5224 9716
rect 8024 9664 8076 9716
rect 16028 9664 16080 9716
rect 17684 9707 17736 9716
rect 17684 9673 17693 9707
rect 17693 9673 17727 9707
rect 17727 9673 17736 9707
rect 17684 9664 17736 9673
rect 21180 9664 21232 9716
rect 25044 9664 25096 9716
rect 28356 9664 28408 9716
rect 2504 9528 2556 9580
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 2228 9460 2280 9512
rect 2688 9460 2740 9512
rect 5448 9596 5500 9648
rect 7748 9639 7800 9648
rect 7748 9605 7757 9639
rect 7757 9605 7791 9639
rect 7791 9605 7800 9639
rect 7748 9596 7800 9605
rect 12532 9596 12584 9648
rect 3424 9460 3476 9512
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 3700 9460 3752 9512
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 9036 9528 9088 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 16764 9596 16816 9648
rect 24676 9596 24728 9648
rect 26792 9596 26844 9648
rect 32220 9596 32272 9648
rect 18604 9528 18656 9580
rect 20720 9528 20772 9580
rect 29092 9528 29144 9580
rect 30472 9528 30524 9580
rect 31484 9528 31536 9580
rect 32680 9528 32732 9580
rect 33048 9528 33100 9580
rect 34336 9596 34388 9648
rect 36176 9664 36228 9716
rect 37280 9707 37332 9716
rect 37280 9673 37289 9707
rect 37289 9673 37323 9707
rect 37323 9673 37332 9707
rect 37280 9664 37332 9673
rect 36084 9596 36136 9648
rect 38752 9596 38804 9648
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 3976 9392 4028 9444
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 8392 9460 8444 9512
rect 8668 9503 8720 9512
rect 8668 9469 8677 9503
rect 8677 9469 8711 9503
rect 8711 9469 8720 9503
rect 8668 9460 8720 9469
rect 3240 9324 3292 9376
rect 7472 9324 7524 9376
rect 8116 9324 8168 9376
rect 10416 9460 10468 9512
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 23020 9460 23072 9512
rect 23756 9503 23808 9512
rect 23756 9469 23765 9503
rect 23765 9469 23799 9503
rect 23799 9469 23808 9503
rect 23756 9460 23808 9469
rect 26332 9460 26384 9512
rect 29920 9503 29972 9512
rect 29920 9469 29929 9503
rect 29929 9469 29963 9503
rect 29963 9469 29972 9503
rect 29920 9460 29972 9469
rect 30564 9460 30616 9512
rect 31208 9503 31260 9512
rect 31208 9469 31217 9503
rect 31217 9469 31251 9503
rect 31251 9469 31260 9503
rect 31208 9460 31260 9469
rect 31300 9460 31352 9512
rect 15108 9392 15160 9444
rect 16672 9392 16724 9444
rect 18512 9392 18564 9444
rect 31668 9392 31720 9444
rect 36820 9503 36872 9512
rect 36820 9469 36829 9503
rect 36829 9469 36863 9503
rect 36863 9469 36872 9503
rect 36820 9460 36872 9469
rect 37832 9503 37884 9512
rect 37832 9469 37841 9503
rect 37841 9469 37875 9503
rect 37875 9469 37884 9503
rect 37832 9460 37884 9469
rect 38016 9460 38068 9512
rect 8944 9324 8996 9376
rect 11244 9324 11296 9376
rect 12164 9324 12216 9376
rect 18420 9367 18472 9376
rect 18420 9333 18429 9367
rect 18429 9333 18463 9367
rect 18463 9333 18472 9367
rect 18420 9324 18472 9333
rect 23204 9367 23256 9376
rect 23204 9333 23213 9367
rect 23213 9333 23247 9367
rect 23247 9333 23256 9367
rect 23204 9324 23256 9333
rect 25504 9367 25556 9376
rect 25504 9333 25513 9367
rect 25513 9333 25547 9367
rect 25547 9333 25556 9367
rect 25504 9324 25556 9333
rect 27160 9367 27212 9376
rect 27160 9333 27169 9367
rect 27169 9333 27203 9367
rect 27203 9333 27212 9367
rect 27160 9324 27212 9333
rect 29000 9324 29052 9376
rect 30564 9367 30616 9376
rect 30564 9333 30573 9367
rect 30573 9333 30607 9367
rect 30607 9333 30616 9367
rect 30564 9324 30616 9333
rect 30656 9367 30708 9376
rect 30656 9333 30665 9367
rect 30665 9333 30699 9367
rect 30699 9333 30708 9367
rect 30656 9324 30708 9333
rect 31024 9324 31076 9376
rect 31484 9324 31536 9376
rect 32956 9367 33008 9376
rect 32956 9333 32965 9367
rect 32965 9333 32999 9367
rect 32999 9333 33008 9367
rect 32956 9324 33008 9333
rect 33324 9367 33376 9376
rect 33324 9333 33333 9367
rect 33333 9333 33367 9367
rect 33367 9333 33376 9367
rect 33324 9324 33376 9333
rect 34520 9324 34572 9376
rect 38936 9324 38988 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 664 9120 716 9172
rect 19432 9120 19484 9172
rect 22744 9120 22796 9172
rect 23296 9120 23348 9172
rect 24676 9163 24728 9172
rect 24676 9129 24685 9163
rect 24685 9129 24719 9163
rect 24719 9129 24728 9163
rect 24676 9120 24728 9129
rect 30840 9120 30892 9172
rect 31300 9120 31352 9172
rect 34336 9163 34388 9172
rect 34336 9129 34345 9163
rect 34345 9129 34379 9163
rect 34379 9129 34388 9163
rect 34336 9120 34388 9129
rect 35348 9163 35400 9172
rect 35348 9129 35357 9163
rect 35357 9129 35391 9163
rect 35391 9129 35400 9163
rect 35348 9120 35400 9129
rect 37740 9163 37792 9172
rect 37740 9129 37749 9163
rect 37749 9129 37783 9163
rect 37783 9129 37792 9163
rect 37740 9120 37792 9129
rect 3608 9095 3660 9104
rect 3608 9061 3617 9095
rect 3617 9061 3651 9095
rect 3651 9061 3660 9095
rect 3608 9052 3660 9061
rect 2688 8984 2740 9036
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4712 9052 4764 9104
rect 7656 9052 7708 9104
rect 8944 8984 8996 9036
rect 26608 9052 26660 9104
rect 12164 8984 12216 9036
rect 16212 8984 16264 9036
rect 16672 8984 16724 9036
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4804 8916 4856 8968
rect 5080 8848 5132 8900
rect 2872 8780 2924 8832
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 3700 8780 3752 8832
rect 8116 8848 8168 8900
rect 8484 8959 8536 8968
rect 8484 8925 8502 8959
rect 8502 8925 8536 8959
rect 8484 8916 8536 8925
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 15936 8959 15988 8968
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 16948 8916 17000 8968
rect 17500 8916 17552 8968
rect 21088 8959 21140 8968
rect 21088 8925 21097 8959
rect 21097 8925 21131 8959
rect 21131 8925 21140 8959
rect 21088 8916 21140 8925
rect 8668 8848 8720 8900
rect 10508 8848 10560 8900
rect 18052 8848 18104 8900
rect 18788 8848 18840 8900
rect 24676 8916 24728 8968
rect 27068 8959 27120 8968
rect 27068 8925 27077 8959
rect 27077 8925 27111 8959
rect 27111 8925 27120 8959
rect 27068 8916 27120 8925
rect 27620 8916 27672 8968
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 30564 8916 30616 8968
rect 31944 8916 31996 8968
rect 34520 8984 34572 9036
rect 35900 9027 35952 9036
rect 35900 8993 35909 9027
rect 35909 8993 35943 9027
rect 35943 8993 35952 9027
rect 35900 8984 35952 8993
rect 37464 8984 37516 9036
rect 32772 8916 32824 8968
rect 33968 8959 34020 8968
rect 33968 8925 33977 8959
rect 33977 8925 34011 8959
rect 34011 8925 34020 8959
rect 33968 8916 34020 8925
rect 36636 8959 36688 8968
rect 36636 8925 36645 8959
rect 36645 8925 36679 8959
rect 36679 8925 36688 8959
rect 36636 8916 36688 8925
rect 37372 8959 37424 8968
rect 37372 8925 37381 8959
rect 37381 8925 37415 8959
rect 37415 8925 37424 8959
rect 37372 8916 37424 8925
rect 23204 8848 23256 8900
rect 24400 8848 24452 8900
rect 25504 8848 25556 8900
rect 28172 8848 28224 8900
rect 8944 8780 8996 8832
rect 9036 8780 9088 8832
rect 9312 8823 9364 8832
rect 9312 8789 9321 8823
rect 9321 8789 9355 8823
rect 9355 8789 9364 8823
rect 9312 8780 9364 8789
rect 9680 8780 9732 8832
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11336 8780 11388 8789
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 20904 8780 20956 8832
rect 21732 8780 21784 8832
rect 22192 8780 22244 8832
rect 22468 8780 22520 8832
rect 22744 8780 22796 8832
rect 26516 8823 26568 8832
rect 26516 8789 26525 8823
rect 26525 8789 26559 8823
rect 26559 8789 26568 8823
rect 26516 8780 26568 8789
rect 27252 8823 27304 8832
rect 27252 8789 27261 8823
rect 27261 8789 27295 8823
rect 27295 8789 27304 8823
rect 27252 8780 27304 8789
rect 27528 8780 27580 8832
rect 27988 8780 28040 8832
rect 30748 8848 30800 8900
rect 29092 8780 29144 8832
rect 29368 8823 29420 8832
rect 29368 8789 29377 8823
rect 29377 8789 29411 8823
rect 29411 8789 29420 8823
rect 29368 8780 29420 8789
rect 29552 8780 29604 8832
rect 31116 8823 31168 8832
rect 31116 8789 31125 8823
rect 31125 8789 31159 8823
rect 31159 8789 31168 8823
rect 31116 8780 31168 8789
rect 32680 8823 32732 8832
rect 32680 8789 32689 8823
rect 32689 8789 32723 8823
rect 32723 8789 32732 8823
rect 32680 8780 32732 8789
rect 34152 8780 34204 8832
rect 35900 8780 35952 8832
rect 36820 8823 36872 8832
rect 36820 8789 36829 8823
rect 36829 8789 36863 8823
rect 36863 8789 36872 8823
rect 36820 8780 36872 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3240 8576 3292 8628
rect 4160 8576 4212 8628
rect 8116 8576 8168 8628
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 11336 8576 11388 8628
rect 12900 8576 12952 8628
rect 13452 8576 13504 8628
rect 16580 8576 16632 8628
rect 17684 8576 17736 8628
rect 18420 8576 18472 8628
rect 2872 8440 2924 8492
rect 4528 8440 4580 8492
rect 6736 8483 6788 8492
rect 6736 8449 6770 8483
rect 6770 8449 6788 8483
rect 6736 8440 6788 8449
rect 7196 8440 7248 8492
rect 12440 8508 12492 8560
rect 14372 8508 14424 8560
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 8944 8483 8996 8492
rect 8944 8449 8978 8483
rect 8978 8449 8996 8483
rect 8944 8440 8996 8449
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 6184 8347 6236 8356
rect 6184 8313 6193 8347
rect 6193 8313 6227 8347
rect 6227 8313 6236 8347
rect 6184 8304 6236 8313
rect 3700 8236 3752 8288
rect 6000 8236 6052 8288
rect 9496 8372 9548 8424
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 11612 8415 11664 8424
rect 11612 8381 11621 8415
rect 11621 8381 11655 8415
rect 11655 8381 11664 8415
rect 11612 8372 11664 8381
rect 6828 8236 6880 8288
rect 8668 8304 8720 8356
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 15384 8483 15436 8492
rect 15384 8449 15418 8483
rect 15418 8449 15436 8483
rect 15384 8440 15436 8449
rect 16672 8440 16724 8492
rect 22192 8576 22244 8628
rect 22376 8576 22428 8628
rect 21088 8508 21140 8560
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 18696 8372 18748 8424
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 21732 8372 21784 8424
rect 21916 8372 21968 8424
rect 22744 8483 22796 8492
rect 22744 8449 22753 8483
rect 22753 8449 22787 8483
rect 22787 8449 22796 8483
rect 22744 8440 22796 8449
rect 26424 8576 26476 8628
rect 27068 8576 27120 8628
rect 30656 8576 30708 8628
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 23848 8372 23900 8424
rect 24584 8372 24636 8424
rect 26240 8372 26292 8424
rect 31208 8576 31260 8628
rect 32680 8576 32732 8628
rect 32772 8576 32824 8628
rect 32956 8576 33008 8628
rect 33968 8576 34020 8628
rect 34428 8576 34480 8628
rect 36176 8576 36228 8628
rect 36636 8576 36688 8628
rect 37372 8576 37424 8628
rect 38384 8619 38436 8628
rect 38384 8585 38393 8619
rect 38393 8585 38427 8619
rect 38427 8585 38436 8619
rect 38384 8576 38436 8585
rect 31668 8508 31720 8560
rect 33048 8508 33100 8560
rect 27160 8372 27212 8424
rect 22376 8304 22428 8356
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 10692 8279 10744 8288
rect 10692 8245 10701 8279
rect 10701 8245 10735 8279
rect 10735 8245 10744 8279
rect 10692 8236 10744 8245
rect 11796 8236 11848 8288
rect 13268 8236 13320 8288
rect 16948 8236 17000 8288
rect 17132 8236 17184 8288
rect 17776 8236 17828 8288
rect 18328 8236 18380 8288
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 23664 8347 23716 8356
rect 23664 8313 23673 8347
rect 23673 8313 23707 8347
rect 23707 8313 23716 8347
rect 23664 8304 23716 8313
rect 23204 8236 23256 8288
rect 23480 8236 23532 8288
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 29460 8415 29512 8424
rect 29460 8381 29469 8415
rect 29469 8381 29503 8415
rect 29503 8381 29512 8415
rect 29460 8372 29512 8381
rect 31484 8372 31536 8424
rect 32588 8415 32640 8424
rect 32588 8381 32597 8415
rect 32597 8381 32631 8415
rect 32631 8381 32640 8415
rect 32588 8372 32640 8381
rect 33048 8372 33100 8424
rect 33324 8372 33376 8424
rect 34336 8483 34388 8492
rect 34336 8449 34345 8483
rect 34345 8449 34379 8483
rect 34379 8449 34388 8483
rect 34336 8440 34388 8449
rect 34520 8440 34572 8492
rect 34704 8483 34756 8492
rect 34704 8449 34738 8483
rect 34738 8449 34756 8483
rect 34704 8440 34756 8449
rect 35992 8508 36044 8560
rect 36084 8415 36136 8424
rect 36084 8381 36093 8415
rect 36093 8381 36127 8415
rect 36127 8381 36136 8415
rect 36084 8372 36136 8381
rect 36452 8440 36504 8492
rect 37188 8440 37240 8492
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 38292 8440 38344 8492
rect 27344 8236 27396 8288
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 30196 8236 30248 8288
rect 31576 8236 31628 8288
rect 31852 8236 31904 8288
rect 32680 8236 32732 8288
rect 34060 8304 34112 8356
rect 34244 8304 34296 8356
rect 37280 8304 37332 8356
rect 37648 8304 37700 8356
rect 37740 8347 37792 8356
rect 37740 8313 37749 8347
rect 37749 8313 37783 8347
rect 37783 8313 37792 8347
rect 37740 8304 37792 8313
rect 38292 8304 38344 8356
rect 36544 8236 36596 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 3976 8032 4028 8084
rect 5448 8032 5500 8084
rect 6736 8032 6788 8084
rect 11060 8032 11112 8084
rect 12072 8032 12124 8084
rect 2596 7828 2648 7880
rect 3884 7760 3936 7812
rect 9496 7964 9548 8016
rect 10048 7964 10100 8016
rect 5264 7896 5316 7948
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 4068 7871 4120 7880
rect 4068 7837 4091 7871
rect 4091 7837 4120 7871
rect 4068 7828 4120 7837
rect 5908 7828 5960 7880
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 9404 7828 9456 7880
rect 9680 7828 9732 7880
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 11612 7896 11664 7948
rect 13728 8032 13780 8084
rect 14740 8032 14792 8084
rect 13820 7964 13872 8016
rect 13912 7964 13964 8016
rect 15936 8032 15988 8084
rect 18144 8032 18196 8084
rect 18236 8032 18288 8084
rect 19616 8032 19668 8084
rect 23756 8032 23808 8084
rect 23848 8032 23900 8084
rect 15108 7964 15160 8016
rect 17132 7964 17184 8016
rect 26240 8032 26292 8084
rect 16212 7896 16264 7948
rect 16948 7896 17000 7948
rect 18328 7896 18380 7948
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 21180 7939 21232 7948
rect 21180 7905 21189 7939
rect 21189 7905 21223 7939
rect 21223 7905 21232 7939
rect 21180 7896 21232 7905
rect 23020 7939 23072 7948
rect 23020 7905 23029 7939
rect 23029 7905 23063 7939
rect 23063 7905 23072 7939
rect 23020 7896 23072 7905
rect 23480 7896 23532 7948
rect 25044 7939 25096 7948
rect 25044 7905 25053 7939
rect 25053 7905 25087 7939
rect 25087 7905 25096 7939
rect 25044 7896 25096 7905
rect 26148 7896 26200 7948
rect 26424 7896 26476 7948
rect 26608 7939 26660 7948
rect 26608 7905 26617 7939
rect 26617 7905 26651 7939
rect 26651 7905 26660 7939
rect 26608 7896 26660 7905
rect 26792 7896 26844 7948
rect 28356 8032 28408 8084
rect 29920 8032 29972 8084
rect 31116 7964 31168 8016
rect 9772 7828 9824 7837
rect 2872 7692 2924 7744
rect 3056 7735 3108 7744
rect 3056 7701 3065 7735
rect 3065 7701 3099 7735
rect 3099 7701 3108 7735
rect 3056 7692 3108 7701
rect 3516 7692 3568 7744
rect 3608 7692 3660 7744
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 4712 7760 4764 7812
rect 8300 7760 8352 7812
rect 8392 7760 8444 7812
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 16120 7828 16172 7880
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 10140 7760 10192 7812
rect 10692 7803 10744 7812
rect 10692 7769 10726 7803
rect 10726 7769 10744 7803
rect 10692 7760 10744 7769
rect 12164 7803 12216 7812
rect 12164 7769 12198 7803
rect 12198 7769 12216 7803
rect 12164 7760 12216 7769
rect 4896 7692 4948 7744
rect 8116 7692 8168 7744
rect 9680 7692 9732 7744
rect 10048 7692 10100 7744
rect 10968 7692 11020 7744
rect 12808 7760 12860 7812
rect 14464 7760 14516 7812
rect 16212 7692 16264 7744
rect 16948 7735 17000 7744
rect 16948 7701 16957 7735
rect 16957 7701 16991 7735
rect 16991 7701 17000 7735
rect 16948 7692 17000 7701
rect 18144 7692 18196 7744
rect 18420 7692 18472 7744
rect 21364 7735 21416 7744
rect 21364 7701 21373 7735
rect 21373 7701 21407 7735
rect 21407 7701 21416 7735
rect 21364 7692 21416 7701
rect 21916 7692 21968 7744
rect 22192 7828 22244 7880
rect 27620 7896 27672 7948
rect 30288 7896 30340 7948
rect 30656 7939 30708 7948
rect 30656 7905 30665 7939
rect 30665 7905 30699 7939
rect 30699 7905 30708 7939
rect 30656 7896 30708 7905
rect 30840 7939 30892 7948
rect 30840 7905 30849 7939
rect 30849 7905 30883 7939
rect 30883 7905 30892 7939
rect 30840 7896 30892 7905
rect 31208 7896 31260 7948
rect 31668 7939 31720 7948
rect 31668 7905 31702 7939
rect 31702 7905 31720 7939
rect 31668 7896 31720 7905
rect 31852 7939 31904 7948
rect 31852 7905 31861 7939
rect 31861 7905 31895 7939
rect 31895 7905 31904 7939
rect 31852 7896 31904 7905
rect 32588 8075 32640 8084
rect 32588 8041 32597 8075
rect 32597 8041 32631 8075
rect 32631 8041 32640 8075
rect 32588 8032 32640 8041
rect 33876 8032 33928 8084
rect 36084 8075 36136 8084
rect 34152 7896 34204 7948
rect 36084 8041 36093 8075
rect 36093 8041 36127 8075
rect 36127 8041 36136 8075
rect 36084 8032 36136 8041
rect 34520 7896 34572 7948
rect 23480 7760 23532 7812
rect 22928 7692 22980 7744
rect 24216 7692 24268 7744
rect 25136 7735 25188 7744
rect 25136 7701 25145 7735
rect 25145 7701 25179 7735
rect 25179 7701 25188 7735
rect 25136 7692 25188 7701
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 26516 7692 26568 7744
rect 29460 7828 29512 7880
rect 29920 7828 29972 7880
rect 30196 7871 30248 7880
rect 30196 7837 30205 7871
rect 30205 7837 30239 7871
rect 30239 7837 30248 7871
rect 30196 7828 30248 7837
rect 29184 7760 29236 7812
rect 34244 7828 34296 7880
rect 34428 7828 34480 7880
rect 37188 7896 37240 7948
rect 38292 7939 38344 7948
rect 38292 7905 38301 7939
rect 38301 7905 38335 7939
rect 38335 7905 38344 7939
rect 38292 7896 38344 7905
rect 36820 7828 36872 7880
rect 29000 7692 29052 7744
rect 30748 7692 30800 7744
rect 32496 7735 32548 7744
rect 32496 7701 32505 7735
rect 32505 7701 32539 7735
rect 32539 7701 32548 7735
rect 32496 7692 32548 7701
rect 34152 7735 34204 7744
rect 34152 7701 34161 7735
rect 34161 7701 34195 7735
rect 34195 7701 34204 7735
rect 34152 7692 34204 7701
rect 34520 7735 34572 7744
rect 34520 7701 34529 7735
rect 34529 7701 34563 7735
rect 34563 7701 34572 7735
rect 34520 7692 34572 7701
rect 35164 7760 35216 7812
rect 36728 7760 36780 7812
rect 37556 7735 37608 7744
rect 37556 7701 37565 7735
rect 37565 7701 37599 7735
rect 37599 7701 37608 7735
rect 37556 7692 37608 7701
rect 37924 7692 37976 7744
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2596 7488 2648 7540
rect 3332 7488 3384 7540
rect 3516 7420 3568 7472
rect 3700 7352 3752 7404
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 4436 7488 4488 7540
rect 4712 7488 4764 7540
rect 4896 7488 4948 7540
rect 4804 7420 4856 7472
rect 5448 7463 5500 7472
rect 5448 7429 5457 7463
rect 5457 7429 5491 7463
rect 5491 7429 5500 7463
rect 5448 7420 5500 7429
rect 7288 7488 7340 7540
rect 9588 7488 9640 7540
rect 14372 7531 14424 7540
rect 14372 7497 14381 7531
rect 14381 7497 14415 7531
rect 14415 7497 14424 7531
rect 14372 7488 14424 7497
rect 15108 7488 15160 7540
rect 15476 7488 15528 7540
rect 17684 7488 17736 7540
rect 18604 7488 18656 7540
rect 18972 7488 19024 7540
rect 21180 7488 21232 7540
rect 24400 7531 24452 7540
rect 24400 7497 24409 7531
rect 24409 7497 24443 7531
rect 24443 7497 24452 7531
rect 24400 7488 24452 7497
rect 27252 7531 27304 7540
rect 27252 7497 27261 7531
rect 27261 7497 27295 7531
rect 27295 7497 27304 7531
rect 27252 7488 27304 7497
rect 28264 7531 28316 7540
rect 28264 7497 28273 7531
rect 28273 7497 28307 7531
rect 28307 7497 28316 7531
rect 28264 7488 28316 7497
rect 30656 7488 30708 7540
rect 31208 7488 31260 7540
rect 31852 7488 31904 7540
rect 32588 7488 32640 7540
rect 9404 7420 9456 7472
rect 2688 7327 2740 7336
rect 2688 7293 2697 7327
rect 2697 7293 2731 7327
rect 2731 7293 2740 7327
rect 2688 7284 2740 7293
rect 3148 7284 3200 7336
rect 2136 7216 2188 7268
rect 3516 7148 3568 7200
rect 4896 7148 4948 7200
rect 7472 7395 7524 7404
rect 7472 7361 7506 7395
rect 7506 7361 7524 7395
rect 7472 7352 7524 7361
rect 9036 7395 9088 7404
rect 9036 7361 9045 7395
rect 9045 7361 9079 7395
rect 9079 7361 9088 7395
rect 9036 7352 9088 7361
rect 12808 7395 12860 7404
rect 12808 7361 12826 7395
rect 12826 7361 12860 7395
rect 12808 7352 12860 7361
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 13912 7420 13964 7472
rect 14556 7420 14608 7472
rect 7196 7327 7248 7336
rect 7196 7293 7205 7327
rect 7205 7293 7239 7327
rect 7239 7293 7248 7327
rect 7196 7284 7248 7293
rect 8944 7284 8996 7336
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 10968 7284 11020 7336
rect 12256 7284 12308 7336
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 13728 7284 13780 7336
rect 5540 7216 5592 7268
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 15384 7352 15436 7404
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 16764 7352 16816 7404
rect 14464 7284 14516 7293
rect 18052 7420 18104 7472
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 25320 7352 25372 7404
rect 26240 7420 26292 7472
rect 27160 7352 27212 7404
rect 27252 7352 27304 7404
rect 29644 7352 29696 7404
rect 29736 7352 29788 7404
rect 18880 7284 18932 7336
rect 19524 7327 19576 7336
rect 19524 7293 19533 7327
rect 19533 7293 19567 7327
rect 19567 7293 19576 7327
rect 19524 7284 19576 7293
rect 23756 7284 23808 7336
rect 27068 7327 27120 7336
rect 27068 7293 27077 7327
rect 27077 7293 27111 7327
rect 27111 7293 27120 7327
rect 27068 7284 27120 7293
rect 29000 7284 29052 7336
rect 32680 7395 32732 7404
rect 32680 7361 32689 7395
rect 32689 7361 32723 7395
rect 32723 7361 32732 7395
rect 32680 7352 32732 7361
rect 31944 7284 31996 7336
rect 34152 7488 34204 7540
rect 35164 7531 35216 7540
rect 35164 7497 35173 7531
rect 35173 7497 35207 7531
rect 35207 7497 35216 7531
rect 35164 7488 35216 7497
rect 36268 7488 36320 7540
rect 37280 7531 37332 7540
rect 37280 7497 37289 7531
rect 37289 7497 37323 7531
rect 37323 7497 37332 7531
rect 37280 7488 37332 7497
rect 37556 7488 37608 7540
rect 34428 7352 34480 7404
rect 34520 7395 34572 7404
rect 34520 7361 34529 7395
rect 34529 7361 34563 7395
rect 34563 7361 34572 7395
rect 34520 7352 34572 7361
rect 36084 7395 36136 7404
rect 36084 7361 36102 7395
rect 36102 7361 36136 7395
rect 36084 7352 36136 7361
rect 36176 7395 36228 7404
rect 36176 7361 36185 7395
rect 36185 7361 36219 7395
rect 36219 7361 36228 7395
rect 36176 7352 36228 7361
rect 38108 7352 38160 7404
rect 37004 7284 37056 7336
rect 38292 7284 38344 7336
rect 22192 7216 22244 7268
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 10416 7148 10468 7200
rect 11060 7148 11112 7200
rect 13084 7148 13136 7200
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 17960 7148 18012 7200
rect 18696 7148 18748 7200
rect 22100 7148 22152 7200
rect 26148 7148 26200 7200
rect 27988 7216 28040 7268
rect 29368 7216 29420 7268
rect 36544 7216 36596 7268
rect 27620 7148 27672 7200
rect 27712 7191 27764 7200
rect 27712 7157 27721 7191
rect 27721 7157 27755 7191
rect 27755 7157 27764 7191
rect 27712 7148 27764 7157
rect 29276 7148 29328 7200
rect 29828 7148 29880 7200
rect 32404 7148 32456 7200
rect 35808 7148 35860 7200
rect 38844 7148 38896 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3700 6944 3752 6996
rect 5264 6944 5316 6996
rect 5908 6987 5960 6996
rect 5908 6953 5917 6987
rect 5917 6953 5951 6987
rect 5951 6953 5960 6987
rect 5908 6944 5960 6953
rect 10968 6987 11020 6996
rect 10968 6953 10977 6987
rect 10977 6953 11011 6987
rect 11011 6953 11020 6987
rect 10968 6944 11020 6953
rect 12164 6944 12216 6996
rect 13728 6944 13780 6996
rect 14464 6944 14516 6996
rect 16304 6944 16356 6996
rect 16764 6944 16816 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 3516 6740 3568 6792
rect 2688 6672 2740 6724
rect 3056 6672 3108 6724
rect 3884 6808 3936 6860
rect 8116 6808 8168 6860
rect 9312 6808 9364 6860
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 11888 6808 11940 6860
rect 3700 6740 3752 6792
rect 4436 6740 4488 6792
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5816 6740 5868 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 8576 6740 8628 6792
rect 9220 6740 9272 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 3700 6604 3752 6656
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 8760 6604 8812 6656
rect 9956 6604 10008 6656
rect 11060 6604 11112 6656
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 13820 6808 13872 6860
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 16948 6808 17000 6860
rect 12900 6740 12952 6792
rect 12992 6740 13044 6792
rect 18420 6808 18472 6860
rect 18696 6851 18748 6860
rect 18696 6817 18705 6851
rect 18705 6817 18739 6851
rect 18739 6817 18748 6851
rect 18696 6808 18748 6817
rect 20720 6808 20772 6860
rect 22008 6851 22060 6860
rect 22008 6817 22017 6851
rect 22017 6817 22051 6851
rect 22051 6817 22060 6851
rect 22008 6808 22060 6817
rect 22100 6851 22152 6860
rect 22100 6817 22109 6851
rect 22109 6817 22143 6851
rect 22143 6817 22152 6851
rect 22100 6808 22152 6817
rect 23296 6944 23348 6996
rect 23480 6987 23532 6996
rect 23480 6953 23489 6987
rect 23489 6953 23523 6987
rect 23523 6953 23532 6987
rect 23480 6944 23532 6953
rect 23756 6944 23808 6996
rect 25044 6987 25096 6996
rect 25044 6953 25053 6987
rect 25053 6953 25087 6987
rect 25087 6953 25096 6987
rect 25044 6944 25096 6953
rect 25320 6987 25372 6996
rect 25320 6953 25329 6987
rect 25329 6953 25363 6987
rect 25363 6953 25372 6987
rect 25320 6944 25372 6953
rect 23572 6876 23624 6928
rect 22928 6851 22980 6860
rect 22928 6817 22937 6851
rect 22937 6817 22971 6851
rect 22971 6817 22980 6851
rect 22928 6808 22980 6817
rect 19524 6740 19576 6792
rect 22284 6740 22336 6792
rect 13176 6672 13228 6724
rect 15476 6672 15528 6724
rect 17224 6672 17276 6724
rect 25044 6808 25096 6860
rect 25228 6808 25280 6860
rect 27160 6987 27212 6996
rect 27160 6953 27169 6987
rect 27169 6953 27203 6987
rect 27203 6953 27212 6987
rect 27160 6944 27212 6953
rect 27988 6944 28040 6996
rect 26608 6808 26660 6860
rect 27712 6851 27764 6860
rect 27712 6817 27721 6851
rect 27721 6817 27755 6851
rect 27755 6817 27764 6851
rect 27712 6808 27764 6817
rect 30288 6944 30340 6996
rect 33968 6944 34020 6996
rect 36084 6944 36136 6996
rect 29460 6876 29512 6928
rect 29920 6808 29972 6860
rect 30748 6851 30800 6860
rect 30748 6817 30757 6851
rect 30757 6817 30791 6851
rect 30791 6817 30800 6851
rect 30748 6808 30800 6817
rect 31116 6808 31168 6860
rect 31392 6808 31444 6860
rect 31944 6808 31996 6860
rect 12256 6604 12308 6656
rect 13728 6604 13780 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14464 6604 14516 6656
rect 15384 6604 15436 6656
rect 16212 6604 16264 6656
rect 17684 6647 17736 6656
rect 17684 6613 17693 6647
rect 17693 6613 17727 6647
rect 17727 6613 17736 6647
rect 17684 6604 17736 6613
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 21272 6647 21324 6656
rect 21272 6613 21281 6647
rect 21281 6613 21315 6647
rect 21315 6613 21324 6647
rect 21272 6604 21324 6613
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 25136 6740 25188 6792
rect 26148 6740 26200 6792
rect 28448 6783 28500 6792
rect 28448 6749 28457 6783
rect 28457 6749 28491 6783
rect 28491 6749 28500 6783
rect 28448 6740 28500 6749
rect 29000 6740 29052 6792
rect 23572 6672 23624 6724
rect 24584 6715 24636 6724
rect 24584 6681 24593 6715
rect 24593 6681 24627 6715
rect 24627 6681 24636 6715
rect 24584 6672 24636 6681
rect 30104 6783 30156 6792
rect 30104 6749 30113 6783
rect 30113 6749 30147 6783
rect 30147 6749 30156 6783
rect 30104 6740 30156 6749
rect 32404 6740 32456 6792
rect 30380 6672 30432 6724
rect 33232 6783 33284 6792
rect 33232 6749 33241 6783
rect 33241 6749 33275 6783
rect 33275 6749 33284 6783
rect 33232 6740 33284 6749
rect 34060 6740 34112 6792
rect 35164 6740 35216 6792
rect 33508 6672 33560 6724
rect 34796 6672 34848 6724
rect 35532 6851 35584 6860
rect 35532 6817 35541 6851
rect 35541 6817 35575 6851
rect 35575 6817 35584 6851
rect 35532 6808 35584 6817
rect 35900 6808 35952 6860
rect 36452 6808 36504 6860
rect 38660 6808 38712 6860
rect 38752 6808 38804 6860
rect 23756 6604 23808 6656
rect 25964 6604 26016 6656
rect 26332 6647 26384 6656
rect 26332 6613 26341 6647
rect 26341 6613 26375 6647
rect 26375 6613 26384 6647
rect 26332 6604 26384 6613
rect 29000 6604 29052 6656
rect 33048 6647 33100 6656
rect 33048 6613 33057 6647
rect 33057 6613 33091 6647
rect 33091 6613 33100 6647
rect 33048 6604 33100 6613
rect 34060 6647 34112 6656
rect 34060 6613 34069 6647
rect 34069 6613 34103 6647
rect 34103 6613 34112 6647
rect 34060 6604 34112 6613
rect 34244 6604 34296 6656
rect 34980 6647 35032 6656
rect 34980 6613 34989 6647
rect 34989 6613 35023 6647
rect 35023 6613 35032 6647
rect 34980 6604 35032 6613
rect 36820 6672 36872 6724
rect 37004 6672 37056 6724
rect 37280 6715 37332 6724
rect 37280 6681 37298 6715
rect 37298 6681 37332 6715
rect 37280 6672 37332 6681
rect 35992 6604 36044 6656
rect 37464 6740 37516 6792
rect 37648 6740 37700 6792
rect 37648 6604 37700 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2136 6443 2188 6452
rect 2136 6409 2145 6443
rect 2145 6409 2179 6443
rect 2179 6409 2188 6443
rect 2136 6400 2188 6409
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 4528 6400 4580 6452
rect 5172 6400 5224 6452
rect 5540 6400 5592 6452
rect 7012 6400 7064 6452
rect 2780 6332 2832 6384
rect 2596 6307 2648 6316
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 2412 6196 2464 6248
rect 3884 6332 3936 6384
rect 3700 6264 3752 6316
rect 4436 6264 4488 6316
rect 3240 6196 3292 6248
rect 4896 6264 4948 6316
rect 5356 6264 5408 6316
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 7380 6332 7432 6384
rect 8576 6375 8628 6384
rect 8576 6341 8585 6375
rect 8585 6341 8619 6375
rect 8619 6341 8628 6375
rect 8576 6332 8628 6341
rect 9036 6400 9088 6452
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 11428 6400 11480 6452
rect 11520 6400 11572 6452
rect 12440 6400 12492 6452
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 14096 6400 14148 6452
rect 15384 6400 15436 6452
rect 15844 6400 15896 6452
rect 20628 6400 20680 6452
rect 6000 6264 6052 6316
rect 6368 6264 6420 6316
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 5172 6196 5224 6248
rect 2688 6060 2740 6112
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 3056 6060 3108 6112
rect 9680 6128 9732 6180
rect 10140 6128 10192 6180
rect 10876 6128 10928 6180
rect 4896 6060 4948 6112
rect 7472 6060 7524 6112
rect 8668 6060 8720 6112
rect 8760 6060 8812 6112
rect 9956 6060 10008 6112
rect 10968 6060 11020 6112
rect 11244 6239 11296 6248
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 14648 6332 14700 6384
rect 13912 6264 13964 6316
rect 15476 6307 15528 6316
rect 15476 6273 15485 6307
rect 15485 6273 15519 6307
rect 15519 6273 15528 6307
rect 15476 6264 15528 6273
rect 19248 6332 19300 6384
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 17592 6239 17644 6248
rect 17592 6205 17601 6239
rect 17601 6205 17635 6239
rect 17635 6205 17644 6239
rect 17592 6196 17644 6205
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 18604 6196 18656 6248
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 21364 6264 21416 6316
rect 23020 6400 23072 6452
rect 23112 6400 23164 6452
rect 24492 6400 24544 6452
rect 25964 6400 26016 6452
rect 23388 6375 23440 6384
rect 23388 6341 23397 6375
rect 23397 6341 23431 6375
rect 23431 6341 23440 6375
rect 23388 6332 23440 6341
rect 24124 6332 24176 6384
rect 27252 6332 27304 6384
rect 21732 6196 21784 6248
rect 24676 6307 24728 6316
rect 24676 6273 24685 6307
rect 24685 6273 24719 6307
rect 24719 6273 24728 6307
rect 24676 6264 24728 6273
rect 26056 6264 26108 6316
rect 26332 6264 26384 6316
rect 27160 6264 27212 6316
rect 24400 6196 24452 6248
rect 19432 6128 19484 6180
rect 22376 6128 22428 6180
rect 24584 6196 24636 6248
rect 25872 6196 25924 6248
rect 25964 6239 26016 6248
rect 25964 6205 25973 6239
rect 25973 6205 26007 6239
rect 26007 6205 26016 6239
rect 25964 6196 26016 6205
rect 27528 6239 27580 6248
rect 27528 6205 27537 6239
rect 27537 6205 27571 6239
rect 27571 6205 27580 6239
rect 27528 6196 27580 6205
rect 27804 6400 27856 6452
rect 28632 6400 28684 6452
rect 30196 6443 30248 6452
rect 30196 6409 30205 6443
rect 30205 6409 30239 6443
rect 30239 6409 30248 6443
rect 30196 6400 30248 6409
rect 32312 6400 32364 6452
rect 33048 6400 33100 6452
rect 34336 6400 34388 6452
rect 34704 6400 34756 6452
rect 34980 6400 35032 6452
rect 35900 6400 35952 6452
rect 36084 6400 36136 6452
rect 38016 6400 38068 6452
rect 29552 6332 29604 6384
rect 30656 6332 30708 6384
rect 29092 6264 29144 6316
rect 29184 6307 29236 6316
rect 29184 6273 29193 6307
rect 29193 6273 29227 6307
rect 29227 6273 29236 6307
rect 29184 6264 29236 6273
rect 32312 6264 32364 6316
rect 32404 6264 32456 6316
rect 26700 6128 26752 6180
rect 30104 6196 30156 6248
rect 30840 6239 30892 6248
rect 30840 6205 30849 6239
rect 30849 6205 30883 6239
rect 30883 6205 30892 6239
rect 30840 6196 30892 6205
rect 31576 6239 31628 6248
rect 31576 6205 31585 6239
rect 31585 6205 31619 6239
rect 31619 6205 31628 6239
rect 31576 6196 31628 6205
rect 32680 6239 32732 6248
rect 32680 6205 32689 6239
rect 32689 6205 32723 6239
rect 32723 6205 32732 6239
rect 32680 6196 32732 6205
rect 33140 6307 33192 6316
rect 33140 6273 33149 6307
rect 33149 6273 33183 6307
rect 33183 6273 33192 6307
rect 33140 6264 33192 6273
rect 34520 6264 34572 6316
rect 32404 6128 32456 6180
rect 33416 6128 33468 6180
rect 34704 6239 34756 6248
rect 34704 6205 34713 6239
rect 34713 6205 34747 6239
rect 34747 6205 34756 6239
rect 34704 6196 34756 6205
rect 35624 6264 35676 6316
rect 37004 6264 37056 6316
rect 38200 6307 38252 6316
rect 38200 6273 38209 6307
rect 38209 6273 38243 6307
rect 38243 6273 38252 6307
rect 38200 6264 38252 6273
rect 35256 6128 35308 6180
rect 35992 6196 36044 6248
rect 36912 6239 36964 6248
rect 36912 6205 36921 6239
rect 36921 6205 36955 6239
rect 36955 6205 36964 6239
rect 36912 6196 36964 6205
rect 38292 6196 38344 6248
rect 38660 6196 38712 6248
rect 13452 6060 13504 6112
rect 15108 6103 15160 6112
rect 15108 6069 15117 6103
rect 15117 6069 15151 6103
rect 15151 6069 15160 6103
rect 15108 6060 15160 6069
rect 15200 6060 15252 6112
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 16672 6060 16724 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 20628 6060 20680 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 22008 6060 22060 6112
rect 25044 6060 25096 6112
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 25136 6060 25188 6069
rect 26148 6060 26200 6112
rect 26332 6060 26384 6112
rect 27620 6060 27672 6112
rect 27712 6103 27764 6112
rect 27712 6069 27721 6103
rect 27721 6069 27755 6103
rect 27755 6069 27764 6103
rect 27712 6060 27764 6069
rect 29736 6060 29788 6112
rect 30288 6103 30340 6112
rect 30288 6069 30297 6103
rect 30297 6069 30331 6103
rect 30331 6069 30340 6103
rect 30288 6060 30340 6069
rect 31208 6060 31260 6112
rect 32036 6060 32088 6112
rect 32128 6103 32180 6112
rect 32128 6069 32137 6103
rect 32137 6069 32171 6103
rect 32171 6069 32180 6103
rect 32128 6060 32180 6069
rect 34152 6103 34204 6112
rect 34152 6069 34161 6103
rect 34161 6069 34195 6103
rect 34195 6069 34204 6103
rect 34152 6060 34204 6069
rect 34612 6060 34664 6112
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 38384 6060 38436 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4068 5856 4120 5908
rect 2780 5720 2832 5772
rect 4068 5720 4120 5772
rect 5356 5856 5408 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6276 5856 6328 5908
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 12164 5856 12216 5908
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 7196 5720 7248 5772
rect 3056 5652 3108 5704
rect 3516 5652 3568 5704
rect 3792 5652 3844 5704
rect 4896 5695 4948 5704
rect 4896 5661 4914 5695
rect 4914 5661 4948 5695
rect 4896 5652 4948 5661
rect 6000 5652 6052 5704
rect 9680 5720 9732 5772
rect 10876 5788 10928 5840
rect 12072 5788 12124 5840
rect 11428 5720 11480 5772
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 3884 5584 3936 5636
rect 3240 5516 3292 5568
rect 4252 5516 4304 5568
rect 5908 5516 5960 5568
rect 7288 5584 7340 5636
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 8484 5584 8536 5636
rect 9128 5584 9180 5636
rect 11336 5652 11388 5704
rect 12440 5856 12492 5908
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 13728 5856 13780 5908
rect 14556 5856 14608 5908
rect 15844 5856 15896 5908
rect 17592 5856 17644 5908
rect 20812 5856 20864 5908
rect 13636 5788 13688 5840
rect 12072 5584 12124 5636
rect 15108 5720 15160 5772
rect 16856 5720 16908 5772
rect 20260 5788 20312 5840
rect 23480 5856 23532 5908
rect 24216 5899 24268 5908
rect 24216 5865 24225 5899
rect 24225 5865 24259 5899
rect 24259 5865 24268 5899
rect 24216 5856 24268 5865
rect 24400 5899 24452 5908
rect 24400 5865 24409 5899
rect 24409 5865 24443 5899
rect 24443 5865 24452 5899
rect 24400 5856 24452 5865
rect 26240 5856 26292 5908
rect 30656 5856 30708 5908
rect 24952 5788 25004 5840
rect 33232 5788 33284 5840
rect 12808 5584 12860 5636
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 15384 5652 15436 5704
rect 15752 5652 15804 5704
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 17868 5652 17920 5704
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 9772 5559 9824 5568
rect 9772 5525 9781 5559
rect 9781 5525 9815 5559
rect 9815 5525 9824 5559
rect 9772 5516 9824 5525
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 11704 5516 11756 5568
rect 15476 5584 15528 5636
rect 20628 5584 20680 5636
rect 21732 5652 21784 5704
rect 23296 5652 23348 5704
rect 23756 5652 23808 5704
rect 26792 5720 26844 5772
rect 13728 5559 13780 5568
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 15384 5516 15436 5568
rect 15660 5516 15712 5568
rect 16212 5516 16264 5568
rect 17132 5516 17184 5568
rect 17960 5516 18012 5568
rect 21456 5516 21508 5568
rect 23572 5516 23624 5568
rect 24308 5652 24360 5704
rect 24492 5584 24544 5636
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 25320 5652 25372 5704
rect 25780 5652 25832 5704
rect 25872 5695 25924 5704
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 27068 5652 27120 5704
rect 28632 5652 28684 5704
rect 30196 5695 30248 5704
rect 30196 5661 30205 5695
rect 30205 5661 30239 5695
rect 30239 5661 30248 5695
rect 30196 5652 30248 5661
rect 25228 5584 25280 5636
rect 29276 5584 29328 5636
rect 31944 5695 31996 5704
rect 31944 5661 31953 5695
rect 31953 5661 31987 5695
rect 31987 5661 31996 5695
rect 31944 5652 31996 5661
rect 32772 5652 32824 5704
rect 34244 5720 34296 5772
rect 34520 5720 34572 5772
rect 25044 5516 25096 5568
rect 25412 5559 25464 5568
rect 25412 5525 25421 5559
rect 25421 5525 25455 5559
rect 25455 5525 25464 5559
rect 25412 5516 25464 5525
rect 25504 5559 25556 5568
rect 25504 5525 25513 5559
rect 25513 5525 25547 5559
rect 25547 5525 25556 5559
rect 25504 5516 25556 5525
rect 27896 5559 27948 5568
rect 27896 5525 27905 5559
rect 27905 5525 27939 5559
rect 27939 5525 27948 5559
rect 27896 5516 27948 5525
rect 28540 5516 28592 5568
rect 29552 5516 29604 5568
rect 30564 5559 30616 5568
rect 30564 5525 30573 5559
rect 30573 5525 30607 5559
rect 30607 5525 30616 5559
rect 30564 5516 30616 5525
rect 32128 5516 32180 5568
rect 32220 5559 32272 5568
rect 32220 5525 32229 5559
rect 32229 5525 32263 5559
rect 32263 5525 32272 5559
rect 32220 5516 32272 5525
rect 32864 5584 32916 5636
rect 34796 5652 34848 5704
rect 34428 5584 34480 5636
rect 36912 5856 36964 5908
rect 37096 5788 37148 5840
rect 35808 5720 35860 5772
rect 36176 5720 36228 5772
rect 37740 5720 37792 5772
rect 37372 5652 37424 5704
rect 38292 5695 38344 5704
rect 38292 5661 38301 5695
rect 38301 5661 38335 5695
rect 38335 5661 38344 5695
rect 38292 5652 38344 5661
rect 35532 5584 35584 5636
rect 37556 5584 37608 5636
rect 34244 5516 34296 5568
rect 34520 5559 34572 5568
rect 34520 5525 34529 5559
rect 34529 5525 34563 5559
rect 34563 5525 34572 5559
rect 34520 5516 34572 5525
rect 35808 5559 35860 5568
rect 35808 5525 35817 5559
rect 35817 5525 35851 5559
rect 35851 5525 35860 5559
rect 35808 5516 35860 5525
rect 36084 5516 36136 5568
rect 36636 5559 36688 5568
rect 36636 5525 36645 5559
rect 36645 5525 36679 5559
rect 36679 5525 36688 5559
rect 36636 5516 36688 5525
rect 37004 5559 37056 5568
rect 37004 5525 37013 5559
rect 37013 5525 37047 5559
rect 37047 5525 37056 5559
rect 37004 5516 37056 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3332 5312 3384 5364
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 4068 5312 4120 5364
rect 4252 5312 4304 5364
rect 4344 5312 4396 5364
rect 4804 5312 4856 5364
rect 5632 5312 5684 5364
rect 6000 5312 6052 5364
rect 6276 5312 6328 5364
rect 3056 5176 3108 5228
rect 3332 5219 3384 5228
rect 3332 5185 3345 5219
rect 3345 5185 3384 5219
rect 3332 5176 3384 5185
rect 3700 5176 3752 5228
rect 7564 5312 7616 5364
rect 9220 5312 9272 5364
rect 10876 5312 10928 5364
rect 10968 5312 11020 5364
rect 12440 5312 12492 5364
rect 13176 5312 13228 5364
rect 13452 5312 13504 5364
rect 17960 5312 18012 5364
rect 18236 5312 18288 5364
rect 18512 5312 18564 5364
rect 21824 5355 21876 5364
rect 21824 5321 21833 5355
rect 21833 5321 21867 5355
rect 21867 5321 21876 5355
rect 21824 5312 21876 5321
rect 24952 5312 25004 5364
rect 25320 5312 25372 5364
rect 26424 5312 26476 5364
rect 27068 5312 27120 5364
rect 28632 5312 28684 5364
rect 29828 5312 29880 5364
rect 30012 5312 30064 5364
rect 4804 5176 4856 5228
rect 5264 5176 5316 5228
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 2688 5151 2740 5160
rect 2688 5117 2697 5151
rect 2697 5117 2731 5151
rect 2731 5117 2740 5151
rect 2688 5108 2740 5117
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 10140 5176 10192 5228
rect 11336 5176 11388 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 3976 5040 4028 5092
rect 4712 5040 4764 5092
rect 5908 5040 5960 5092
rect 7932 5083 7984 5092
rect 7932 5049 7941 5083
rect 7941 5049 7975 5083
rect 7975 5049 7984 5083
rect 7932 5040 7984 5049
rect 9956 5108 10008 5160
rect 10416 5108 10468 5160
rect 12900 5244 12952 5296
rect 14740 5287 14792 5296
rect 14740 5253 14749 5287
rect 14749 5253 14783 5287
rect 14783 5253 14792 5287
rect 14740 5244 14792 5253
rect 15200 5244 15252 5296
rect 12256 5176 12308 5228
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 13176 5108 13228 5160
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 3516 4972 3568 5024
rect 4344 4972 4396 5024
rect 5356 4972 5408 5024
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 7748 4972 7800 5024
rect 10048 4972 10100 5024
rect 11060 4972 11112 5024
rect 11704 4972 11756 5024
rect 12440 4972 12492 5024
rect 12716 4972 12768 5024
rect 17960 5176 18012 5228
rect 16580 5108 16632 5160
rect 17868 5108 17920 5160
rect 18972 5176 19024 5228
rect 21456 5244 21508 5296
rect 22284 5244 22336 5296
rect 22468 5244 22520 5296
rect 23112 5244 23164 5296
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 23480 5219 23532 5228
rect 23480 5185 23489 5219
rect 23489 5185 23523 5219
rect 23523 5185 23532 5219
rect 23480 5176 23532 5185
rect 19248 5151 19300 5160
rect 19248 5117 19257 5151
rect 19257 5117 19291 5151
rect 19291 5117 19300 5151
rect 19248 5108 19300 5117
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 21640 5108 21692 5160
rect 21732 5108 21784 5160
rect 23848 5108 23900 5160
rect 24124 5108 24176 5160
rect 24492 5108 24544 5160
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 24952 5176 25004 5228
rect 25136 5219 25188 5228
rect 25136 5185 25170 5219
rect 25170 5185 25188 5219
rect 25136 5176 25188 5185
rect 26240 5176 26292 5228
rect 26516 5219 26568 5228
rect 26516 5185 26525 5219
rect 26525 5185 26559 5219
rect 26559 5185 26568 5219
rect 26516 5176 26568 5185
rect 26700 5219 26752 5228
rect 26700 5185 26709 5219
rect 26709 5185 26743 5219
rect 26743 5185 26752 5219
rect 26700 5176 26752 5185
rect 29000 5244 29052 5296
rect 29184 5244 29236 5296
rect 30288 5244 30340 5296
rect 29460 5219 29512 5228
rect 29460 5185 29469 5219
rect 29469 5185 29503 5219
rect 29503 5185 29512 5219
rect 29460 5176 29512 5185
rect 31576 5312 31628 5364
rect 31668 5355 31720 5364
rect 31668 5321 31677 5355
rect 31677 5321 31711 5355
rect 31711 5321 31720 5355
rect 31668 5312 31720 5321
rect 32496 5312 32548 5364
rect 32864 5355 32916 5364
rect 32864 5321 32873 5355
rect 32873 5321 32907 5355
rect 32907 5321 32916 5355
rect 32864 5312 32916 5321
rect 33416 5312 33468 5364
rect 30564 5244 30616 5296
rect 27068 5151 27120 5160
rect 27068 5117 27077 5151
rect 27077 5117 27111 5151
rect 27111 5117 27120 5151
rect 27068 5108 27120 5117
rect 27160 5108 27212 5160
rect 27620 5108 27672 5160
rect 29000 5108 29052 5160
rect 17040 4972 17092 5024
rect 18052 4972 18104 5024
rect 18788 4972 18840 5024
rect 19708 4972 19760 5024
rect 21272 4972 21324 5024
rect 22468 4972 22520 5024
rect 24492 5015 24544 5024
rect 24492 4981 24501 5015
rect 24501 4981 24535 5015
rect 24535 4981 24544 5015
rect 24492 4972 24544 4981
rect 26884 5040 26936 5092
rect 27436 5040 27488 5092
rect 30656 5108 30708 5160
rect 31392 5108 31444 5160
rect 31944 5219 31996 5228
rect 31944 5185 31953 5219
rect 31953 5185 31987 5219
rect 31987 5185 31996 5219
rect 31944 5176 31996 5185
rect 32036 5176 32088 5228
rect 30472 5040 30524 5092
rect 32220 5151 32272 5160
rect 32220 5117 32229 5151
rect 32229 5117 32263 5151
rect 32263 5117 32272 5151
rect 32220 5108 32272 5117
rect 32496 5219 32548 5228
rect 32496 5185 32505 5219
rect 32505 5185 32539 5219
rect 32539 5185 32548 5219
rect 32496 5176 32548 5185
rect 32588 5176 32640 5228
rect 33324 5176 33376 5228
rect 33876 5219 33928 5228
rect 33876 5185 33885 5219
rect 33885 5185 33919 5219
rect 33919 5185 33928 5219
rect 33876 5176 33928 5185
rect 34152 5312 34204 5364
rect 37280 5312 37332 5364
rect 36176 5244 36228 5296
rect 34244 5176 34296 5228
rect 32864 5040 32916 5092
rect 26332 5015 26384 5024
rect 26332 4981 26341 5015
rect 26341 4981 26375 5015
rect 26375 4981 26384 5015
rect 26332 4972 26384 4981
rect 26700 4972 26752 5024
rect 28908 4972 28960 5024
rect 31852 4972 31904 5024
rect 32220 4972 32272 5024
rect 32588 4972 32640 5024
rect 32956 5015 33008 5024
rect 32956 4981 32965 5015
rect 32965 4981 32999 5015
rect 32999 4981 33008 5015
rect 32956 4972 33008 4981
rect 33048 4972 33100 5024
rect 37280 5219 37332 5228
rect 37280 5185 37289 5219
rect 37289 5185 37323 5219
rect 37323 5185 37332 5219
rect 37280 5176 37332 5185
rect 38016 5176 38068 5228
rect 34888 4972 34940 5024
rect 36452 5040 36504 5092
rect 37740 5040 37792 5092
rect 37924 5040 37976 5092
rect 36084 4972 36136 5024
rect 37832 4972 37884 5024
rect 38292 5015 38344 5024
rect 38292 4981 38301 5015
rect 38301 4981 38335 5015
rect 38335 4981 38344 5015
rect 38292 4972 38344 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4528 4768 4580 4820
rect 6460 4768 6512 4820
rect 3056 4700 3108 4752
rect 7012 4700 7064 4752
rect 3240 4564 3292 4616
rect 4528 4564 4580 4616
rect 6276 4632 6328 4684
rect 7380 4768 7432 4820
rect 8668 4768 8720 4820
rect 9956 4768 10008 4820
rect 12164 4768 12216 4820
rect 13452 4768 13504 4820
rect 11244 4700 11296 4752
rect 8300 4632 8352 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 11520 4632 11572 4684
rect 11704 4632 11756 4684
rect 12164 4675 12216 4684
rect 12164 4641 12198 4675
rect 12198 4641 12216 4675
rect 12164 4632 12216 4641
rect 13084 4632 13136 4684
rect 17500 4768 17552 4820
rect 19340 4811 19392 4820
rect 19340 4777 19349 4811
rect 19349 4777 19383 4811
rect 19383 4777 19392 4811
rect 19340 4768 19392 4777
rect 20260 4768 20312 4820
rect 14740 4700 14792 4752
rect 4712 4496 4764 4548
rect 4804 4496 4856 4548
rect 2964 4428 3016 4480
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 4896 4428 4948 4480
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 5448 4564 5500 4616
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 5908 4564 5960 4616
rect 6828 4564 6880 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 6276 4496 6328 4548
rect 6552 4496 6604 4548
rect 7104 4496 7156 4548
rect 7932 4496 7984 4548
rect 9772 4564 9824 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 14740 4564 14792 4616
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 17776 4675 17828 4684
rect 17776 4641 17785 4675
rect 17785 4641 17819 4675
rect 17819 4641 17828 4675
rect 17776 4632 17828 4641
rect 18328 4632 18380 4684
rect 19248 4632 19300 4684
rect 16580 4564 16632 4616
rect 17408 4564 17460 4616
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 10600 4496 10652 4548
rect 15384 4539 15436 4548
rect 15384 4505 15418 4539
rect 15418 4505 15436 4539
rect 15384 4496 15436 4505
rect 18236 4496 18288 4548
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 19708 4564 19760 4616
rect 20168 4564 20220 4616
rect 22284 4768 22336 4820
rect 23112 4811 23164 4820
rect 23112 4777 23121 4811
rect 23121 4777 23155 4811
rect 23155 4777 23164 4811
rect 23112 4768 23164 4777
rect 23296 4700 23348 4752
rect 23388 4632 23440 4684
rect 24124 4768 24176 4820
rect 24492 4768 24544 4820
rect 24768 4768 24820 4820
rect 23664 4675 23716 4684
rect 23664 4641 23673 4675
rect 23673 4641 23707 4675
rect 23707 4641 23716 4675
rect 23664 4632 23716 4641
rect 21732 4607 21784 4616
rect 21732 4573 21741 4607
rect 21741 4573 21775 4607
rect 21775 4573 21784 4607
rect 21732 4564 21784 4573
rect 22928 4607 22980 4616
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 22928 4564 22980 4573
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 28448 4768 28500 4820
rect 28908 4811 28960 4820
rect 28908 4777 28917 4811
rect 28917 4777 28951 4811
rect 28951 4777 28960 4811
rect 28908 4768 28960 4777
rect 29276 4811 29328 4820
rect 29276 4777 29285 4811
rect 29285 4777 29319 4811
rect 29319 4777 29328 4811
rect 29276 4768 29328 4777
rect 30196 4768 30248 4820
rect 30472 4768 30524 4820
rect 31116 4768 31168 4820
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 19984 4496 20036 4548
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 6460 4471 6512 4480
rect 6460 4437 6469 4471
rect 6469 4437 6503 4471
rect 6503 4437 6512 4471
rect 6460 4428 6512 4437
rect 10416 4428 10468 4480
rect 10508 4428 10560 4480
rect 14924 4428 14976 4480
rect 16212 4428 16264 4480
rect 18512 4428 18564 4480
rect 18880 4471 18932 4480
rect 18880 4437 18889 4471
rect 18889 4437 18923 4471
rect 18923 4437 18932 4471
rect 18880 4428 18932 4437
rect 18972 4428 19024 4480
rect 23848 4496 23900 4548
rect 26240 4564 26292 4616
rect 26424 4607 26476 4616
rect 26424 4573 26433 4607
rect 26433 4573 26467 4607
rect 26467 4573 26476 4607
rect 26424 4564 26476 4573
rect 27436 4632 27488 4684
rect 27528 4632 27580 4684
rect 30012 4632 30064 4684
rect 30196 4675 30248 4684
rect 30196 4641 30205 4675
rect 30205 4641 30239 4675
rect 30239 4641 30248 4675
rect 30196 4632 30248 4641
rect 30564 4632 30616 4684
rect 31576 4768 31628 4820
rect 32220 4768 32272 4820
rect 32496 4768 32548 4820
rect 32680 4768 32732 4820
rect 28540 4607 28592 4616
rect 28540 4573 28558 4607
rect 28558 4573 28592 4607
rect 28540 4564 28592 4573
rect 29000 4564 29052 4616
rect 29828 4564 29880 4616
rect 24124 4471 24176 4480
rect 24124 4437 24133 4471
rect 24133 4437 24167 4471
rect 24167 4437 24176 4471
rect 24124 4428 24176 4437
rect 24768 4428 24820 4480
rect 27344 4428 27396 4480
rect 27436 4471 27488 4480
rect 27436 4437 27445 4471
rect 27445 4437 27479 4471
rect 27479 4437 27488 4471
rect 27436 4428 27488 4437
rect 29368 4539 29420 4548
rect 29368 4505 29377 4539
rect 29377 4505 29411 4539
rect 29411 4505 29420 4539
rect 29368 4496 29420 4505
rect 29460 4428 29512 4480
rect 30472 4607 30524 4616
rect 30472 4573 30481 4607
rect 30481 4573 30515 4607
rect 30515 4573 30524 4607
rect 30472 4564 30524 4573
rect 31484 4564 31536 4616
rect 32956 4768 33008 4820
rect 33692 4811 33744 4820
rect 33692 4777 33701 4811
rect 33701 4777 33735 4811
rect 33735 4777 33744 4811
rect 33692 4768 33744 4777
rect 34796 4768 34848 4820
rect 36636 4768 36688 4820
rect 32864 4675 32916 4684
rect 32864 4641 32873 4675
rect 32873 4641 32907 4675
rect 32907 4641 32916 4675
rect 32864 4632 32916 4641
rect 33232 4632 33284 4684
rect 33324 4632 33376 4684
rect 33508 4632 33560 4684
rect 33600 4675 33652 4684
rect 33600 4641 33609 4675
rect 33609 4641 33643 4675
rect 33643 4641 33652 4675
rect 33600 4632 33652 4641
rect 33876 4675 33928 4684
rect 33876 4641 33885 4675
rect 33885 4641 33919 4675
rect 33919 4641 33928 4675
rect 33876 4632 33928 4641
rect 34060 4675 34112 4684
rect 34060 4641 34069 4675
rect 34069 4641 34103 4675
rect 34103 4641 34112 4675
rect 34060 4632 34112 4641
rect 34336 4632 34388 4684
rect 35164 4632 35216 4684
rect 36452 4700 36504 4752
rect 35992 4675 36044 4684
rect 35992 4641 36010 4675
rect 36010 4641 36044 4675
rect 35992 4632 36044 4641
rect 37464 4768 37516 4820
rect 33416 4607 33468 4616
rect 33416 4573 33425 4607
rect 33425 4573 33459 4607
rect 33459 4573 33468 4607
rect 33416 4564 33468 4573
rect 32588 4496 32640 4548
rect 33968 4564 34020 4616
rect 34612 4564 34664 4616
rect 34888 4607 34940 4616
rect 34888 4573 34897 4607
rect 34897 4573 34931 4607
rect 34931 4573 34940 4607
rect 34888 4564 34940 4573
rect 36084 4607 36136 4616
rect 36084 4573 36093 4607
rect 36093 4573 36127 4607
rect 36127 4573 36136 4607
rect 36084 4564 36136 4573
rect 32128 4428 32180 4480
rect 34336 4428 34388 4480
rect 37188 4564 37240 4616
rect 36912 4496 36964 4548
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2504 4156 2556 4208
rect 3792 4224 3844 4276
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 2872 4088 2924 4140
rect 3332 4088 3384 4140
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 1768 4020 1820 4072
rect 4804 4224 4856 4276
rect 5816 4224 5868 4276
rect 6828 4267 6880 4276
rect 6828 4233 6837 4267
rect 6837 4233 6871 4267
rect 6871 4233 6880 4267
rect 6828 4224 6880 4233
rect 7472 4224 7524 4276
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4988 4088 5040 4140
rect 6276 4156 6328 4208
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 6368 4156 6420 4165
rect 7748 4156 7800 4208
rect 11060 4224 11112 4276
rect 11336 4224 11388 4276
rect 14188 4224 14240 4276
rect 14924 4224 14976 4276
rect 16764 4224 16816 4276
rect 18328 4224 18380 4276
rect 18512 4267 18564 4276
rect 18512 4233 18521 4267
rect 18521 4233 18555 4267
rect 18555 4233 18564 4267
rect 18512 4224 18564 4233
rect 18696 4224 18748 4276
rect 6460 4088 6512 4140
rect 7564 4088 7616 4140
rect 8300 4088 8352 4140
rect 9496 4156 9548 4208
rect 9588 4156 9640 4208
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 9772 4088 9824 4140
rect 10048 4156 10100 4208
rect 12532 4156 12584 4208
rect 12716 4199 12768 4208
rect 12716 4165 12734 4199
rect 12734 4165 12768 4199
rect 12716 4156 12768 4165
rect 14740 4156 14792 4208
rect 15384 4156 15436 4208
rect 5356 4020 5408 4072
rect 6184 4020 6236 4072
rect 7104 4020 7156 4072
rect 9496 4063 9548 4072
rect 9496 4029 9505 4063
rect 9505 4029 9539 4063
rect 9539 4029 9548 4063
rect 9496 4020 9548 4029
rect 12164 4088 12216 4140
rect 12900 4088 12952 4140
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 14372 4088 14424 4140
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 16580 4088 16632 4140
rect 16948 4131 17000 4140
rect 16948 4097 16982 4131
rect 16982 4097 17000 4131
rect 16948 4088 17000 4097
rect 17316 4088 17368 4140
rect 18972 4156 19024 4208
rect 20168 4224 20220 4276
rect 23112 4224 23164 4276
rect 24124 4224 24176 4276
rect 24860 4224 24912 4276
rect 26516 4224 26568 4276
rect 27344 4267 27396 4276
rect 27344 4233 27353 4267
rect 27353 4233 27387 4267
rect 27387 4233 27396 4267
rect 27344 4224 27396 4233
rect 29368 4224 29420 4276
rect 32036 4224 32088 4276
rect 32128 4267 32180 4276
rect 32128 4233 32137 4267
rect 32137 4233 32171 4267
rect 32171 4233 32180 4267
rect 32128 4224 32180 4233
rect 32864 4224 32916 4276
rect 33416 4224 33468 4276
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 18512 4088 18564 4140
rect 19248 4088 19300 4140
rect 2964 3952 3016 4004
rect 3608 3952 3660 4004
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 3332 3884 3384 3936
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 3976 3927 4028 3936
rect 3976 3893 3985 3927
rect 3985 3893 4019 3927
rect 4019 3893 4028 3927
rect 3976 3884 4028 3893
rect 4068 3884 4120 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 5172 3952 5224 4004
rect 8300 3952 8352 4004
rect 11244 4020 11296 4072
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6000 3884 6052 3936
rect 8760 3884 8812 3936
rect 9956 3952 10008 4004
rect 13544 3952 13596 4004
rect 15108 4020 15160 4072
rect 15568 4020 15620 4072
rect 18052 4020 18104 4072
rect 20536 4088 20588 4140
rect 21364 4131 21416 4140
rect 21364 4097 21382 4131
rect 21382 4097 21416 4131
rect 21364 4088 21416 4097
rect 23112 4088 23164 4140
rect 24032 4156 24084 4208
rect 15752 3995 15804 4004
rect 15752 3961 15761 3995
rect 15761 3961 15795 3995
rect 15795 3961 15804 3995
rect 15752 3952 15804 3961
rect 20260 4020 20312 4072
rect 20536 3952 20588 4004
rect 12716 3884 12768 3936
rect 13912 3927 13964 3936
rect 13912 3893 13921 3927
rect 13921 3893 13955 3927
rect 13955 3893 13964 3927
rect 13912 3884 13964 3893
rect 14832 3927 14884 3936
rect 14832 3893 14841 3927
rect 14841 3893 14875 3927
rect 14875 3893 14884 3927
rect 14832 3884 14884 3893
rect 16856 3884 16908 3936
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 20168 3927 20220 3936
rect 20168 3893 20177 3927
rect 20177 3893 20211 3927
rect 20211 3893 20220 3927
rect 20168 3884 20220 3893
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 24492 4131 24544 4140
rect 24492 4097 24501 4131
rect 24501 4097 24535 4131
rect 24535 4097 24544 4131
rect 24492 4088 24544 4097
rect 25136 4156 25188 4208
rect 27160 4156 27212 4208
rect 29184 4156 29236 4208
rect 30012 4156 30064 4208
rect 25412 4088 25464 4140
rect 27804 4088 27856 4140
rect 27988 4131 28040 4140
rect 27988 4097 27997 4131
rect 27997 4097 28031 4131
rect 28031 4097 28040 4131
rect 27988 4088 28040 4097
rect 29552 4131 29604 4140
rect 29552 4097 29586 4131
rect 29586 4097 29604 4131
rect 29552 4088 29604 4097
rect 30656 4156 30708 4208
rect 31484 4156 31536 4208
rect 35900 4224 35952 4276
rect 37096 4224 37148 4276
rect 37464 4224 37516 4276
rect 38384 4224 38436 4276
rect 31208 4131 31260 4140
rect 31208 4097 31217 4131
rect 31217 4097 31251 4131
rect 31251 4097 31260 4131
rect 31208 4088 31260 4097
rect 31760 4131 31812 4140
rect 31760 4097 31769 4131
rect 31769 4097 31803 4131
rect 31803 4097 31812 4131
rect 31760 4088 31812 4097
rect 32404 4088 32456 4140
rect 32680 4131 32732 4140
rect 32680 4097 32689 4131
rect 32689 4097 32723 4131
rect 32723 4097 32732 4131
rect 32680 4088 32732 4097
rect 34244 4156 34296 4208
rect 26884 4020 26936 4072
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 27620 4020 27672 4072
rect 27896 4020 27948 4072
rect 29000 4020 29052 4072
rect 26240 3952 26292 4004
rect 29092 3952 29144 4004
rect 22100 3884 22152 3936
rect 23296 3927 23348 3936
rect 23296 3893 23305 3927
rect 23305 3893 23339 3927
rect 23339 3893 23348 3927
rect 23296 3884 23348 3893
rect 23388 3884 23440 3936
rect 24124 3927 24176 3936
rect 24124 3893 24133 3927
rect 24133 3893 24167 3927
rect 24167 3893 24176 3927
rect 24124 3884 24176 3893
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 27436 3884 27488 3936
rect 31024 4020 31076 4072
rect 30288 3952 30340 4004
rect 32220 4020 32272 4072
rect 34428 4088 34480 4140
rect 37740 4156 37792 4208
rect 38200 4156 38252 4208
rect 35624 4131 35676 4140
rect 35624 4097 35658 4131
rect 35658 4097 35676 4131
rect 35624 4088 35676 4097
rect 35900 4088 35952 4140
rect 36820 4088 36872 4140
rect 38568 4088 38620 4140
rect 38660 4088 38712 4140
rect 37924 4063 37976 4072
rect 37924 4029 37933 4063
rect 37933 4029 37967 4063
rect 37967 4029 37976 4063
rect 37924 4020 37976 4029
rect 29920 3884 29972 3936
rect 30656 3927 30708 3936
rect 30656 3893 30665 3927
rect 30665 3893 30699 3927
rect 30699 3893 30708 3927
rect 30656 3884 30708 3893
rect 30840 3884 30892 3936
rect 30932 3884 30984 3936
rect 31944 3884 31996 3936
rect 37188 3952 37240 4004
rect 33232 3884 33284 3936
rect 35992 3884 36044 3936
rect 36268 3884 36320 3936
rect 37924 3884 37976 3936
rect 38108 3927 38160 3936
rect 38108 3893 38117 3927
rect 38117 3893 38151 3927
rect 38151 3893 38160 3927
rect 38108 3884 38160 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2688 3680 2740 3732
rect 2872 3723 2924 3732
rect 2872 3689 2881 3723
rect 2881 3689 2915 3723
rect 2915 3689 2924 3723
rect 2872 3680 2924 3689
rect 2412 3655 2464 3664
rect 2412 3621 2421 3655
rect 2421 3621 2455 3655
rect 2455 3621 2464 3655
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 3700 3680 3752 3732
rect 4160 3680 4212 3732
rect 4252 3680 4304 3732
rect 6000 3680 6052 3732
rect 2412 3612 2464 3621
rect 5448 3612 5500 3664
rect 3700 3544 3752 3596
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 2872 3476 2924 3528
rect 3884 3519 3936 3528
rect 3884 3485 3893 3519
rect 3893 3485 3927 3519
rect 3927 3485 3936 3519
rect 3884 3476 3936 3485
rect 3976 3476 4028 3528
rect 4252 3476 4304 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 5448 3476 5500 3528
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 7380 3655 7432 3664
rect 7380 3621 7389 3655
rect 7389 3621 7423 3655
rect 7423 3621 7432 3655
rect 7380 3612 7432 3621
rect 7196 3544 7248 3596
rect 4160 3408 4212 3460
rect 5172 3451 5224 3460
rect 5172 3417 5181 3451
rect 5181 3417 5215 3451
rect 5215 3417 5224 3451
rect 5172 3408 5224 3417
rect 5264 3408 5316 3460
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 2320 3340 2372 3392
rect 2596 3340 2648 3392
rect 3332 3340 3384 3392
rect 3516 3340 3568 3392
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 6092 3408 6144 3460
rect 7472 3340 7524 3392
rect 9404 3680 9456 3732
rect 12164 3680 12216 3732
rect 9956 3612 10008 3664
rect 10140 3612 10192 3664
rect 11152 3612 11204 3664
rect 12624 3655 12676 3664
rect 12624 3621 12633 3655
rect 12633 3621 12667 3655
rect 12667 3621 12676 3655
rect 12624 3612 12676 3621
rect 13912 3612 13964 3664
rect 8300 3476 8352 3528
rect 8484 3544 8536 3596
rect 10508 3544 10560 3596
rect 12532 3544 12584 3596
rect 12900 3587 12952 3596
rect 12900 3553 12909 3587
rect 12909 3553 12943 3587
rect 12943 3553 12952 3587
rect 12900 3544 12952 3553
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9404 3476 9456 3528
rect 10232 3476 10284 3528
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 12716 3476 12768 3528
rect 16856 3680 16908 3732
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 19248 3680 19300 3732
rect 22008 3680 22060 3732
rect 22928 3680 22980 3732
rect 17224 3587 17276 3596
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 17224 3544 17276 3553
rect 17684 3544 17736 3596
rect 24032 3680 24084 3732
rect 24768 3680 24820 3732
rect 25044 3680 25096 3732
rect 27528 3680 27580 3732
rect 29184 3723 29236 3732
rect 29184 3689 29193 3723
rect 29193 3689 29227 3723
rect 29227 3689 29236 3723
rect 29184 3680 29236 3689
rect 29644 3723 29696 3732
rect 29644 3689 29653 3723
rect 29653 3689 29687 3723
rect 29687 3689 29696 3723
rect 29644 3680 29696 3689
rect 30012 3680 30064 3732
rect 30932 3680 30984 3732
rect 31576 3680 31628 3732
rect 32036 3680 32088 3732
rect 33048 3680 33100 3732
rect 34704 3723 34756 3732
rect 34704 3689 34713 3723
rect 34713 3689 34747 3723
rect 34747 3689 34756 3723
rect 34704 3680 34756 3689
rect 35348 3680 35400 3732
rect 37280 3680 37332 3732
rect 22376 3587 22428 3596
rect 22376 3553 22385 3587
rect 22385 3553 22419 3587
rect 22419 3553 22428 3587
rect 22376 3544 22428 3553
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 10876 3408 10928 3460
rect 10324 3340 10376 3392
rect 12624 3408 12676 3460
rect 13820 3340 13872 3392
rect 14004 3408 14056 3460
rect 14924 3476 14976 3528
rect 17316 3476 17368 3528
rect 17868 3476 17920 3528
rect 18972 3476 19024 3528
rect 14556 3408 14608 3460
rect 14648 3451 14700 3460
rect 14648 3417 14657 3451
rect 14657 3417 14691 3451
rect 14691 3417 14700 3451
rect 14648 3408 14700 3417
rect 16580 3408 16632 3460
rect 16672 3408 16724 3460
rect 17408 3408 17460 3460
rect 17960 3408 18012 3460
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 22100 3476 22152 3528
rect 23020 3476 23072 3528
rect 23112 3476 23164 3528
rect 14188 3383 14240 3392
rect 14188 3349 14197 3383
rect 14197 3349 14231 3383
rect 14231 3349 14240 3383
rect 14188 3340 14240 3349
rect 15108 3340 15160 3392
rect 22744 3408 22796 3460
rect 19064 3383 19116 3392
rect 19064 3349 19073 3383
rect 19073 3349 19107 3383
rect 19107 3349 19116 3383
rect 19064 3340 19116 3349
rect 19432 3340 19484 3392
rect 22100 3340 22152 3392
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 23204 3340 23256 3392
rect 23480 3340 23532 3392
rect 31944 3612 31996 3664
rect 24860 3544 24912 3596
rect 27436 3587 27488 3596
rect 27436 3553 27445 3587
rect 27445 3553 27479 3587
rect 27479 3553 27488 3587
rect 27436 3544 27488 3553
rect 25964 3476 26016 3528
rect 26700 3408 26752 3460
rect 26976 3408 27028 3460
rect 29368 3519 29420 3528
rect 29368 3485 29377 3519
rect 29377 3485 29411 3519
rect 29411 3485 29420 3519
rect 29368 3476 29420 3485
rect 31668 3544 31720 3596
rect 32956 3544 33008 3596
rect 35440 3612 35492 3664
rect 33232 3544 33284 3596
rect 35532 3587 35584 3596
rect 35532 3553 35541 3587
rect 35541 3553 35575 3587
rect 35575 3553 35584 3587
rect 35532 3544 35584 3553
rect 29920 3476 29972 3528
rect 31392 3476 31444 3528
rect 32036 3476 32088 3528
rect 34428 3519 34480 3528
rect 34428 3485 34437 3519
rect 34437 3485 34471 3519
rect 34471 3485 34480 3519
rect 34428 3476 34480 3485
rect 35808 3612 35860 3664
rect 36360 3612 36412 3664
rect 38108 3680 38160 3732
rect 35900 3587 35952 3596
rect 35900 3553 35909 3587
rect 35909 3553 35943 3587
rect 35943 3553 35952 3587
rect 35900 3544 35952 3553
rect 35716 3519 35768 3528
rect 35716 3485 35725 3519
rect 35725 3485 35759 3519
rect 35759 3485 35768 3519
rect 35716 3476 35768 3485
rect 38292 3544 38344 3596
rect 24492 3340 24544 3392
rect 28264 3383 28316 3392
rect 28264 3349 28273 3383
rect 28273 3349 28307 3383
rect 28307 3349 28316 3383
rect 28264 3340 28316 3349
rect 30472 3408 30524 3460
rect 30656 3408 30708 3460
rect 33600 3451 33652 3460
rect 33600 3417 33609 3451
rect 33609 3417 33643 3451
rect 33643 3417 33652 3451
rect 33600 3408 33652 3417
rect 35992 3408 36044 3460
rect 36544 3408 36596 3460
rect 37832 3476 37884 3528
rect 30104 3340 30156 3392
rect 34152 3340 34204 3392
rect 35164 3383 35216 3392
rect 35164 3349 35173 3383
rect 35173 3349 35207 3383
rect 35207 3349 35216 3383
rect 35164 3340 35216 3349
rect 36360 3340 36412 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 1860 3136 1912 3188
rect 2320 3111 2372 3120
rect 2320 3077 2329 3111
rect 2329 3077 2363 3111
rect 2363 3077 2372 3111
rect 2320 3068 2372 3077
rect 2780 3068 2832 3120
rect 1032 3000 1084 3052
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 3424 3043 3476 3052
rect 3424 3009 3433 3043
rect 3433 3009 3467 3043
rect 3467 3009 3476 3043
rect 3424 3000 3476 3009
rect 2964 2932 3016 2984
rect 3056 2975 3108 2984
rect 3056 2941 3065 2975
rect 3065 2941 3099 2975
rect 3099 2941 3108 2975
rect 3056 2932 3108 2941
rect 4252 3136 4304 3188
rect 4804 3136 4856 3188
rect 6276 3136 6328 3188
rect 7564 3136 7616 3188
rect 8760 3136 8812 3188
rect 6644 3068 6696 3120
rect 4068 3000 4120 3052
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 9220 3068 9272 3120
rect 10784 3068 10836 3120
rect 3608 2932 3660 2984
rect 2504 2907 2556 2916
rect 2504 2873 2513 2907
rect 2513 2873 2547 2907
rect 2547 2873 2556 2907
rect 2504 2864 2556 2873
rect 2688 2864 2740 2916
rect 5356 2932 5408 2984
rect 6184 2975 6236 2984
rect 6184 2941 6193 2975
rect 6193 2941 6227 2975
rect 6227 2941 6236 2975
rect 6184 2932 6236 2941
rect 7012 2932 7064 2984
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7748 3000 7800 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 9036 3000 9088 3052
rect 10416 3000 10468 3052
rect 8208 2932 8260 2984
rect 9588 2932 9640 2984
rect 3792 2796 3844 2848
rect 6000 2796 6052 2848
rect 6092 2796 6144 2848
rect 11244 3179 11296 3188
rect 11244 3145 11253 3179
rect 11253 3145 11287 3179
rect 11287 3145 11296 3179
rect 11244 3136 11296 3145
rect 14188 3136 14240 3188
rect 14556 3136 14608 3188
rect 18788 3136 18840 3188
rect 19064 3136 19116 3188
rect 19984 3136 20036 3188
rect 20536 3136 20588 3188
rect 22100 3179 22152 3188
rect 22100 3145 22109 3179
rect 22109 3145 22143 3179
rect 22143 3145 22152 3179
rect 22100 3136 22152 3145
rect 23572 3136 23624 3188
rect 11428 3000 11480 3052
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 16580 3068 16632 3120
rect 16764 3068 16816 3120
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 11980 2932 12032 2984
rect 11428 2864 11480 2916
rect 12900 2864 12952 2916
rect 14464 3000 14516 3052
rect 15476 3000 15528 3052
rect 17040 3000 17092 3052
rect 22376 3068 22428 3120
rect 19984 3000 20036 3052
rect 20260 3000 20312 3052
rect 20904 3000 20956 3052
rect 23296 3000 23348 3052
rect 24124 3043 24176 3052
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14188 2932 14240 2984
rect 15016 2932 15068 2984
rect 17224 2932 17276 2984
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 13176 2796 13228 2848
rect 13820 2796 13872 2848
rect 19340 2796 19392 2848
rect 21088 2975 21140 2984
rect 21088 2941 21097 2975
rect 21097 2941 21131 2975
rect 21131 2941 21140 2975
rect 21088 2932 21140 2941
rect 22744 2932 22796 2984
rect 24952 3179 25004 3188
rect 24952 3145 24961 3179
rect 24961 3145 24995 3179
rect 24995 3145 25004 3179
rect 24952 3136 25004 3145
rect 26608 3179 26660 3188
rect 26608 3145 26617 3179
rect 26617 3145 26651 3179
rect 26651 3145 26660 3179
rect 26608 3136 26660 3145
rect 26792 3136 26844 3188
rect 27712 3136 27764 3188
rect 28264 3136 28316 3188
rect 30196 3179 30248 3188
rect 30196 3145 30205 3179
rect 30205 3145 30239 3179
rect 30239 3145 30248 3179
rect 30196 3136 30248 3145
rect 30840 3136 30892 3188
rect 34520 3136 34572 3188
rect 35164 3136 35216 3188
rect 36820 3136 36872 3188
rect 37004 3136 37056 3188
rect 25320 3068 25372 3120
rect 24952 2932 25004 2984
rect 26332 3043 26384 3052
rect 26332 3009 26341 3043
rect 26341 3009 26375 3043
rect 26375 3009 26384 3043
rect 26332 3000 26384 3009
rect 26424 2932 26476 2984
rect 30288 3000 30340 3052
rect 30656 3068 30708 3120
rect 31392 3068 31444 3120
rect 31944 3068 31996 3120
rect 32312 3068 32364 3120
rect 35808 3068 35860 3120
rect 31852 3000 31904 3052
rect 27344 2932 27396 2984
rect 28264 2932 28316 2984
rect 30472 2932 30524 2984
rect 31208 2932 31260 2984
rect 26884 2864 26936 2916
rect 29184 2864 29236 2916
rect 22008 2796 22060 2848
rect 24032 2796 24084 2848
rect 24308 2796 24360 2848
rect 26516 2796 26568 2848
rect 28632 2796 28684 2848
rect 32036 2796 32088 2848
rect 34060 3000 34112 3052
rect 34336 3000 34388 3052
rect 37556 3068 37608 3120
rect 38660 3000 38712 3052
rect 32956 2975 33008 2984
rect 32956 2941 32965 2975
rect 32965 2941 32999 2975
rect 32999 2941 33008 2975
rect 32956 2932 33008 2941
rect 32220 2907 32272 2916
rect 32220 2873 32229 2907
rect 32229 2873 32263 2907
rect 32263 2873 32272 2907
rect 32220 2864 32272 2873
rect 34796 2932 34848 2984
rect 36084 2932 36136 2984
rect 37924 2975 37976 2984
rect 37924 2941 37933 2975
rect 37933 2941 37967 2975
rect 37967 2941 37976 2975
rect 37924 2932 37976 2941
rect 32588 2839 32640 2848
rect 32588 2805 32597 2839
rect 32597 2805 32631 2839
rect 32631 2805 32640 2839
rect 32588 2796 32640 2805
rect 33416 2796 33468 2848
rect 36084 2796 36136 2848
rect 36636 2796 36688 2848
rect 37832 2796 37884 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2872 2592 2924 2644
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 3148 2592 3200 2644
rect 8392 2592 8444 2644
rect 9496 2592 9548 2644
rect 12808 2592 12860 2644
rect 13084 2592 13136 2644
rect 14372 2635 14424 2644
rect 14372 2601 14381 2635
rect 14381 2601 14415 2635
rect 14415 2601 14424 2635
rect 14372 2592 14424 2601
rect 16580 2592 16632 2644
rect 18512 2592 18564 2644
rect 19156 2592 19208 2644
rect 20444 2592 20496 2644
rect 22652 2592 22704 2644
rect 24216 2635 24268 2644
rect 24216 2601 24225 2635
rect 24225 2601 24259 2635
rect 24259 2601 24268 2635
rect 24216 2592 24268 2601
rect 25228 2592 25280 2644
rect 26608 2635 26660 2644
rect 26608 2601 26617 2635
rect 26617 2601 26651 2635
rect 26651 2601 26660 2635
rect 26608 2592 26660 2601
rect 29368 2592 29420 2644
rect 29828 2592 29880 2644
rect 30380 2592 30432 2644
rect 33140 2592 33192 2644
rect 33692 2592 33744 2644
rect 35532 2592 35584 2644
rect 36084 2592 36136 2644
rect 36912 2635 36964 2644
rect 36912 2601 36921 2635
rect 36921 2601 36955 2635
rect 36955 2601 36964 2635
rect 36912 2592 36964 2601
rect 37648 2592 37700 2644
rect 38016 2635 38068 2644
rect 38016 2601 38025 2635
rect 38025 2601 38059 2635
rect 38059 2601 38068 2635
rect 38016 2592 38068 2601
rect 1400 2456 1452 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3240 2388 3292 2440
rect 5632 2456 5684 2508
rect 6828 2456 6880 2508
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5540 2388 5592 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7656 2388 7708 2440
rect 5080 2363 5132 2372
rect 5080 2329 5089 2363
rect 5089 2329 5123 2363
rect 5123 2329 5132 2363
rect 5080 2320 5132 2329
rect 12072 2524 12124 2576
rect 23940 2524 23992 2576
rect 9772 2456 9824 2508
rect 10600 2499 10652 2508
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 12992 2499 13044 2508
rect 12992 2465 13001 2499
rect 13001 2465 13035 2499
rect 13035 2465 13044 2499
rect 12992 2456 13044 2465
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 12348 2388 12400 2440
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 17316 2456 17368 2508
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19248 2456 19300 2508
rect 20720 2499 20772 2508
rect 20720 2465 20729 2499
rect 20729 2465 20763 2499
rect 20763 2465 20772 2499
rect 20720 2456 20772 2465
rect 23388 2456 23440 2508
rect 26148 2456 26200 2508
rect 29368 2456 29420 2508
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 15752 2320 15804 2372
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 16856 2388 16908 2440
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 18696 2320 18748 2372
rect 11152 2252 11204 2304
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 23480 2388 23532 2440
rect 24032 2431 24084 2440
rect 24032 2397 24041 2431
rect 24041 2397 24075 2431
rect 24075 2397 24084 2431
rect 24032 2388 24084 2397
rect 25504 2388 25556 2440
rect 26424 2431 26476 2440
rect 26424 2397 26433 2431
rect 26433 2397 26467 2431
rect 26467 2397 26476 2431
rect 26424 2388 26476 2397
rect 26516 2388 26568 2440
rect 27252 2388 27304 2440
rect 21916 2320 21968 2372
rect 24124 2320 24176 2372
rect 24768 2320 24820 2372
rect 29184 2431 29236 2440
rect 29184 2397 29193 2431
rect 29193 2397 29227 2431
rect 29227 2397 29236 2431
rect 29184 2388 29236 2397
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 29000 2320 29052 2372
rect 31944 2431 31996 2440
rect 31944 2397 31953 2431
rect 31953 2397 31987 2431
rect 31987 2397 31996 2431
rect 31944 2388 31996 2397
rect 34060 2456 34112 2508
rect 35808 2456 35860 2508
rect 37832 2499 37884 2508
rect 37832 2465 37841 2499
rect 37841 2465 37875 2499
rect 37875 2465 37884 2499
rect 37832 2456 37884 2465
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 34520 2431 34572 2440
rect 34520 2397 34529 2431
rect 34529 2397 34563 2431
rect 34563 2397 34572 2431
rect 34520 2388 34572 2397
rect 34612 2388 34664 2440
rect 38476 2456 38528 2508
rect 38660 2456 38712 2508
rect 31668 2320 31720 2372
rect 34428 2320 34480 2372
rect 29276 2252 29328 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 6368 2048 6420 2100
rect 9864 2048 9916 2100
rect 33600 1708 33652 1760
rect 39304 1708 39356 1760
rect 11520 1504 11572 1556
rect 16488 1504 16540 1556
<< metal2 >>
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 37372 32428 37424 32434
rect 37372 32370 37424 32376
rect 14096 32360 14148 32366
rect 14096 32302 14148 32308
rect 15016 32360 15068 32366
rect 15016 32302 15068 32308
rect 24584 32360 24636 32366
rect 24584 32302 24636 32308
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 28816 32360 28868 32366
rect 28816 32302 28868 32308
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 10060 31958 10088 32166
rect 10048 31952 10100 31958
rect 10048 31894 10100 31900
rect 9680 31680 9732 31686
rect 9680 31622 9732 31628
rect 9692 31482 9720 31622
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 10060 31278 10088 31894
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 11244 31816 11296 31822
rect 11244 31758 11296 31764
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 8760 31136 8812 31142
rect 8760 31078 8812 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 8772 30326 8800 31078
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 8760 30320 8812 30326
rect 8760 30262 8812 30268
rect 7840 30184 7892 30190
rect 7840 30126 7892 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 6000 29640 6052 29646
rect 6000 29582 6052 29588
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5080 29232 5132 29238
rect 5080 29174 5132 29180
rect 4620 28960 4672 28966
rect 4620 28902 4672 28908
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3792 28552 3844 28558
rect 4632 28506 4660 28902
rect 4724 28558 4752 28902
rect 3792 28494 3844 28500
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 3608 28008 3660 28014
rect 3608 27950 3660 27956
rect 2792 27674 2820 27950
rect 2964 27872 3016 27878
rect 2964 27814 3016 27820
rect 3056 27872 3108 27878
rect 3056 27814 3108 27820
rect 2780 27668 2832 27674
rect 2780 27610 2832 27616
rect 2044 27328 2096 27334
rect 2044 27270 2096 27276
rect 2056 26790 2084 27270
rect 2976 27062 3004 27814
rect 2964 27056 3016 27062
rect 2964 26998 3016 27004
rect 2044 26784 2096 26790
rect 2044 26726 2096 26732
rect 2320 26784 2372 26790
rect 2320 26726 2372 26732
rect 2056 26586 2084 26726
rect 2044 26580 2096 26586
rect 2044 26522 2096 26528
rect 2332 26382 2360 26726
rect 3068 26382 3096 27814
rect 3620 27130 3648 27950
rect 3712 27334 3740 28018
rect 3700 27328 3752 27334
rect 3700 27270 3752 27276
rect 3608 27124 3660 27130
rect 3608 27066 3660 27072
rect 3712 26994 3740 27270
rect 3700 26988 3752 26994
rect 3700 26930 3752 26936
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 2320 26376 2372 26382
rect 2320 26318 2372 26324
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 2332 25974 2360 26318
rect 2320 25968 2372 25974
rect 2320 25910 2372 25916
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 2056 25498 2084 25842
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 2872 24064 2924 24070
rect 2872 24006 2924 24012
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 2044 23112 2096 23118
rect 2044 23054 2096 23060
rect 2056 22642 2084 23054
rect 2516 22710 2544 23462
rect 2504 22704 2556 22710
rect 2504 22646 2556 22652
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 2056 22030 2084 22578
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 2056 19922 2084 21966
rect 2884 21962 2912 24006
rect 3436 23866 3464 24142
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 2872 21956 2924 21962
rect 2872 21898 2924 21904
rect 3068 21690 3096 23598
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 3620 21486 3648 26862
rect 3712 26246 3740 26930
rect 3804 26450 3832 28494
rect 4540 28478 4660 28506
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4540 28014 4568 28478
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4712 28416 4764 28422
rect 4712 28358 4764 28364
rect 4528 28008 4580 28014
rect 4528 27950 4580 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27130 4660 28358
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4724 26926 4752 28358
rect 4988 27600 5040 27606
rect 4988 27542 5040 27548
rect 4712 26920 4764 26926
rect 4712 26862 4764 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 3700 26240 3752 26246
rect 3700 26182 3752 26188
rect 3712 25158 3740 26182
rect 3988 25974 4016 26318
rect 4724 26058 4752 26318
rect 4724 26030 4844 26058
rect 3976 25968 4028 25974
rect 3976 25910 4028 25916
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 25424 4028 25430
rect 3976 25366 4028 25372
rect 3884 25356 3936 25362
rect 3884 25298 3936 25304
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3896 24614 3924 25298
rect 3988 24818 4016 25366
rect 4724 24954 4752 25842
rect 4816 25770 4844 26030
rect 4804 25764 4856 25770
rect 4804 25706 4856 25712
rect 4816 25362 4844 25706
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4908 25498 4936 25638
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3792 24064 3844 24070
rect 3792 24006 3844 24012
rect 3804 23118 3832 24006
rect 3896 23662 3924 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3988 22574 4016 23598
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 4080 23304 4108 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 24142
rect 4908 23746 4936 25094
rect 5000 23866 5028 27542
rect 5092 27470 5120 29174
rect 5368 28218 5396 29446
rect 5816 29164 5868 29170
rect 5816 29106 5868 29112
rect 5448 28484 5500 28490
rect 5448 28426 5500 28432
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5460 27878 5488 28426
rect 5540 28416 5592 28422
rect 5540 28358 5592 28364
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 5460 27538 5488 27814
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 5448 27532 5500 27538
rect 5448 27474 5500 27480
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 5080 25424 5132 25430
rect 5080 25366 5132 25372
rect 5092 24954 5120 25366
rect 5276 24954 5304 27474
rect 5552 27470 5580 28358
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5356 27056 5408 27062
rect 5356 26998 5408 27004
rect 5368 25906 5396 26998
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 5552 25498 5580 26386
rect 5632 26240 5684 26246
rect 5632 26182 5684 26188
rect 5644 26042 5672 26182
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 5092 24410 5120 24890
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 4712 23724 4764 23730
rect 4908 23718 5028 23746
rect 4712 23666 4764 23672
rect 4724 23322 4752 23666
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4620 23316 4672 23322
rect 4080 23276 4200 23304
rect 4172 23118 4200 23276
rect 4620 23258 4672 23264
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4252 23248 4304 23254
rect 4250 23216 4252 23225
rect 4344 23248 4396 23254
rect 4304 23216 4306 23225
rect 4344 23190 4396 23196
rect 4710 23216 4766 23225
rect 4250 23151 4306 23160
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4356 22642 4384 23190
rect 4710 23151 4766 23160
rect 4436 23044 4488 23050
rect 4436 22986 4488 22992
rect 4448 22642 4476 22986
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4540 22778 4568 22918
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4344 22636 4396 22642
rect 4172 22596 4344 22624
rect 3976 22568 4028 22574
rect 4172 22522 4200 22596
rect 4344 22578 4396 22584
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 3976 22510 4028 22516
rect 3884 22500 3936 22506
rect 3884 22442 3936 22448
rect 3896 22166 3924 22442
rect 3988 22234 4016 22510
rect 4080 22494 4200 22522
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3884 22160 3936 22166
rect 3884 22102 3936 22108
rect 4080 21962 4108 22494
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 21956 4120 21962
rect 4068 21898 4120 21904
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3436 21146 3464 21422
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3620 21078 3648 21422
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3608 21072 3660 21078
rect 3608 21014 3660 21020
rect 4632 21010 4660 22374
rect 4724 22094 4752 23151
rect 4816 23050 4844 23598
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4724 22066 4844 22094
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20398 4568 20742
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2056 19514 2084 19858
rect 2516 19854 2544 20198
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 2056 18834 2084 19450
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2044 18828 2096 18834
rect 2044 18770 2096 18776
rect 2056 18290 2084 18770
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2976 17882 3004 19314
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3436 18902 3464 19246
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3804 18766 3832 19654
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3344 17882 3372 18226
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3804 17746 3832 18566
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2148 15706 2176 16526
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 15094 1624 15506
rect 2332 15502 2360 15982
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2424 15366 2452 16458
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 15434 2636 16390
rect 2792 16182 2820 16934
rect 3160 16794 3188 16934
rect 3436 16794 3464 17070
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2596 15428 2648 15434
rect 2596 15370 2648 15376
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 1596 14006 1624 15030
rect 1688 14074 1716 15302
rect 2424 15094 2452 15302
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2792 14958 2820 15438
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14618 1992 14758
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2792 14414 2820 14894
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10810 1716 10950
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1780 9994 1808 11766
rect 1872 11354 1900 11766
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1964 10742 1992 12786
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2332 11898 2360 12174
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2056 10810 2084 11086
rect 2332 10810 2360 11562
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 1952 10736 2004 10742
rect 2424 10724 2452 12038
rect 2516 11762 2544 12310
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2792 11558 2820 14350
rect 2884 13530 2912 14962
rect 2976 13870 3004 16594
rect 3896 16590 3924 20334
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 20058 4660 20334
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4264 19378 4292 19994
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4080 18358 4108 19178
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18970 4660 19790
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4632 18578 4660 18770
rect 4724 18766 4752 19654
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4816 18578 4844 22066
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 4908 20262 4936 21014
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4908 19922 4936 20198
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 4172 18170 4200 18362
rect 4264 18222 4292 18566
rect 4632 18550 4844 18578
rect 4080 18142 4200 18170
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4080 17762 4108 18142
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4080 17734 4200 17762
rect 4172 17542 4200 17734
rect 4632 17610 4660 18550
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4724 17746 4752 18090
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4172 17082 4200 17478
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4080 17054 4200 17082
rect 4080 16776 4108 17054
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4080 16748 4200 16776
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 16250 3832 16390
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 4172 15994 4200 16748
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4540 16182 4568 16594
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4632 16114 4660 17206
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4080 15966 4200 15994
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15094 3096 15846
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 4080 15586 4108 15966
rect 4724 15910 4752 17070
rect 4816 16697 4844 17138
rect 4802 16688 4858 16697
rect 4802 16623 4858 16632
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 3344 13938 3372 15302
rect 3620 14618 3648 15574
rect 4080 15558 4292 15586
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15162 4200 15302
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 14822 4292 15558
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4448 15162 4476 15506
rect 4724 15502 4752 15846
rect 4816 15706 4844 16458
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4908 15094 4936 19858
rect 5000 17338 5028 23718
rect 5092 23225 5120 24346
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5078 23216 5134 23225
rect 5184 23186 5212 23802
rect 5276 23662 5304 24006
rect 5736 23866 5764 28086
rect 5828 26314 5856 29106
rect 6012 28218 6040 29582
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 6196 29306 6224 29446
rect 6184 29300 6236 29306
rect 6184 29242 6236 29248
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 6000 28212 6052 28218
rect 6000 28154 6052 28160
rect 5908 27532 5960 27538
rect 5908 27474 5960 27480
rect 5920 26586 5948 27474
rect 6012 27452 6040 28154
rect 6196 28014 6224 28494
rect 6380 28422 6408 29582
rect 6460 29096 6512 29102
rect 6460 29038 6512 29044
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6184 28008 6236 28014
rect 6184 27950 6236 27956
rect 6092 27464 6144 27470
rect 6012 27424 6092 27452
rect 6092 27406 6144 27412
rect 6196 27062 6224 27950
rect 6472 27520 6500 29038
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 6932 27674 6960 28018
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 6552 27532 6604 27538
rect 6472 27492 6552 27520
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 5908 26580 5960 26586
rect 5908 26522 5960 26528
rect 5816 26308 5868 26314
rect 5816 26250 5868 26256
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5078 23151 5134 23160
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 5184 23066 5212 23122
rect 5092 23038 5212 23066
rect 5092 20618 5120 23038
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5184 21690 5212 22034
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5276 21010 5304 23598
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 5368 23050 5396 23530
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5460 23118 5488 23462
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 5368 22930 5396 22986
rect 5368 22902 5488 22930
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5368 21962 5396 22374
rect 5460 21962 5488 22902
rect 5920 22234 5948 26522
rect 6104 25702 6132 26930
rect 6380 26450 6408 27406
rect 6472 27130 6500 27492
rect 6552 27474 6604 27480
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 6460 27124 6512 27130
rect 6460 27066 6512 27072
rect 6368 26444 6420 26450
rect 6368 26386 6420 26392
rect 7024 26042 7052 27270
rect 7116 26382 7144 28358
rect 7208 28218 7236 28494
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 7668 28218 7696 28358
rect 7196 28212 7248 28218
rect 7196 28154 7248 28160
rect 7656 28212 7708 28218
rect 7656 28154 7708 28160
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 26994 7696 27270
rect 7852 26994 7880 30126
rect 9324 29646 9352 30670
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9508 29850 9536 29990
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 8760 29640 8812 29646
rect 8760 29582 8812 29588
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 8208 29504 8260 29510
rect 8208 29446 8260 29452
rect 7932 29028 7984 29034
rect 7932 28970 7984 28976
rect 7656 26988 7708 26994
rect 7656 26930 7708 26936
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7012 26036 7064 26042
rect 7012 25978 7064 25984
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 6736 25696 6788 25702
rect 6736 25638 6788 25644
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5644 22094 5672 22170
rect 5552 22066 5672 22094
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5092 20590 5304 20618
rect 5276 20534 5304 20590
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5092 19718 5120 20402
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 19446 5120 19654
rect 5184 19514 5212 19790
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5080 19440 5132 19446
rect 5080 19382 5132 19388
rect 5092 18630 5120 19382
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5184 18970 5212 19110
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5276 18850 5304 20470
rect 5552 20262 5580 22066
rect 5908 21956 5960 21962
rect 5908 21898 5960 21904
rect 5920 21622 5948 21898
rect 5908 21616 5960 21622
rect 5908 21558 5960 21564
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5368 19514 5396 19654
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5552 19360 5580 20198
rect 5632 19372 5684 19378
rect 5552 19332 5632 19360
rect 5552 19174 5580 19332
rect 5632 19314 5684 19320
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5184 18822 5304 18850
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 16250 5028 16526
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4896 15088 4948 15094
rect 4434 15056 4490 15065
rect 4896 15030 4948 15036
rect 4434 14991 4436 15000
rect 4488 14991 4490 15000
rect 4436 14962 4488 14968
rect 4448 14906 4476 14962
rect 4448 14878 4660 14906
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14618 4660 14878
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12442 2912 12718
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 3068 11830 3096 12582
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2504 11552 2556 11558
rect 2780 11552 2832 11558
rect 2556 11512 2728 11540
rect 2504 11494 2556 11500
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2424 10696 2544 10724
rect 1952 10678 2004 10684
rect 2516 10606 2544 10696
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 2240 9518 2268 10542
rect 2424 9722 2452 10542
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9586 2544 10542
rect 2608 10266 2636 11018
rect 2700 10606 2728 11512
rect 2780 11494 2832 11500
rect 2792 11150 2820 11494
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 3160 10674 3188 12786
rect 3252 10810 3280 12786
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3344 10810 3372 11018
rect 3436 11014 3464 13874
rect 3620 13394 3648 14554
rect 3974 13968 4030 13977
rect 3974 13903 3976 13912
rect 4028 13903 4030 13912
rect 4632 13920 4660 14554
rect 4632 13892 4752 13920
rect 3976 13874 4028 13880
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3988 12442 4016 12786
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 13738
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2884 9586 2912 10474
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9722 3096 9862
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 664 9172 716 9178
rect 664 9114 716 9120
rect 676 800 704 9114
rect 2700 9042 2728 9454
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2608 7546 2636 7822
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2700 7426 2728 8978
rect 2884 8838 2912 9522
rect 3252 9382 3280 10746
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3436 10062 3464 10678
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3436 8974 3464 9454
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 3240 8832 3292 8838
rect 3528 8820 3556 12310
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3620 11898 3648 12174
rect 3608 11892 3660 11898
rect 3660 11852 3740 11880
rect 3608 11834 3660 11840
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 10198 3648 10950
rect 3712 10674 3740 11852
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4724 10810 4752 13892
rect 4816 12374 4844 14758
rect 5092 13802 5120 18566
rect 5184 17542 5212 18822
rect 5644 18426 5672 19110
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 16998 5304 17478
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5276 16182 5304 16934
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11694 4844 12174
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 11014 4844 11630
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4816 10674 4844 10950
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4724 10198 4752 10474
rect 4804 10464 4856 10470
rect 4908 10452 4936 11290
rect 4856 10424 4936 10452
rect 4804 10406 4856 10412
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 3620 9722 3648 10134
rect 4816 10130 4844 10406
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 3700 9988 3752 9994
rect 3700 9930 3752 9936
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3712 9518 3740 9930
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3620 9110 3648 9454
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3712 8838 3740 9454
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3988 8974 4016 9386
rect 3976 8968 4028 8974
rect 4080 8956 4108 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4160 8968 4212 8974
rect 4080 8928 4160 8956
rect 3976 8910 4028 8916
rect 4160 8910 4212 8916
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 3240 8774 3292 8780
rect 3436 8792 3556 8820
rect 3700 8832 3752 8838
rect 3252 8634 3280 8774
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2884 7750 2912 8434
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3146 7712 3202 7721
rect 2608 7398 2728 7426
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2148 6458 2176 7210
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2608 6322 2636 7398
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2700 6914 2728 7278
rect 2700 6886 2820 6914
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 1044 800 1072 2994
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 800 1440 2450
rect 1688 2446 1716 3334
rect 1780 3194 1808 4014
rect 2424 3670 2452 6190
rect 2700 6118 2728 6666
rect 2792 6390 2820 6886
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2792 6118 2820 6326
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2700 5166 2728 6054
rect 2792 5778 2820 6054
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 2228 3528 2280 3534
rect 2516 3482 2544 4150
rect 2884 4146 2912 7686
rect 3068 6730 3096 7686
rect 3146 7647 3202 7656
rect 3160 7342 3188 7647
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3160 6458 3188 7278
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3252 6254 3280 8570
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 6248 3292 6254
rect 3146 6216 3202 6225
rect 3068 6174 3146 6202
rect 3068 6118 3096 6174
rect 3240 6190 3292 6196
rect 3146 6151 3202 6160
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5710 3096 6054
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3068 5234 3096 5646
rect 3252 5574 3280 6190
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3056 5228 3108 5234
rect 3252 5216 3280 5510
rect 3344 5370 3372 7482
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3332 5228 3384 5234
rect 3252 5188 3332 5216
rect 3056 5170 3108 5176
rect 3332 5170 3384 5176
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3641 2636 3878
rect 2700 3738 2728 4082
rect 2870 4040 2926 4049
rect 2976 4010 3004 4422
rect 2870 3975 2926 3984
rect 2964 4004 3016 4010
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2594 3632 2650 3641
rect 2594 3567 2650 3576
rect 2228 3470 2280 3476
rect 1872 3194 1900 3470
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1964 1850 1992 3470
rect 2240 1850 2268 3470
rect 2424 3454 2544 3482
rect 2686 3496 2742 3505
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3126 2360 3334
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2424 2774 2452 3454
rect 2686 3431 2742 3440
rect 2596 3392 2648 3398
rect 2502 3360 2558 3369
rect 2596 3334 2648 3340
rect 2502 3295 2558 3304
rect 2516 2922 2544 3295
rect 2608 3058 2636 3334
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2700 2922 2728 3431
rect 2792 3126 2820 3878
rect 2884 3738 2912 3975
rect 2964 3946 3016 3952
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2962 3632 3018 3641
rect 2962 3567 3018 3576
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2424 2746 2544 2774
rect 1780 1822 1992 1850
rect 2148 1822 2268 1850
rect 1780 800 1808 1822
rect 2148 800 2176 1822
rect 2516 800 2544 2746
rect 2884 2650 2912 3470
rect 2976 3233 3004 3567
rect 2962 3224 3018 3233
rect 2962 3159 3018 3168
rect 3068 2990 3096 4694
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2976 2650 3004 2926
rect 3160 2650 3188 2994
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3252 2530 3280 4558
rect 3344 4146 3372 5170
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3641 3372 3878
rect 3330 3632 3386 3641
rect 3330 3567 3386 3576
rect 3344 3398 3372 3567
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3436 3058 3464 8792
rect 3700 8774 3752 8780
rect 3712 8294 3740 8774
rect 4172 8634 4200 8910
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4540 8498 4568 8910
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3528 7478 3556 7686
rect 3516 7472 3568 7478
rect 3516 7414 3568 7420
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6798 3556 7142
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3620 6610 3648 7686
rect 3712 7410 3740 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3896 7818 3924 8026
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3988 7528 4016 8026
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3804 7500 4016 7528
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3712 6798 3740 6938
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3528 6582 3648 6610
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3528 5710 3556 6582
rect 3712 6322 3740 6598
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 5370 3556 5646
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3712 5234 3740 6258
rect 3804 5710 3832 7500
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3896 6390 3924 6802
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 3398 3556 4966
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4282 3832 4422
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3620 3738 3648 3946
rect 3712 3738 3740 4082
rect 3896 4026 3924 5578
rect 3988 5098 4016 7346
rect 4080 5914 4108 7822
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7546 4476 7686
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 7313 4200 7346
rect 4158 7304 4214 7313
rect 4158 7239 4214 7248
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4448 6322 4476 6734
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6458 4568 6598
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5370 4108 5714
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5370 4292 5510
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 4356 5030 4384 5306
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 4622 4568 4762
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 3804 3998 3924 4026
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3712 3602 3740 3674
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3160 2502 3280 2530
rect 2884 870 3004 898
rect 2884 800 2912 870
rect 662 0 718 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 2976 762 3004 870
rect 3160 762 3188 2502
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3252 800 3280 2382
rect 3620 800 3648 2926
rect 3804 2854 3832 3998
rect 4632 3942 4660 9522
rect 4724 9110 4752 9862
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4816 8974 4844 10066
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4724 7721 4752 7754
rect 4896 7744 4948 7750
rect 4710 7712 4766 7721
rect 4766 7670 4844 7698
rect 4896 7686 4948 7692
rect 4710 7647 4766 7656
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4724 5098 4752 7482
rect 4816 7478 4844 7670
rect 4908 7546 4936 7686
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4802 7304 4858 7313
rect 4802 7239 4858 7248
rect 4816 6225 4844 7239
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6322 4936 7142
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4802 6216 4858 6225
rect 4802 6151 4858 6160
rect 4816 5370 4844 6151
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 5710 4936 6054
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4816 4554 4844 5170
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 3896 3534 3924 3878
rect 3988 3534 4016 3878
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4080 3058 4108 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4172 3466 4200 3674
rect 4264 3534 4292 3674
rect 4618 3632 4674 3641
rect 4540 3590 4618 3618
rect 4540 3534 4568 3590
rect 4618 3567 4674 3576
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4264 3194 4292 3470
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 4724 2774 4752 4490
rect 4816 4282 4844 4490
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3194 4844 4082
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4908 3058 4936 4422
rect 5000 4298 5028 12106
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5184 11558 5212 11766
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5092 10198 5120 10746
rect 5184 10606 5212 11494
rect 5276 11286 5304 11834
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5276 10810 5304 11222
rect 5368 10810 5396 16050
rect 5460 16046 5488 16390
rect 5552 16250 5580 16934
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5092 8906 5120 10134
rect 5184 9722 5212 10542
rect 5276 10266 5304 10746
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5460 9654 5488 15982
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5644 15162 5672 15302
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5552 10198 5580 11222
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5276 7002 5304 7890
rect 5460 7478 5488 8026
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 6458 5212 6734
rect 5552 6458 5580 7210
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5184 5778 5212 6190
rect 5368 5914 5396 6258
rect 5644 5914 5672 13670
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5644 5370 5672 5850
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5276 4622 5304 5170
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5000 4270 5120 4298
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 3602 5028 4082
rect 5092 4049 5120 4270
rect 5078 4040 5134 4049
rect 5078 3975 5134 3984
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5184 3466 5212 3946
rect 5276 3466 5304 4558
rect 5368 4078 5396 4966
rect 5644 4622 5672 5306
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5184 3233 5212 3402
rect 5170 3224 5226 3233
rect 5170 3159 5226 3168
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5368 2990 5396 3878
rect 5460 3670 5488 4558
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5736 3534 5764 18566
rect 5920 12442 5948 21558
rect 6104 21350 6132 25638
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6196 21894 6224 22442
rect 6288 21962 6316 23598
rect 6380 23225 6408 24142
rect 6366 23216 6422 23225
rect 6366 23151 6422 23160
rect 6380 22778 6408 23151
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 19334 6132 19858
rect 6012 19306 6132 19334
rect 6012 15978 6040 19306
rect 6196 18850 6224 21830
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6380 19922 6408 20334
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6288 19446 6316 19722
rect 6276 19440 6328 19446
rect 6276 19382 6328 19388
rect 6092 18828 6144 18834
rect 6196 18822 6316 18850
rect 6092 18770 6144 18776
rect 6104 18086 6132 18770
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6104 14958 6132 18022
rect 6196 17746 6224 18566
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 16046 6224 16526
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6012 10470 6040 14010
rect 6104 13734 6132 14894
rect 6196 14890 6224 15982
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6196 14414 6224 14826
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6196 12306 6224 14350
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7002 5948 7822
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 6322 5856 6734
rect 6012 6322 6040 8230
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5920 5234 5948 5510
rect 6012 5370 6040 5646
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6012 5234 6040 5306
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 5920 5098 5948 5170
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5920 4622 5948 5034
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 4282 5856 4422
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 6012 3942 6040 4966
rect 6196 4078 6224 8298
rect 6288 5914 6316 18822
rect 6380 18766 6408 19858
rect 6472 19718 6500 20810
rect 6656 20058 6684 20878
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6380 18290 6408 18702
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6656 17882 6684 18226
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6380 13852 6408 15914
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 15162 6500 15302
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6656 14074 6684 15098
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6380 13824 6592 13852
rect 6564 13394 6592 13824
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6380 11354 6408 12786
rect 6564 12434 6592 13330
rect 6564 12406 6684 12434
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6288 5370 6316 5850
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6288 4690 6316 5306
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 4214 6316 4490
rect 6380 4214 6408 6258
rect 6472 4826 6500 11834
rect 6656 11626 6684 12406
rect 6748 11898 6776 25638
rect 7668 25498 7696 26182
rect 7852 25906 7880 26930
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7656 25492 7708 25498
rect 7656 25434 7708 25440
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 7024 24954 7052 25230
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6840 23322 6868 24074
rect 7024 23730 7052 24686
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 6932 23066 6960 23122
rect 6840 23038 6960 23066
rect 6840 22658 6868 23038
rect 7024 22982 7052 23666
rect 7116 23662 7144 24142
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7104 23520 7156 23526
rect 7208 23508 7236 24618
rect 7392 24410 7420 24754
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7156 23480 7236 23508
rect 7104 23462 7156 23468
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6932 22778 6960 22918
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6840 22630 6960 22658
rect 6932 22234 6960 22630
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7024 22094 7052 22918
rect 7392 22556 7420 23122
rect 7576 22710 7604 25094
rect 7668 23322 7696 25434
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7760 23866 7788 25094
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 7654 23216 7710 23225
rect 7654 23151 7710 23160
rect 7668 23118 7696 23151
rect 7665 23112 7717 23118
rect 7665 23054 7717 23060
rect 7564 22704 7616 22710
rect 7564 22646 7616 22652
rect 7852 22642 7880 23462
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7392 22528 7604 22556
rect 7024 22066 7144 22094
rect 7116 22030 7144 22066
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7208 20534 7236 20742
rect 7196 20528 7248 20534
rect 7196 20470 7248 20476
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6932 19446 6960 19654
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6932 18970 6960 19246
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 17814 6868 18566
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 16182 6960 16934
rect 7024 16794 7052 17070
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 7024 15586 7052 16730
rect 7116 16658 7144 19110
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 6932 15570 7052 15586
rect 6920 15564 7052 15570
rect 6972 15558 7052 15564
rect 6920 15506 6972 15512
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7116 15366 7144 15438
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7392 14618 7420 15438
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 7024 14006 7052 14282
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6932 12434 6960 13194
rect 6840 12406 6960 12434
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6564 11354 6592 11494
rect 6748 11354 6776 11630
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 10810 6868 12406
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 10810 6960 11698
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6748 8090 6776 8434
rect 6840 8294 6868 10406
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 7024 6798 7052 13942
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7300 11898 7328 12718
rect 7484 12434 7512 20402
rect 7576 19310 7604 22528
rect 7852 22098 7880 22578
rect 7944 22098 7972 28970
rect 8024 28960 8076 28966
rect 8024 28902 8076 28908
rect 8036 28014 8064 28902
rect 8220 28218 8248 29446
rect 8772 29102 8800 29582
rect 9864 29504 9916 29510
rect 9864 29446 9916 29452
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9784 28218 9812 28494
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 8036 26994 8064 27950
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 8404 26586 8432 27406
rect 9048 27062 9076 27814
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 9036 27056 9088 27062
rect 9036 26998 9088 27004
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8760 26308 8812 26314
rect 8760 26250 8812 26256
rect 8116 26036 8168 26042
rect 8116 25978 8168 25984
rect 8128 22574 8156 25978
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8220 23866 8248 24550
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8404 23662 8432 25230
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8404 23254 8432 23598
rect 8392 23248 8444 23254
rect 8392 23190 8444 23196
rect 8588 23186 8616 23802
rect 8680 23186 8708 24006
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8576 22704 8628 22710
rect 8496 22664 8576 22692
rect 8116 22568 8168 22574
rect 8116 22510 8168 22516
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8036 22273 8064 22374
rect 8022 22264 8078 22273
rect 8022 22199 8078 22208
rect 7840 22092 7892 22098
rect 7840 22034 7892 22040
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 8312 21894 8340 22374
rect 8496 22098 8524 22664
rect 8576 22646 8628 22652
rect 8680 22642 8708 23122
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7760 20262 7788 20878
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 19378 7788 20198
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7576 18426 7604 19246
rect 7852 18426 7880 19246
rect 7944 18970 7972 21626
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8312 20806 8340 21286
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8312 19242 8340 20742
rect 8404 20466 8432 20810
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7852 17746 7880 18362
rect 8312 18086 8340 19178
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16794 7604 17070
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7668 15094 7696 16934
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 16250 7788 16390
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7852 15638 7880 17206
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7852 15162 7880 15574
rect 8220 15570 8248 15914
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8220 15162 8248 15506
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14278 8248 14758
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7392 12406 7512 12434
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 8498 7236 11086
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 7342 7236 8434
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7546 7328 7822
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7024 6458 7052 6734
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7208 5778 7236 7278
rect 7392 6390 7420 12406
rect 7668 12238 7696 12582
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7746 12200 7802 12209
rect 7746 12135 7802 12144
rect 7760 11880 7788 12135
rect 7668 11852 7788 11880
rect 7668 10198 7696 11852
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7760 9654 7788 11698
rect 7852 10198 7880 13738
rect 7944 12986 7972 13806
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7944 11642 7972 12922
rect 8128 11898 8156 13126
rect 8220 12209 8248 14214
rect 8312 14006 8340 18022
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16250 8432 17070
rect 8496 17066 8524 22034
rect 8588 21690 8616 22510
rect 8772 22506 8800 26250
rect 9232 26042 9260 27338
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9416 27130 9444 27270
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9600 26586 9628 26862
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 8852 24744 8904 24750
rect 8852 24686 8904 24692
rect 8864 23322 8892 24686
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9048 23866 9076 24142
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 9324 23118 9352 24006
rect 9508 23304 9536 26318
rect 9692 26042 9720 27950
rect 9876 26926 9904 29446
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9968 27674 9996 28494
rect 9956 27668 10008 27674
rect 9956 27610 10008 27616
rect 9968 27130 9996 27610
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9876 26518 9904 26862
rect 9864 26512 9916 26518
rect 9864 26454 9916 26460
rect 10060 26058 10088 31214
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 10152 30190 10180 30534
rect 10140 30184 10192 30190
rect 10140 30126 10192 30132
rect 10152 26874 10180 30126
rect 10336 29646 10364 31078
rect 10428 30258 10456 31758
rect 10600 31680 10652 31686
rect 10600 31622 10652 31628
rect 10612 30734 10640 31622
rect 11060 31340 11112 31346
rect 11060 31282 11112 31288
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 10888 30938 10916 31214
rect 10876 30932 10928 30938
rect 10876 30874 10928 30880
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 11072 30598 11100 31282
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 11152 30252 11204 30258
rect 11152 30194 11204 30200
rect 10428 30054 10456 30194
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 10416 30048 10468 30054
rect 10416 29990 10468 29996
rect 10324 29640 10376 29646
rect 10324 29582 10376 29588
rect 10612 29306 10640 30126
rect 10784 30116 10836 30122
rect 10784 30058 10836 30064
rect 10796 29510 10824 30058
rect 11164 29850 11192 30194
rect 11256 30190 11284 31758
rect 13268 31680 13320 31686
rect 13268 31622 13320 31628
rect 13280 31482 13308 31622
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11348 30802 11376 31078
rect 11532 30938 11560 31214
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11336 30796 11388 30802
rect 11336 30738 11388 30744
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 11152 29844 11204 29850
rect 11152 29786 11204 29792
rect 11244 29776 11296 29782
rect 11244 29718 11296 29724
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 11152 29504 11204 29510
rect 11152 29446 11204 29452
rect 10600 29300 10652 29306
rect 10600 29242 10652 29248
rect 10796 28762 10824 29446
rect 11072 29170 11100 29446
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10428 27470 10456 28358
rect 10520 28218 10548 28358
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 11060 28008 11112 28014
rect 11060 27950 11112 27956
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10416 27464 10468 27470
rect 10416 27406 10468 27412
rect 10416 27328 10468 27334
rect 10416 27270 10468 27276
rect 10428 27130 10456 27270
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10428 26994 10456 27066
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10152 26858 10272 26874
rect 10152 26852 10284 26858
rect 10152 26846 10232 26852
rect 10232 26794 10284 26800
rect 10244 26314 10272 26794
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 9680 26036 9732 26042
rect 10060 26030 10180 26058
rect 9680 25978 9732 25984
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 23866 9628 24550
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9588 23316 9640 23322
rect 9508 23276 9588 23304
rect 9588 23258 9640 23264
rect 9600 23186 9628 23258
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 8760 22500 8812 22506
rect 8760 22442 8812 22448
rect 9600 22438 9628 23122
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8576 19712 8628 19718
rect 8628 19660 8708 19666
rect 8576 19654 8708 19660
rect 8588 19638 8708 19654
rect 8680 19378 8708 19638
rect 8864 19378 8892 19994
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9508 19514 9536 19790
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8852 19372 8904 19378
rect 9600 19334 9628 22374
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20398 9720 20742
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9692 19922 9720 20334
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 8852 19314 8904 19320
rect 8588 18970 8616 19314
rect 9508 19310 9628 19334
rect 9496 19306 9628 19310
rect 9496 19304 9548 19306
rect 9496 19246 9548 19252
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8864 18834 8892 19110
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8496 16250 8524 16526
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8404 15162 8432 15982
rect 8496 15570 8524 16186
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8588 14958 8616 18702
rect 9508 18630 9536 19246
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8680 16658 8708 17002
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 9232 16046 9260 18566
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8496 14618 8524 14894
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8588 14346 8616 14894
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12442 8340 12786
rect 8772 12442 8800 13262
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8392 12232 8444 12238
rect 8206 12200 8262 12209
rect 8392 12174 8444 12180
rect 8206 12135 8262 12144
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11642 8064 11698
rect 7944 11614 8064 11642
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 10810 7972 11494
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 7410 7512 9318
rect 7668 9110 7696 9522
rect 7852 9518 7880 10134
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8036 9722 8064 9998
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 8128 8906 8156 9318
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8634 8156 8842
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8128 7750 8156 8366
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 8128 6866 8156 7686
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7392 6225 7420 6326
rect 7378 6216 7434 6225
rect 7378 6151 7434 6160
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6564 4554 6592 4966
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 4146 6500 4422
rect 6840 4282 6868 4558
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5460 3369 5488 3470
rect 5540 3392 5592 3398
rect 5446 3360 5502 3369
rect 5540 3334 5592 3340
rect 5446 3295 5502 3304
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2746 4752 2774
rect 4356 870 4476 898
rect 4356 800 4384 870
rect 2976 734 3188 762
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4448 762 4476 870
rect 4632 762 4660 2746
rect 5552 2446 5580 3334
rect 6012 2854 6040 3674
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6104 2854 6132 3402
rect 6288 3194 6316 3470
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 4724 800 4752 2382
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 5092 800 5120 2314
rect 5644 1306 5672 2450
rect 5644 1278 5856 1306
rect 5828 800 5856 1278
rect 6196 800 6224 2926
rect 6656 2446 6684 3062
rect 7024 2990 7052 4694
rect 7208 4622 7236 5714
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4078 7144 4490
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7208 3602 7236 4558
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6380 2106 6408 2382
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6564 870 6684 898
rect 6564 800 6592 870
rect 4448 734 4660 762
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6656 762 6684 870
rect 6840 762 6868 2450
rect 7300 800 7328 5578
rect 7392 4826 7420 6151
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5166 7512 6054
rect 8220 5914 8248 12038
rect 8404 11830 8432 12174
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8392 11688 8444 11694
rect 8298 11656 8354 11665
rect 8392 11630 8444 11636
rect 8298 11591 8354 11600
rect 8312 11354 8340 11591
rect 8404 11354 8432 11630
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8312 7818 8340 11290
rect 8496 10810 8524 12106
rect 8772 11694 8800 12378
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8588 10470 8616 11562
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8772 10674 8800 11290
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8864 10146 8892 15846
rect 9232 15366 9260 15982
rect 9324 15434 9352 16934
rect 9784 15706 9812 25774
rect 10060 25498 10088 25842
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10152 24818 10180 26030
rect 10520 25770 10548 26930
rect 10612 26042 10640 27814
rect 10704 26790 10732 27950
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10704 25906 10732 26726
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10508 25764 10560 25770
rect 10508 25706 10560 25712
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9876 22778 9904 22918
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9876 20330 9904 22714
rect 10152 22094 10180 24754
rect 10324 23792 10376 23798
rect 10324 23734 10376 23740
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 10244 23118 10272 23598
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10244 22642 10272 23054
rect 10336 22778 10364 23734
rect 10692 23044 10744 23050
rect 10692 22986 10744 22992
rect 10704 22778 10732 22986
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 9968 22066 10180 22094
rect 9968 21962 9996 22066
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 20534 9996 21286
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9876 20058 9904 20266
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 10060 18970 10088 22066
rect 10244 20806 10272 22578
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10232 19712 10284 19718
rect 10336 19700 10364 21830
rect 10600 21480 10652 21486
rect 10600 21422 10652 21428
rect 10612 21146 10640 21422
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10284 19672 10364 19700
rect 10232 19654 10284 19660
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10060 18426 10088 18906
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 10060 17678 10088 18362
rect 10244 18086 10272 19654
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 17202 10088 17478
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9876 16250 9904 17002
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9968 16794 9996 16934
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9324 15026 9352 15370
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9048 14618 9076 14758
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8956 10674 8984 11222
rect 9048 10810 9076 13806
rect 9140 12186 9168 14282
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9232 12918 9260 13670
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9232 12356 9260 12854
rect 9324 12628 9352 14962
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9416 13734 9444 14010
rect 9496 13864 9548 13870
rect 9494 13832 9496 13841
rect 9548 13832 9550 13841
rect 9494 13767 9550 13776
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 12850 9444 13670
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9508 12764 9536 13767
rect 9508 12736 9628 12764
rect 9324 12600 9536 12628
rect 9232 12328 9352 12356
rect 9140 12170 9260 12186
rect 9140 12164 9272 12170
rect 9140 12158 9220 12164
rect 9140 11558 9168 12158
rect 9220 12106 9272 12112
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9232 11354 9260 11630
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8668 10124 8720 10130
rect 8864 10118 8984 10146
rect 8668 10066 8720 10072
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 7818 8432 9454
rect 8496 8974 8524 9862
rect 8680 9518 8708 10066
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8680 8906 8708 9454
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7576 5370 7604 5646
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7392 3670 7420 4762
rect 7484 4282 7512 5102
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7760 4214 7788 4966
rect 7944 4554 7972 5034
rect 8312 4690 8340 6598
rect 8588 6390 8616 6734
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8680 6202 8708 8298
rect 8772 7954 8800 8910
rect 8864 8498 8892 9998
rect 8956 9382 8984 10118
rect 9048 9586 9076 10406
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 9042 8984 9318
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 9048 8838 9076 9522
rect 9324 8922 9352 12328
rect 9404 11688 9456 11694
rect 9508 11676 9536 12600
rect 9600 12238 9628 12736
rect 9692 12306 9720 15302
rect 9876 12850 9904 16186
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9692 11898 9720 12242
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9456 11648 9536 11676
rect 9588 11688 9640 11694
rect 9404 11630 9456 11636
rect 9588 11630 9640 11636
rect 9416 11354 9444 11630
rect 9404 11348 9456 11354
rect 9456 11308 9536 11336
rect 9404 11290 9456 11296
rect 9232 8894 9352 8922
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8956 8498 8984 8774
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 6662 8800 7890
rect 8956 7342 8984 8434
rect 9048 7410 9076 8774
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 9048 6458 9076 7346
rect 9232 7342 9260 8894
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9232 6798 9260 7278
rect 9324 6866 9352 8774
rect 9508 8430 9536 11308
rect 9600 10538 9628 11630
rect 9876 10606 9904 12786
rect 9968 10690 9996 15370
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10152 12782 10180 14350
rect 10244 13394 10272 18022
rect 10428 13938 10456 20538
rect 10704 19854 10732 21286
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 16590 10548 18566
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10704 17746 10732 18022
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 13802 10456 13874
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10520 13530 10548 13670
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10336 12434 10364 13126
rect 10612 12850 10640 13670
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10796 12434 10824 27270
rect 10888 26382 10916 27610
rect 10968 27124 11020 27130
rect 11072 27112 11100 27950
rect 11164 27418 11192 29446
rect 11256 27538 11284 29718
rect 11348 29594 11376 30738
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11440 30394 11468 30670
rect 11428 30388 11480 30394
rect 11428 30330 11480 30336
rect 11532 30258 11560 30874
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11612 30252 11664 30258
rect 11716 30240 11744 30534
rect 12176 30394 12204 31078
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12164 30388 12216 30394
rect 12164 30330 12216 30336
rect 12636 30258 12664 30670
rect 12912 30326 12940 31078
rect 13464 30666 13492 32166
rect 14108 32026 14136 32302
rect 14280 32224 14332 32230
rect 14280 32166 14332 32172
rect 14292 32026 14320 32166
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 13912 31816 13964 31822
rect 13912 31758 13964 31764
rect 13636 31680 13688 31686
rect 13636 31622 13688 31628
rect 13648 31278 13676 31622
rect 13636 31272 13688 31278
rect 13636 31214 13688 31220
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13452 30660 13504 30666
rect 13452 30602 13504 30608
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 11664 30212 11744 30240
rect 12624 30252 12676 30258
rect 11612 30194 11664 30200
rect 12624 30194 12676 30200
rect 11348 29566 11468 29594
rect 11336 29504 11388 29510
rect 11336 29446 11388 29452
rect 11348 28082 11376 29446
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 11164 27390 11284 27418
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11164 27130 11192 27270
rect 11020 27084 11100 27112
rect 11152 27124 11204 27130
rect 10968 27066 11020 27072
rect 11152 27066 11204 27072
rect 11256 27010 11284 27390
rect 11072 26982 11284 27010
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 25362 11008 26182
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 11072 24750 11100 26982
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11256 26314 11284 26862
rect 11440 26602 11468 29566
rect 11624 29510 11652 30194
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11612 29504 11664 29510
rect 11612 29446 11664 29452
rect 11808 29306 11836 29650
rect 12636 29306 12664 30194
rect 13648 30138 13676 31214
rect 13740 30802 13768 31214
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13924 30394 13952 31758
rect 14740 31748 14792 31754
rect 14740 31690 14792 31696
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 13912 30388 13964 30394
rect 13912 30330 13964 30336
rect 13648 30110 13768 30138
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12912 29714 12940 29990
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 11520 28008 11572 28014
rect 11520 27950 11572 27956
rect 11348 26574 11468 26602
rect 11532 26586 11560 27950
rect 12164 27872 12216 27878
rect 12164 27814 12216 27820
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11624 27130 11652 27270
rect 12176 27130 12204 27814
rect 12544 27470 12572 27814
rect 12636 27674 12664 29242
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12268 27130 12296 27406
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 12256 27124 12308 27130
rect 12256 27066 12308 27072
rect 11704 26920 11756 26926
rect 11704 26862 11756 26868
rect 11520 26580 11572 26586
rect 11348 26518 11376 26574
rect 11520 26522 11572 26528
rect 11336 26512 11388 26518
rect 11336 26454 11388 26460
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11164 26042 11192 26182
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 11244 25968 11296 25974
rect 11244 25910 11296 25916
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 11164 25226 11192 25774
rect 11256 25362 11284 25910
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10888 24206 10916 24550
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10888 22098 10916 24142
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21146 11100 21830
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11060 20868 11112 20874
rect 11164 20856 11192 25162
rect 11440 25158 11468 26386
rect 11612 26240 11664 26246
rect 11612 26182 11664 26188
rect 11624 25838 11652 26182
rect 11716 26042 11744 26862
rect 11796 26784 11848 26790
rect 11796 26726 11848 26732
rect 11808 26314 11836 26726
rect 12544 26518 12572 27406
rect 12636 27130 12664 27610
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 12728 27130 12756 27270
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12820 26586 12848 27270
rect 12808 26580 12860 26586
rect 12808 26522 12860 26528
rect 12532 26512 12584 26518
rect 12532 26454 12584 26460
rect 13004 26450 13032 27814
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13096 26586 13124 27406
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 12992 26444 13044 26450
rect 12992 26386 13044 26392
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 13096 26042 13124 26182
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 11612 25832 11664 25838
rect 11612 25774 11664 25780
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11348 22234 11376 22510
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11440 21350 11468 25094
rect 12728 24954 12756 25094
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 12084 24342 12112 24550
rect 12072 24336 12124 24342
rect 12072 24278 12124 24284
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11624 22710 11652 24006
rect 11808 22710 11836 24006
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11440 21010 11468 21286
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11112 20828 11192 20856
rect 11060 20810 11112 20816
rect 11072 20602 11100 20810
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11440 20466 11468 20946
rect 11624 20602 11652 21966
rect 12452 21894 12480 22646
rect 12544 22642 12572 23734
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12728 23322 12756 23666
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12728 23118 12756 23258
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11716 21146 11744 21558
rect 12452 21554 12480 21830
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11716 20466 11744 21082
rect 12360 20618 12388 21422
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 12452 20942 12480 21354
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12268 20590 12388 20618
rect 12268 20466 12296 20590
rect 12544 20482 12572 22578
rect 12728 22094 12756 23054
rect 12912 22098 12940 23054
rect 13004 22778 13032 24686
rect 13280 23322 13308 25230
rect 13372 24070 13400 29650
rect 13740 29646 13768 30110
rect 13728 29640 13780 29646
rect 13728 29582 13780 29588
rect 13740 29238 13768 29582
rect 14108 29306 14136 31282
rect 14660 30734 14688 31622
rect 14752 31414 14780 31690
rect 14740 31408 14792 31414
rect 14740 31350 14792 31356
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 14752 30666 14780 31350
rect 15028 30938 15056 32302
rect 23940 32292 23992 32298
rect 23940 32234 23992 32240
rect 23952 32026 23980 32234
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 24044 32026 24072 32166
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 19064 31816 19116 31822
rect 19064 31758 19116 31764
rect 19248 31816 19300 31822
rect 19248 31758 19300 31764
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 14740 30660 14792 30666
rect 14740 30602 14792 30608
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14568 29850 14596 30126
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14752 29510 14780 30602
rect 14924 30388 14976 30394
rect 14924 30330 14976 30336
rect 14936 30258 14964 30330
rect 15028 30258 15056 30874
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15200 30116 15252 30122
rect 15200 30058 15252 30064
rect 15212 30002 15240 30058
rect 15028 29974 15240 30002
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14096 29300 14148 29306
rect 14096 29242 14148 29248
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 13820 28960 13872 28966
rect 13820 28902 13872 28908
rect 13832 28490 13860 28902
rect 14464 28552 14516 28558
rect 14464 28494 14516 28500
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 14476 28218 14504 28494
rect 14648 28484 14700 28490
rect 14648 28426 14700 28432
rect 14464 28212 14516 28218
rect 14464 28154 14516 28160
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 14004 28008 14056 28014
rect 14004 27950 14056 27956
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13556 27470 13584 27814
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 13832 27130 13860 27950
rect 14016 27402 14044 27950
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14004 27396 14056 27402
rect 14004 27338 14056 27344
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 13820 27124 13872 27130
rect 13820 27066 13872 27072
rect 13924 26926 13952 27270
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 14016 26246 14044 27338
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14096 26852 14148 26858
rect 14096 26794 14148 26800
rect 14108 26586 14136 26794
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 13544 25968 13596 25974
rect 13544 25910 13596 25916
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13464 23798 13492 24550
rect 13556 24206 13584 25910
rect 14200 25498 14228 26862
rect 14292 25838 14320 27814
rect 14660 26858 14688 28426
rect 14752 28150 14780 29446
rect 15028 28762 15056 29974
rect 15304 29714 15332 31078
rect 15580 30938 15608 31758
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 16120 31476 16172 31482
rect 16120 31418 16172 31424
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15568 30932 15620 30938
rect 15568 30874 15620 30880
rect 15752 30864 15804 30870
rect 15752 30806 15804 30812
rect 15764 30258 15792 30806
rect 15856 30258 15884 31214
rect 16132 30802 16160 31418
rect 18524 31346 18552 31622
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18236 31272 18288 31278
rect 18236 31214 18288 31220
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 16132 30598 16160 30738
rect 18248 30734 18276 31214
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 16120 30592 16172 30598
rect 16120 30534 16172 30540
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16132 30394 16160 30534
rect 16120 30388 16172 30394
rect 16120 30330 16172 30336
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 15120 29102 15148 29446
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 14740 28144 14792 28150
rect 14740 28086 14792 28092
rect 15028 28014 15056 28358
rect 15212 28218 15240 29106
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15200 28212 15252 28218
rect 15200 28154 15252 28160
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14648 26852 14700 26858
rect 14648 26794 14700 26800
rect 14660 26314 14688 26794
rect 14752 26382 14780 27610
rect 14832 27124 14884 27130
rect 14832 27066 14884 27072
rect 14844 26994 14872 27066
rect 14936 26994 14964 27814
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14556 26240 14608 26246
rect 14556 26182 14608 26188
rect 14568 25906 14596 26182
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14740 25832 14792 25838
rect 14740 25774 14792 25780
rect 14752 25498 14780 25774
rect 14936 25770 14964 26930
rect 14924 25764 14976 25770
rect 14924 25706 14976 25712
rect 15028 25498 15056 27950
rect 14188 25492 14240 25498
rect 14188 25434 14240 25440
rect 14464 25492 14516 25498
rect 14464 25434 14516 25440
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13648 23730 13676 24754
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13924 24410 13952 24686
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12728 22066 12848 22094
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12636 20874 12664 21490
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12360 20454 12572 20482
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11992 20058 12020 20198
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12256 19508 12308 19514
rect 12360 19496 12388 20454
rect 12544 20398 12572 20454
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12452 19718 12480 20334
rect 12636 19854 12664 20810
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12308 19468 12388 19496
rect 12256 19450 12308 19456
rect 12636 19378 12664 19790
rect 12728 19514 12756 21286
rect 12820 21026 12848 22066
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12820 20998 13124 21026
rect 13188 21010 13216 22918
rect 13280 22574 13308 23258
rect 13360 23248 13412 23254
rect 13360 23190 13412 23196
rect 13372 22642 13400 23190
rect 13648 22710 13676 23666
rect 13740 23662 13768 24006
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13832 23662 13860 23802
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13820 23656 13872 23662
rect 13820 23598 13872 23604
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13740 23186 13768 23462
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 13924 23118 13952 24346
rect 14200 23730 14228 25434
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14292 23866 14320 24550
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22778 14136 22918
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13740 21010 13768 21626
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 11888 19304 11940 19310
rect 11518 19272 11574 19281
rect 12256 19304 12308 19310
rect 11940 19252 12256 19258
rect 11888 19246 12308 19252
rect 11900 19230 12296 19246
rect 11518 19207 11520 19216
rect 11572 19207 11574 19216
rect 11520 19178 11572 19184
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12268 18834 12296 19110
rect 12820 18970 12848 20810
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12912 20466 12940 20538
rect 13096 20466 13124 20998
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 19378 12940 19654
rect 13096 19514 13124 20402
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11532 18426 11560 18702
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12360 18170 12388 18362
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11072 17134 11100 17478
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 15162 11008 17002
rect 11072 16114 11100 17070
rect 11348 16998 11376 18158
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11716 16590 11744 17070
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 12268 16250 12296 18158
rect 12360 18142 12480 18170
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12360 17678 12388 18022
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12452 17542 12480 18142
rect 12728 17746 12756 18906
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12452 16946 12480 17478
rect 12624 17128 12676 17134
rect 12676 17076 12756 17082
rect 12624 17070 12756 17076
rect 12636 17054 12756 17070
rect 12452 16918 12572 16946
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11256 14278 11284 15438
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11624 15026 11652 15302
rect 12452 15094 12480 16730
rect 12544 16114 12572 16918
rect 12728 16454 12756 17054
rect 12912 16794 12940 17478
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12544 15502 12572 16050
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11348 14618 11376 14894
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 12268 14482 12296 14758
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10244 12406 10364 12434
rect 10612 12406 10824 12434
rect 10244 12238 10272 12406
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10060 10810 10088 11018
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9968 10662 10088 10690
rect 10152 10674 10180 11494
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9876 10198 9904 10542
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 8022 9536 8366
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 7478 9444 7822
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 8680 6174 8800 6202
rect 8772 6118 8800 6174
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8576 5704 8628 5710
rect 8680 5681 8708 6054
rect 8576 5646 8628 5652
rect 8666 5672 8722 5681
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 3058 7512 3334
rect 7576 3194 7604 4082
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7760 3058 7788 4150
rect 8312 4146 8340 4626
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 8300 4004 8352 4010
rect 7852 3058 7880 3975
rect 8300 3946 8352 3952
rect 8312 3534 8340 3946
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7668 800 7696 2382
rect 8220 1578 8248 2926
rect 8404 2650 8432 5646
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8496 3602 8524 5578
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 2774 8616 5646
rect 8666 5607 8722 5616
rect 9128 5636 9180 5642
rect 8680 5234 8708 5607
rect 9128 5578 9180 5584
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8680 4826 8708 5170
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8772 3942 8800 5510
rect 9140 4622 9168 5578
rect 9232 5370 9260 6258
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 9140 3618 9168 4558
rect 9508 4214 9536 7958
rect 9600 7546 9628 9862
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 7886 9720 8774
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 10060 8242 10088 10662
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10244 10266 10272 12174
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10336 8634 10364 11562
rect 10520 10606 10548 11698
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10428 8430 10456 9454
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9680 7744 9732 7750
rect 9784 7732 9812 7822
rect 9732 7704 9812 7732
rect 9680 7686 9732 7692
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6186 9720 7142
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5778 9720 6122
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9692 4298 9720 4626
rect 9784 4622 9812 5510
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9600 4270 9720 4298
rect 9600 4214 9628 4270
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9772 4140 9824 4146
rect 9876 4128 9904 8230
rect 10060 8214 10364 8242
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7750 10088 7958
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6118 9996 6598
rect 10152 6186 10180 7754
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4826 9996 5102
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10060 4214 10088 4966
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9876 4100 9996 4128
rect 9772 4082 9824 4088
rect 9416 3738 9444 4082
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9048 3590 9168 3618
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3194 8800 3334
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9048 3058 9076 3590
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9232 3126 9260 3470
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9416 2774 9444 3470
rect 8588 2746 8800 2774
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8036 1550 8248 1578
rect 8036 800 8064 1550
rect 8772 800 8800 2746
rect 9140 2746 9444 2774
rect 9140 800 9168 2746
rect 9508 2650 9536 4014
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9600 1578 9628 2926
rect 9784 2514 9812 4082
rect 9968 4010 9996 4100
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 10152 3670 10180 5170
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9968 2446 9996 3606
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 9508 1550 9628 1578
rect 9508 800 9536 1550
rect 9876 800 9904 2042
rect 10244 800 10272 3470
rect 10336 3398 10364 8214
rect 10428 7206 10456 8366
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 5166 10456 6734
rect 10520 6458 10548 8842
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10612 4554 10640 12406
rect 10980 11898 11008 13738
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11348 12986 11376 13194
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11440 12442 11468 14282
rect 11980 14068 12032 14074
rect 12452 14056 12480 15030
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12532 14068 12584 14074
rect 12452 14028 12532 14056
rect 11980 14010 12032 14016
rect 12532 14010 12584 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11808 12714 11836 13874
rect 11992 13326 12020 14010
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11992 11762 12020 13262
rect 12544 12918 12572 13806
rect 12636 13530 12664 14350
rect 12728 14278 12756 14418
rect 12820 14278 12848 15370
rect 12912 15162 12940 15438
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 13004 14482 13032 14826
rect 13096 14822 13124 17070
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12728 12918 12756 14214
rect 12820 13938 12848 14214
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12306 12204 12582
rect 12452 12442 12480 12718
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 11354 12020 11698
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11532 10810 11560 11018
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 7818 10732 8230
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7342 11008 7686
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 7002 11008 7278
rect 11072 7206 11100 8026
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11072 6662 11100 7142
rect 11256 6866 11284 9318
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11348 8634 11376 8774
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11624 7954 11652 8366
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5846 10916 6122
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10888 5370 10916 5510
rect 10980 5370 11008 6054
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11072 5030 11100 6598
rect 11532 6458 11560 6734
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11440 6361 11468 6394
rect 11426 6352 11482 6361
rect 11426 6287 11482 6296
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11256 4758 11284 6190
rect 11440 5778 11468 6287
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11348 5234 11376 5646
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11058 4584 11114 4593
rect 10600 4548 10652 4554
rect 11058 4519 11114 4528
rect 10600 4490 10652 4496
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10428 3058 10456 4422
rect 10520 3602 10548 4422
rect 11072 4282 11100 4519
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11164 3670 11192 4626
rect 11256 4078 11284 4694
rect 11532 4690 11560 6190
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11716 5234 11744 5510
rect 11808 5234 11836 8230
rect 12084 8090 12112 9862
rect 12176 9382 12204 12106
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10674 12480 10950
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12544 9654 12572 12854
rect 13188 12434 13216 20742
rect 13464 19922 13492 20878
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20602 13584 20742
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13832 20262 13860 20878
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 14016 19718 14044 20334
rect 14004 19712 14056 19718
rect 14056 19660 14136 19666
rect 14004 19654 14136 19660
rect 14016 19638 14136 19654
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17270 13308 17478
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13280 16522 13308 17002
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13372 15162 13400 16934
rect 13648 16590 13676 18158
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13832 15570 13860 19246
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13372 14618 13400 14962
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13556 14414 13584 15438
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13464 13530 13492 14350
rect 13740 13818 13768 14758
rect 13556 13790 13768 13818
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13188 12406 13308 12434
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12728 10606 12756 12038
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13004 10606 13032 11290
rect 13096 10810 13124 12038
rect 13188 11762 13216 12038
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 9994 12848 10474
rect 13188 10266 13216 10542
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12912 9674 12940 10066
rect 12532 9648 12584 9654
rect 12912 9646 13032 9674
rect 12532 9590 12584 9596
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 9042 12204 9318
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8566 12480 8774
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 6866 11928 7822
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 7002 12204 7754
rect 12256 7336 12308 7342
rect 12308 7296 12388 7324
rect 12256 7278 12308 7284
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12176 5914 12204 6190
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12084 5642 12112 5782
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12268 5234 12296 6598
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4690 11744 4966
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12176 4690 12204 4762
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12360 4622 12388 7296
rect 12452 6458 12480 8502
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12452 5914 12480 6394
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12452 5370 12480 5850
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11348 4282 11376 4558
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3126 10824 3470
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10888 2774 10916 3402
rect 11256 3194 11284 3839
rect 12176 3738 12204 4082
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11440 2922 11468 2994
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 10888 2746 11008 2774
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10612 800 10640 2450
rect 10980 800 11008 2746
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 1306 11192 2246
rect 11532 1562 11560 2994
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11164 1278 11376 1306
rect 11348 800 11376 1278
rect 11716 870 11836 898
rect 11716 800 11744 870
rect 6656 734 6868 762
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 11808 762 11836 870
rect 11992 762 12020 2926
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 12084 800 12112 2518
rect 12360 2446 12388 4558
rect 12452 2564 12480 4966
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12544 3602 12572 4150
rect 12636 3670 12664 9522
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12820 7410 12848 7754
rect 12912 7410 12940 8570
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13004 6798 13032 9646
rect 13280 8294 13308 12406
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 11898 13492 12174
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13464 11082 13492 11834
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12728 4214 12756 4966
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12728 3534 12756 3878
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12452 2536 12572 2564
rect 12544 2446 12572 2536
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12636 1306 12664 3402
rect 12820 2650 12848 5578
rect 12912 5302 12940 6734
rect 13004 6254 13032 6734
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 5914 13032 6190
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12912 4146 12940 5238
rect 13096 4690 13124 7142
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13188 6458 13216 6666
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5370 13492 6054
rect 13556 5710 13584 13790
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13326 13676 13670
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13740 12918 13768 13262
rect 13728 12912 13780 12918
rect 13648 12860 13728 12866
rect 13648 12854 13780 12860
rect 13648 12838 13768 12854
rect 13648 11694 13676 12838
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 11830 13768 12582
rect 13832 12102 13860 15506
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13924 12306 13952 15302
rect 14108 14822 14136 19638
rect 14200 19514 14228 20402
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14292 19854 14320 20334
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14482 14136 14758
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 14074 14136 14214
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13924 11558 13952 12242
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 14016 11218 14044 12038
rect 14108 11898 14136 12038
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11286 14136 11494
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14200 11098 14228 14282
rect 14292 14006 14320 19790
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14384 19281 14412 19382
rect 14476 19310 14504 25434
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14568 23798 14596 24142
rect 14660 23866 14688 24142
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14568 23594 14596 23734
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 15212 23322 15240 28154
rect 15304 26314 15332 28358
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15384 27396 15436 27402
rect 15384 27338 15436 27344
rect 15396 27130 15424 27338
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15384 27124 15436 27130
rect 15384 27066 15436 27072
rect 15488 26450 15516 27270
rect 15580 26586 15608 27950
rect 16040 27538 16068 29990
rect 16592 29850 16620 30534
rect 17236 30258 17264 30670
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 17224 30252 17276 30258
rect 17224 30194 17276 30200
rect 17408 30252 17460 30258
rect 17408 30194 17460 30200
rect 17420 29850 17448 30194
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 17408 29844 17460 29850
rect 17408 29786 17460 29792
rect 16028 27532 16080 27538
rect 16028 27474 16080 27480
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15568 26580 15620 26586
rect 15568 26522 15620 26528
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15580 26042 15608 26182
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 14556 20256 14608 20262
rect 14556 20198 14608 20204
rect 14568 19854 14596 20198
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19304 14516 19310
rect 14370 19272 14426 19281
rect 14464 19246 14516 19252
rect 14370 19207 14426 19216
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14752 17746 14780 18090
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14752 17542 14780 17682
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14476 13530 14504 14214
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14292 11898 14320 12718
rect 14752 12306 14780 17478
rect 15028 16572 15056 18022
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 15120 16794 15148 17070
rect 15212 16794 15240 17138
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15108 16584 15160 16590
rect 15028 16544 15108 16572
rect 15108 16526 15160 16532
rect 15304 14618 15332 25842
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 15396 23730 15424 24550
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15396 23254 15424 23462
rect 15580 23322 15608 24006
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15384 23248 15436 23254
rect 15384 23190 15436 23196
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15672 19446 15700 23054
rect 15856 22094 15884 27270
rect 15948 27130 15976 27270
rect 16592 27130 16620 29786
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 16132 26382 16160 26726
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16408 25838 16436 26862
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 16132 24410 16160 24686
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 16224 23526 16252 24278
rect 16408 24206 16436 25094
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16776 24138 16804 25230
rect 16868 24750 16896 29514
rect 17972 29306 18000 30602
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18156 29306 18184 29582
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18064 27674 18092 28494
rect 18248 28218 18276 30670
rect 19076 29850 19104 31758
rect 19156 31136 19208 31142
rect 19156 31078 19208 31084
rect 19168 30190 19196 31078
rect 19260 30938 19288 31758
rect 23940 31748 23992 31754
rect 23940 31690 23992 31696
rect 19340 31680 19392 31686
rect 19340 31622 19392 31628
rect 20352 31680 20404 31686
rect 20352 31622 20404 31628
rect 23664 31680 23716 31686
rect 23664 31622 23716 31628
rect 19352 31482 19380 31622
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 20364 31482 20392 31622
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 20352 31476 20404 31482
rect 20352 31418 20404 31424
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 19984 31272 20036 31278
rect 19984 31214 20036 31220
rect 19616 31136 19668 31142
rect 19616 31078 19668 31084
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19260 30394 19288 30874
rect 19628 30802 19656 31078
rect 19616 30796 19668 30802
rect 19616 30738 19668 30744
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19352 30394 19380 30534
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19352 30190 19380 30330
rect 19444 30274 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19444 30258 19840 30274
rect 19444 30252 19852 30258
rect 19444 30246 19800 30252
rect 19800 30194 19852 30200
rect 19156 30184 19208 30190
rect 19156 30126 19208 30132
rect 19340 30184 19392 30190
rect 19340 30126 19392 30132
rect 19616 30184 19668 30190
rect 19616 30126 19668 30132
rect 19628 30054 19656 30126
rect 19616 30048 19668 30054
rect 19444 29996 19616 30002
rect 19444 29990 19668 29996
rect 19708 30048 19760 30054
rect 19708 29990 19760 29996
rect 19444 29974 19656 29990
rect 19064 29844 19116 29850
rect 19064 29786 19116 29792
rect 18880 29708 18932 29714
rect 18880 29650 18932 29656
rect 18892 29578 18920 29650
rect 18880 29572 18932 29578
rect 18880 29514 18932 29520
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 18340 29306 18368 29446
rect 19352 29306 19380 29446
rect 19444 29306 19472 29974
rect 19720 29866 19748 29990
rect 19628 29838 19748 29866
rect 19628 29646 19656 29838
rect 19616 29640 19668 29646
rect 19616 29582 19668 29588
rect 19812 29578 19840 30194
rect 19800 29572 19852 29578
rect 19800 29514 19852 29520
rect 19996 29510 20024 31214
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 20548 30734 20576 31078
rect 21928 30802 21956 31078
rect 21916 30796 21968 30802
rect 21916 30738 21968 30744
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20720 30592 20772 30598
rect 20720 30534 20772 30540
rect 20732 29714 20760 30534
rect 22296 30394 22324 31282
rect 22468 30728 22520 30734
rect 22468 30670 22520 30676
rect 22284 30388 22336 30394
rect 22284 30330 22336 30336
rect 21088 30116 21140 30122
rect 21088 30058 21140 30064
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19352 28506 19380 29242
rect 19260 28478 19380 28506
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18972 28416 19024 28422
rect 18972 28358 19024 28364
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17696 26790 17724 27270
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17512 26382 17540 26522
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16776 23866 16804 24074
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 15856 22066 15976 22094
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 20602 15884 21422
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19854 15884 20198
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15856 19174 15884 19790
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15672 17882 15700 18158
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15488 17270 15516 17478
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15396 15706 15424 17138
rect 15856 16250 15884 18022
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15706 15792 15846
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15488 15162 15516 15370
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14936 12434 14964 13874
rect 14936 12406 15056 12434
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 14016 11070 14228 11098
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 13832 10588 13860 11018
rect 13912 10600 13964 10606
rect 13832 10560 13912 10588
rect 13912 10542 13964 10548
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13740 8090 13768 8366
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13832 7410 13860 7958
rect 13924 7478 13952 7958
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 7002 13768 7278
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13832 6866 13860 7346
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 5914 13768 6598
rect 13924 6322 13952 7142
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13188 5166 13216 5306
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13464 4826 13492 5306
rect 13452 4820 13504 4826
rect 13188 4780 13452 4808
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13188 4570 13216 4780
rect 13452 4762 13504 4768
rect 13096 4542 13216 4570
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12912 2922 12940 3538
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 13096 2650 13124 4542
rect 13648 4146 13676 5782
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 12452 1278 12664 1306
rect 12452 800 12480 1278
rect 13004 1170 13032 2450
rect 12820 1142 13032 1170
rect 12820 800 12848 1142
rect 13188 800 13216 2790
rect 13556 800 13584 3946
rect 13740 3058 13768 5510
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13924 3670 13952 3878
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14016 3466 14044 11070
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10606 14136 10950
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 10266 14228 10542
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14292 10062 14320 11086
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14384 7546 14412 8502
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14476 7818 14504 8366
rect 14752 8090 14780 12242
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14936 11354 14964 11630
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14936 10266 14964 10406
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14476 7002 14504 7278
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14108 6458 14136 6598
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14372 5228 14424 5234
rect 14292 5188 14372 5216
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4282 14228 5102
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 13820 3392 13872 3398
rect 14188 3392 14240 3398
rect 13820 3334 13872 3340
rect 14186 3360 14188 3369
rect 14240 3360 14242 3369
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13832 2854 13860 3334
rect 14186 3295 14242 3304
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14200 2990 14228 3130
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14108 2774 14136 2926
rect 13924 2746 14136 2774
rect 13924 800 13952 2746
rect 14292 800 14320 5188
rect 14372 5170 14424 5176
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14384 2650 14412 4082
rect 14476 3058 14504 6598
rect 14568 5914 14596 7414
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14660 5710 14688 6326
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14740 5296 14792 5302
rect 14740 5238 14792 5244
rect 14752 4758 14780 5238
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14752 4214 14780 4558
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 4282 14964 4422
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14830 4040 14886 4049
rect 14830 3975 14886 3984
rect 14844 3942 14872 3975
rect 14832 3936 14884 3942
rect 15028 3913 15056 12406
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15304 11558 15332 12038
rect 15396 11762 15424 12038
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15120 10674 15148 11290
rect 15396 11082 15424 11698
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15396 10606 15424 11018
rect 15580 10606 15608 14418
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15384 10600 15436 10606
rect 15568 10600 15620 10606
rect 15436 10548 15516 10554
rect 15384 10542 15516 10548
rect 15568 10542 15620 10548
rect 15396 10526 15516 10542
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15120 9450 15148 9998
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15120 8498 15148 9386
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15396 8498 15424 8774
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15120 7546 15148 7958
rect 15488 7546 15516 10526
rect 15580 9926 15608 10542
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15396 6662 15424 7346
rect 15672 6866 15700 12854
rect 15764 12442 15792 13262
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15856 11082 15884 12582
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15856 10266 15884 11018
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 9058 15976 22066
rect 16224 20874 16252 23462
rect 16316 23322 16344 23734
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16316 22642 16344 23258
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16868 22234 16896 24686
rect 17040 24064 17092 24070
rect 17040 24006 17092 24012
rect 17052 23662 17080 24006
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 17144 21434 17172 25638
rect 17316 24404 17368 24410
rect 17512 24392 17540 26318
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17972 26042 18000 26250
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 18064 25378 18092 27066
rect 18156 25838 18184 27950
rect 18248 27130 18276 28154
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18248 26382 18276 27066
rect 18524 26994 18552 28358
rect 18984 28014 19012 28358
rect 19260 28098 19288 28478
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19352 28218 19380 28358
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19260 28082 19380 28098
rect 19260 28076 19392 28082
rect 19260 28070 19340 28076
rect 19340 28018 19392 28024
rect 18972 28008 19024 28014
rect 18972 27950 19024 27956
rect 19352 27334 19380 28018
rect 19444 27674 19472 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 18972 27328 19024 27334
rect 18972 27270 19024 27276
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18880 26852 18932 26858
rect 18880 26794 18932 26800
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18064 25350 18184 25378
rect 18052 25288 18104 25294
rect 18052 25230 18104 25236
rect 18064 24682 18092 25230
rect 18052 24676 18104 24682
rect 18052 24618 18104 24624
rect 17368 24364 17540 24392
rect 17316 24346 17368 24352
rect 17512 23594 17540 24364
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23730 17908 24006
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17972 23322 18000 24142
rect 18064 23866 18092 24618
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 18156 23746 18184 25350
rect 18248 24818 18276 26318
rect 18892 26314 18920 26794
rect 18880 26308 18932 26314
rect 18880 26250 18932 26256
rect 18984 25906 19012 27270
rect 19444 27130 19472 27610
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 20088 26926 20116 29514
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 27470 20760 27814
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 21100 27130 21128 30058
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21284 26926 21312 27338
rect 21376 27130 21404 27406
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 19708 26920 19760 26926
rect 19444 26880 19708 26908
rect 19340 26852 19392 26858
rect 19340 26794 19392 26800
rect 19352 26586 19380 26794
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19444 26450 19472 26880
rect 19708 26862 19760 26868
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18708 25498 18736 25842
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 18696 25492 18748 25498
rect 18696 25434 18748 25440
rect 18984 25430 19012 25706
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18524 23866 18552 24210
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18064 23730 18368 23746
rect 18052 23724 18368 23730
rect 18104 23718 18368 23724
rect 18052 23666 18104 23672
rect 18236 23656 18288 23662
rect 18236 23598 18288 23604
rect 17960 23316 18012 23322
rect 18012 23276 18092 23304
rect 17960 23258 18012 23264
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17880 22778 17908 23122
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17696 22234 17724 22578
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17236 21554 17264 21830
rect 17972 21554 18000 22918
rect 18064 22234 18092 23276
rect 18248 22778 18276 23598
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17868 21480 17920 21486
rect 17144 21418 17264 21434
rect 17868 21422 17920 21428
rect 17144 21412 17276 21418
rect 17144 21406 17224 21412
rect 17224 21354 17276 21360
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 21146 16804 21286
rect 17880 21146 17908 21422
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16132 20534 16160 20742
rect 16500 20534 16528 20742
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 17144 20466 17172 21082
rect 18064 20806 18092 22170
rect 18156 22098 18184 22374
rect 18144 22092 18196 22098
rect 18340 22094 18368 23718
rect 18524 22982 18552 23802
rect 18616 23322 18644 24142
rect 18708 23866 18736 25094
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18892 23866 18920 24686
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18708 23254 18736 23598
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 18984 22094 19012 25366
rect 19444 25362 19472 26386
rect 20260 26240 20312 26246
rect 20260 26182 20312 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20272 25906 20300 26182
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20260 25764 20312 25770
rect 20260 25706 20312 25712
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 18340 22066 18460 22094
rect 18144 22034 18196 22040
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18248 20806 18276 21422
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18340 21146 18368 21354
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18248 20602 18276 20742
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18156 20466 18184 20538
rect 17132 20460 17184 20466
rect 18052 20460 18104 20466
rect 17132 20402 17184 20408
rect 17972 20420 18052 20448
rect 17972 20058 18000 20420
rect 18052 20402 18104 20408
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16040 17678 16068 19110
rect 16500 18970 16528 19722
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16960 18834 16988 19110
rect 17420 18970 17448 19246
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 17604 18630 17632 19246
rect 17972 18834 18000 19994
rect 18064 19718 18092 20198
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19378 18092 19654
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 16040 16658 16068 17614
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16224 16794 16252 17070
rect 16500 17066 16528 18158
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16794 16344 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16592 16250 16620 17478
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 12434 16252 15982
rect 16684 15570 16712 16934
rect 17236 16590 17264 18022
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17307 17196 17359 17202
rect 17307 17138 17359 17144
rect 17328 16794 17356 17138
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15026 16528 15302
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16316 13870 16344 14350
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16500 13530 16528 14282
rect 16684 14074 16712 14758
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16132 12406 16252 12434
rect 16132 11268 16160 12406
rect 16212 11824 16264 11830
rect 16316 11812 16344 13262
rect 16684 12306 16712 13806
rect 16776 12782 16804 15982
rect 16960 15570 16988 16118
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17052 15570 17080 15642
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 15162 16896 15302
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 17052 14822 17080 15506
rect 17328 15450 17356 16730
rect 17512 16590 17540 17546
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17604 16522 17632 18566
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17788 17882 17816 18158
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17880 17066 17908 18022
rect 18156 17898 18184 20198
rect 18248 19378 18276 20538
rect 18328 20460 18380 20466
rect 18432 20448 18460 22066
rect 18800 22066 19012 22094
rect 18800 21894 18828 22066
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 21010 18828 21830
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18380 20420 18460 20448
rect 18328 20402 18380 20408
rect 18340 20262 18368 20402
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18616 19922 18644 20878
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18708 19514 18736 20742
rect 18800 19854 18828 20946
rect 19168 20602 19196 21422
rect 19352 21010 19380 23462
rect 19628 23118 19656 23462
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20168 22432 20220 22438
rect 19996 22392 20168 22420
rect 19996 22030 20024 22392
rect 20168 22374 20220 22380
rect 20272 22094 20300 25706
rect 20180 22066 20300 22094
rect 19984 22024 20036 22030
rect 19984 21966 20036 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19248 20800 19300 20806
rect 19246 20768 19248 20777
rect 19340 20800 19392 20806
rect 19300 20768 19302 20777
rect 19340 20742 19392 20748
rect 19246 20703 19302 20712
rect 19352 20602 19380 20742
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18984 20058 19012 20334
rect 18972 20052 19024 20058
rect 18892 20012 18972 20040
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18892 19378 18920 20012
rect 18972 19994 19024 20000
rect 19444 19922 19472 21014
rect 19904 21010 19932 21286
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 21490
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18064 17870 18184 17898
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 17144 15422 17356 15450
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16264 11784 16344 11812
rect 16212 11766 16264 11772
rect 16684 11762 16712 12242
rect 16868 12238 16896 12582
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 17144 11898 17172 15422
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17328 13682 17356 15302
rect 17420 15162 17448 15302
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17406 14920 17462 14929
rect 17406 14855 17408 14864
rect 17460 14855 17462 14864
rect 17408 14826 17460 14832
rect 17420 14414 17448 14826
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17236 13654 17356 13682
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16212 11280 16264 11286
rect 16132 11240 16212 11268
rect 16212 11222 16264 11228
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 9722 16068 10474
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15856 9030 15976 9058
rect 16224 9042 16252 11222
rect 16212 9036 16264 9042
rect 15660 6860 15712 6866
rect 15580 6820 15660 6848
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15120 5778 15148 6054
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15212 5302 15240 6054
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14832 3878 14884 3884
rect 15014 3904 15070 3913
rect 15014 3839 15070 3848
rect 14924 3528 14976 3534
rect 14646 3496 14702 3505
rect 14556 3460 14608 3466
rect 14924 3470 14976 3476
rect 14646 3431 14648 3440
rect 14556 3402 14608 3408
rect 14700 3431 14702 3440
rect 14648 3402 14700 3408
rect 14568 3194 14596 3402
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14936 2774 14964 3470
rect 15120 3398 15148 4014
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14660 2746 14964 2774
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14660 800 14688 2746
rect 15028 800 15056 2926
rect 15304 2446 15332 6054
rect 15396 5710 15424 6394
rect 15488 6322 15516 6666
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 4554 15424 5510
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15396 800 15424 4150
rect 15488 3058 15516 5578
rect 15580 4078 15608 6820
rect 15660 6802 15712 6808
rect 15856 6458 15884 9030
rect 16212 8978 16264 8984
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8090 15976 8910
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 16132 7886 16160 8774
rect 16224 7954 16252 8978
rect 16592 8634 16620 11290
rect 16684 11218 16712 11698
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16684 10674 16712 11154
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16684 10130 16712 10610
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16684 9450 16712 10066
rect 16776 9654 16804 11494
rect 17144 11354 17172 11834
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16684 9042 16712 9386
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16684 8498 16712 8978
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16224 7834 16252 7890
rect 16224 7806 16344 7834
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 6662 16252 7686
rect 16316 7002 16344 7806
rect 16684 7410 16712 8434
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16776 7002 16804 7346
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15856 5914 15884 6190
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16224 5710 16252 6598
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 15752 5704 15804 5710
rect 16212 5704 16264 5710
rect 15752 5646 15804 5652
rect 16132 5652 16212 5658
rect 16132 5646 16264 5652
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 4146 15700 5510
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15764 4010 15792 5646
rect 16132 5630 16252 5646
rect 16132 4146 16160 5630
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16224 4593 16252 5510
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16592 4622 16620 5102
rect 16580 4616 16632 4622
rect 16210 4584 16266 4593
rect 16580 4558 16632 4564
rect 16210 4519 16266 4528
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4146 16252 4422
rect 16592 4146 16620 4558
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 16592 3466 16620 4082
rect 16684 3466 16712 6054
rect 16868 5778 16896 9862
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8294 16988 8910
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 16960 7954 16988 8230
rect 17144 8022 17172 8230
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 6866 16988 7686
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17236 6730 17264 13654
rect 17512 13326 17540 15574
rect 17604 14498 17632 16458
rect 17880 15314 17908 17002
rect 17788 15286 17908 15314
rect 17788 14929 17816 15286
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 15008 18000 15098
rect 18064 15026 18092 17870
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 18156 17202 18184 17750
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16114 18184 17138
rect 18248 16674 18276 19314
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17270 18644 17546
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18340 16794 18368 17138
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18248 16646 18368 16674
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18052 15020 18104 15026
rect 17972 14980 18052 15008
rect 17868 14952 17920 14958
rect 17774 14920 17830 14929
rect 17868 14894 17920 14900
rect 17774 14855 17830 14864
rect 17604 14470 17724 14498
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17500 13320 17552 13326
rect 17328 13268 17500 13274
rect 17328 13262 17552 13268
rect 17328 13246 17540 13262
rect 17328 8956 17356 13246
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12102 17540 12786
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17512 11898 17540 12038
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17420 11762 17448 11834
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17512 11150 17540 11834
rect 17604 11558 17632 14350
rect 17696 13394 17724 14470
rect 17880 14074 17908 14894
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17696 12986 17724 13330
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17604 10810 17632 11494
rect 17592 10804 17644 10810
rect 17644 10764 17816 10792
rect 17592 10746 17644 10752
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17696 9722 17724 9930
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17500 8968 17552 8974
rect 17328 8928 17500 8956
rect 17500 8910 17552 8916
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17696 7886 17724 8570
rect 17788 8294 17816 10764
rect 17972 9674 18000 14980
rect 18052 14962 18104 14968
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18156 14074 18184 14554
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18340 12918 18368 16646
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18708 16250 18736 16526
rect 18892 16250 18920 19314
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 18290 20116 18566
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18432 15570 18460 16118
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18432 13870 18460 15302
rect 18512 14952 18564 14958
rect 18604 14952 18656 14958
rect 18512 14894 18564 14900
rect 18602 14920 18604 14929
rect 18656 14920 18658 14929
rect 18524 14278 18552 14894
rect 18602 14855 18658 14864
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18524 13394 18552 14214
rect 18800 14074 18828 14282
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18248 12442 18276 12854
rect 18236 12436 18288 12442
rect 18984 12434 19012 17478
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19260 14618 19288 14894
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19352 13938 19380 15302
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 18984 12406 19288 12434
rect 18236 12378 18288 12384
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18616 11898 18644 12310
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 19260 11694 19288 12406
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 18064 10266 18092 11630
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10266 18184 10950
rect 18432 10810 18460 11630
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 17880 9646 18000 9674
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17696 6662 17724 7482
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17222 6352 17278 6361
rect 17278 6310 17356 6338
rect 17222 6287 17278 6296
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16776 3126 16804 4218
rect 16960 4146 16988 6054
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3738 16896 3878
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 16592 2650 16620 3062
rect 17052 3058 17080 4966
rect 17144 4672 17172 5510
rect 17224 4684 17276 4690
rect 17144 4644 17224 4672
rect 17224 4626 17276 4632
rect 17328 4570 17356 6310
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17604 5914 17632 6190
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17512 4622 17540 4762
rect 17236 4542 17356 4570
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17236 3602 17264 4542
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17328 3534 17356 4082
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17420 3466 17448 4558
rect 17696 3602 17724 6054
rect 17788 4690 17816 8230
rect 17880 7018 17908 9646
rect 18616 9586 18644 10950
rect 18708 10674 18736 11494
rect 19260 11082 19288 11630
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17972 7206 18000 7822
rect 18064 7478 18092 8842
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8090 18276 8774
rect 18432 8634 18460 9318
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18156 7834 18184 8026
rect 18340 7954 18368 8230
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18156 7806 18368 7834
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17880 6990 18000 7018
rect 18156 7002 18184 7686
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17880 5166 17908 5646
rect 17972 5574 18000 6990
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18248 5370 18276 6190
rect 18340 5896 18368 7806
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 6866 18460 7686
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18340 5868 18460 5896
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 17960 5364 18012 5370
rect 18236 5364 18288 5370
rect 18012 5324 18092 5352
rect 17960 5306 18012 5312
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17880 3534 17908 5102
rect 17972 3738 18000 5170
rect 18064 5030 18092 5324
rect 18236 5306 18288 5312
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4078 18092 4966
rect 18248 4554 18276 5306
rect 18340 4690 18368 5646
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18340 4282 18368 4626
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18432 4146 18460 5868
rect 18524 5370 18552 9386
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 7546 18644 8230
rect 18708 7954 18736 8366
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18708 6866 18736 7142
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18602 6352 18658 6361
rect 18602 6287 18658 6296
rect 18616 6254 18644 6287
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18800 5114 18828 8842
rect 18892 7342 18920 11018
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 7546 19012 9454
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 18972 5228 19024 5234
rect 19024 5188 19196 5216
rect 18972 5170 19024 5176
rect 18616 5086 18828 5114
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 4282 18552 4422
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15764 800 15792 2314
rect 16132 800 16160 2314
rect 16488 1556 16540 1562
rect 16488 1498 16540 1504
rect 16500 800 16528 1498
rect 16868 800 16896 2382
rect 17236 800 17264 2926
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 11808 734 12020 762
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17328 762 17356 2450
rect 17512 870 17632 898
rect 17512 762 17540 870
rect 17604 800 17632 870
rect 17972 800 18000 3402
rect 18524 2650 18552 4082
rect 18616 4049 18644 5086
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18708 4282 18736 4558
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18602 4040 18658 4049
rect 18602 3975 18658 3984
rect 18800 3194 18828 4966
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 18892 3074 18920 4422
rect 18984 4214 19012 4422
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 18970 4040 19026 4049
rect 18970 3975 19026 3984
rect 18984 3534 19012 3975
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19076 3194 19104 3334
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18800 3046 18920 3074
rect 18800 2774 18828 3046
rect 18880 2984 18932 2990
rect 18932 2944 19104 2972
rect 18880 2926 18932 2932
rect 18800 2746 18920 2774
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18340 800 18368 2450
rect 18892 2446 18920 2746
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 18708 800 18736 2314
rect 19076 800 19104 2944
rect 19168 2650 19196 5188
rect 19260 5166 19288 6326
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19260 4690 19288 5102
rect 19352 4826 19380 12786
rect 19444 9178 19472 17546
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 20180 16794 20208 22066
rect 20258 21040 20314 21049
rect 20258 20975 20260 20984
rect 20312 20975 20314 20984
rect 20260 20946 20312 20952
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19536 14482 19564 15098
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19720 14482 19748 14758
rect 19996 14618 20024 15438
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 20088 15162 20116 15370
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 20088 14074 20116 14554
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 14074 20208 14214
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 8090 19656 8366
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19536 6798 19564 7278
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19430 6216 19486 6225
rect 19430 6151 19432 6160
rect 19484 6151 19486 6160
rect 19432 6122 19484 6128
rect 20272 5846 20300 20946
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 15026 20484 15302
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20640 12434 20668 26726
rect 21928 26382 21956 27270
rect 22112 26586 22140 27406
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 27130 22324 27270
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22388 26926 22416 27814
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21916 26376 21968 26382
rect 21916 26318 21968 26324
rect 21284 26042 21312 26318
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 22480 24818 22508 30670
rect 23572 30660 23624 30666
rect 23572 30602 23624 30608
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22756 29850 22784 30126
rect 23584 29850 23612 30602
rect 23676 30598 23704 31622
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23664 30592 23716 30598
rect 23664 30534 23716 30540
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 23676 29578 23704 30534
rect 23768 30258 23796 30874
rect 23860 30258 23888 31418
rect 23952 30938 23980 31690
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 24412 30734 24440 31622
rect 24596 30938 24624 32302
rect 25412 32224 25464 32230
rect 25412 32166 25464 32172
rect 26608 32224 26660 32230
rect 26608 32166 26660 32172
rect 27068 32224 27120 32230
rect 27068 32166 27120 32172
rect 27528 32224 27580 32230
rect 27528 32166 27580 32172
rect 28264 32224 28316 32230
rect 28264 32166 28316 32172
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24780 31346 24808 31826
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25136 31680 25188 31686
rect 25136 31622 25188 31628
rect 25148 31414 25176 31622
rect 25136 31408 25188 31414
rect 25136 31350 25188 31356
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24124 30592 24176 30598
rect 24124 30534 24176 30540
rect 23756 30252 23808 30258
rect 23756 30194 23808 30200
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23664 29572 23716 29578
rect 23664 29514 23716 29520
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22744 28212 22796 28218
rect 22744 28154 22796 28160
rect 22756 26994 22784 28154
rect 22848 27470 22876 28358
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 22836 27464 22888 27470
rect 22836 27406 22888 27412
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22560 25696 22612 25702
rect 22664 25684 22692 26862
rect 23124 25974 23152 27610
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23308 26926 23336 27406
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23296 26920 23348 26926
rect 23296 26862 23348 26868
rect 23400 26858 23428 27270
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 23204 26580 23256 26586
rect 23204 26522 23256 26528
rect 23112 25968 23164 25974
rect 23112 25910 23164 25916
rect 23216 25838 23244 26522
rect 23400 26450 23428 26794
rect 23492 26586 23520 27814
rect 23584 26586 23612 28494
rect 23676 28150 23704 28494
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23664 28144 23716 28150
rect 23664 28086 23716 28092
rect 23768 27538 23796 28358
rect 23860 27538 23888 29990
rect 24136 29714 24164 30534
rect 24596 30394 24624 30874
rect 24584 30388 24636 30394
rect 24584 30330 24636 30336
rect 24584 30048 24636 30054
rect 24584 29990 24636 29996
rect 23940 29708 23992 29714
rect 23940 29650 23992 29656
rect 24124 29708 24176 29714
rect 24124 29650 24176 29656
rect 23952 29034 23980 29650
rect 24124 29504 24176 29510
rect 24124 29446 24176 29452
rect 23940 29028 23992 29034
rect 23940 28970 23992 28976
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23664 26920 23716 26926
rect 23664 26862 23716 26868
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23572 26580 23624 26586
rect 23572 26522 23624 26528
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23676 26382 23704 26862
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 22612 25656 22692 25684
rect 22560 25638 22612 25644
rect 22664 25362 22692 25656
rect 23768 25498 23796 27270
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23860 26586 23888 26726
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23952 25362 23980 28970
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 24044 27674 24072 27814
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 24032 26920 24084 26926
rect 24032 26862 24084 26868
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 23940 25356 23992 25362
rect 23940 25298 23992 25304
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22480 23866 22508 24754
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 21622 20760 22918
rect 21284 22778 21312 23054
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22778 21956 22918
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 21376 22574 21404 22714
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 21690 21220 21830
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 20942 20944 21286
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20732 17270 20760 18634
rect 20824 18290 20852 19654
rect 21284 19514 21312 19790
rect 21376 19718 21404 22510
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21836 22030 21864 22170
rect 22112 22030 22140 23054
rect 22204 22438 22232 23802
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22480 23186 22508 23462
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22388 22710 22416 22918
rect 22480 22778 22508 22918
rect 22468 22772 22520 22778
rect 22468 22714 22520 22720
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22192 22432 22244 22438
rect 22244 22380 22324 22386
rect 22192 22374 22324 22380
rect 22204 22358 22324 22374
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22112 21894 22140 21966
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21376 19378 21404 19654
rect 21560 19378 21588 20878
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21928 20602 21956 20810
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21732 19712 21784 19718
rect 21732 19654 21784 19660
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20916 17882 20944 18294
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 21376 17610 21404 19314
rect 21560 18834 21588 19314
rect 21744 19310 21772 19654
rect 22204 19514 22232 19654
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22112 18358 22140 18702
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 21468 17270 21496 17478
rect 21928 17270 21956 17478
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 21456 17264 21508 17270
rect 21456 17206 21508 17212
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 14550 20760 14962
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20548 12406 20668 12434
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11898 20484 12038
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20260 5840 20312 5846
rect 20260 5782 20312 5788
rect 19616 5704 19668 5710
rect 19614 5672 19616 5681
rect 20168 5704 20220 5710
rect 19668 5672 19670 5681
rect 20168 5646 20220 5652
rect 19614 5607 19670 5616
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19260 4146 19288 4626
rect 19720 4622 19748 4966
rect 20180 4622 20208 5646
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20272 4826 20300 5102
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19260 3738 19288 4082
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19352 2938 19380 3878
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19260 2910 19380 2938
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19260 2514 19288 2910
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19352 1442 19380 2790
rect 19444 2446 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3194 20024 4490
rect 20180 4282 20208 4558
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20548 4162 20576 12406
rect 20732 12306 20760 13806
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20916 11898 20944 12718
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21192 9722 21220 11290
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21284 9674 21312 16458
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 15026 21680 15438
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21928 15162 21956 15370
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21732 13864 21784 13870
rect 21732 13806 21784 13812
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21560 12434 21588 12582
rect 21560 12406 21680 12434
rect 21652 12238 21680 12406
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21744 11694 21772 13806
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21824 12232 21876 12238
rect 21928 12220 21956 12786
rect 21876 12192 21956 12220
rect 21824 12174 21876 12180
rect 21836 11694 21864 12174
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21744 11354 21772 11630
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 22020 11150 22048 17478
rect 22296 15042 22324 22358
rect 22572 22166 22600 22510
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22572 21842 22600 22102
rect 22756 22098 22784 23122
rect 23400 23118 23428 23598
rect 23768 23526 23796 24686
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23860 23866 23888 24550
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22388 21814 22600 21842
rect 22388 21690 22416 21814
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22388 18766 22416 18906
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22388 17202 22416 18702
rect 22480 17746 22508 21558
rect 22572 20942 22600 21626
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22560 19848 22612 19854
rect 22558 19816 22560 19825
rect 22612 19816 22614 19825
rect 22558 19751 22614 19760
rect 22664 19446 22692 20198
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22756 19334 22784 22034
rect 22848 20874 22876 22374
rect 23020 22160 23072 22166
rect 23020 22102 23072 22108
rect 23032 21978 23060 22102
rect 23308 22098 23336 22986
rect 23400 22642 23428 23054
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 22940 21950 23060 21978
rect 23204 21956 23256 21962
rect 22940 21026 22968 21950
rect 23204 21898 23256 21904
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23032 21146 23060 21830
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 22940 20998 23060 21026
rect 22836 20868 22888 20874
rect 22836 20810 22888 20816
rect 22928 20324 22980 20330
rect 22928 20266 22980 20272
rect 22940 19922 22968 20266
rect 22928 19916 22980 19922
rect 22928 19858 22980 19864
rect 22756 19306 22968 19334
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22572 18850 22600 19110
rect 22848 18902 22876 19110
rect 22836 18896 22888 18902
rect 22572 18822 22784 18850
rect 22836 18838 22888 18844
rect 22756 18630 22784 18822
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22664 17610 22692 18566
rect 22848 18358 22876 18838
rect 22940 18766 22968 19306
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16658 22600 16934
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22756 15042 22784 17478
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22204 15014 22324 15042
rect 22388 15014 22784 15042
rect 22204 14006 22232 15014
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14278 22324 14894
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22296 13394 22324 14214
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22100 13320 22152 13326
rect 22152 13280 22232 13308
rect 22100 13262 22152 13268
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 12918 22140 13126
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22204 10810 22232 13280
rect 22388 12434 22416 15014
rect 22744 14952 22796 14958
rect 22848 14906 22876 15506
rect 22796 14900 22876 14906
rect 22744 14894 22876 14900
rect 22652 14884 22704 14890
rect 22652 14826 22704 14832
rect 22756 14878 22876 14894
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22388 12406 22508 12434
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22296 11286 22324 11834
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22388 10742 22416 11766
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 22480 10690 22508 12406
rect 22572 12306 22600 12582
rect 22664 12322 22692 14826
rect 22756 14278 22784 14878
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 23032 13308 23060 20998
rect 23124 20466 23152 21830
rect 23216 21078 23244 21898
rect 23400 21690 23428 22578
rect 23492 22506 23520 22918
rect 23480 22500 23532 22506
rect 23480 22442 23532 22448
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23308 20058 23336 20334
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23124 19825 23152 19858
rect 23110 19816 23166 19825
rect 23110 19751 23166 19760
rect 23216 19718 23244 19994
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23308 19310 23336 19790
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23308 18970 23336 19246
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23308 18290 23336 18702
rect 23400 18358 23428 20198
rect 23492 19922 23520 21830
rect 23584 21146 23612 21830
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23676 18426 23704 18906
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23216 16114 23244 18158
rect 23676 17746 23704 18362
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23308 16250 23336 16934
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23400 16130 23428 17070
rect 23768 16538 23796 23462
rect 23952 22982 23980 25298
rect 24044 24410 24072 26862
rect 24136 24682 24164 29446
rect 24596 29034 24624 29990
rect 24688 29714 24716 31214
rect 24860 31204 24912 31210
rect 24860 31146 24912 31152
rect 24872 30258 24900 31146
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24964 30734 24992 31078
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24964 30394 24992 30670
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 25240 29850 25268 31758
rect 25424 30666 25452 32166
rect 26620 31890 26648 32166
rect 27080 31890 27108 32166
rect 26608 31884 26660 31890
rect 26608 31826 26660 31832
rect 27068 31884 27120 31890
rect 27068 31826 27120 31832
rect 26332 31816 26384 31822
rect 26332 31758 26384 31764
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 25872 31136 25924 31142
rect 25872 31078 25924 31084
rect 25412 30660 25464 30666
rect 25412 30602 25464 30608
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 24676 29708 24728 29714
rect 24676 29650 24728 29656
rect 24768 29708 24820 29714
rect 24768 29650 24820 29656
rect 24780 29510 24808 29650
rect 25884 29646 25912 31078
rect 26160 30734 26188 31282
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26160 29714 26188 30670
rect 26344 30666 26372 31758
rect 26620 30938 26648 31826
rect 26608 30932 26660 30938
rect 26608 30874 26660 30880
rect 26332 30660 26384 30666
rect 26332 30602 26384 30608
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 26240 30116 26292 30122
rect 26240 30058 26292 30064
rect 26148 29708 26200 29714
rect 26148 29650 26200 29656
rect 25872 29640 25924 29646
rect 25872 29582 25924 29588
rect 26252 29510 26280 30058
rect 26436 29510 26464 30194
rect 27080 29782 27108 31826
rect 27540 31414 27568 32166
rect 28276 32026 28304 32166
rect 28460 32026 28488 32302
rect 28264 32020 28316 32026
rect 28264 31962 28316 31968
rect 28448 32020 28500 32026
rect 28448 31962 28500 31968
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28540 31680 28592 31686
rect 28540 31622 28592 31628
rect 28080 31476 28132 31482
rect 28080 31418 28132 31424
rect 27528 31408 27580 31414
rect 27528 31350 27580 31356
rect 27988 30932 28040 30938
rect 27988 30874 28040 30880
rect 28000 30258 28028 30874
rect 28092 30258 28120 31418
rect 28460 31346 28488 31622
rect 28448 31340 28500 31346
rect 28448 31282 28500 31288
rect 28552 30734 28580 31622
rect 28828 31482 28856 32302
rect 36360 32224 36412 32230
rect 36360 32166 36412 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 29184 31816 29236 31822
rect 29184 31758 29236 31764
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 29196 31482 29224 31758
rect 29276 31748 29328 31754
rect 29276 31690 29328 31696
rect 29288 31482 29316 31690
rect 29736 31680 29788 31686
rect 29736 31622 29788 31628
rect 28816 31476 28868 31482
rect 28816 31418 28868 31424
rect 29184 31476 29236 31482
rect 29184 31418 29236 31424
rect 29276 31476 29328 31482
rect 29276 31418 29328 31424
rect 29460 31340 29512 31346
rect 29460 31282 29512 31288
rect 28632 31272 28684 31278
rect 28632 31214 28684 31220
rect 28644 30938 28672 31214
rect 28632 30932 28684 30938
rect 28632 30874 28684 30880
rect 29000 30932 29052 30938
rect 29000 30874 29052 30880
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 27804 30252 27856 30258
rect 27804 30194 27856 30200
rect 27988 30252 28040 30258
rect 27988 30194 28040 30200
rect 28080 30252 28132 30258
rect 28080 30194 28132 30200
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 27068 29776 27120 29782
rect 27068 29718 27120 29724
rect 26976 29708 27028 29714
rect 26976 29650 27028 29656
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24492 28008 24544 28014
rect 24492 27950 24544 27956
rect 24504 27674 24532 27950
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24400 27328 24452 27334
rect 24400 27270 24452 27276
rect 24216 26444 24268 26450
rect 24216 26386 24268 26392
rect 24228 25498 24256 26386
rect 24412 26353 24440 27270
rect 24596 26994 24624 28970
rect 24676 27940 24728 27946
rect 24676 27882 24728 27888
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24688 26926 24716 27882
rect 24964 27334 24992 29446
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24780 27130 24808 27270
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24964 26926 24992 27270
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24398 26344 24454 26353
rect 24398 26279 24454 26288
rect 24964 26246 24992 26862
rect 25056 26858 25084 28494
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 26056 27872 26108 27878
rect 26056 27814 26108 27820
rect 25332 27130 25360 27814
rect 25688 27600 25740 27606
rect 25688 27542 25740 27548
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25320 27124 25372 27130
rect 25320 27066 25372 27072
rect 25044 26852 25096 26858
rect 25044 26794 25096 26800
rect 25424 26314 25452 27406
rect 25412 26308 25464 26314
rect 25412 26250 25464 26256
rect 24952 26240 25004 26246
rect 24952 26182 25004 26188
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24216 25492 24268 25498
rect 24216 25434 24268 25440
rect 24124 24676 24176 24682
rect 24124 24618 24176 24624
rect 24032 24404 24084 24410
rect 24032 24346 24084 24352
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 24044 22166 24072 24346
rect 24780 24206 24808 25638
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24032 22160 24084 22166
rect 24032 22102 24084 22108
rect 24044 21690 24072 22102
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24136 21894 24164 22034
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23952 20058 23980 20334
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 24032 18692 24084 18698
rect 24032 18634 24084 18640
rect 24044 18358 24072 18634
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 23860 16794 23888 17070
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23308 16102 23428 16130
rect 23492 16510 23796 16538
rect 23308 15910 23336 16102
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 23124 15162 23152 15302
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23216 14328 23244 15438
rect 23308 14958 23336 15846
rect 23400 15570 23428 15846
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23296 14340 23348 14346
rect 23216 14300 23296 14328
rect 23296 14282 23348 14288
rect 23308 13530 23336 14282
rect 23492 13802 23520 16510
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23584 15570 23612 16390
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23584 14090 23612 15506
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23768 15026 23796 15098
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23664 14952 23716 14958
rect 23860 14906 23888 15302
rect 23716 14900 23888 14906
rect 23664 14894 23888 14900
rect 23676 14878 23888 14894
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23768 14618 23796 14758
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23860 14482 23888 14878
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23584 14062 23704 14090
rect 23952 14074 23980 15302
rect 24228 14498 24256 22442
rect 24308 21684 24360 21690
rect 24308 21626 24360 21632
rect 24320 18970 24348 21626
rect 24872 21350 24900 25638
rect 24964 23746 24992 26182
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25240 24750 25268 25434
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 25056 23866 25084 24346
rect 25240 24154 25268 24686
rect 25148 24126 25268 24154
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 24964 23718 25084 23746
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24964 20874 24992 23462
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24596 18970 24624 19246
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24320 16998 24348 17682
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 24320 14618 24348 15438
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24136 14470 24256 14498
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 24044 14074 24072 14282
rect 23676 14006 23704 14062
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23204 13320 23256 13326
rect 23032 13280 23204 13308
rect 23020 12912 23072 12918
rect 23020 12854 23072 12860
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22664 12306 22784 12322
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22652 12300 22784 12306
rect 22704 12294 22784 12300
rect 22652 12242 22704 12248
rect 22572 11354 22600 12242
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22664 10810 22692 11766
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22480 10662 22692 10690
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 6866 20760 9522
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20916 7886 20944 8774
rect 21100 8566 21128 8910
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 21192 7954 21220 9658
rect 21284 9646 21864 9674
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21744 8430 21772 8774
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 21192 7546 21220 7890
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 20640 6458 20668 6598
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5642 20668 6054
rect 20824 5914 20852 6190
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 21284 5030 21312 6598
rect 21376 6322 21404 7686
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 20456 4146 20576 4162
rect 21376 4146 21404 6054
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 5302 21496 5510
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21652 5166 21680 6598
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21744 5710 21772 6190
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21836 5370 21864 9646
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22204 8634 22232 8774
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21928 7750 21956 8366
rect 22204 7886 22232 8570
rect 22388 8362 22416 8570
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 22204 7274 22232 7822
rect 22480 7410 22508 8774
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6866 22140 7142
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22020 6118 22048 6802
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21744 4622 21772 5102
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 20456 4140 20588 4146
rect 20456 4134 20536 4140
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 1442 20024 2994
rect 19352 1414 19472 1442
rect 19444 800 19472 1414
rect 19812 1414 20024 1442
rect 19812 800 19840 1414
rect 20088 1034 20116 3470
rect 20180 2774 20208 3878
rect 20272 3058 20300 4014
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20180 2746 20300 2774
rect 20272 2446 20300 2746
rect 20456 2650 20484 4134
rect 20536 4082 20588 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20548 3194 20576 3946
rect 22020 3738 22048 5170
rect 22100 3936 22152 3942
rect 22204 3924 22232 7210
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22664 6746 22692 10662
rect 22756 9178 22784 12294
rect 22848 12102 22876 12582
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22940 11558 22968 12174
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 23032 11150 23060 12854
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23020 10600 23072 10606
rect 23124 10554 23152 13280
rect 23204 13262 23256 13268
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23216 12102 23244 12786
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23216 11898 23244 12038
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23308 11694 23336 13466
rect 23584 12986 23612 13874
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23676 12434 23704 13942
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23860 13530 23888 13738
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23584 12406 23704 12434
rect 23584 11830 23612 12406
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 11150 23244 11494
rect 23308 11218 23336 11630
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23400 11014 23428 11698
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23492 10810 23520 11494
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23388 10736 23440 10742
rect 23584 10690 23612 11766
rect 23860 11694 23888 13466
rect 24136 12850 24164 14470
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24228 14006 24256 14214
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 24308 13796 24360 13802
rect 24308 13738 24360 13744
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23440 10684 23612 10690
rect 23388 10678 23612 10684
rect 23072 10548 23152 10554
rect 23020 10542 23152 10548
rect 23032 10526 23152 10542
rect 23400 10662 23612 10678
rect 23032 9926 23060 10526
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 23032 9518 23060 9862
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22756 8498 22784 8774
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 23032 7954 23060 9454
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23216 8906 23244 9318
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23204 8900 23256 8906
rect 23204 8842 23256 8848
rect 23204 8288 23256 8294
rect 23308 8276 23336 9114
rect 23256 8248 23336 8276
rect 23204 8230 23256 8236
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22940 6866 22968 7686
rect 23308 7002 23336 8248
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 22296 5302 22324 6734
rect 22664 6718 22784 6746
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22296 4826 22324 5238
rect 22388 5137 22416 6122
rect 22468 5296 22520 5302
rect 22468 5238 22520 5244
rect 22374 5128 22430 5137
rect 22374 5063 22430 5072
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22152 3896 22232 3924
rect 22100 3878 22152 3884
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22112 3534 22140 3878
rect 22388 3602 22416 5063
rect 22480 5030 22508 5238
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22756 3466 22784 6718
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23032 6458 23060 6598
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5302 23152 6394
rect 23308 5710 23336 6938
rect 23400 6390 23428 10662
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23492 7954 23520 8230
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23492 7002 23520 7754
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23572 6928 23624 6934
rect 23572 6870 23624 6876
rect 23584 6730 23612 6870
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22940 3738 22968 4558
rect 23124 4282 23152 4762
rect 23308 4758 23336 5646
rect 23492 5234 23520 5850
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23112 4276 23164 4282
rect 23032 4236 23112 4264
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23032 3534 23060 4236
rect 23112 4218 23164 4224
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 23124 3618 23152 4082
rect 23400 3942 23428 4626
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23124 3590 23244 3618
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22112 3194 22140 3334
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20732 1442 20760 2450
rect 20548 1414 20760 1442
rect 20088 1006 20208 1034
rect 20180 800 20208 1006
rect 20548 800 20576 1414
rect 20916 800 20944 2994
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 21100 2774 21128 2926
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21100 2746 21312 2774
rect 21284 800 21312 2746
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21652 870 21772 898
rect 21652 800 21680 870
rect 17328 734 17540 762
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 21744 762 21772 870
rect 21928 762 21956 2314
rect 22020 800 22048 2790
rect 22388 800 22416 3062
rect 22664 2650 22692 3334
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22756 800 22784 2926
rect 23124 800 23152 3470
rect 23216 3398 23244 3590
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23308 3058 23336 3878
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23400 2514 23428 3878
rect 23584 3505 23612 5510
rect 23676 4690 23704 8298
rect 23768 8090 23796 9454
rect 23860 8430 23888 10746
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23860 8090 23888 8366
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23768 7002 23796 7278
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23768 5710 23796 6598
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23768 4434 23796 5646
rect 23860 5166 23888 8026
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23860 4554 23888 5102
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23768 4406 23888 4434
rect 23860 4078 23888 4406
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23570 3496 23626 3505
rect 23570 3431 23626 3440
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23492 2446 23520 3334
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23584 1578 23612 3130
rect 23860 2774 23888 4014
rect 23952 3505 23980 11018
rect 24228 10810 24256 12242
rect 24216 10804 24268 10810
rect 24216 10746 24268 10752
rect 24216 7744 24268 7750
rect 24214 7712 24216 7721
rect 24268 7712 24270 7721
rect 24214 7647 24270 7656
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24136 5166 24164 6326
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24124 5160 24176 5166
rect 24124 5102 24176 5108
rect 24136 4826 24164 5102
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 24136 4282 24164 4422
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 24044 3738 24072 4150
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 23938 3496 23994 3505
rect 23938 3431 23994 3440
rect 24136 3058 24164 3878
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 23860 2746 23980 2774
rect 23952 2582 23980 2746
rect 23940 2576 23992 2582
rect 23940 2518 23992 2524
rect 24044 2446 24072 2790
rect 24228 2650 24256 5850
rect 24320 5710 24348 13738
rect 24412 12238 24440 14758
rect 24504 13784 24532 17546
rect 24596 17066 24624 18226
rect 24964 17882 24992 20810
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 24596 13802 24624 17002
rect 24964 16794 24992 17818
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 25056 16590 25084 23718
rect 25148 23526 25176 24126
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 25240 23730 25268 24006
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25240 22778 25268 23666
rect 25424 23526 25452 26250
rect 25700 26042 25728 27542
rect 26068 27402 26096 27814
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 26160 27130 26188 27950
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25700 24138 25728 25094
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25792 23730 25820 24686
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 25424 23322 25452 23462
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 25688 23180 25740 23186
rect 25688 23122 25740 23128
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25700 22234 25728 23122
rect 25780 22976 25832 22982
rect 25884 22964 25912 23598
rect 25832 22936 25912 22964
rect 25780 22918 25832 22924
rect 25688 22228 25740 22234
rect 25688 22170 25740 22176
rect 25700 21962 25728 22170
rect 25792 22098 25820 22918
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25688 21956 25740 21962
rect 25608 21916 25688 21944
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25148 19378 25176 19790
rect 25240 19514 25268 20198
rect 25504 19712 25556 19718
rect 25504 19654 25556 19660
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25148 18834 25176 19314
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 25424 18970 25452 19110
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25516 18766 25544 19654
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25608 18630 25636 21916
rect 25688 21898 25740 21904
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18222 25636 18566
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25700 17678 25728 20198
rect 25792 18426 25820 20334
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25884 20058 25912 20198
rect 25872 20052 25924 20058
rect 25872 19994 25924 20000
rect 25976 19718 26004 24210
rect 26068 23730 26096 26930
rect 26252 26314 26280 29446
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26436 25702 26464 29446
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26804 27130 26832 28358
rect 26988 28082 27016 29650
rect 27816 29034 27844 30194
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 27804 29028 27856 29034
rect 27804 28970 27856 28976
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 26988 27538 27016 28018
rect 27356 27674 27384 28494
rect 27344 27668 27396 27674
rect 27344 27610 27396 27616
rect 26976 27532 27028 27538
rect 26976 27474 27028 27480
rect 26792 27124 26844 27130
rect 26792 27066 26844 27072
rect 26988 26994 27016 27474
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 26976 26988 27028 26994
rect 26976 26930 27028 26936
rect 26516 26920 26568 26926
rect 26516 26862 26568 26868
rect 26528 26586 26556 26862
rect 26516 26580 26568 26586
rect 26568 26540 26648 26568
rect 26516 26522 26568 26528
rect 26424 25696 26476 25702
rect 26424 25638 26476 25644
rect 26424 25288 26476 25294
rect 26424 25230 26476 25236
rect 26240 24880 26292 24886
rect 26240 24822 26292 24828
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 26160 24410 26188 24686
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 26252 24070 26280 24822
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26344 24070 26372 24550
rect 26436 24410 26464 25230
rect 26516 24608 26568 24614
rect 26516 24550 26568 24556
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26528 24206 26556 24550
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 26252 23882 26280 24006
rect 26252 23866 26372 23882
rect 26252 23860 26384 23866
rect 26252 23854 26332 23860
rect 26056 23724 26108 23730
rect 26108 23684 26188 23712
rect 26056 23666 26108 23672
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 26068 22778 26096 22986
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 26160 22098 26188 23684
rect 26252 23186 26280 23854
rect 26332 23802 26384 23808
rect 26620 23322 26648 26540
rect 27080 26518 27108 27406
rect 27068 26512 27120 26518
rect 27068 26454 27120 26460
rect 27448 26042 27476 28494
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27540 28218 27568 28358
rect 28000 28218 28028 29990
rect 28828 29850 28856 30194
rect 29012 30190 29040 30874
rect 29472 30802 29500 31282
rect 29748 31142 29776 31622
rect 29920 31272 29972 31278
rect 29920 31214 29972 31220
rect 29736 31136 29788 31142
rect 29736 31078 29788 31084
rect 29932 30938 29960 31214
rect 31116 31136 31168 31142
rect 31116 31078 31168 31084
rect 29920 30932 29972 30938
rect 29920 30874 29972 30880
rect 29460 30796 29512 30802
rect 29460 30738 29512 30744
rect 29368 30592 29420 30598
rect 29368 30534 29420 30540
rect 29000 30184 29052 30190
rect 29000 30126 29052 30132
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29104 29850 29132 29990
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 29092 29844 29144 29850
rect 29092 29786 29144 29792
rect 28540 29028 28592 29034
rect 28540 28970 28592 28976
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 27712 27872 27764 27878
rect 27712 27814 27764 27820
rect 27724 27538 27752 27814
rect 27712 27532 27764 27538
rect 27712 27474 27764 27480
rect 27804 27532 27856 27538
rect 27804 27474 27856 27480
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 27436 26036 27488 26042
rect 27436 25978 27488 25984
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27632 24410 27660 25774
rect 27620 24404 27672 24410
rect 27620 24346 27672 24352
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27356 23866 27384 24006
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 27724 23662 27752 26726
rect 27816 26314 27844 27474
rect 28092 27470 28120 28018
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 28092 27130 28120 27406
rect 28080 27124 28132 27130
rect 28080 27066 28132 27072
rect 27804 26308 27856 26314
rect 27804 26250 27856 26256
rect 28276 26042 28304 28358
rect 28368 27946 28396 28494
rect 28356 27940 28408 27946
rect 28356 27882 28408 27888
rect 28552 27538 28580 28970
rect 28632 28416 28684 28422
rect 28632 28358 28684 28364
rect 28644 28014 28672 28358
rect 29000 28076 29052 28082
rect 29000 28018 29052 28024
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 28632 28008 28684 28014
rect 28632 27950 28684 27956
rect 28540 27532 28592 27538
rect 28540 27474 28592 27480
rect 28644 27334 28672 27950
rect 28724 27940 28776 27946
rect 28724 27882 28776 27888
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28264 26036 28316 26042
rect 28264 25978 28316 25984
rect 28448 26036 28500 26042
rect 28448 25978 28500 25984
rect 28460 25498 28488 25978
rect 28644 25974 28672 27270
rect 28736 27130 28764 27882
rect 29012 27674 29040 28018
rect 29000 27668 29052 27674
rect 29000 27610 29052 27616
rect 29196 27606 29224 28018
rect 29276 27872 29328 27878
rect 29276 27814 29328 27820
rect 29288 27713 29316 27814
rect 29274 27704 29330 27713
rect 29274 27639 29330 27648
rect 28908 27600 28960 27606
rect 28908 27542 28960 27548
rect 29184 27600 29236 27606
rect 29380 27554 29408 30534
rect 29184 27542 29236 27548
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28920 26926 28948 27542
rect 29000 27532 29052 27538
rect 29000 27474 29052 27480
rect 29288 27526 29408 27554
rect 28908 26920 28960 26926
rect 28908 26862 28960 26868
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 28632 25968 28684 25974
rect 28632 25910 28684 25916
rect 28448 25492 28500 25498
rect 28448 25434 28500 25440
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28368 23866 28396 24550
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28172 23792 28224 23798
rect 28172 23734 28224 23740
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 26976 23520 27028 23526
rect 26976 23462 27028 23468
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 26988 23186 27016 23462
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26332 23044 26384 23050
rect 26332 22986 26384 22992
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26252 22234 26280 22918
rect 26344 22778 26372 22986
rect 26608 22976 26660 22982
rect 26608 22918 26660 22924
rect 26620 22778 26648 22918
rect 27632 22778 27660 23530
rect 27724 23322 27752 23598
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26528 20602 26556 20742
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25976 19514 26004 19654
rect 26712 19514 26740 19858
rect 26988 19786 27016 20198
rect 27264 20058 27292 20878
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 26976 19780 27028 19786
rect 26976 19722 27028 19728
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 26332 18352 26384 18358
rect 26332 18294 26384 18300
rect 26344 17882 26372 18294
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24688 14074 24716 14758
rect 24780 14346 24808 14962
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24964 14074 24992 15982
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24584 13796 24636 13802
rect 24504 13756 24552 13784
rect 24524 13546 24552 13756
rect 24584 13738 24636 13744
rect 24504 13518 24552 13546
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24412 10674 24440 12038
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24412 7546 24440 8842
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24504 6458 24532 13518
rect 25056 13258 25084 16050
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25240 14958 25268 15302
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 14074 25268 14214
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24780 12306 24808 12786
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24780 11830 24808 12038
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24596 11529 24624 11630
rect 24582 11520 24638 11529
rect 24582 11455 24638 11464
rect 24596 8430 24624 11455
rect 24872 11354 24900 12038
rect 24964 11762 24992 12582
rect 25332 12434 25360 16526
rect 25332 12406 25452 12434
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25240 11082 25268 12242
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24688 9654 24716 10406
rect 25056 9722 25084 10406
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24688 9178 24716 9590
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24688 8498 24716 8910
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24596 6730 24624 8366
rect 25056 7954 25084 9658
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 25056 7002 25084 7890
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 24674 6896 24730 6905
rect 24674 6831 24730 6840
rect 25044 6860 25096 6866
rect 24584 6724 24636 6730
rect 24584 6666 24636 6672
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24688 6322 24716 6831
rect 25044 6802 25096 6808
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24412 5914 24440 6190
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 24490 5672 24546 5681
rect 24490 5607 24492 5616
rect 24544 5607 24546 5616
rect 24492 5578 24544 5584
rect 24490 5264 24546 5273
rect 24490 5199 24546 5208
rect 24504 5166 24532 5199
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 24504 4826 24532 4966
rect 24492 4820 24544 4826
rect 24492 4762 24544 4768
rect 24596 4706 24624 6190
rect 25056 6118 25084 6802
rect 25148 6798 25176 7686
rect 25240 6866 25268 11018
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25332 7002 25360 7346
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 25228 6860 25280 6866
rect 25228 6802 25280 6808
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 4826 24808 5646
rect 24964 5370 24992 5782
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24504 4678 24624 4706
rect 24504 4146 24532 4678
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24504 3398 24532 4082
rect 24780 3738 24808 4422
rect 24872 4282 24900 5170
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24872 3602 24900 4218
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24964 3194 24992 5170
rect 25056 3738 25084 5510
rect 25148 5234 25176 6054
rect 25332 5710 25360 6938
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25424 5658 25452 12406
rect 25516 12306 25544 16934
rect 25700 15570 25728 17614
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26252 16726 26280 16934
rect 26436 16794 26464 19450
rect 27080 19378 27108 19994
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26528 17134 26556 18158
rect 26792 17876 26844 17882
rect 26792 17818 26844 17824
rect 26804 17338 26832 17818
rect 26896 17746 26924 19246
rect 27172 18630 27200 19314
rect 27356 18970 27384 20878
rect 27448 20398 27476 20878
rect 27724 20534 27752 23258
rect 28000 23118 28028 23462
rect 27896 23112 27948 23118
rect 27896 23054 27948 23060
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 27908 22710 27936 23054
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 28184 22094 28212 23734
rect 28540 23520 28592 23526
rect 28540 23462 28592 23468
rect 28552 22778 28580 23462
rect 28540 22772 28592 22778
rect 28540 22714 28592 22720
rect 28644 22642 28672 25910
rect 28736 24614 28764 26318
rect 28920 26042 28948 26862
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 28724 24608 28776 24614
rect 28724 24550 28776 24556
rect 28736 23594 28764 24550
rect 29012 23662 29040 27474
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 29196 27130 29224 27406
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 29092 26988 29144 26994
rect 29092 26930 29144 26936
rect 29104 25906 29132 26930
rect 29092 25900 29144 25906
rect 29092 25842 29144 25848
rect 29000 23656 29052 23662
rect 29000 23598 29052 23604
rect 28724 23588 28776 23594
rect 28724 23530 28776 23536
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28540 22432 28592 22438
rect 28540 22374 28592 22380
rect 28448 22160 28500 22166
rect 28448 22102 28500 22108
rect 28184 22066 28396 22094
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28000 20806 28028 21286
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27540 19718 27568 20402
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27632 20058 27660 20334
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 27528 19712 27580 19718
rect 27528 19654 27580 19660
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 27540 18630 27568 19654
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27448 18222 27476 18566
rect 27540 18426 27568 18566
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27724 18154 27752 20470
rect 27908 19922 27936 20742
rect 28000 20466 28028 20742
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27908 18970 27936 19314
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 27712 18148 27764 18154
rect 27712 18090 27764 18096
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 27724 17678 27752 18090
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26516 17128 26568 17134
rect 26516 17070 26568 17076
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26240 16720 26292 16726
rect 26240 16662 26292 16668
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25700 14482 25728 15506
rect 26068 15094 26096 16594
rect 26252 16538 26280 16662
rect 26160 16510 26280 16538
rect 26344 16522 26556 16538
rect 26332 16516 26556 16522
rect 26160 16114 26188 16510
rect 26384 16510 26556 16516
rect 26332 16458 26384 16464
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26252 15706 26280 16118
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 26056 15088 26108 15094
rect 25976 15036 26056 15042
rect 25976 15030 26108 15036
rect 25976 15014 26096 15030
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 25700 13954 25728 14418
rect 25976 14074 26004 15014
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 25700 13926 25820 13954
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25700 12850 25728 13806
rect 25792 13394 25820 13926
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25516 11150 25544 12242
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25608 11218 25636 11494
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25516 8906 25544 9318
rect 25504 8900 25556 8906
rect 25504 8842 25556 8848
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25228 5636 25280 5642
rect 25424 5630 25636 5658
rect 25228 5578 25280 5584
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25148 4214 25176 4558
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 23492 1550 23612 1578
rect 23492 800 23520 1550
rect 23860 870 23980 898
rect 23860 800 23888 870
rect 21744 734 21956 762
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 23952 762 23980 870
rect 24136 762 24164 2314
rect 24320 1442 24348 2790
rect 24768 2372 24820 2378
rect 24228 1414 24348 1442
rect 24596 2332 24768 2360
rect 24228 800 24256 1414
rect 24596 800 24624 2332
rect 24768 2314 24820 2320
rect 24964 800 24992 2926
rect 25240 2650 25268 5578
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 25332 4690 25360 5306
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25424 4146 25452 5510
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25320 3120 25372 3126
rect 25320 3062 25372 3068
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25332 800 25360 3062
rect 25516 2446 25544 5510
rect 25608 3913 25636 5630
rect 25700 4049 25728 7686
rect 25792 5710 25820 12038
rect 25976 6662 26004 14010
rect 26068 13530 26096 14894
rect 26252 14482 26280 15642
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 26252 12238 26280 14418
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26344 13530 26372 14214
rect 26436 13938 26464 16390
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26528 13802 26556 16510
rect 26804 15502 26832 16934
rect 27080 16658 27108 16934
rect 27448 16658 27476 17070
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26712 14074 26740 15098
rect 27068 14952 27120 14958
rect 27448 14906 27476 16594
rect 27632 16454 27660 17070
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27068 14894 27120 14900
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26988 14074 27016 14214
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 26516 13796 26568 13802
rect 26516 13738 26568 13744
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26528 13190 26556 13738
rect 27080 13530 27108 14894
rect 27172 14890 27476 14906
rect 27160 14884 27476 14890
rect 27212 14878 27476 14884
rect 27160 14826 27212 14832
rect 27448 14006 27476 14878
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27540 13870 27568 14350
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 26608 13524 26660 13530
rect 26608 13466 26660 13472
rect 27068 13524 27120 13530
rect 27068 13466 27120 13472
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26056 11144 26108 11150
rect 26054 11112 26056 11121
rect 26108 11112 26110 11121
rect 26054 11047 26110 11056
rect 26160 10810 26188 11698
rect 26240 11144 26292 11150
rect 26344 11132 26372 12582
rect 26292 11104 26372 11132
rect 26240 11086 26292 11092
rect 26620 10962 26648 13466
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26712 12170 26740 12582
rect 26804 12434 26832 13126
rect 26804 12406 26924 12434
rect 26700 12164 26752 12170
rect 26700 12106 26752 12112
rect 26792 11008 26844 11014
rect 26620 10956 26792 10962
rect 26620 10950 26844 10956
rect 26620 10934 26832 10950
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26804 9926 26832 10934
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 26804 9654 26832 9862
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26252 8090 26280 8366
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26148 7948 26200 7954
rect 26148 7890 26200 7896
rect 26160 7206 26188 7890
rect 26240 7472 26292 7478
rect 26240 7414 26292 7420
rect 26148 7200 26200 7206
rect 26148 7142 26200 7148
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25976 6458 26004 6598
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25976 6254 26004 6394
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 25884 5710 25912 6190
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25686 4040 25742 4049
rect 25686 3975 25742 3984
rect 26068 3942 26096 6258
rect 26160 6118 26188 6734
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26252 5914 26280 7414
rect 26344 6662 26372 9454
rect 26608 9104 26660 9110
rect 26608 9046 26660 9052
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 26436 7954 26464 8570
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26528 7750 26556 8774
rect 26620 7954 26648 9046
rect 26804 7954 26832 9590
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 26620 6866 26648 7890
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26332 6316 26384 6322
rect 26332 6258 26384 6264
rect 26344 6118 26372 6258
rect 26700 6180 26752 6186
rect 26700 6122 26752 6128
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26240 5908 26292 5914
rect 26240 5850 26292 5856
rect 26252 5234 26280 5850
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 26252 4010 26280 4558
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26056 3936 26108 3942
rect 25594 3904 25650 3913
rect 26056 3878 26108 3884
rect 25594 3839 25650 3848
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25700 870 25820 898
rect 25700 800 25728 870
rect 23952 734 24164 762
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 25792 762 25820 870
rect 25976 762 26004 3470
rect 26344 3058 26372 4966
rect 26436 4622 26464 5306
rect 26712 5234 26740 6122
rect 26792 5772 26844 5778
rect 26792 5714 26844 5720
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 26424 4616 26476 4622
rect 26424 4558 26476 4564
rect 26528 4282 26556 5170
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 26606 3496 26662 3505
rect 26712 3466 26740 4966
rect 26606 3431 26662 3440
rect 26700 3460 26752 3466
rect 26620 3194 26648 3431
rect 26700 3402 26752 3408
rect 26804 3194 26832 5714
rect 26896 5098 26924 12406
rect 27080 12170 27108 13466
rect 27344 13184 27396 13190
rect 27344 13126 27396 13132
rect 27356 12986 27384 13126
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27448 12782 27476 13806
rect 27528 13184 27580 13190
rect 27528 13126 27580 13132
rect 27540 12782 27568 13126
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27068 12164 27120 12170
rect 27068 12106 27120 12112
rect 27080 11830 27108 12106
rect 27448 12102 27476 12718
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27068 11824 27120 11830
rect 27068 11766 27120 11772
rect 27080 10266 27108 11766
rect 27448 10674 27476 12038
rect 27632 10810 27660 14758
rect 27724 14074 27752 16050
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27816 15026 27844 15642
rect 27908 15638 27936 17070
rect 28000 16726 28028 20402
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28092 19514 28120 19790
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28092 18834 28120 19450
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 28184 17746 28212 19246
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28276 18426 28304 18702
rect 28264 18420 28316 18426
rect 28264 18362 28316 18368
rect 28172 17740 28224 17746
rect 28172 17682 28224 17688
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 27988 16720 28040 16726
rect 27988 16662 28040 16668
rect 28276 16658 28304 17614
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 27988 16448 28040 16454
rect 27988 16390 28040 16396
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 27896 15632 27948 15638
rect 27896 15574 27948 15580
rect 27804 15020 27856 15026
rect 27804 14962 27856 14968
rect 28000 14482 28028 16390
rect 28092 14618 28120 16390
rect 28080 14612 28132 14618
rect 28080 14554 28132 14560
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 28368 13530 28396 22066
rect 28460 21962 28488 22102
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28552 20482 28580 22374
rect 28736 20584 28764 23530
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 28816 22228 28868 22234
rect 28816 22170 28868 22176
rect 28828 21894 28856 22170
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28736 20556 28856 20584
rect 28552 20454 28764 20482
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28552 18426 28580 19722
rect 28736 18902 28764 20454
rect 28828 19224 28856 20556
rect 28920 20262 28948 22646
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 28908 20256 28960 20262
rect 28908 20198 28960 20204
rect 28920 19514 28948 20198
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28908 19236 28960 19242
rect 28828 19196 28908 19224
rect 28828 18970 28856 19196
rect 28908 19178 28960 19184
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 28724 18896 28776 18902
rect 28724 18838 28776 18844
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28828 18714 28856 18770
rect 28736 18686 28856 18714
rect 28540 18420 28592 18426
rect 28540 18362 28592 18368
rect 28736 18086 28764 18686
rect 29012 18222 29040 22510
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28540 16652 28592 16658
rect 28540 16594 28592 16600
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28460 14958 28488 15846
rect 28552 15706 28580 16594
rect 28644 16182 28672 17614
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28632 14952 28684 14958
rect 28632 14894 28684 14900
rect 28644 14550 28672 14894
rect 28632 14544 28684 14550
rect 28632 14486 28684 14492
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 28736 13462 28764 18022
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29012 17338 29040 17478
rect 29104 17338 29132 25842
rect 29288 25294 29316 27526
rect 29472 26994 29500 30738
rect 31024 30728 31076 30734
rect 31024 30670 31076 30676
rect 30472 30660 30524 30666
rect 30472 30602 30524 30608
rect 29552 30592 29604 30598
rect 29552 30534 29604 30540
rect 29564 30258 29592 30534
rect 30484 30394 30512 30602
rect 31036 30394 31064 30670
rect 30472 30388 30524 30394
rect 30472 30330 30524 30336
rect 31024 30388 31076 30394
rect 31024 30330 31076 30336
rect 29552 30252 29604 30258
rect 29552 30194 29604 30200
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30668 29850 30696 30194
rect 30656 29844 30708 29850
rect 30656 29786 30708 29792
rect 31128 29034 31156 31078
rect 31300 30660 31352 30666
rect 31300 30602 31352 30608
rect 31312 29306 31340 30602
rect 31772 29646 31800 31758
rect 32048 30054 32076 31758
rect 33324 31408 33376 31414
rect 33324 31350 33376 31356
rect 32312 31136 32364 31142
rect 32312 31078 32364 31084
rect 32324 30734 32352 31078
rect 33140 30932 33192 30938
rect 33140 30874 33192 30880
rect 32312 30728 32364 30734
rect 32312 30670 32364 30676
rect 32324 30394 32352 30670
rect 33048 30592 33100 30598
rect 33048 30534 33100 30540
rect 32312 30388 32364 30394
rect 32312 30330 32364 30336
rect 32324 30274 32352 30330
rect 32324 30246 32444 30274
rect 33060 30258 33088 30534
rect 32036 30048 32088 30054
rect 32036 29990 32088 29996
rect 32048 29850 32076 29990
rect 32036 29844 32088 29850
rect 32036 29786 32088 29792
rect 31760 29640 31812 29646
rect 31760 29582 31812 29588
rect 32220 29504 32272 29510
rect 32220 29446 32272 29452
rect 32232 29306 32260 29446
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32220 29096 32272 29102
rect 32218 29064 32220 29073
rect 32272 29064 32274 29073
rect 30748 29028 30800 29034
rect 30748 28970 30800 28976
rect 31116 29028 31168 29034
rect 32218 28999 32274 29008
rect 31116 28970 31168 28976
rect 30564 27464 30616 27470
rect 30564 27406 30616 27412
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 29564 27130 29592 27270
rect 29552 27124 29604 27130
rect 29552 27066 29604 27072
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29656 26586 29684 26930
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 30012 26784 30064 26790
rect 30012 26726 30064 26732
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 30024 26382 30052 26726
rect 30300 26586 30328 26862
rect 30576 26790 30604 27406
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30668 27130 30696 27270
rect 30656 27124 30708 27130
rect 30656 27066 30708 27072
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30288 26580 30340 26586
rect 30288 26522 30340 26528
rect 30576 26450 30604 26726
rect 30564 26444 30616 26450
rect 30564 26386 30616 26392
rect 30012 26376 30064 26382
rect 30012 26318 30064 26324
rect 30760 25362 30788 28970
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 29644 25356 29696 25362
rect 29644 25298 29696 25304
rect 30748 25356 30800 25362
rect 30748 25298 30800 25304
rect 29276 25288 29328 25294
rect 29276 25230 29328 25236
rect 29288 24750 29316 25230
rect 29552 25152 29604 25158
rect 29552 25094 29604 25100
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29288 24070 29316 24686
rect 29276 24064 29328 24070
rect 29276 24006 29328 24012
rect 29380 23730 29408 24754
rect 29564 24206 29592 25094
rect 29656 24274 29684 25298
rect 30196 25288 30248 25294
rect 30196 25230 30248 25236
rect 29828 24744 29880 24750
rect 29828 24686 29880 24692
rect 29736 24676 29788 24682
rect 29736 24618 29788 24624
rect 29748 24274 29776 24618
rect 29840 24410 29868 24686
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29828 24404 29880 24410
rect 29828 24346 29880 24352
rect 29644 24268 29696 24274
rect 29644 24210 29696 24216
rect 29736 24268 29788 24274
rect 29736 24210 29788 24216
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29748 23866 29776 24210
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29380 23322 29408 23666
rect 29840 23662 29868 24346
rect 29932 24274 29960 24550
rect 30208 24410 30236 25230
rect 30748 24608 30800 24614
rect 30748 24550 30800 24556
rect 30196 24404 30248 24410
rect 30196 24346 30248 24352
rect 29920 24268 29972 24274
rect 29920 24210 29972 24216
rect 30760 24206 30788 24550
rect 30748 24200 30800 24206
rect 30748 24142 30800 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 30288 24132 30340 24138
rect 30288 24074 30340 24080
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 30208 23769 30236 24006
rect 30194 23760 30250 23769
rect 30300 23730 30328 24074
rect 30380 24064 30432 24070
rect 30380 24006 30432 24012
rect 30194 23695 30250 23704
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 29368 23316 29420 23322
rect 29368 23258 29420 23264
rect 30116 22778 30144 23598
rect 30300 23322 30328 23666
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30104 22772 30156 22778
rect 30104 22714 30156 22720
rect 30392 22710 30420 24006
rect 30944 23866 30972 24142
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 30472 23656 30524 23662
rect 30472 23598 30524 23604
rect 30380 22704 30432 22710
rect 30380 22646 30432 22652
rect 30484 22522 30512 23598
rect 30392 22494 30512 22522
rect 30392 22438 30420 22494
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 29380 21894 29408 22170
rect 30392 22166 30420 22374
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 29368 21888 29420 21894
rect 29368 21830 29420 21836
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 29104 15706 29132 16390
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 28816 15428 28868 15434
rect 28816 15370 28868 15376
rect 28828 14958 28856 15370
rect 28816 14952 28868 14958
rect 28816 14894 28868 14900
rect 28724 13456 28776 13462
rect 28724 13398 28776 13404
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27724 12306 27752 13262
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 28000 11898 28028 12038
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27724 11744 27752 11834
rect 27804 11756 27856 11762
rect 27724 11716 27804 11744
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27356 10266 27384 10610
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 27528 10192 27580 10198
rect 27528 10134 27580 10140
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27080 8634 27108 8910
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 27172 8430 27200 9318
rect 27540 8838 27568 10134
rect 27724 10130 27752 11716
rect 27804 11698 27856 11704
rect 27896 11688 27948 11694
rect 27896 11630 27948 11636
rect 27804 11280 27856 11286
rect 27908 11268 27936 11630
rect 28080 11620 28132 11626
rect 28080 11562 28132 11568
rect 27856 11240 27936 11268
rect 27804 11222 27856 11228
rect 28092 11082 28120 11562
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27712 10124 27764 10130
rect 27712 10066 27764 10072
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 27066 7712 27122 7721
rect 27066 7647 27122 7656
rect 27080 7342 27108 7647
rect 27264 7546 27292 8774
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 27252 7404 27304 7410
rect 27356 7392 27384 8230
rect 27632 7954 27660 8910
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27304 7364 27384 7392
rect 27252 7346 27304 7352
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27172 7002 27200 7346
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 27264 6882 27292 7346
rect 27632 7206 27660 7890
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27712 7200 27764 7206
rect 27712 7142 27764 7148
rect 27172 6854 27292 6882
rect 27724 6866 27752 7142
rect 27712 6860 27764 6866
rect 27172 6322 27200 6854
rect 27712 6802 27764 6808
rect 27816 6458 27844 10406
rect 28184 8906 28212 13330
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28448 12912 28500 12918
rect 28448 12854 28500 12860
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 28368 12442 28396 12718
rect 28460 12442 28488 12854
rect 28540 12640 28592 12646
rect 28540 12582 28592 12588
rect 28356 12436 28408 12442
rect 28356 12378 28408 12384
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 28552 12306 28580 12582
rect 28540 12300 28592 12306
rect 28540 12242 28592 12248
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28460 11762 28488 12106
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28276 10810 28304 11494
rect 28354 11112 28410 11121
rect 28354 11047 28410 11056
rect 28264 10804 28316 10810
rect 28264 10746 28316 10752
rect 28368 10606 28396 11047
rect 28264 10600 28316 10606
rect 28264 10542 28316 10548
rect 28356 10600 28408 10606
rect 28356 10542 28408 10548
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 28000 7274 28028 8774
rect 28276 7546 28304 10542
rect 28368 10198 28396 10542
rect 28356 10192 28408 10198
rect 28356 10134 28408 10140
rect 28368 9722 28396 10134
rect 28356 9716 28408 9722
rect 28356 9658 28408 9664
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28368 8090 28396 8366
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 27988 7268 28040 7274
rect 27988 7210 28040 7216
rect 28000 7002 28028 7210
rect 27988 6996 28040 7002
rect 27988 6938 28040 6944
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27252 6384 27304 6390
rect 27252 6326 27304 6332
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 27068 5704 27120 5710
rect 27068 5646 27120 5652
rect 27080 5370 27108 5646
rect 27068 5364 27120 5370
rect 27068 5306 27120 5312
rect 27172 5166 27200 6258
rect 27068 5160 27120 5166
rect 27066 5128 27068 5137
rect 27160 5160 27212 5166
rect 27120 5128 27122 5137
rect 26884 5092 26936 5098
rect 27160 5102 27212 5108
rect 27066 5063 27122 5072
rect 26884 5034 26936 5040
rect 26896 4078 26924 5034
rect 27172 4214 27200 5102
rect 27160 4208 27212 4214
rect 27160 4150 27212 4156
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 26160 898 26188 2450
rect 26436 2446 26464 2926
rect 26884 2916 26936 2922
rect 26884 2858 26936 2864
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26528 2446 26556 2790
rect 26896 2774 26924 2858
rect 26712 2746 26924 2774
rect 26606 2680 26662 2689
rect 26606 2615 26608 2624
rect 26660 2615 26662 2624
rect 26608 2586 26660 2592
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 26068 870 26188 898
rect 26436 870 26556 898
rect 26068 800 26096 870
rect 26436 800 26464 870
rect 25792 734 26004 762
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26528 762 26556 870
rect 26712 762 26740 2746
rect 26988 1850 27016 3402
rect 27264 2446 27292 6326
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27436 5092 27488 5098
rect 27436 5034 27488 5040
rect 27448 4690 27476 5034
rect 27540 4690 27568 6190
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27712 6112 27764 6118
rect 27712 6054 27764 6060
rect 27632 5166 27660 6054
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27618 4992 27674 5001
rect 27618 4927 27674 4936
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27448 4486 27476 4626
rect 27344 4480 27396 4486
rect 27344 4422 27396 4428
rect 27436 4480 27488 4486
rect 27436 4422 27488 4428
rect 27356 4282 27384 4422
rect 27344 4276 27396 4282
rect 27344 4218 27396 4224
rect 27436 4072 27488 4078
rect 27434 4040 27436 4049
rect 27488 4040 27490 4049
rect 27434 3975 27490 3984
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27448 3602 27476 3878
rect 27540 3738 27568 4626
rect 27632 4078 27660 4927
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27436 3596 27488 3602
rect 27436 3538 27488 3544
rect 27724 3194 27752 6054
rect 27896 5568 27948 5574
rect 27896 5510 27948 5516
rect 27908 4162 27936 5510
rect 27816 4146 27936 4162
rect 28000 4146 28028 6938
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 28460 4826 28488 6734
rect 28644 6458 28672 13194
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 28828 12374 28856 12718
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28828 11762 28856 12310
rect 29092 12096 29144 12102
rect 29092 12038 29144 12044
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 29000 11688 29052 11694
rect 29000 11630 29052 11636
rect 28736 11370 28764 11630
rect 29012 11529 29040 11630
rect 28998 11520 29054 11529
rect 28998 11455 29054 11464
rect 28736 11354 28856 11370
rect 29012 11354 29040 11455
rect 28736 11348 28868 11354
rect 28736 11342 28816 11348
rect 28736 10674 28764 11342
rect 28816 11290 28868 11296
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29104 11150 29132 12038
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 29196 10198 29224 17478
rect 29288 13190 29316 21286
rect 29380 21146 29408 21830
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29380 19922 29408 21082
rect 29368 19916 29420 19922
rect 29368 19858 29420 19864
rect 29380 19514 29408 19858
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29368 19508 29420 19514
rect 29368 19450 29420 19456
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18426 29592 18566
rect 29932 18426 29960 19654
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30024 18426 30052 19110
rect 30208 18630 30236 21490
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 30484 20602 30512 21422
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30392 19854 30420 19994
rect 30484 19922 30512 20538
rect 30944 20534 30972 21286
rect 31036 20806 31064 28358
rect 31128 27146 31156 28970
rect 32416 28422 32444 30246
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 32772 30184 32824 30190
rect 32824 30144 32904 30172
rect 32772 30126 32824 30132
rect 32770 29744 32826 29753
rect 32770 29679 32772 29688
rect 32824 29679 32826 29688
rect 32772 29650 32824 29656
rect 32588 29504 32640 29510
rect 32588 29446 32640 29452
rect 32680 29504 32732 29510
rect 32680 29446 32732 29452
rect 32600 29170 32628 29446
rect 32692 29306 32720 29446
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 32588 29164 32640 29170
rect 32588 29106 32640 29112
rect 32404 28416 32456 28422
rect 32404 28358 32456 28364
rect 31392 27872 31444 27878
rect 31392 27814 31444 27820
rect 31128 27118 31248 27146
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 31128 24410 31156 24890
rect 31116 24404 31168 24410
rect 31116 24346 31168 24352
rect 31220 24290 31248 27118
rect 31404 26382 31432 27814
rect 31576 27668 31628 27674
rect 31576 27610 31628 27616
rect 31588 26926 31616 27610
rect 32416 27470 32444 28358
rect 32600 28082 32628 29106
rect 32784 29034 32812 29650
rect 32772 29028 32824 29034
rect 32772 28970 32824 28976
rect 32588 28076 32640 28082
rect 32588 28018 32640 28024
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32600 27334 32628 28018
rect 32128 27328 32180 27334
rect 32128 27270 32180 27276
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 31576 26920 31628 26926
rect 31576 26862 31628 26868
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31588 26042 31616 26862
rect 32140 26042 32168 27270
rect 31576 26036 31628 26042
rect 31576 25978 31628 25984
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32600 25974 32628 27270
rect 32772 26988 32824 26994
rect 32876 26976 32904 30144
rect 32968 29850 32996 30194
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32956 29572 33008 29578
rect 32956 29514 33008 29520
rect 32968 29170 32996 29514
rect 33060 29170 33088 30194
rect 33152 29714 33180 30874
rect 33232 30660 33284 30666
rect 33232 30602 33284 30608
rect 33244 29850 33272 30602
rect 33336 30394 33364 31350
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 33784 31204 33836 31210
rect 33784 31146 33836 31152
rect 33324 30388 33376 30394
rect 33324 30330 33376 30336
rect 33600 30388 33652 30394
rect 33600 30330 33652 30336
rect 33336 30122 33364 30330
rect 33324 30116 33376 30122
rect 33324 30058 33376 30064
rect 33416 30048 33468 30054
rect 33416 29990 33468 29996
rect 33232 29844 33284 29850
rect 33232 29786 33284 29792
rect 33140 29708 33192 29714
rect 33140 29650 33192 29656
rect 33152 29617 33180 29650
rect 33138 29608 33194 29617
rect 33138 29543 33194 29552
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 33152 29102 33180 29543
rect 33140 29096 33192 29102
rect 33140 29038 33192 29044
rect 33140 28552 33192 28558
rect 33140 28494 33192 28500
rect 32956 28416 33008 28422
rect 32956 28358 33008 28364
rect 32968 28218 32996 28358
rect 32956 28212 33008 28218
rect 32956 28154 33008 28160
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32824 26948 32904 26976
rect 32772 26930 32824 26936
rect 32968 26042 32996 27814
rect 33152 27010 33180 28494
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 33244 27130 33272 27950
rect 33324 27600 33376 27606
rect 33324 27542 33376 27548
rect 33232 27124 33284 27130
rect 33232 27066 33284 27072
rect 33060 26994 33180 27010
rect 33048 26988 33180 26994
rect 33100 26982 33180 26988
rect 33048 26930 33100 26936
rect 33152 26382 33180 26982
rect 33244 26926 33272 27066
rect 33232 26920 33284 26926
rect 33232 26862 33284 26868
rect 33232 26784 33284 26790
rect 33232 26726 33284 26732
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 33244 26042 33272 26726
rect 32956 26036 33008 26042
rect 32956 25978 33008 25984
rect 33232 26036 33284 26042
rect 33232 25978 33284 25984
rect 32588 25968 32640 25974
rect 32588 25910 32640 25916
rect 32864 25900 32916 25906
rect 32864 25842 32916 25848
rect 31944 25696 31996 25702
rect 31944 25638 31996 25644
rect 31128 24262 31248 24290
rect 31128 23662 31156 24262
rect 31852 24064 31904 24070
rect 31852 24006 31904 24012
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31128 23254 31156 23598
rect 31116 23248 31168 23254
rect 31116 23190 31168 23196
rect 31864 23050 31892 24006
rect 31852 23044 31904 23050
rect 31852 22986 31904 22992
rect 31956 21962 31984 25638
rect 32876 25498 32904 25842
rect 32864 25492 32916 25498
rect 32864 25434 32916 25440
rect 33336 24342 33364 27542
rect 33428 25838 33456 29990
rect 33612 26858 33640 30330
rect 33796 30258 33824 31146
rect 33968 30796 34020 30802
rect 33968 30738 34020 30744
rect 33876 30592 33928 30598
rect 33876 30534 33928 30540
rect 33784 30252 33836 30258
rect 33784 30194 33836 30200
rect 33888 29306 33916 30534
rect 33980 30258 34008 30738
rect 33968 30252 34020 30258
rect 33968 30194 34020 30200
rect 34164 29850 34192 31214
rect 34336 31136 34388 31142
rect 34336 31078 34388 31084
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 34348 29646 34376 31078
rect 34428 30388 34480 30394
rect 34428 30330 34480 30336
rect 34440 29730 34468 30330
rect 34716 30326 34744 31826
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 35348 31680 35400 31686
rect 35348 31622 35400 31628
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30666 35388 31622
rect 35348 30660 35400 30666
rect 35348 30602 35400 30608
rect 34704 30320 34756 30326
rect 34704 30262 34756 30268
rect 34612 30184 34664 30190
rect 34612 30126 34664 30132
rect 34704 30184 34756 30190
rect 34704 30126 34756 30132
rect 34440 29702 34560 29730
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 34428 29640 34480 29646
rect 34428 29582 34480 29588
rect 34440 29306 34468 29582
rect 34532 29306 34560 29702
rect 34624 29510 34652 30126
rect 34716 29578 34744 30126
rect 35452 30122 35480 31758
rect 36372 31414 36400 32166
rect 36452 31816 36504 31822
rect 36452 31758 36504 31764
rect 36360 31408 36412 31414
rect 36360 31350 36412 31356
rect 35808 31136 35860 31142
rect 35808 31078 35860 31084
rect 36176 31136 36228 31142
rect 36176 31078 36228 31084
rect 35820 30734 35848 31078
rect 35808 30728 35860 30734
rect 35808 30670 35860 30676
rect 34796 30116 34848 30122
rect 34796 30058 34848 30064
rect 35440 30116 35492 30122
rect 35440 30058 35492 30064
rect 34704 29572 34756 29578
rect 34704 29514 34756 29520
rect 34612 29504 34664 29510
rect 34612 29446 34664 29452
rect 33876 29300 33928 29306
rect 33876 29242 33928 29248
rect 34428 29300 34480 29306
rect 34428 29242 34480 29248
rect 34520 29300 34572 29306
rect 34520 29242 34572 29248
rect 34244 28552 34296 28558
rect 34244 28494 34296 28500
rect 33692 28416 33744 28422
rect 33692 28358 33744 28364
rect 33704 27538 33732 28358
rect 33784 28008 33836 28014
rect 33784 27950 33836 27956
rect 33692 27532 33744 27538
rect 33692 27474 33744 27480
rect 33796 26926 33824 27950
rect 34256 27538 34284 28494
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34336 27872 34388 27878
rect 34336 27814 34388 27820
rect 34244 27532 34296 27538
rect 34244 27474 34296 27480
rect 34152 27328 34204 27334
rect 34152 27270 34204 27276
rect 33784 26920 33836 26926
rect 33784 26862 33836 26868
rect 34164 26874 34192 27270
rect 34256 26994 34284 27474
rect 34348 27130 34376 27814
rect 34532 27334 34560 27950
rect 34520 27328 34572 27334
rect 34520 27270 34572 27276
rect 34336 27124 34388 27130
rect 34336 27066 34388 27072
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 33600 26852 33652 26858
rect 33600 26794 33652 26800
rect 33612 26246 33640 26794
rect 33796 26586 33824 26862
rect 34164 26858 34284 26874
rect 34164 26852 34296 26858
rect 34164 26846 34244 26852
rect 34244 26794 34296 26800
rect 33784 26580 33836 26586
rect 33784 26522 33836 26528
rect 33968 26308 34020 26314
rect 33968 26250 34020 26256
rect 33600 26240 33652 26246
rect 33600 26182 33652 26188
rect 33612 26042 33640 26182
rect 33980 26042 34008 26250
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33968 26036 34020 26042
rect 33968 25978 34020 25984
rect 33416 25832 33468 25838
rect 33416 25774 33468 25780
rect 33692 25696 33744 25702
rect 33692 25638 33744 25644
rect 32588 24336 32640 24342
rect 32588 24278 32640 24284
rect 33324 24336 33376 24342
rect 33324 24278 33376 24284
rect 32600 23322 32628 24278
rect 33324 23520 33376 23526
rect 33324 23462 33376 23468
rect 32588 23316 32640 23322
rect 32588 23258 32640 23264
rect 32600 23186 32628 23258
rect 32588 23180 32640 23186
rect 32588 23122 32640 23128
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 32324 22642 32352 23054
rect 32588 22976 32640 22982
rect 32588 22918 32640 22924
rect 32600 22642 32628 22918
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32588 22636 32640 22642
rect 32588 22578 32640 22584
rect 32220 22094 32272 22098
rect 32324 22094 32352 22578
rect 32220 22092 32352 22094
rect 32272 22066 32352 22092
rect 32220 22034 32272 22040
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31956 21554 31984 21898
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 32416 21146 32444 21830
rect 32784 21690 32812 23054
rect 33048 22976 33100 22982
rect 33048 22918 33100 22924
rect 33060 22030 33088 22918
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33336 21690 33364 23462
rect 33600 23044 33652 23050
rect 33600 22986 33652 22992
rect 33612 21690 33640 22986
rect 32772 21684 32824 21690
rect 32772 21626 32824 21632
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 33600 21684 33652 21690
rect 33600 21626 33652 21632
rect 33416 21412 33468 21418
rect 33416 21354 33468 21360
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 31220 20602 31248 20810
rect 31208 20596 31260 20602
rect 31208 20538 31260 20544
rect 30932 20528 30984 20534
rect 30932 20470 30984 20476
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31128 19990 31156 20402
rect 31312 19990 31340 21082
rect 31392 20936 31444 20942
rect 31392 20878 31444 20884
rect 31404 20398 31432 20878
rect 33428 20602 33456 21354
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 33428 20466 33456 20538
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 31760 20392 31812 20398
rect 31760 20334 31812 20340
rect 30656 19984 30708 19990
rect 30656 19926 30708 19932
rect 31116 19984 31168 19990
rect 31116 19926 31168 19932
rect 31300 19984 31352 19990
rect 31300 19926 31352 19932
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30392 19514 30420 19654
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30668 18970 30696 19926
rect 31312 19854 31340 19926
rect 31024 19848 31076 19854
rect 31024 19790 31076 19796
rect 31300 19848 31352 19854
rect 31300 19790 31352 19796
rect 31036 19446 31064 19790
rect 31024 19440 31076 19446
rect 31024 19382 31076 19388
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 30748 19304 30800 19310
rect 30748 19246 30800 19252
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 29552 18420 29604 18426
rect 29552 18362 29604 18368
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29748 17542 29776 18158
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29920 17196 29972 17202
rect 29920 17138 29972 17144
rect 29552 16720 29604 16726
rect 29552 16662 29604 16668
rect 29564 16250 29592 16662
rect 29552 16244 29604 16250
rect 29552 16186 29604 16192
rect 29564 15094 29592 16186
rect 29736 16040 29788 16046
rect 29736 15982 29788 15988
rect 29748 15502 29776 15982
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29932 15450 29960 17138
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29564 14074 29592 15030
rect 29748 14278 29776 15438
rect 29932 15422 30052 15450
rect 29920 15360 29972 15366
rect 29920 15302 29972 15308
rect 29736 14272 29788 14278
rect 29788 14232 29868 14260
rect 29736 14214 29788 14220
rect 29552 14068 29604 14074
rect 29552 14010 29604 14016
rect 29276 13184 29328 13190
rect 29276 13126 29328 13132
rect 29564 12434 29592 14010
rect 29736 13252 29788 13258
rect 29736 13194 29788 13200
rect 29564 12406 29684 12434
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29288 10810 29316 11698
rect 29276 10804 29328 10810
rect 29276 10746 29328 10752
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29184 10192 29236 10198
rect 29184 10134 29236 10140
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 29012 7750 29040 9318
rect 29104 8838 29132 9522
rect 29380 8838 29408 10406
rect 29656 10146 29684 12406
rect 29748 11626 29776 13194
rect 29840 11694 29868 14232
rect 29932 13938 29960 15302
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29932 11830 29960 12582
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29736 11620 29788 11626
rect 29736 11562 29788 11568
rect 29840 11218 29868 11630
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29656 10130 29868 10146
rect 29656 10124 29880 10130
rect 29656 10118 29828 10124
rect 29828 10066 29880 10072
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 29552 8832 29604 8838
rect 29552 8774 29604 8780
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7342 29040 7686
rect 29000 7336 29052 7342
rect 29000 7278 29052 7284
rect 29012 6798 29040 7278
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 29000 6656 29052 6662
rect 29104 6644 29132 8774
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29196 7818 29224 8230
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 29380 7274 29408 8774
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 29472 7886 29500 8366
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29368 7268 29420 7274
rect 29368 7210 29420 7216
rect 29276 7200 29328 7206
rect 29276 7142 29328 7148
rect 29182 6896 29238 6905
rect 29182 6831 29238 6840
rect 29052 6616 29132 6644
rect 29000 6598 29052 6604
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 28552 4622 28580 5510
rect 28644 5370 28672 5646
rect 28632 5364 28684 5370
rect 28632 5306 28684 5312
rect 29012 5302 29040 6598
rect 29196 6322 29224 6831
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29000 5160 29052 5166
rect 29000 5102 29052 5108
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 28920 4826 28948 4966
rect 28908 4820 28960 4826
rect 28908 4762 28960 4768
rect 29012 4622 29040 5102
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 27804 4140 27936 4146
rect 27856 4134 27936 4140
rect 27988 4140 28040 4146
rect 27804 4082 27856 4088
rect 27988 4082 28040 4088
rect 29012 4078 29040 4558
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 26804 1822 27016 1850
rect 26804 800 26832 1822
rect 27356 1578 27384 2926
rect 27526 2816 27582 2825
rect 27526 2751 27582 2760
rect 27172 1550 27384 1578
rect 27172 800 27200 1550
rect 27540 800 27568 2751
rect 27908 800 27936 4014
rect 29104 4010 29132 6258
rect 29288 5642 29316 7142
rect 29276 5636 29328 5642
rect 29276 5578 29328 5584
rect 29184 5296 29236 5302
rect 29184 5238 29236 5244
rect 29196 4457 29224 5238
rect 29380 5114 29408 7210
rect 29472 6934 29500 7822
rect 29460 6928 29512 6934
rect 29460 6870 29512 6876
rect 29472 5234 29500 6870
rect 29564 6390 29592 8774
rect 29748 7410 29776 8910
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 29552 6384 29604 6390
rect 29552 6326 29604 6332
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29460 5228 29512 5234
rect 29460 5170 29512 5176
rect 29380 5086 29500 5114
rect 29276 4820 29328 4826
rect 29276 4762 29328 4768
rect 29182 4448 29238 4457
rect 29182 4383 29238 4392
rect 29184 4208 29236 4214
rect 29184 4150 29236 4156
rect 29092 4004 29144 4010
rect 29092 3946 29144 3952
rect 29196 3738 29224 4150
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 28276 3194 28304 3334
rect 28264 3188 28316 3194
rect 28264 3130 28316 3136
rect 28264 2984 28316 2990
rect 28264 2926 28316 2932
rect 28276 800 28304 2926
rect 29184 2916 29236 2922
rect 29184 2858 29236 2864
rect 28632 2848 28684 2854
rect 28632 2790 28684 2796
rect 28644 800 28672 2790
rect 29196 2446 29224 2858
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29012 800 29040 2314
rect 29288 2310 29316 4762
rect 29368 4548 29420 4554
rect 29368 4490 29420 4496
rect 29380 4282 29408 4490
rect 29472 4486 29500 5086
rect 29460 4480 29512 4486
rect 29460 4422 29512 4428
rect 29368 4276 29420 4282
rect 29368 4218 29420 4224
rect 29564 4146 29592 5510
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29656 3738 29684 7346
rect 29840 7206 29868 10066
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 29932 8090 29960 9454
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 29932 7018 29960 7822
rect 29840 6990 29960 7018
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 29368 3528 29420 3534
rect 29368 3470 29420 3476
rect 29380 2650 29408 3470
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29368 2508 29420 2514
rect 29368 2450 29420 2456
rect 29276 2304 29328 2310
rect 29276 2246 29328 2252
rect 29380 800 29408 2450
rect 29748 2446 29776 6054
rect 29840 5370 29868 6990
rect 29920 6860 29972 6866
rect 30024 6848 30052 15422
rect 30116 15366 30144 15642
rect 30104 15360 30156 15366
rect 30104 15302 30156 15308
rect 30104 14340 30156 14346
rect 30104 14282 30156 14288
rect 30116 14074 30144 14282
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 30116 11898 30144 12174
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 30208 10810 30236 18566
rect 30760 18086 30788 19246
rect 30840 18828 30892 18834
rect 30840 18770 30892 18776
rect 30380 18080 30432 18086
rect 30380 18022 30432 18028
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30392 16674 30420 18022
rect 30392 16646 30512 16674
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 30392 16046 30420 16526
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30288 15564 30340 15570
rect 30288 15506 30340 15512
rect 30300 15162 30328 15506
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 30484 14226 30512 16646
rect 30564 15428 30616 15434
rect 30564 15370 30616 15376
rect 30392 14198 30512 14226
rect 30288 14000 30340 14006
rect 30288 13942 30340 13948
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30300 10470 30328 13942
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30392 8956 30420 14198
rect 30576 14074 30604 15370
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 30668 13954 30696 14758
rect 30760 14618 30788 18022
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30576 13926 30696 13954
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30484 12918 30512 13670
rect 30576 13258 30604 13926
rect 30746 13832 30802 13841
rect 30852 13818 30880 18770
rect 30944 18630 30972 19314
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 31312 18698 31340 19110
rect 31772 18970 31800 20334
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 31864 19378 31892 19994
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 32048 19446 32076 19790
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 32956 19712 33008 19718
rect 32956 19654 33008 19660
rect 32232 19514 32260 19654
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 32036 19440 32088 19446
rect 32036 19382 32088 19388
rect 31852 19372 31904 19378
rect 31852 19314 31904 19320
rect 31760 18964 31812 18970
rect 31760 18906 31812 18912
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31300 18692 31352 18698
rect 31300 18634 31352 18640
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 30944 15570 30972 16934
rect 31404 15978 31616 15994
rect 31404 15972 31628 15978
rect 31404 15966 31576 15972
rect 31404 15570 31432 15966
rect 31576 15914 31628 15920
rect 30932 15564 30984 15570
rect 30932 15506 30984 15512
rect 31392 15564 31444 15570
rect 31392 15506 31444 15512
rect 31576 15564 31628 15570
rect 31576 15506 31628 15512
rect 30802 13790 30880 13818
rect 30746 13767 30802 13776
rect 30944 13734 30972 15506
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31024 14816 31076 14822
rect 31024 14758 31076 14764
rect 31036 14414 31064 14758
rect 31220 14618 31248 15438
rect 31484 15156 31536 15162
rect 31484 15098 31536 15104
rect 31208 14612 31260 14618
rect 31208 14554 31260 14560
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 31220 13938 31248 14554
rect 31496 14278 31524 15098
rect 31588 14890 31616 15506
rect 31576 14884 31628 14890
rect 31576 14826 31628 14832
rect 31484 14272 31536 14278
rect 31484 14214 31536 14220
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30564 13252 30616 13258
rect 30564 13194 30616 13200
rect 30668 12986 30696 13262
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30472 12912 30524 12918
rect 30472 12854 30524 12860
rect 30472 12776 30524 12782
rect 30472 12718 30524 12724
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 30484 10810 30512 12718
rect 30576 12102 30604 12718
rect 30944 12374 30972 13670
rect 31208 13184 31260 13190
rect 31208 13126 31260 13132
rect 31300 13184 31352 13190
rect 31300 13126 31352 13132
rect 31024 12844 31076 12850
rect 31024 12786 31076 12792
rect 30932 12368 30984 12374
rect 30932 12310 30984 12316
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30472 10532 30524 10538
rect 30472 10474 30524 10480
rect 30484 9586 30512 10474
rect 30472 9580 30524 9586
rect 30472 9522 30524 9528
rect 30576 9518 30604 12038
rect 30944 10266 30972 12310
rect 31036 10810 31064 12786
rect 31116 12096 31168 12102
rect 31116 12038 31168 12044
rect 31128 11354 31156 12038
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 31220 11150 31248 13126
rect 31312 12986 31340 13126
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31208 11144 31260 11150
rect 31208 11086 31260 11092
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 31036 10470 31064 10746
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 31312 10266 31340 11290
rect 31392 10464 31444 10470
rect 31392 10406 31444 10412
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 31300 10260 31352 10266
rect 31300 10202 31352 10208
rect 30944 10062 30972 10202
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 30748 9920 30800 9926
rect 30748 9862 30800 9868
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 30656 9376 30708 9382
rect 30656 9318 30708 9324
rect 30576 8974 30604 9318
rect 30564 8968 30616 8974
rect 30392 8928 30512 8956
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30208 7886 30236 8230
rect 30288 7948 30340 7954
rect 30288 7890 30340 7896
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 30300 7002 30328 7890
rect 30288 6996 30340 7002
rect 30288 6938 30340 6944
rect 29972 6820 30052 6848
rect 29920 6802 29972 6808
rect 30104 6792 30156 6798
rect 30300 6769 30328 6938
rect 30104 6734 30156 6740
rect 30286 6760 30342 6769
rect 30116 6361 30144 6734
rect 30286 6695 30342 6704
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30194 6488 30250 6497
rect 30194 6423 30196 6432
rect 30248 6423 30250 6432
rect 30196 6394 30248 6400
rect 30102 6352 30158 6361
rect 30102 6287 30158 6296
rect 30104 6248 30156 6254
rect 30104 6190 30156 6196
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 30024 4690 30052 5306
rect 30012 4684 30064 4690
rect 30012 4626 30064 4632
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 29840 2650 29868 4558
rect 30024 4214 30052 4626
rect 30012 4208 30064 4214
rect 30012 4150 30064 4156
rect 30116 4049 30144 6190
rect 30288 6112 30340 6118
rect 30288 6054 30340 6060
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 30208 4826 30236 5646
rect 30300 5302 30328 6054
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30194 4720 30250 4729
rect 30194 4655 30196 4664
rect 30248 4655 30250 4664
rect 30196 4626 30248 4632
rect 30102 4040 30158 4049
rect 30102 3975 30158 3984
rect 30288 4004 30340 4010
rect 30288 3946 30340 3952
rect 29920 3936 29972 3942
rect 29920 3878 29972 3884
rect 30194 3904 30250 3913
rect 29932 3534 29960 3878
rect 30194 3839 30250 3848
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 29748 870 29868 898
rect 29748 800 29776 870
rect 26528 734 26740 762
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 29840 762 29868 870
rect 30024 762 30052 3674
rect 30104 3392 30156 3398
rect 30104 3334 30156 3340
rect 30116 800 30144 3334
rect 30208 3194 30236 3839
rect 30196 3188 30248 3194
rect 30196 3130 30248 3136
rect 30300 3058 30328 3946
rect 30288 3052 30340 3058
rect 30288 2994 30340 3000
rect 30392 2650 30420 6666
rect 30484 5545 30512 8928
rect 30564 8910 30616 8916
rect 30668 8634 30696 9318
rect 30760 8906 30788 9862
rect 31208 9512 31260 9518
rect 31208 9454 31260 9460
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31024 9376 31076 9382
rect 31024 9318 31076 9324
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30852 7954 30880 9114
rect 30656 7948 30708 7954
rect 30656 7890 30708 7896
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 30668 7546 30696 7890
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30656 7540 30708 7546
rect 30656 7482 30708 7488
rect 30760 6866 30788 7686
rect 30748 6860 30800 6866
rect 30748 6802 30800 6808
rect 30656 6384 30708 6390
rect 30656 6326 30708 6332
rect 30668 5914 30696 6326
rect 30840 6248 30892 6254
rect 30840 6190 30892 6196
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30564 5568 30616 5574
rect 30470 5536 30526 5545
rect 30564 5510 30616 5516
rect 30470 5471 30526 5480
rect 30576 5302 30604 5510
rect 30564 5296 30616 5302
rect 30564 5238 30616 5244
rect 30472 5092 30524 5098
rect 30472 5034 30524 5040
rect 30484 4826 30512 5034
rect 30472 4820 30524 4826
rect 30472 4762 30524 4768
rect 30576 4690 30604 5238
rect 30668 5166 30696 5850
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 30564 4684 30616 4690
rect 30564 4626 30616 4632
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30484 3466 30512 4558
rect 30656 4208 30708 4214
rect 30656 4150 30708 4156
rect 30668 3942 30696 4150
rect 30852 3942 30880 6190
rect 31036 4078 31064 9318
rect 31116 8832 31168 8838
rect 31116 8774 31168 8780
rect 31128 8022 31156 8774
rect 31220 8634 31248 9454
rect 31312 9178 31340 9454
rect 31300 9172 31352 9178
rect 31300 9114 31352 9120
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 31116 8016 31168 8022
rect 31116 7958 31168 7964
rect 31128 6866 31156 7958
rect 31208 7948 31260 7954
rect 31208 7890 31260 7896
rect 31220 7546 31248 7890
rect 31208 7540 31260 7546
rect 31208 7482 31260 7488
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31220 6644 31248 7482
rect 31404 6866 31432 10406
rect 31496 9586 31524 14214
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31680 12102 31708 12174
rect 31668 12096 31720 12102
rect 31668 12038 31720 12044
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31576 10056 31628 10062
rect 31576 9998 31628 10004
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 31496 9382 31524 9522
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31496 8430 31524 9318
rect 31484 8424 31536 8430
rect 31484 8366 31536 8372
rect 31588 8294 31616 9998
rect 31680 9450 31708 10202
rect 31668 9444 31720 9450
rect 31668 9386 31720 9392
rect 31668 8560 31720 8566
rect 31668 8502 31720 8508
rect 31576 8288 31628 8294
rect 31576 8230 31628 8236
rect 31680 7954 31708 8502
rect 31668 7948 31720 7954
rect 31668 7890 31720 7896
rect 31392 6860 31444 6866
rect 31392 6802 31444 6808
rect 31128 6616 31248 6644
rect 31128 5137 31156 6616
rect 31576 6248 31628 6254
rect 31576 6190 31628 6196
rect 31208 6112 31260 6118
rect 31208 6054 31260 6060
rect 31114 5128 31170 5137
rect 31114 5063 31170 5072
rect 31128 4826 31156 5063
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31220 4146 31248 6054
rect 31588 5370 31616 6190
rect 31576 5364 31628 5370
rect 31576 5306 31628 5312
rect 31668 5364 31720 5370
rect 31668 5306 31720 5312
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 31404 4706 31432 5102
rect 31588 4826 31616 5306
rect 31576 4820 31628 4826
rect 31576 4762 31628 4768
rect 31404 4678 31616 4706
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31496 4214 31524 4558
rect 31484 4208 31536 4214
rect 31482 4176 31484 4185
rect 31536 4176 31538 4185
rect 31208 4140 31260 4146
rect 31482 4111 31538 4120
rect 31208 4082 31260 4088
rect 31024 4072 31076 4078
rect 31024 4014 31076 4020
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30932 3936 30984 3942
rect 30932 3878 30984 3884
rect 30944 3738 30972 3878
rect 31588 3738 31616 4678
rect 30932 3732 30984 3738
rect 30932 3674 30984 3680
rect 31576 3732 31628 3738
rect 31576 3674 31628 3680
rect 31680 3602 31708 5306
rect 31772 4146 31800 18770
rect 32968 18766 32996 19654
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 33416 19168 33468 19174
rect 33416 19110 33468 19116
rect 32956 18760 33008 18766
rect 32956 18702 33008 18708
rect 33232 18760 33284 18766
rect 33232 18702 33284 18708
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 33060 17270 33088 18566
rect 33244 18358 33272 18702
rect 33336 18698 33364 19110
rect 33324 18692 33376 18698
rect 33324 18634 33376 18640
rect 33232 18352 33284 18358
rect 33232 18294 33284 18300
rect 33324 17536 33376 17542
rect 33324 17478 33376 17484
rect 33048 17264 33100 17270
rect 33048 17206 33100 17212
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 33152 16658 33180 17070
rect 33140 16652 33192 16658
rect 33140 16594 33192 16600
rect 32588 16584 32640 16590
rect 32588 16526 32640 16532
rect 31852 16448 31904 16454
rect 31852 16390 31904 16396
rect 31864 16182 31892 16390
rect 31852 16176 31904 16182
rect 31852 16118 31904 16124
rect 31864 15638 31892 16118
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 31852 15632 31904 15638
rect 31852 15574 31904 15580
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 32036 13320 32088 13326
rect 32036 13262 32088 13268
rect 31852 12300 31904 12306
rect 31852 12242 31904 12248
rect 31864 11558 31892 12242
rect 31956 12102 31984 13262
rect 32048 12306 32076 13262
rect 32140 12986 32168 15302
rect 32324 14618 32352 15438
rect 32416 15162 32444 15982
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 32508 15042 32536 15302
rect 32416 15026 32536 15042
rect 32404 15020 32536 15026
rect 32456 15014 32536 15020
rect 32404 14962 32456 14968
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 32128 12776 32180 12782
rect 32128 12718 32180 12724
rect 32036 12300 32088 12306
rect 32036 12242 32088 12248
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 32048 11830 32076 12242
rect 32036 11824 32088 11830
rect 32036 11766 32088 11772
rect 31852 11552 31904 11558
rect 31852 11494 31904 11500
rect 31864 10674 31892 11494
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31852 10192 31904 10198
rect 31852 10134 31904 10140
rect 31864 8786 31892 10134
rect 31956 8974 31984 11086
rect 32048 9926 32076 11766
rect 32140 10198 32168 12718
rect 32416 12186 32444 14962
rect 32600 14822 32628 16526
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 32680 15564 32732 15570
rect 32680 15506 32732 15512
rect 32588 14816 32640 14822
rect 32588 14758 32640 14764
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32508 12442 32536 12786
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32416 12158 32536 12186
rect 32508 12102 32536 12158
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32496 12096 32548 12102
rect 32496 12038 32548 12044
rect 32416 11150 32444 12038
rect 32404 11144 32456 11150
rect 32404 11086 32456 11092
rect 32508 10962 32536 12038
rect 32416 10934 32536 10962
rect 32312 10736 32364 10742
rect 32312 10678 32364 10684
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 32128 10192 32180 10198
rect 32128 10134 32180 10140
rect 32140 9926 32168 10134
rect 32232 10062 32260 10542
rect 32220 10056 32272 10062
rect 32220 9998 32272 10004
rect 32036 9920 32088 9926
rect 32036 9862 32088 9868
rect 32128 9920 32180 9926
rect 32128 9862 32180 9868
rect 32232 9654 32260 9998
rect 32220 9648 32272 9654
rect 32220 9590 32272 9596
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 31864 8758 31984 8786
rect 31852 8288 31904 8294
rect 31852 8230 31904 8236
rect 31864 7954 31892 8230
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 31864 7546 31892 7890
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 31956 7426 31984 8758
rect 31864 7398 31984 7426
rect 31864 5273 31892 7398
rect 31944 7336 31996 7342
rect 31944 7278 31996 7284
rect 31956 6866 31984 7278
rect 31944 6860 31996 6866
rect 31944 6802 31996 6808
rect 31956 5710 31984 6802
rect 32324 6458 32352 10678
rect 32416 10606 32444 10934
rect 32404 10600 32456 10606
rect 32404 10542 32456 10548
rect 32416 7206 32444 10542
rect 32692 9586 32720 15506
rect 32876 15162 32904 15846
rect 32864 15156 32916 15162
rect 32864 15098 32916 15104
rect 32772 14884 32824 14890
rect 32968 14872 32996 15846
rect 33140 15632 33192 15638
rect 33140 15574 33192 15580
rect 32824 14844 32996 14872
rect 32772 14826 32824 14832
rect 32784 14074 32812 14826
rect 33152 14482 33180 15574
rect 33336 15570 33364 17478
rect 33324 15564 33376 15570
rect 33324 15506 33376 15512
rect 33232 15360 33284 15366
rect 33232 15302 33284 15308
rect 33244 14618 33272 15302
rect 33232 14612 33284 14618
rect 33232 14554 33284 14560
rect 33140 14476 33192 14482
rect 33140 14418 33192 14424
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32784 12714 32812 14010
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 32772 12708 32824 12714
rect 32772 12650 32824 12656
rect 32784 12442 32812 12650
rect 32956 12640 33008 12646
rect 32956 12582 33008 12588
rect 32772 12436 32824 12442
rect 32772 12378 32824 12384
rect 32784 11354 32812 12378
rect 32968 12306 32996 12582
rect 33152 12306 33180 12718
rect 32956 12300 33008 12306
rect 32956 12242 33008 12248
rect 33140 12300 33192 12306
rect 33140 12242 33192 12248
rect 33152 11898 33180 12242
rect 33232 12096 33284 12102
rect 33232 12038 33284 12044
rect 33140 11892 33192 11898
rect 33140 11834 33192 11840
rect 33244 11762 33272 12038
rect 33232 11756 33284 11762
rect 33232 11698 33284 11704
rect 33428 11665 33456 19110
rect 33600 15904 33652 15910
rect 33600 15846 33652 15852
rect 33612 15162 33640 15846
rect 33600 15156 33652 15162
rect 33600 15098 33652 15104
rect 33704 12918 33732 25638
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33796 22778 33824 24142
rect 33876 23656 33928 23662
rect 33876 23598 33928 23604
rect 33784 22772 33836 22778
rect 33784 22714 33836 22720
rect 33796 21554 33824 22714
rect 33888 22438 33916 23598
rect 33968 22976 34020 22982
rect 33968 22918 34020 22924
rect 33876 22432 33928 22438
rect 33876 22374 33928 22380
rect 33876 22160 33928 22166
rect 33876 22102 33928 22108
rect 33784 21548 33836 21554
rect 33784 21490 33836 21496
rect 33888 21350 33916 22102
rect 33876 21344 33928 21350
rect 33876 21286 33928 21292
rect 33980 20602 34008 22918
rect 34152 21480 34204 21486
rect 34152 21422 34204 21428
rect 34164 21146 34192 21422
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33796 18290 33824 19654
rect 33784 18284 33836 18290
rect 33784 18226 33836 18232
rect 33782 17640 33838 17649
rect 33782 17575 33838 17584
rect 33796 17542 33824 17575
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33876 17536 33928 17542
rect 33876 17478 33928 17484
rect 33796 14278 33824 17478
rect 33888 17338 33916 17478
rect 33876 17332 33928 17338
rect 33876 17274 33928 17280
rect 33876 16516 33928 16522
rect 33876 16458 33928 16464
rect 33888 15706 33916 16458
rect 33876 15700 33928 15706
rect 33876 15642 33928 15648
rect 34256 15162 34284 26794
rect 34520 26784 34572 26790
rect 34520 26726 34572 26732
rect 34532 25906 34560 26726
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34336 24608 34388 24614
rect 34336 24550 34388 24556
rect 34348 23730 34376 24550
rect 34624 24410 34652 29446
rect 34808 29238 34836 30058
rect 35716 30048 35768 30054
rect 35716 29990 35768 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35348 28008 35400 28014
rect 35348 27950 35400 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27464 34848 27470
rect 34796 27406 34848 27412
rect 34808 26926 34836 27406
rect 34704 26920 34756 26926
rect 34704 26862 34756 26868
rect 34796 26920 34848 26926
rect 34796 26862 34848 26868
rect 34716 26382 34744 26862
rect 34808 26450 34836 26862
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26586 35388 27950
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 35532 26444 35584 26450
rect 35532 26386 35584 26392
rect 34704 26376 34756 26382
rect 34704 26318 34756 26324
rect 34808 25906 34836 26386
rect 35348 26308 35400 26314
rect 35348 26250 35400 26256
rect 35360 26042 35388 26250
rect 35348 26036 35400 26042
rect 35348 25978 35400 25984
rect 35440 25968 35492 25974
rect 35440 25910 35492 25916
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35452 25498 35480 25910
rect 35544 25770 35572 26386
rect 35532 25764 35584 25770
rect 35532 25706 35584 25712
rect 35440 25492 35492 25498
rect 35440 25434 35492 25440
rect 35728 25226 35756 29990
rect 35820 29646 35848 30670
rect 36188 30258 36216 31078
rect 36464 30938 36492 31758
rect 36648 31226 36676 32302
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 36912 31816 36964 31822
rect 36912 31758 36964 31764
rect 36556 31198 36676 31226
rect 36556 31142 36584 31198
rect 36544 31136 36596 31142
rect 36544 31078 36596 31084
rect 36452 30932 36504 30938
rect 36372 30892 36452 30920
rect 36176 30252 36228 30258
rect 36176 30194 36228 30200
rect 36372 30190 36400 30892
rect 36452 30874 36504 30880
rect 36360 30184 36412 30190
rect 36360 30126 36412 30132
rect 35900 30048 35952 30054
rect 35900 29990 35952 29996
rect 35808 29640 35860 29646
rect 35808 29582 35860 29588
rect 35912 29238 35940 29990
rect 36636 29640 36688 29646
rect 36636 29582 36688 29588
rect 36452 29504 36504 29510
rect 36452 29446 36504 29452
rect 35900 29232 35952 29238
rect 35900 29174 35952 29180
rect 36464 29170 36492 29446
rect 36084 29164 36136 29170
rect 36084 29106 36136 29112
rect 36452 29164 36504 29170
rect 36452 29106 36504 29112
rect 35898 29064 35954 29073
rect 35898 28999 35900 29008
rect 35952 28999 35954 29008
rect 35900 28970 35952 28976
rect 36096 28082 36124 29106
rect 36268 29028 36320 29034
rect 36268 28970 36320 28976
rect 36280 28218 36308 28970
rect 36648 28422 36676 29582
rect 36740 29306 36768 31758
rect 36820 31272 36872 31278
rect 36820 31214 36872 31220
rect 36832 29306 36860 31214
rect 36924 30666 36952 31758
rect 36912 30660 36964 30666
rect 36912 30602 36964 30608
rect 36924 30394 36952 30602
rect 36912 30388 36964 30394
rect 36912 30330 36964 30336
rect 37384 30122 37412 32370
rect 37740 32224 37792 32230
rect 37740 32166 37792 32172
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37476 30258 37504 31758
rect 37752 30326 37780 32166
rect 38108 31816 38160 31822
rect 38108 31758 38160 31764
rect 37924 31136 37976 31142
rect 37924 31078 37976 31084
rect 37936 30938 37964 31078
rect 37924 30932 37976 30938
rect 37924 30874 37976 30880
rect 37740 30320 37792 30326
rect 37740 30262 37792 30268
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 37648 30252 37700 30258
rect 37648 30194 37700 30200
rect 37372 30116 37424 30122
rect 37372 30058 37424 30064
rect 37476 29850 37504 30194
rect 37464 29844 37516 29850
rect 37464 29786 37516 29792
rect 37280 29708 37332 29714
rect 37280 29650 37332 29656
rect 37292 29617 37320 29650
rect 37278 29608 37334 29617
rect 37278 29543 37334 29552
rect 37660 29510 37688 30194
rect 37832 30184 37884 30190
rect 37832 30126 37884 30132
rect 37844 29753 37872 30126
rect 37830 29744 37886 29753
rect 37830 29679 37886 29688
rect 38120 29646 38148 31758
rect 38108 29640 38160 29646
rect 38108 29582 38160 29588
rect 37648 29504 37700 29510
rect 37648 29446 37700 29452
rect 36728 29300 36780 29306
rect 36728 29242 36780 29248
rect 36820 29300 36872 29306
rect 36820 29242 36872 29248
rect 37648 29096 37700 29102
rect 37648 29038 37700 29044
rect 36636 28416 36688 28422
rect 36636 28358 36688 28364
rect 36912 28416 36964 28422
rect 36912 28358 36964 28364
rect 36268 28212 36320 28218
rect 36268 28154 36320 28160
rect 36084 28076 36136 28082
rect 36084 28018 36136 28024
rect 35900 28008 35952 28014
rect 35900 27950 35952 27956
rect 35808 27872 35860 27878
rect 35808 27814 35860 27820
rect 35820 27062 35848 27814
rect 35912 27674 35940 27950
rect 35900 27668 35952 27674
rect 35900 27610 35952 27616
rect 35808 27056 35860 27062
rect 35808 26998 35860 27004
rect 36096 26994 36124 28018
rect 36648 27470 36676 28358
rect 36636 27464 36688 27470
rect 36636 27406 36688 27412
rect 36924 27402 36952 28358
rect 37372 27872 37424 27878
rect 37372 27814 37424 27820
rect 36912 27396 36964 27402
rect 36912 27338 36964 27344
rect 36636 27328 36688 27334
rect 37096 27328 37148 27334
rect 36688 27276 36768 27282
rect 36636 27270 36768 27276
rect 37096 27270 37148 27276
rect 36648 27254 36768 27270
rect 36084 26988 36136 26994
rect 36084 26930 36136 26936
rect 36096 26450 36124 26930
rect 36268 26920 36320 26926
rect 36268 26862 36320 26868
rect 36084 26444 36136 26450
rect 36084 26386 36136 26392
rect 35900 26308 35952 26314
rect 35900 26250 35952 26256
rect 35912 25294 35940 26250
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35716 25220 35768 25226
rect 35716 25162 35768 25168
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 35900 24744 35952 24750
rect 35900 24686 35952 24692
rect 34612 24404 34664 24410
rect 34612 24346 34664 24352
rect 34336 23724 34388 23730
rect 34336 23666 34388 23672
rect 34624 23186 34652 24346
rect 34716 23322 34744 24686
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 23316 34756 23322
rect 34704 23258 34756 23264
rect 34796 23316 34848 23322
rect 34796 23258 34848 23264
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34428 22092 34480 22098
rect 34428 22034 34480 22040
rect 34440 20942 34468 22034
rect 34532 21468 34560 22374
rect 34624 21865 34652 23122
rect 34808 22234 34836 23258
rect 35360 23118 35388 24550
rect 35624 24268 35676 24274
rect 35624 24210 35676 24216
rect 35636 23730 35664 24210
rect 35716 24200 35768 24206
rect 35768 24148 35848 24154
rect 35716 24142 35848 24148
rect 35728 24126 35848 24142
rect 35716 24064 35768 24070
rect 35716 24006 35768 24012
rect 35624 23724 35676 23730
rect 35624 23666 35676 23672
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35348 22772 35400 22778
rect 35348 22714 35400 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22228 34848 22234
rect 34716 22188 34796 22216
rect 34610 21856 34666 21865
rect 34610 21791 34666 21800
rect 34716 21536 34744 22188
rect 34796 22170 34848 22176
rect 35360 22030 35388 22714
rect 35544 22710 35572 22918
rect 35636 22778 35664 23666
rect 35624 22772 35676 22778
rect 35624 22714 35676 22720
rect 35532 22704 35584 22710
rect 35532 22646 35584 22652
rect 35440 22568 35492 22574
rect 35440 22510 35492 22516
rect 35452 22438 35480 22510
rect 35728 22506 35756 24006
rect 35716 22500 35768 22506
rect 35716 22442 35768 22448
rect 35440 22432 35492 22438
rect 35440 22374 35492 22380
rect 35624 22432 35676 22438
rect 35624 22374 35676 22380
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35256 22024 35308 22030
rect 35256 21966 35308 21972
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 34980 21888 35032 21894
rect 34980 21830 35032 21836
rect 34796 21548 34848 21554
rect 34716 21508 34796 21536
rect 34796 21490 34848 21496
rect 34992 21486 35020 21830
rect 34612 21480 34664 21486
rect 34532 21440 34612 21468
rect 34612 21422 34664 21428
rect 34980 21480 35032 21486
rect 34980 21422 35032 21428
rect 35268 21418 35296 21966
rect 35452 21554 35480 22170
rect 35530 21856 35586 21865
rect 35530 21791 35586 21800
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35256 21412 35308 21418
rect 35256 21354 35308 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34612 21140 34664 21146
rect 34612 21082 34664 21088
rect 34428 20936 34480 20942
rect 34428 20878 34480 20884
rect 34624 20466 34652 21082
rect 34704 20868 34756 20874
rect 34704 20810 34756 20816
rect 34716 20602 34744 20810
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 34612 20460 34664 20466
rect 34612 20402 34664 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34888 19848 34940 19854
rect 34888 19790 34940 19796
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34716 19514 34744 19654
rect 34900 19514 34928 19790
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34888 19508 34940 19514
rect 34888 19450 34940 19456
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 34612 19168 34664 19174
rect 34612 19110 34664 19116
rect 34624 18630 34652 19110
rect 34612 18624 34664 18630
rect 34612 18566 34664 18572
rect 34336 15904 34388 15910
rect 34336 15846 34388 15852
rect 34348 15706 34376 15846
rect 34336 15700 34388 15706
rect 34336 15642 34388 15648
rect 34244 15156 34296 15162
rect 34244 15098 34296 15104
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 33876 15020 33928 15026
rect 33876 14962 33928 14968
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33784 13184 33836 13190
rect 33784 13126 33836 13132
rect 33692 12912 33744 12918
rect 33692 12854 33744 12860
rect 33796 12238 33824 13126
rect 33784 12232 33836 12238
rect 33784 12174 33836 12180
rect 33508 11756 33560 11762
rect 33508 11698 33560 11704
rect 33414 11656 33470 11665
rect 33414 11591 33470 11600
rect 33520 11354 33548 11698
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 33508 11348 33560 11354
rect 33508 11290 33560 11296
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32968 10742 32996 11018
rect 33048 11008 33100 11014
rect 33048 10950 33100 10956
rect 33060 10810 33088 10950
rect 33048 10804 33100 10810
rect 33048 10746 33100 10752
rect 32956 10736 33008 10742
rect 32956 10678 33008 10684
rect 33048 10532 33100 10538
rect 33048 10474 33100 10480
rect 33060 10130 33088 10474
rect 33796 10130 33824 12174
rect 33048 10124 33100 10130
rect 33048 10066 33100 10072
rect 33784 10124 33836 10130
rect 33784 10066 33836 10072
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 33048 9580 33100 9586
rect 33048 9522 33100 9528
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32772 8968 32824 8974
rect 32772 8910 32824 8916
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 32692 8634 32720 8774
rect 32784 8634 32812 8910
rect 32968 8634 32996 9318
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32956 8628 33008 8634
rect 32956 8570 33008 8576
rect 33060 8566 33088 9522
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 33060 8430 33088 8502
rect 33336 8430 33364 9318
rect 32588 8424 32640 8430
rect 32588 8366 32640 8372
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 33324 8424 33376 8430
rect 33324 8366 33376 8372
rect 32600 8090 32628 8366
rect 32680 8288 32732 8294
rect 32680 8230 32732 8236
rect 32588 8084 32640 8090
rect 32588 8026 32640 8032
rect 32496 7744 32548 7750
rect 32496 7686 32548 7692
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32416 6322 32444 6734
rect 32312 6316 32364 6322
rect 32312 6258 32364 6264
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 32128 6112 32180 6118
rect 32128 6054 32180 6060
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 32048 5409 32076 6054
rect 32140 5574 32168 6054
rect 32218 5672 32274 5681
rect 32218 5607 32274 5616
rect 32232 5574 32260 5607
rect 32128 5568 32180 5574
rect 32128 5510 32180 5516
rect 32220 5568 32272 5574
rect 32220 5510 32272 5516
rect 32034 5400 32090 5409
rect 32034 5335 32090 5344
rect 31850 5264 31906 5273
rect 32218 5264 32274 5273
rect 31850 5199 31906 5208
rect 31944 5228 31996 5234
rect 31944 5170 31996 5176
rect 32036 5228 32088 5234
rect 32218 5199 32274 5208
rect 32036 5170 32088 5176
rect 31852 5024 31904 5030
rect 31852 4966 31904 4972
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 31668 3596 31720 3602
rect 31668 3538 31720 3544
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 30472 3460 30524 3466
rect 30472 3402 30524 3408
rect 30656 3460 30708 3466
rect 30656 3402 30708 3408
rect 30668 3126 30696 3402
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 30656 3120 30708 3126
rect 30656 3062 30708 3068
rect 30472 2984 30524 2990
rect 30472 2926 30524 2932
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30484 800 30512 2926
rect 30852 800 30880 3130
rect 31404 3126 31432 3470
rect 31392 3120 31444 3126
rect 31392 3062 31444 3068
rect 31864 3058 31892 4966
rect 31956 3942 31984 5170
rect 32048 5137 32076 5170
rect 32232 5166 32260 5199
rect 32220 5160 32272 5166
rect 32034 5128 32090 5137
rect 32220 5102 32272 5108
rect 32034 5063 32090 5072
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 32232 4826 32260 4966
rect 32220 4820 32272 4826
rect 32220 4762 32272 4768
rect 32128 4480 32180 4486
rect 32128 4422 32180 4428
rect 32140 4282 32168 4422
rect 32036 4276 32088 4282
rect 32036 4218 32088 4224
rect 32128 4276 32180 4282
rect 32128 4218 32180 4224
rect 31944 3936 31996 3942
rect 31944 3878 31996 3884
rect 32048 3738 32076 4218
rect 32220 4072 32272 4078
rect 32140 4032 32220 4060
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 31944 3664 31996 3670
rect 31944 3606 31996 3612
rect 31956 3126 31984 3606
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 31944 3120 31996 3126
rect 31944 3062 31996 3068
rect 31852 3052 31904 3058
rect 31852 2994 31904 3000
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31220 800 31248 2926
rect 32048 2854 32076 3470
rect 32036 2848 32088 2854
rect 31942 2816 31998 2825
rect 32036 2790 32088 2796
rect 31942 2751 31998 2760
rect 32140 2774 32168 4032
rect 32220 4014 32272 4020
rect 32218 3632 32274 3641
rect 32218 3567 32274 3576
rect 32232 2922 32260 3567
rect 32324 3233 32352 6258
rect 32404 6180 32456 6186
rect 32404 6122 32456 6128
rect 32416 4146 32444 6122
rect 32508 5370 32536 7686
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 32496 5364 32548 5370
rect 32496 5306 32548 5312
rect 32600 5234 32628 7482
rect 32692 7410 32720 8230
rect 33888 8090 33916 14962
rect 34336 13252 34388 13258
rect 34336 13194 34388 13200
rect 34244 12708 34296 12714
rect 34244 12650 34296 12656
rect 34256 11286 34284 12650
rect 34244 11280 34296 11286
rect 34244 11222 34296 11228
rect 33968 11212 34020 11218
rect 33968 11154 34020 11160
rect 33980 11121 34008 11154
rect 33966 11112 34022 11121
rect 33966 11047 34022 11056
rect 33980 10810 34008 11047
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 34348 10198 34376 13194
rect 34336 10192 34388 10198
rect 34336 10134 34388 10140
rect 34348 9654 34376 10134
rect 34336 9648 34388 9654
rect 34336 9590 34388 9596
rect 34348 9178 34376 9590
rect 34336 9172 34388 9178
rect 34336 9114 34388 9120
rect 33968 8968 34020 8974
rect 33968 8910 34020 8916
rect 33980 8634 34008 8910
rect 34152 8832 34204 8838
rect 34152 8774 34204 8780
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34060 8356 34112 8362
rect 34060 8298 34112 8304
rect 34164 8344 34192 8774
rect 34440 8634 34468 15098
rect 34520 14816 34572 14822
rect 34520 14758 34572 14764
rect 34532 13938 34560 14758
rect 34624 13977 34652 18566
rect 34716 17542 34744 19314
rect 35360 19174 35388 19790
rect 35440 19712 35492 19718
rect 35440 19654 35492 19660
rect 35452 19514 35480 19654
rect 35440 19508 35492 19514
rect 35440 19450 35492 19456
rect 35348 19168 35400 19174
rect 35348 19110 35400 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18970 35388 19110
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 35440 18964 35492 18970
rect 35440 18906 35492 18912
rect 35452 18426 35480 18906
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35256 17740 35308 17746
rect 35176 17700 35256 17728
rect 34980 17604 35032 17610
rect 35176 17592 35204 17700
rect 35256 17682 35308 17688
rect 35348 17740 35400 17746
rect 35544 17728 35572 21791
rect 35636 19334 35664 22374
rect 35820 22094 35848 24126
rect 35912 23526 35940 24686
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35912 23186 35940 23462
rect 35992 23248 36044 23254
rect 35992 23190 36044 23196
rect 35900 23180 35952 23186
rect 35900 23122 35952 23128
rect 36004 22642 36032 23190
rect 35992 22636 36044 22642
rect 35992 22578 36044 22584
rect 35820 22066 35940 22094
rect 35912 21962 35940 22066
rect 35992 22092 36044 22098
rect 35992 22034 36044 22040
rect 35900 21956 35952 21962
rect 35900 21898 35952 21904
rect 35808 21140 35860 21146
rect 35808 21082 35860 21088
rect 35636 19306 35756 19334
rect 35624 18828 35676 18834
rect 35624 18770 35676 18776
rect 35636 18358 35664 18770
rect 35624 18352 35676 18358
rect 35624 18294 35676 18300
rect 35400 17700 35572 17728
rect 35348 17682 35400 17688
rect 35032 17564 35204 17592
rect 35254 17640 35310 17649
rect 35360 17626 35388 17682
rect 35310 17598 35388 17626
rect 35254 17575 35310 17584
rect 34980 17546 35032 17552
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 34716 16250 34744 17478
rect 35256 17264 35308 17270
rect 35308 17212 35388 17218
rect 35256 17206 35388 17212
rect 35268 17190 35388 17206
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16454 35388 17190
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 35624 17128 35676 17134
rect 35624 17070 35676 17076
rect 35452 16590 35480 17070
rect 35440 16584 35492 16590
rect 35440 16526 35492 16532
rect 35636 16522 35664 17070
rect 35624 16516 35676 16522
rect 35624 16458 35676 16464
rect 35348 16448 35400 16454
rect 35348 16390 35400 16396
rect 34704 16244 34756 16250
rect 34704 16186 34756 16192
rect 35360 16114 35388 16390
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34808 15706 34836 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35636 15706 35664 16458
rect 35728 16046 35756 19306
rect 35820 18970 35848 21082
rect 36004 20534 36032 22034
rect 35992 20528 36044 20534
rect 35992 20470 36044 20476
rect 36096 19334 36124 26386
rect 36176 24200 36228 24206
rect 36176 24142 36228 24148
rect 36188 21894 36216 24142
rect 36280 22166 36308 26862
rect 36544 26784 36596 26790
rect 36544 26726 36596 26732
rect 36452 26444 36504 26450
rect 36556 26432 36584 26726
rect 36504 26404 36584 26432
rect 36452 26386 36504 26392
rect 36360 24608 36412 24614
rect 36360 24550 36412 24556
rect 36372 22574 36400 24550
rect 36464 23526 36492 26386
rect 36740 26382 36768 27254
rect 37108 26450 37136 27270
rect 37280 26784 37332 26790
rect 37280 26726 37332 26732
rect 37292 26518 37320 26726
rect 37280 26512 37332 26518
rect 37280 26454 37332 26460
rect 37004 26444 37056 26450
rect 37004 26386 37056 26392
rect 37096 26444 37148 26450
rect 37096 26386 37148 26392
rect 36728 26376 36780 26382
rect 36728 26318 36780 26324
rect 37016 25906 37044 26386
rect 36820 25900 36872 25906
rect 36820 25842 36872 25848
rect 37004 25900 37056 25906
rect 37004 25842 37056 25848
rect 36636 24064 36688 24070
rect 36636 24006 36688 24012
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 36452 23520 36504 23526
rect 36452 23462 36504 23468
rect 36464 23322 36492 23462
rect 36452 23316 36504 23322
rect 36452 23258 36504 23264
rect 36464 23118 36492 23258
rect 36452 23112 36504 23118
rect 36452 23054 36504 23060
rect 36556 22778 36584 23598
rect 36648 22778 36676 24006
rect 36832 23338 36860 25842
rect 37108 25430 37136 26386
rect 37188 26240 37240 26246
rect 37188 26182 37240 26188
rect 37200 25498 37228 26182
rect 37384 25974 37412 27814
rect 37660 26450 37688 29038
rect 37924 28552 37976 28558
rect 37924 28494 37976 28500
rect 37740 28144 37792 28150
rect 37740 28086 37792 28092
rect 37752 27062 37780 28086
rect 37936 27130 37964 28494
rect 38016 27396 38068 27402
rect 38016 27338 38068 27344
rect 37924 27124 37976 27130
rect 37924 27066 37976 27072
rect 37740 27056 37792 27062
rect 37740 26998 37792 27004
rect 37924 26988 37976 26994
rect 37924 26930 37976 26936
rect 37648 26444 37700 26450
rect 37648 26386 37700 26392
rect 37372 25968 37424 25974
rect 37372 25910 37424 25916
rect 37660 25838 37688 26386
rect 37936 26382 37964 26930
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 37924 26376 37976 26382
rect 37924 26318 37976 26324
rect 37740 26240 37792 26246
rect 37740 26182 37792 26188
rect 37648 25832 37700 25838
rect 37648 25774 37700 25780
rect 37188 25492 37240 25498
rect 37188 25434 37240 25440
rect 37096 25424 37148 25430
rect 37096 25366 37148 25372
rect 37752 25362 37780 26182
rect 37844 25906 37872 26318
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 38028 25498 38056 27338
rect 38200 26444 38252 26450
rect 38200 26386 38252 26392
rect 38212 26042 38240 26386
rect 38200 26036 38252 26042
rect 38200 25978 38252 25984
rect 38016 25492 38068 25498
rect 38016 25434 38068 25440
rect 37740 25356 37792 25362
rect 37740 25298 37792 25304
rect 38292 25152 38344 25158
rect 38292 25094 38344 25100
rect 37004 24744 37056 24750
rect 37004 24686 37056 24692
rect 37096 24744 37148 24750
rect 37096 24686 37148 24692
rect 36912 24608 36964 24614
rect 36912 24550 36964 24556
rect 36924 24206 36952 24550
rect 36912 24200 36964 24206
rect 36912 24142 36964 24148
rect 37016 23866 37044 24686
rect 37004 23860 37056 23866
rect 37004 23802 37056 23808
rect 36832 23310 36952 23338
rect 37016 23322 37044 23802
rect 36924 23202 36952 23310
rect 37004 23316 37056 23322
rect 37004 23258 37056 23264
rect 36924 23186 37044 23202
rect 36924 23180 37056 23186
rect 36924 23174 37004 23180
rect 37004 23122 37056 23128
rect 36912 22976 36964 22982
rect 36912 22918 36964 22924
rect 36544 22772 36596 22778
rect 36544 22714 36596 22720
rect 36636 22772 36688 22778
rect 36636 22714 36688 22720
rect 36924 22710 36952 22918
rect 37108 22778 37136 24686
rect 37740 24404 37792 24410
rect 37740 24346 37792 24352
rect 37186 23760 37242 23769
rect 37186 23695 37242 23704
rect 37200 23474 37228 23695
rect 37200 23446 37320 23474
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 37096 22772 37148 22778
rect 37096 22714 37148 22720
rect 36452 22704 36504 22710
rect 36452 22646 36504 22652
rect 36912 22704 36964 22710
rect 36912 22646 36964 22652
rect 36360 22568 36412 22574
rect 36360 22510 36412 22516
rect 36268 22160 36320 22166
rect 36268 22102 36320 22108
rect 36360 22024 36412 22030
rect 36360 21966 36412 21972
rect 36176 21888 36228 21894
rect 36176 21830 36228 21836
rect 36372 21146 36400 21966
rect 36464 21962 36492 22646
rect 36728 22568 36780 22574
rect 36728 22510 36780 22516
rect 36452 21956 36504 21962
rect 36452 21898 36504 21904
rect 36740 21146 36768 22510
rect 37200 22030 37228 22918
rect 37292 22574 37320 23446
rect 37752 23186 37780 24346
rect 37740 23180 37792 23186
rect 37740 23122 37792 23128
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 37280 22568 37332 22574
rect 37280 22510 37332 22516
rect 37188 22024 37240 22030
rect 37188 21966 37240 21972
rect 37292 21146 37320 22510
rect 37476 22234 37504 23054
rect 37556 22704 37608 22710
rect 37556 22646 37608 22652
rect 37464 22228 37516 22234
rect 37464 22170 37516 22176
rect 37568 21690 37596 22646
rect 37648 22636 37700 22642
rect 37648 22578 37700 22584
rect 37660 22234 37688 22578
rect 37740 22568 37792 22574
rect 37740 22510 37792 22516
rect 37648 22228 37700 22234
rect 37648 22170 37700 22176
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 37464 21480 37516 21486
rect 37464 21422 37516 21428
rect 36360 21140 36412 21146
rect 36360 21082 36412 21088
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 37280 21140 37332 21146
rect 37280 21082 37332 21088
rect 36452 19848 36504 19854
rect 36452 19790 36504 19796
rect 36176 19712 36228 19718
rect 36176 19654 36228 19660
rect 36188 19514 36216 19654
rect 36176 19508 36228 19514
rect 36176 19450 36228 19456
rect 35992 19304 36044 19310
rect 36096 19306 36400 19334
rect 35992 19246 36044 19252
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 35808 18964 35860 18970
rect 35808 18906 35860 18912
rect 35912 18834 35940 19110
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 36004 17626 36032 19246
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 36096 18086 36124 18702
rect 36176 18352 36228 18358
rect 36176 18294 36228 18300
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 36188 17678 36216 18294
rect 35912 17598 36032 17626
rect 36176 17672 36228 17678
rect 36176 17614 36228 17620
rect 36084 17604 36136 17610
rect 35716 16040 35768 16046
rect 35716 15982 35768 15988
rect 35728 15706 35756 15982
rect 34796 15700 34848 15706
rect 34796 15642 34848 15648
rect 35624 15700 35676 15706
rect 35624 15642 35676 15648
rect 35716 15700 35768 15706
rect 35716 15642 35768 15648
rect 35912 15065 35940 17598
rect 36084 17546 36136 17552
rect 36096 17490 36124 17546
rect 36004 17462 36124 17490
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 36004 16250 36032 17462
rect 36084 17332 36136 17338
rect 36084 17274 36136 17280
rect 36096 17202 36124 17274
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36176 16652 36228 16658
rect 36176 16594 36228 16600
rect 36084 16516 36136 16522
rect 36084 16458 36136 16464
rect 36096 16250 36124 16458
rect 35992 16244 36044 16250
rect 35992 16186 36044 16192
rect 36084 16244 36136 16250
rect 36084 16186 36136 16192
rect 35898 15056 35954 15065
rect 35898 14991 35954 15000
rect 34796 14952 34848 14958
rect 34796 14894 34848 14900
rect 35900 14952 35952 14958
rect 35900 14894 35952 14900
rect 34808 14618 34836 14894
rect 35348 14816 35400 14822
rect 35348 14758 35400 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14618 35388 14758
rect 34796 14612 34848 14618
rect 34796 14554 34848 14560
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 35912 14074 35940 14894
rect 36188 14414 36216 16594
rect 36280 16114 36308 17478
rect 36268 16108 36320 16114
rect 36268 16050 36320 16056
rect 36372 15706 36400 19306
rect 36464 18086 36492 19790
rect 36544 19440 36596 19446
rect 36544 19382 36596 19388
rect 36556 18358 36584 19382
rect 36740 19334 36768 21082
rect 37292 20754 37320 21082
rect 37476 21078 37504 21422
rect 37464 21072 37516 21078
rect 37462 21040 37464 21049
rect 37516 21040 37518 21049
rect 37462 20975 37518 20984
rect 37200 20726 37320 20754
rect 36820 19848 36872 19854
rect 36820 19790 36872 19796
rect 36648 19306 36768 19334
rect 36544 18352 36596 18358
rect 36544 18294 36596 18300
rect 36452 18080 36504 18086
rect 36452 18022 36504 18028
rect 36544 17740 36596 17746
rect 36648 17728 36676 19306
rect 36832 18902 36860 19790
rect 36820 18896 36872 18902
rect 36820 18838 36872 18844
rect 36728 18828 36780 18834
rect 36728 18770 36780 18776
rect 36740 18086 36768 18770
rect 36832 18426 36860 18838
rect 36820 18420 36872 18426
rect 36820 18362 36872 18368
rect 36728 18080 36780 18086
rect 36728 18022 36780 18028
rect 36596 17700 36676 17728
rect 36544 17682 36596 17688
rect 36452 17672 36504 17678
rect 36452 17614 36504 17620
rect 36464 17134 36492 17614
rect 36452 17128 36504 17134
rect 36452 17070 36504 17076
rect 36740 16998 36768 18022
rect 36912 17672 36964 17678
rect 36912 17614 36964 17620
rect 36924 17338 36952 17614
rect 36912 17332 36964 17338
rect 36912 17274 36964 17280
rect 36728 16992 36780 16998
rect 36728 16934 36780 16940
rect 37200 16250 37228 20726
rect 37752 18714 37780 22510
rect 38016 21344 38068 21350
rect 38016 21286 38068 21292
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 37372 18692 37424 18698
rect 37372 18634 37424 18640
rect 37476 18686 37780 18714
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37292 17746 37320 18022
rect 37384 17882 37412 18634
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37188 16244 37240 16250
rect 37188 16186 37240 16192
rect 37372 16040 37424 16046
rect 37372 15982 37424 15988
rect 36360 15700 36412 15706
rect 36360 15642 36412 15648
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 35900 14068 35952 14074
rect 35900 14010 35952 14016
rect 34610 13968 34666 13977
rect 34520 13932 34572 13938
rect 35912 13954 35940 14010
rect 35912 13938 36032 13954
rect 35912 13932 36044 13938
rect 35912 13926 35992 13932
rect 34610 13903 34666 13912
rect 34520 13874 34572 13880
rect 35992 13874 36044 13880
rect 34796 13864 34848 13870
rect 34796 13806 34848 13812
rect 34808 13394 34836 13806
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 36188 13530 36216 14350
rect 36360 13864 36412 13870
rect 36360 13806 36412 13812
rect 36176 13524 36228 13530
rect 36176 13466 36228 13472
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34520 12912 34572 12918
rect 34518 12880 34520 12889
rect 34572 12880 34574 12889
rect 34808 12850 34836 13330
rect 36372 12986 36400 13806
rect 36360 12980 36412 12986
rect 36360 12922 36412 12928
rect 34518 12815 34574 12824
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34532 11218 34560 12038
rect 34808 11694 34836 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 36372 12322 36400 12922
rect 36464 12424 36492 15370
rect 37384 15162 37412 15982
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 36544 14952 36596 14958
rect 36544 14894 36596 14900
rect 36556 14618 36584 14894
rect 37188 14816 37240 14822
rect 37188 14758 37240 14764
rect 37280 14816 37332 14822
rect 37280 14758 37332 14764
rect 36544 14612 36596 14618
rect 36544 14554 36596 14560
rect 36556 14074 36584 14554
rect 37200 14074 37228 14758
rect 37292 14618 37320 14758
rect 37384 14618 37412 15098
rect 37280 14612 37332 14618
rect 37280 14554 37332 14560
rect 37372 14612 37424 14618
rect 37372 14554 37424 14560
rect 37372 14272 37424 14278
rect 37372 14214 37424 14220
rect 36544 14068 36596 14074
rect 36544 14010 36596 14016
rect 37188 14068 37240 14074
rect 37188 14010 37240 14016
rect 37004 13796 37056 13802
rect 37004 13738 37056 13744
rect 37016 13190 37044 13738
rect 37280 13252 37332 13258
rect 37280 13194 37332 13200
rect 37004 13184 37056 13190
rect 37004 13126 37056 13132
rect 36728 12776 36780 12782
rect 36728 12718 36780 12724
rect 36740 12442 36768 12718
rect 36728 12436 36780 12442
rect 36464 12396 36575 12424
rect 36547 12356 36575 12396
rect 36728 12378 36780 12384
rect 36547 12328 36584 12356
rect 36372 12306 36492 12322
rect 36372 12300 36504 12306
rect 36372 12294 36452 12300
rect 36452 12242 36504 12248
rect 36084 12096 36136 12102
rect 36084 12038 36136 12044
rect 34704 11688 34756 11694
rect 34704 11630 34756 11636
rect 34796 11688 34848 11694
rect 34796 11630 34848 11636
rect 35532 11688 35584 11694
rect 35532 11630 35584 11636
rect 34716 11354 34744 11630
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34532 10674 34560 11154
rect 35360 10742 35388 11494
rect 35348 10736 35400 10742
rect 35348 10678 35400 10684
rect 35544 10674 35572 11630
rect 35716 11280 35768 11286
rect 35716 11222 35768 11228
rect 34520 10668 34572 10674
rect 34520 10610 34572 10616
rect 35532 10668 35584 10674
rect 35532 10610 35584 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34532 9382 34560 9998
rect 35348 9988 35400 9994
rect 35348 9930 35400 9936
rect 34520 9376 34572 9382
rect 34520 9318 34572 9324
rect 34532 9042 34560 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 9178 35388 9930
rect 35348 9172 35400 9178
rect 35348 9114 35400 9120
rect 34520 9036 34572 9042
rect 34520 8978 34572 8984
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34532 8498 34560 8978
rect 34336 8492 34388 8498
rect 34336 8434 34388 8440
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34244 8356 34296 8362
rect 34164 8316 34244 8344
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 33968 6996 34020 7002
rect 33968 6938 34020 6944
rect 33232 6792 33284 6798
rect 33232 6734 33284 6740
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33060 6458 33088 6598
rect 33048 6452 33100 6458
rect 33048 6394 33100 6400
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 32680 6248 32732 6254
rect 32680 6190 32732 6196
rect 32496 5228 32548 5234
rect 32496 5170 32548 5176
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 32508 4826 32536 5170
rect 32600 5030 32628 5170
rect 32588 5024 32640 5030
rect 32588 4966 32640 4972
rect 32692 4826 32720 6190
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32496 4820 32548 4826
rect 32496 4762 32548 4768
rect 32680 4820 32732 4826
rect 32680 4762 32732 4768
rect 32588 4548 32640 4554
rect 32588 4490 32640 4496
rect 32404 4140 32456 4146
rect 32404 4082 32456 4088
rect 32310 3224 32366 3233
rect 32310 3159 32366 3168
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 32220 2916 32272 2922
rect 32220 2858 32272 2864
rect 31956 2446 31984 2751
rect 32140 2746 32260 2774
rect 31944 2440 31996 2446
rect 31588 2378 31708 2394
rect 31944 2382 31996 2388
rect 31588 2372 31720 2378
rect 31588 2366 31668 2372
rect 31588 800 31616 2366
rect 31668 2314 31720 2320
rect 31956 870 32076 898
rect 31956 800 31984 870
rect 29840 734 30052 762
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32048 762 32076 870
rect 32232 762 32260 2746
rect 32324 800 32352 3062
rect 32600 2854 32628 4490
rect 32678 4176 32734 4185
rect 32678 4111 32680 4120
rect 32732 4111 32734 4120
rect 32680 4082 32732 4088
rect 32784 3369 32812 5646
rect 32864 5636 32916 5642
rect 32864 5578 32916 5584
rect 32876 5370 32904 5578
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32864 5092 32916 5098
rect 32864 5034 32916 5040
rect 32876 4690 32904 5034
rect 32956 5024 33008 5030
rect 32956 4966 33008 4972
rect 33048 5024 33100 5030
rect 33048 4966 33100 4972
rect 32968 4826 32996 4966
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 32876 4282 32904 4626
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 33060 3738 33088 4966
rect 33048 3732 33100 3738
rect 33048 3674 33100 3680
rect 32956 3596 33008 3602
rect 33008 3556 33088 3584
rect 32956 3538 33008 3544
rect 32770 3360 32826 3369
rect 32770 3295 32826 3304
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 32588 2848 32640 2854
rect 32588 2790 32640 2796
rect 32968 2774 32996 2926
rect 32876 2746 32996 2774
rect 32876 1578 32904 2746
rect 32692 1550 32904 1578
rect 32692 800 32720 1550
rect 33060 800 33088 3556
rect 33152 2650 33180 6258
rect 33244 5846 33272 6734
rect 33508 6724 33560 6730
rect 33508 6666 33560 6672
rect 33416 6180 33468 6186
rect 33416 6122 33468 6128
rect 33232 5840 33284 5846
rect 33428 5817 33456 6122
rect 33232 5782 33284 5788
rect 33414 5808 33470 5817
rect 33414 5743 33470 5752
rect 33428 5370 33456 5743
rect 33416 5364 33468 5370
rect 33416 5306 33468 5312
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33336 4690 33364 5170
rect 33520 4690 33548 6666
rect 33874 5536 33930 5545
rect 33874 5471 33930 5480
rect 33888 5234 33916 5471
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 33232 4684 33284 4690
rect 33232 4626 33284 4632
rect 33324 4684 33376 4690
rect 33324 4626 33376 4632
rect 33508 4684 33560 4690
rect 33508 4626 33560 4632
rect 33600 4684 33652 4690
rect 33600 4626 33652 4632
rect 33244 4457 33272 4626
rect 33416 4616 33468 4622
rect 33416 4558 33468 4564
rect 33230 4448 33286 4457
rect 33230 4383 33286 4392
rect 33428 4282 33456 4558
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33612 4185 33640 4626
rect 33598 4176 33654 4185
rect 33598 4111 33654 4120
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 33244 3602 33272 3878
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33428 800 33456 2790
rect 33612 1766 33640 3402
rect 33704 2650 33732 4762
rect 33874 4720 33930 4729
rect 33874 4655 33876 4664
rect 33928 4655 33930 4664
rect 33876 4626 33928 4632
rect 33980 4622 34008 6938
rect 34072 6798 34100 8298
rect 34164 7954 34192 8316
rect 34244 8298 34296 8304
rect 34152 7948 34204 7954
rect 34152 7890 34204 7896
rect 34244 7880 34296 7886
rect 34244 7822 34296 7828
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 34164 7546 34192 7686
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 34256 6662 34284 7822
rect 34060 6656 34112 6662
rect 34060 6598 34112 6604
rect 34244 6656 34296 6662
rect 34244 6598 34296 6604
rect 34072 4690 34100 6598
rect 34348 6458 34376 8434
rect 34532 7954 34560 8434
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34440 7410 34468 7822
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34532 7410 34560 7686
rect 34428 7404 34480 7410
rect 34428 7346 34480 7352
rect 34520 7404 34572 7410
rect 34520 7346 34572 7352
rect 34716 6458 34744 8434
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35164 7812 35216 7818
rect 35164 7754 35216 7760
rect 35176 7546 35204 7754
rect 35164 7540 35216 7546
rect 35164 7482 35216 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35532 6860 35584 6866
rect 35532 6802 35584 6808
rect 35164 6792 35216 6798
rect 35544 6769 35572 6802
rect 35164 6734 35216 6740
rect 35530 6760 35586 6769
rect 34796 6724 34848 6730
rect 34796 6666 34848 6672
rect 34336 6452 34388 6458
rect 34336 6394 34388 6400
rect 34704 6452 34756 6458
rect 34704 6394 34756 6400
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 34152 6112 34204 6118
rect 34152 6054 34204 6060
rect 34164 5370 34192 6054
rect 34242 5808 34298 5817
rect 34532 5778 34560 6258
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 34520 5772 34572 5778
rect 34298 5752 34376 5760
rect 34242 5743 34244 5752
rect 34296 5732 34376 5752
rect 34244 5714 34296 5720
rect 34244 5568 34296 5574
rect 34244 5510 34296 5516
rect 34152 5364 34204 5370
rect 34152 5306 34204 5312
rect 34256 5234 34284 5510
rect 34244 5228 34296 5234
rect 34244 5170 34296 5176
rect 34060 4684 34112 4690
rect 34060 4626 34112 4632
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 34256 4214 34284 5170
rect 34348 4690 34376 5732
rect 34520 5714 34572 5720
rect 34428 5636 34480 5642
rect 34428 5578 34480 5584
rect 34336 4684 34388 4690
rect 34336 4626 34388 4632
rect 34336 4480 34388 4486
rect 34336 4422 34388 4428
rect 34244 4208 34296 4214
rect 34244 4150 34296 4156
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 34058 3224 34114 3233
rect 34058 3159 34114 3168
rect 34072 3058 34100 3159
rect 34060 3052 34112 3058
rect 34060 2994 34112 3000
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 34060 2508 34112 2514
rect 34060 2450 34112 2456
rect 33600 1760 33652 1766
rect 33600 1702 33652 1708
rect 33796 870 33916 898
rect 33796 800 33824 870
rect 32048 734 32260 762
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 33888 762 33916 870
rect 34072 762 34100 2450
rect 34164 2446 34192 3334
rect 34348 3058 34376 4422
rect 34440 4146 34468 5578
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34532 4162 34560 5510
rect 34624 4622 34652 6054
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34428 4140 34480 4146
rect 34532 4134 34652 4162
rect 34428 4082 34480 4088
rect 34426 4040 34482 4049
rect 34426 3975 34482 3984
rect 34440 3534 34468 3975
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 34532 2446 34560 3130
rect 34624 2446 34652 4134
rect 34716 3738 34744 6190
rect 34808 5794 34836 6666
rect 34980 6656 35032 6662
rect 34980 6598 35032 6604
rect 34992 6458 35020 6598
rect 34980 6452 35032 6458
rect 34980 6394 35032 6400
rect 35176 6338 35204 6734
rect 35530 6695 35586 6704
rect 35176 6310 35480 6338
rect 35256 6180 35308 6186
rect 35256 6122 35308 6128
rect 35268 6066 35296 6122
rect 35268 6038 35388 6066
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34808 5766 34928 5794
rect 34796 5704 34848 5710
rect 34796 5646 34848 5652
rect 34808 4826 34836 5646
rect 34900 5030 34928 5766
rect 34888 5024 34940 5030
rect 34888 4966 34940 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 4820 34848 4826
rect 35360 4808 35388 6038
rect 34796 4762 34848 4768
rect 34992 4780 35388 4808
rect 34886 4720 34942 4729
rect 34886 4655 34942 4664
rect 34900 4622 34928 4655
rect 34888 4616 34940 4622
rect 34888 4558 34940 4564
rect 34992 3992 35020 4780
rect 35164 4684 35216 4690
rect 35164 4626 35216 4632
rect 35176 4060 35204 4626
rect 35176 4032 35388 4060
rect 34808 3964 35020 3992
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34808 3618 34836 3964
rect 35360 3913 35388 4032
rect 35346 3904 35402 3913
rect 34934 3836 35242 3845
rect 35346 3839 35402 3848
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35348 3732 35400 3738
rect 35348 3674 35400 3680
rect 34716 3590 34836 3618
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34428 2372 34480 2378
rect 34428 2314 34480 2320
rect 34164 870 34284 898
rect 34164 800 34192 870
rect 33888 734 34100 762
rect 34150 0 34206 800
rect 34256 762 34284 870
rect 34440 762 34468 2314
rect 34716 2258 34744 3590
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 35176 3194 35204 3334
rect 35164 3188 35216 3194
rect 35164 3130 35216 3136
rect 34796 2984 34848 2990
rect 34796 2926 34848 2932
rect 34532 2230 34744 2258
rect 34532 800 34560 2230
rect 34808 1578 34836 2926
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1850 35388 3674
rect 35452 3670 35480 6310
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35532 5636 35584 5642
rect 35532 5578 35584 5584
rect 35544 4026 35572 5578
rect 35636 4146 35664 6258
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 35544 3998 35664 4026
rect 35440 3664 35492 3670
rect 35440 3606 35492 3612
rect 35532 3596 35584 3602
rect 35532 3538 35584 3544
rect 35544 2650 35572 3538
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 35268 1822 35388 1850
rect 34808 1550 34928 1578
rect 34900 800 34928 1550
rect 35268 800 35296 1822
rect 35636 800 35664 3998
rect 35728 3534 35756 11222
rect 36096 11014 36124 12038
rect 36360 11144 36412 11150
rect 36358 11112 36360 11121
rect 36452 11144 36504 11150
rect 36412 11112 36414 11121
rect 36452 11086 36504 11092
rect 36358 11047 36414 11056
rect 36084 11008 36136 11014
rect 36084 10950 36136 10956
rect 36096 10810 36124 10950
rect 36084 10804 36136 10810
rect 36084 10746 36136 10752
rect 36176 10600 36228 10606
rect 36176 10542 36228 10548
rect 36268 10600 36320 10606
rect 36268 10542 36320 10548
rect 35900 10464 35952 10470
rect 35900 10406 35952 10412
rect 35912 9042 35940 10406
rect 36188 9722 36216 10542
rect 36280 10266 36308 10542
rect 36268 10260 36320 10266
rect 36268 10202 36320 10208
rect 36464 9926 36492 11086
rect 36452 9920 36504 9926
rect 36452 9862 36504 9868
rect 36176 9716 36228 9722
rect 36176 9658 36228 9664
rect 36084 9648 36136 9654
rect 36084 9590 36136 9596
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 35900 8832 35952 8838
rect 35900 8774 35952 8780
rect 35808 7200 35860 7206
rect 35808 7142 35860 7148
rect 35820 5778 35848 7142
rect 35912 6866 35940 8774
rect 35992 8560 36044 8566
rect 35992 8502 36044 8508
rect 35900 6860 35952 6866
rect 35900 6802 35952 6808
rect 36004 6662 36032 8502
rect 36096 8430 36124 9590
rect 36176 8628 36228 8634
rect 36176 8570 36228 8576
rect 36084 8424 36136 8430
rect 36084 8366 36136 8372
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36096 7410 36124 8026
rect 36188 7410 36216 8570
rect 36452 8492 36504 8498
rect 36452 8434 36504 8440
rect 36268 7540 36320 7546
rect 36268 7482 36320 7488
rect 36084 7404 36136 7410
rect 36084 7346 36136 7352
rect 36176 7404 36228 7410
rect 36176 7346 36228 7352
rect 36084 6996 36136 7002
rect 36084 6938 36136 6944
rect 35992 6656 36044 6662
rect 35992 6598 36044 6604
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 35808 5568 35860 5574
rect 35808 5510 35860 5516
rect 35820 4162 35848 5510
rect 35912 4282 35940 6394
rect 36004 6338 36032 6598
rect 36096 6458 36124 6938
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36004 6310 36124 6338
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 36004 4690 36032 6190
rect 36096 5574 36124 6310
rect 36176 5772 36228 5778
rect 36176 5714 36228 5720
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 36188 5386 36216 5714
rect 36096 5358 36216 5386
rect 36096 5273 36124 5358
rect 36176 5296 36228 5302
rect 36082 5264 36138 5273
rect 36176 5238 36228 5244
rect 36082 5199 36138 5208
rect 36084 5024 36136 5030
rect 36084 4966 36136 4972
rect 35992 4684 36044 4690
rect 35992 4626 36044 4632
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 35820 4146 35940 4162
rect 35820 4140 35952 4146
rect 35820 4134 35900 4140
rect 35820 3670 35848 4134
rect 35900 4082 35952 4088
rect 36004 3942 36032 4626
rect 36096 4622 36124 4966
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 35992 3936 36044 3942
rect 35898 3904 35954 3913
rect 35992 3878 36044 3884
rect 35898 3839 35954 3848
rect 35808 3664 35860 3670
rect 35808 3606 35860 3612
rect 35912 3602 35940 3839
rect 35900 3596 35952 3602
rect 35900 3538 35952 3544
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 35808 3120 35860 3126
rect 35808 3062 35860 3068
rect 35820 2514 35848 3062
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 36004 800 36032 3402
rect 36096 2990 36124 4558
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 36084 2848 36136 2854
rect 36084 2790 36136 2796
rect 36096 2650 36124 2790
rect 36084 2644 36136 2650
rect 36084 2586 36136 2592
rect 36188 2122 36216 5238
rect 36280 3942 36308 7482
rect 36464 6866 36492 8434
rect 36556 8294 36584 12328
rect 37016 11218 37044 13126
rect 37292 12986 37320 13194
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37384 12850 37412 14214
rect 37476 13818 37504 18686
rect 37648 18624 37700 18630
rect 37648 18566 37700 18572
rect 37556 18216 37608 18222
rect 37556 18158 37608 18164
rect 37568 17542 37596 18158
rect 37556 17536 37608 17542
rect 37556 17478 37608 17484
rect 37568 16046 37596 17478
rect 37660 17338 37688 18566
rect 37844 18426 37872 19654
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37844 17814 37872 18158
rect 37832 17808 37884 17814
rect 37832 17750 37884 17756
rect 37648 17332 37700 17338
rect 37648 17274 37700 17280
rect 37740 16584 37792 16590
rect 37740 16526 37792 16532
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37556 16040 37608 16046
rect 37556 15982 37608 15988
rect 37660 15706 37688 16050
rect 37648 15700 37700 15706
rect 37648 15642 37700 15648
rect 37752 15570 37780 16526
rect 37740 15564 37792 15570
rect 37740 15506 37792 15512
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37648 14340 37700 14346
rect 37648 14282 37700 14288
rect 37660 14074 37688 14282
rect 37648 14068 37700 14074
rect 37648 14010 37700 14016
rect 37648 13932 37700 13938
rect 37648 13874 37700 13880
rect 37476 13790 37596 13818
rect 37464 13728 37516 13734
rect 37464 13670 37516 13676
rect 37476 13190 37504 13670
rect 37464 13184 37516 13190
rect 37464 13126 37516 13132
rect 37568 13002 37596 13790
rect 37476 12974 37596 13002
rect 37372 12844 37424 12850
rect 37372 12786 37424 12792
rect 37476 12442 37504 12974
rect 37556 12912 37608 12918
rect 37556 12854 37608 12860
rect 37464 12436 37516 12442
rect 37464 12378 37516 12384
rect 37568 12186 37596 12854
rect 37292 12158 37596 12186
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 37200 11694 37228 12038
rect 37188 11688 37240 11694
rect 37188 11630 37240 11636
rect 37096 11552 37148 11558
rect 37096 11494 37148 11500
rect 37108 11286 37136 11494
rect 37096 11280 37148 11286
rect 37096 11222 37148 11228
rect 36820 11212 36872 11218
rect 36820 11154 36872 11160
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36832 10062 36860 11154
rect 37016 10810 37044 11154
rect 37004 10804 37056 10810
rect 37004 10746 37056 10752
rect 37200 10742 37228 11630
rect 37188 10736 37240 10742
rect 37188 10678 37240 10684
rect 37292 10606 37320 12158
rect 37660 12050 37688 13874
rect 37740 13796 37792 13802
rect 37740 13738 37792 13744
rect 37752 13530 37780 13738
rect 37740 13524 37792 13530
rect 37740 13466 37792 13472
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37476 12022 37688 12050
rect 37476 11694 37504 12022
rect 37752 11914 37780 13126
rect 37844 12442 37872 14350
rect 37936 14074 37964 14894
rect 37924 14068 37976 14074
rect 37924 14010 37976 14016
rect 37924 13524 37976 13530
rect 37924 13466 37976 13472
rect 37832 12436 37884 12442
rect 37832 12378 37884 12384
rect 37936 12306 37964 13466
rect 38028 12434 38056 21286
rect 38108 17128 38160 17134
rect 38108 17070 38160 17076
rect 38120 12918 38148 17070
rect 38200 16992 38252 16998
rect 38200 16934 38252 16940
rect 38108 12912 38160 12918
rect 38108 12854 38160 12860
rect 38028 12406 38148 12434
rect 37924 12300 37976 12306
rect 37924 12242 37976 12248
rect 38016 12164 38068 12170
rect 38016 12106 38068 12112
rect 37568 11886 37780 11914
rect 37464 11688 37516 11694
rect 37464 11630 37516 11636
rect 37372 11620 37424 11626
rect 37372 11562 37424 11568
rect 37384 11218 37412 11562
rect 37372 11212 37424 11218
rect 37372 11154 37424 11160
rect 37280 10600 37332 10606
rect 37280 10542 37332 10548
rect 37384 10130 37412 11154
rect 37464 11144 37516 11150
rect 37464 11086 37516 11092
rect 37476 10266 37504 11086
rect 37568 10810 37596 11886
rect 37740 11824 37792 11830
rect 37740 11766 37792 11772
rect 37648 11348 37700 11354
rect 37648 11290 37700 11296
rect 37660 10810 37688 11290
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 37648 10804 37700 10810
rect 37648 10746 37700 10752
rect 37648 10600 37700 10606
rect 37648 10542 37700 10548
rect 37464 10260 37516 10266
rect 37464 10202 37516 10208
rect 37372 10124 37424 10130
rect 37372 10066 37424 10072
rect 36820 10056 36872 10062
rect 36820 9998 36872 10004
rect 37280 9988 37332 9994
rect 37280 9930 37332 9936
rect 36820 9920 36872 9926
rect 36820 9862 36872 9868
rect 36832 9518 36860 9862
rect 37292 9722 37320 9930
rect 37280 9716 37332 9722
rect 37280 9658 37332 9664
rect 36820 9512 36872 9518
rect 36820 9454 36872 9460
rect 37476 9042 37504 10202
rect 37660 9058 37688 10542
rect 37752 9178 37780 11766
rect 37924 11688 37976 11694
rect 37924 11630 37976 11636
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 9518 37872 11494
rect 37936 11150 37964 11630
rect 37924 11144 37976 11150
rect 37924 11086 37976 11092
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 37936 10266 37964 10950
rect 37924 10260 37976 10266
rect 37924 10202 37976 10208
rect 38028 9518 38056 12106
rect 37832 9512 37884 9518
rect 37832 9454 37884 9460
rect 38016 9512 38068 9518
rect 38016 9454 38068 9460
rect 37740 9172 37792 9178
rect 37740 9114 37792 9120
rect 37464 9036 37516 9042
rect 37660 9030 37780 9058
rect 37464 8978 37516 8984
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 37372 8968 37424 8974
rect 37372 8910 37424 8916
rect 36648 8634 36676 8910
rect 36820 8832 36872 8838
rect 36820 8774 36872 8780
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 36544 8288 36596 8294
rect 36544 8230 36596 8236
rect 36832 7886 36860 8774
rect 37384 8634 37412 8910
rect 37372 8628 37424 8634
rect 37372 8570 37424 8576
rect 37292 8498 37412 8514
rect 37188 8492 37240 8498
rect 37188 8434 37240 8440
rect 37280 8492 37412 8498
rect 37332 8486 37412 8492
rect 37280 8434 37332 8440
rect 37200 7954 37228 8434
rect 37280 8356 37332 8362
rect 37280 8298 37332 8304
rect 37188 7948 37240 7954
rect 37188 7890 37240 7896
rect 36820 7880 36872 7886
rect 36820 7822 36872 7828
rect 36728 7812 36780 7818
rect 36728 7754 36780 7760
rect 36544 7268 36596 7274
rect 36544 7210 36596 7216
rect 36452 6860 36504 6866
rect 36452 6802 36504 6808
rect 36556 6746 36584 7210
rect 36464 6718 36584 6746
rect 36358 5672 36414 5681
rect 36358 5607 36414 5616
rect 36268 3936 36320 3942
rect 36268 3878 36320 3884
rect 36372 3670 36400 5607
rect 36464 5098 36492 6718
rect 36636 5568 36688 5574
rect 36636 5510 36688 5516
rect 36542 5400 36598 5409
rect 36542 5335 36598 5344
rect 36452 5092 36504 5098
rect 36452 5034 36504 5040
rect 36464 4758 36492 5034
rect 36452 4752 36504 4758
rect 36452 4694 36504 4700
rect 36360 3664 36412 3670
rect 36360 3606 36412 3612
rect 36556 3466 36584 5335
rect 36648 4826 36676 5510
rect 36636 4820 36688 4826
rect 36636 4762 36688 4768
rect 36740 3720 36768 7754
rect 37292 7546 37320 8298
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 37004 7336 37056 7342
rect 37004 7278 37056 7284
rect 37016 6730 37044 7278
rect 36820 6724 36872 6730
rect 36820 6666 36872 6672
rect 37004 6724 37056 6730
rect 37004 6666 37056 6672
rect 37280 6724 37332 6730
rect 37280 6666 37332 6672
rect 36832 5114 36860 6666
rect 37016 6322 37044 6666
rect 37004 6316 37056 6322
rect 37004 6258 37056 6264
rect 36912 6248 36964 6254
rect 36912 6190 36964 6196
rect 36924 5914 36952 6190
rect 36912 5908 36964 5914
rect 36912 5850 36964 5856
rect 37096 5840 37148 5846
rect 37096 5782 37148 5788
rect 37004 5568 37056 5574
rect 37004 5510 37056 5516
rect 36832 5086 36952 5114
rect 36924 4554 36952 5086
rect 36912 4548 36964 4554
rect 36912 4490 36964 4496
rect 36910 4176 36966 4185
rect 36820 4140 36872 4146
rect 36910 4111 36966 4120
rect 36820 4082 36872 4088
rect 36648 3692 36768 3720
rect 36544 3460 36596 3466
rect 36544 3402 36596 3408
rect 36360 3392 36412 3398
rect 36360 3334 36412 3340
rect 36372 3233 36400 3334
rect 36358 3224 36414 3233
rect 36358 3159 36414 3168
rect 36648 2854 36676 3692
rect 36726 3632 36782 3641
rect 36726 3567 36782 3576
rect 36636 2848 36688 2854
rect 36636 2790 36688 2796
rect 36188 2094 36400 2122
rect 36372 800 36400 2094
rect 36740 800 36768 3567
rect 36832 3194 36860 4082
rect 36820 3188 36872 3194
rect 36820 3130 36872 3136
rect 36924 2650 36952 4111
rect 37016 3194 37044 5510
rect 37108 4282 37136 5782
rect 37292 5370 37320 6666
rect 37384 6497 37412 8486
rect 37752 8362 37780 9030
rect 37648 8356 37700 8362
rect 37648 8298 37700 8304
rect 37740 8356 37792 8362
rect 37740 8298 37792 8304
rect 37556 7744 37608 7750
rect 37556 7686 37608 7692
rect 37568 7546 37596 7686
rect 37556 7540 37608 7546
rect 37556 7482 37608 7488
rect 37660 6798 37688 8298
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 37648 6792 37700 6798
rect 37648 6734 37700 6740
rect 37370 6488 37426 6497
rect 37370 6423 37426 6432
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37280 5228 37332 5234
rect 37280 5170 37332 5176
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 37096 4276 37148 4282
rect 37096 4218 37148 4224
rect 37200 4010 37228 4558
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 37292 3738 37320 5170
rect 37280 3732 37332 3738
rect 37280 3674 37332 3680
rect 37384 3618 37412 5646
rect 37476 4826 37504 6734
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37556 5636 37608 5642
rect 37556 5578 37608 5584
rect 37464 4820 37516 4826
rect 37464 4762 37516 4768
rect 37476 4282 37504 4762
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37108 3590 37412 3618
rect 37004 3188 37056 3194
rect 37004 3130 37056 3136
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 37108 800 37136 3590
rect 37462 3360 37518 3369
rect 37462 3295 37518 3304
rect 37476 800 37504 3295
rect 37568 3126 37596 5578
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 37660 2650 37688 6598
rect 37752 5778 37780 8298
rect 37924 7744 37976 7750
rect 37924 7686 37976 7692
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 37740 5772 37792 5778
rect 37740 5714 37792 5720
rect 37936 5098 37964 7686
rect 38028 6458 38056 7686
rect 38120 7410 38148 12406
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38016 6452 38068 6458
rect 38016 6394 38068 6400
rect 38212 6322 38240 16934
rect 38304 15162 38332 25094
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38488 18970 38516 19790
rect 38476 18964 38528 18970
rect 38476 18906 38528 18912
rect 38384 16584 38436 16590
rect 38384 16526 38436 16532
rect 38396 16250 38424 16526
rect 38384 16244 38436 16250
rect 38384 16186 38436 16192
rect 38384 16040 38436 16046
rect 38384 15982 38436 15988
rect 38292 15156 38344 15162
rect 38292 15098 38344 15104
rect 38292 14544 38344 14550
rect 38292 14486 38344 14492
rect 38304 12986 38332 14486
rect 38292 12980 38344 12986
rect 38292 12922 38344 12928
rect 38292 11892 38344 11898
rect 38292 11834 38344 11840
rect 38304 11354 38332 11834
rect 38292 11348 38344 11354
rect 38292 11290 38344 11296
rect 38292 10464 38344 10470
rect 38292 10406 38344 10412
rect 38304 8498 38332 10406
rect 38396 8634 38424 15982
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 38476 10532 38528 10538
rect 38476 10474 38528 10480
rect 38384 8628 38436 8634
rect 38384 8570 38436 8576
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38292 8356 38344 8362
rect 38292 8298 38344 8304
rect 38304 7954 38332 8298
rect 38292 7948 38344 7954
rect 38292 7890 38344 7896
rect 38292 7336 38344 7342
rect 38292 7278 38344 7284
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38304 6254 38332 7278
rect 38292 6248 38344 6254
rect 38292 6190 38344 6196
rect 38016 6112 38068 6118
rect 38016 6054 38068 6060
rect 38028 5234 38056 6054
rect 38304 5817 38332 6190
rect 38384 6112 38436 6118
rect 38384 6054 38436 6060
rect 38290 5808 38346 5817
rect 38290 5743 38346 5752
rect 38292 5704 38344 5710
rect 38292 5646 38344 5652
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 38304 5114 38332 5646
rect 37740 5092 37792 5098
rect 37740 5034 37792 5040
rect 37924 5092 37976 5098
rect 37924 5034 37976 5040
rect 38212 5086 38332 5114
rect 37752 4214 37780 5034
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37740 4208 37792 4214
rect 37740 4150 37792 4156
rect 37844 3534 37872 4966
rect 37922 4448 37978 4457
rect 37922 4383 37978 4392
rect 37936 4078 37964 4383
rect 38212 4298 38240 5086
rect 38292 5024 38344 5030
rect 38292 4966 38344 4972
rect 38028 4270 38240 4298
rect 37924 4072 37976 4078
rect 37924 4014 37976 4020
rect 37924 3936 37976 3942
rect 37924 3878 37976 3884
rect 37832 3528 37884 3534
rect 37738 3496 37794 3505
rect 37832 3470 37884 3476
rect 37738 3431 37794 3440
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 37752 1714 37780 3431
rect 37936 2990 37964 3878
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 37832 2848 37884 2854
rect 37832 2790 37884 2796
rect 37844 2514 37872 2790
rect 38028 2650 38056 4270
rect 38200 4208 38252 4214
rect 38200 4150 38252 4156
rect 38108 3936 38160 3942
rect 38108 3878 38160 3884
rect 38120 3738 38148 3878
rect 38108 3732 38160 3738
rect 38108 3674 38160 3680
rect 38016 2644 38068 2650
rect 38016 2586 38068 2592
rect 37832 2508 37884 2514
rect 37832 2450 37884 2456
rect 37752 1686 37872 1714
rect 37844 800 37872 1686
rect 38212 800 38240 4150
rect 38304 3602 38332 4966
rect 38396 4282 38424 6054
rect 38384 4276 38436 4282
rect 38384 4218 38436 4224
rect 38292 3596 38344 3602
rect 38292 3538 38344 3544
rect 38488 2514 38516 10474
rect 38580 4146 38608 15098
rect 38752 13728 38804 13734
rect 38752 13670 38804 13676
rect 38660 11076 38712 11082
rect 38660 11018 38712 11024
rect 38672 6866 38700 11018
rect 38764 9654 38792 13670
rect 38752 9648 38804 9654
rect 38752 9590 38804 9596
rect 38764 6866 38792 9590
rect 38936 9376 38988 9382
rect 38936 9318 38988 9324
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 38660 6860 38712 6866
rect 38660 6802 38712 6808
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38660 6248 38712 6254
rect 38660 6190 38712 6196
rect 38672 4146 38700 6190
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 38566 3088 38622 3097
rect 38672 3058 38700 4082
rect 38856 4049 38884 7142
rect 38842 4040 38898 4049
rect 38842 3975 38898 3984
rect 38566 3023 38622 3032
rect 38660 3052 38712 3058
rect 38476 2508 38528 2514
rect 38476 2450 38528 2456
rect 38580 800 38608 3023
rect 38660 2994 38712 3000
rect 38672 2514 38700 2994
rect 38660 2508 38712 2514
rect 38660 2450 38712 2456
rect 38948 800 38976 9318
rect 39304 1760 39356 1766
rect 39304 1702 39356 1708
rect 39316 800 39344 1702
rect 34256 734 34468 762
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4250 23196 4252 23216
rect 4252 23196 4304 23216
rect 4304 23196 4306 23216
rect 4250 23160 4306 23196
rect 4710 23160 4766 23216
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4802 16632 4858 16688
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 5078 23160 5134 23216
rect 4434 15020 4490 15056
rect 4434 15000 4436 15020
rect 4436 15000 4488 15020
rect 4488 15000 4490 15020
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3974 13932 4030 13968
rect 3974 13912 3976 13932
rect 3976 13912 4028 13932
rect 4028 13912 4030 13932
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3146 7656 3202 7712
rect 3146 6160 3202 6216
rect 2870 3984 2926 4040
rect 2594 3576 2650 3632
rect 2686 3440 2742 3496
rect 2502 3304 2558 3360
rect 2962 3576 3018 3632
rect 2962 3168 3018 3224
rect 3330 3576 3386 3632
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4158 7248 4214 7304
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4710 7656 4766 7712
rect 4802 7248 4858 7304
rect 4802 6160 4858 6216
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 3576 4674 3632
rect 5078 3984 5134 4040
rect 5170 3168 5226 3224
rect 6366 23160 6422 23216
rect 7654 23160 7710 23216
rect 8022 22208 8078 22264
rect 7746 12144 7802 12200
rect 8206 12144 8262 12200
rect 7378 6160 7434 6216
rect 5446 3304 5502 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8298 11600 8354 11656
rect 9494 13812 9496 13832
rect 9496 13812 9548 13832
rect 9548 13812 9550 13832
rect 9494 13776 9550 13812
rect 11518 19236 11574 19272
rect 11518 19216 11520 19236
rect 11520 19216 11572 19236
rect 11572 19216 11574 19236
rect 7838 3984 7894 4040
rect 8666 5616 8722 5672
rect 11426 6296 11482 6352
rect 11058 4528 11114 4584
rect 11242 3848 11298 3904
rect 14370 19216 14426 19272
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 14186 3340 14188 3360
rect 14188 3340 14240 3360
rect 14240 3340 14242 3360
rect 14186 3304 14242 3340
rect 14830 3984 14886 4040
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19246 20748 19248 20768
rect 19248 20748 19300 20768
rect 19300 20748 19302 20768
rect 19246 20712 19302 20748
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 17406 14884 17462 14920
rect 17406 14864 17408 14884
rect 17408 14864 17460 14884
rect 17460 14864 17462 14884
rect 15014 3848 15070 3904
rect 14646 3460 14702 3496
rect 14646 3440 14648 3460
rect 14648 3440 14700 3460
rect 14700 3440 14702 3460
rect 16210 4528 16266 4584
rect 17774 14864 17830 14920
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 18602 14900 18604 14920
rect 18604 14900 18656 14920
rect 18656 14900 18658 14920
rect 18602 14864 18658 14900
rect 17222 6296 17278 6352
rect 18602 6296 18658 6352
rect 18602 3984 18658 4040
rect 18970 3984 19026 4040
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 20258 21004 20314 21040
rect 20258 20984 20260 21004
rect 20260 20984 20312 21004
rect 20312 20984 20314 21004
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19430 6180 19486 6216
rect 19430 6160 19432 6180
rect 19432 6160 19484 6180
rect 19484 6160 19486 6180
rect 19614 5652 19616 5672
rect 19616 5652 19668 5672
rect 19668 5652 19670 5672
rect 19614 5616 19670 5652
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 22558 19796 22560 19816
rect 22560 19796 22612 19816
rect 22612 19796 22614 19816
rect 22558 19760 22614 19796
rect 23110 19760 23166 19816
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 24398 26288 24454 26344
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22374 5072 22430 5128
rect 23570 3440 23626 3496
rect 24214 7692 24216 7712
rect 24216 7692 24268 7712
rect 24268 7692 24270 7712
rect 24214 7656 24270 7692
rect 23938 3440 23994 3496
rect 29274 27648 29330 27704
rect 24582 11464 24638 11520
rect 24674 6840 24730 6896
rect 24490 5636 24546 5672
rect 24490 5616 24492 5636
rect 24492 5616 24544 5636
rect 24544 5616 24546 5636
rect 24490 5208 24546 5264
rect 26054 11092 26056 11112
rect 26056 11092 26108 11112
rect 26108 11092 26110 11112
rect 26054 11056 26110 11092
rect 25686 3984 25742 4040
rect 25594 3848 25650 3904
rect 26606 3440 26662 3496
rect 32218 29044 32220 29064
rect 32220 29044 32272 29064
rect 32272 29044 32274 29064
rect 32218 29008 32274 29044
rect 30194 23704 30250 23760
rect 27066 7656 27122 7712
rect 28354 11056 28410 11112
rect 27066 5108 27068 5128
rect 27068 5108 27120 5128
rect 27120 5108 27122 5128
rect 27066 5072 27122 5108
rect 26606 2644 26662 2680
rect 26606 2624 26608 2644
rect 26608 2624 26660 2644
rect 26660 2624 26662 2644
rect 27618 4936 27674 4992
rect 27434 4020 27436 4040
rect 27436 4020 27488 4040
rect 27488 4020 27490 4040
rect 27434 3984 27490 4020
rect 28998 11464 29054 11520
rect 32770 29708 32826 29744
rect 32770 29688 32772 29708
rect 32772 29688 32824 29708
rect 32824 29688 32826 29708
rect 33138 29552 33194 29608
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 29182 6840 29238 6896
rect 27526 2760 27582 2816
rect 29182 4392 29238 4448
rect 30746 13776 30802 13832
rect 30286 6704 30342 6760
rect 30194 6452 30250 6488
rect 30194 6432 30196 6452
rect 30196 6432 30248 6452
rect 30248 6432 30250 6452
rect 30102 6296 30158 6352
rect 30194 4684 30250 4720
rect 30194 4664 30196 4684
rect 30196 4664 30248 4684
rect 30248 4664 30250 4684
rect 30102 3984 30158 4040
rect 30194 3848 30250 3904
rect 30470 5480 30526 5536
rect 31114 5072 31170 5128
rect 31482 4156 31484 4176
rect 31484 4156 31536 4176
rect 31536 4156 31538 4176
rect 31482 4120 31538 4156
rect 33782 17584 33838 17640
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35898 29028 35954 29064
rect 35898 29008 35900 29028
rect 35900 29008 35952 29028
rect 35952 29008 35954 29028
rect 37278 29552 37334 29608
rect 37830 29688 37886 29744
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34610 21800 34666 21856
rect 35530 21800 35586 21856
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 33414 11600 33470 11656
rect 32218 5616 32274 5672
rect 32034 5344 32090 5400
rect 31850 5208 31906 5264
rect 32218 5208 32274 5264
rect 32034 5072 32090 5128
rect 31942 2760 31998 2816
rect 32218 3576 32274 3632
rect 33966 11056 34022 11112
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35254 17584 35310 17640
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 37186 23704 37242 23760
rect 35898 15000 35954 15056
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 37462 21020 37464 21040
rect 37464 21020 37516 21040
rect 37516 21020 37518 21040
rect 37462 20984 37518 21020
rect 34610 13912 34666 13968
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34518 12860 34520 12880
rect 34520 12860 34572 12880
rect 34572 12860 34574 12880
rect 34518 12824 34574 12860
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 32310 3168 32366 3224
rect 32678 4140 32734 4176
rect 32678 4120 32680 4140
rect 32680 4120 32732 4140
rect 32732 4120 32734 4140
rect 32770 3304 32826 3360
rect 33414 5752 33470 5808
rect 33874 5480 33930 5536
rect 33230 4392 33286 4448
rect 33598 4120 33654 4176
rect 33874 4684 33930 4720
rect 33874 4664 33876 4684
rect 33876 4664 33928 4684
rect 33928 4664 33930 4684
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34242 5772 34298 5808
rect 34242 5752 34244 5772
rect 34244 5752 34296 5772
rect 34296 5752 34298 5772
rect 34058 3168 34114 3224
rect 34426 3984 34482 4040
rect 35530 6704 35586 6760
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34886 4664 34942 4720
rect 35346 3848 35402 3904
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36358 11092 36360 11112
rect 36360 11092 36412 11112
rect 36412 11092 36414 11112
rect 36358 11056 36414 11092
rect 36082 5208 36138 5264
rect 35898 3848 35954 3904
rect 36358 5616 36414 5672
rect 36542 5344 36598 5400
rect 36910 4120 36966 4176
rect 36358 3168 36414 3224
rect 36726 3576 36782 3632
rect 37370 6432 37426 6488
rect 37462 3304 37518 3360
rect 38290 5752 38346 5808
rect 37922 4392 37978 4448
rect 37738 3440 37794 3496
rect 38566 3032 38622 3088
rect 38842 3984 38898 4040
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 32765 29746 32831 29749
rect 37825 29746 37891 29749
rect 32765 29744 37891 29746
rect 32765 29688 32770 29744
rect 32826 29688 37830 29744
rect 37886 29688 37891 29744
rect 32765 29686 37891 29688
rect 32765 29683 32831 29686
rect 37825 29683 37891 29686
rect 33133 29610 33199 29613
rect 37273 29610 37339 29613
rect 33133 29608 37339 29610
rect 33133 29552 33138 29608
rect 33194 29552 37278 29608
rect 37334 29552 37339 29608
rect 33133 29550 37339 29552
rect 33133 29547 33199 29550
rect 37273 29547 37339 29550
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 32213 29066 32279 29069
rect 35893 29066 35959 29069
rect 32213 29064 35959 29066
rect 32213 29008 32218 29064
rect 32274 29008 35898 29064
rect 35954 29008 35959 29064
rect 32213 29006 35959 29008
rect 32213 29003 32279 29006
rect 35893 29003 35959 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 29269 27708 29335 27709
rect 29269 27704 29316 27708
rect 29380 27706 29386 27708
rect 29269 27648 29274 27704
rect 29269 27644 29316 27648
rect 29380 27646 29426 27706
rect 29380 27644 29386 27646
rect 29269 27643 29335 27644
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 24393 26346 24459 26349
rect 24710 26346 24716 26348
rect 24393 26344 24716 26346
rect 24393 26288 24398 26344
rect 24454 26288 24716 26344
rect 24393 26286 24716 26288
rect 24393 26283 24459 26286
rect 24710 26284 24716 26286
rect 24780 26284 24786 26348
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 30189 23762 30255 23765
rect 37181 23762 37247 23765
rect 30189 23760 37247 23762
rect 30189 23704 30194 23760
rect 30250 23704 37186 23760
rect 37242 23704 37247 23760
rect 30189 23702 37247 23704
rect 30189 23699 30255 23702
rect 37181 23699 37247 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4245 23218 4311 23221
rect 4705 23218 4771 23221
rect 5073 23218 5139 23221
rect 4245 23216 5139 23218
rect 4245 23160 4250 23216
rect 4306 23160 4710 23216
rect 4766 23160 5078 23216
rect 5134 23160 5139 23216
rect 4245 23158 5139 23160
rect 4245 23155 4311 23158
rect 4705 23155 4771 23158
rect 5073 23155 5139 23158
rect 6361 23218 6427 23221
rect 7649 23218 7715 23221
rect 6361 23216 7715 23218
rect 6361 23160 6366 23216
rect 6422 23160 7654 23216
rect 7710 23160 7715 23216
rect 6361 23158 7715 23160
rect 6361 23155 6427 23158
rect 7649 23155 7715 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 8017 22268 8083 22269
rect 7966 22266 7972 22268
rect 7926 22206 7972 22266
rect 8036 22264 8083 22268
rect 8078 22208 8083 22264
rect 7966 22204 7972 22206
rect 8036 22204 8083 22208
rect 8017 22203 8083 22204
rect 34605 21858 34671 21861
rect 35525 21858 35591 21861
rect 34605 21856 35591 21858
rect 34605 21800 34610 21856
rect 34666 21800 35530 21856
rect 35586 21800 35591 21856
rect 34605 21798 35591 21800
rect 34605 21795 34671 21798
rect 35525 21795 35591 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 20253 21042 20319 21045
rect 37457 21042 37523 21045
rect 20253 21040 37523 21042
rect 20253 20984 20258 21040
rect 20314 20984 37462 21040
rect 37518 20984 37523 21040
rect 20253 20982 37523 20984
rect 20253 20979 20319 20982
rect 37457 20979 37523 20982
rect 19006 20708 19012 20772
rect 19076 20770 19082 20772
rect 19241 20770 19307 20773
rect 19076 20768 19307 20770
rect 19076 20712 19246 20768
rect 19302 20712 19307 20768
rect 19076 20710 19307 20712
rect 19076 20708 19082 20710
rect 19241 20707 19307 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 22553 19818 22619 19821
rect 23105 19818 23171 19821
rect 22553 19816 23171 19818
rect 22553 19760 22558 19816
rect 22614 19760 23110 19816
rect 23166 19760 23171 19816
rect 22553 19758 23171 19760
rect 22553 19755 22619 19758
rect 23105 19755 23171 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 11513 19274 11579 19277
rect 14365 19274 14431 19277
rect 11513 19272 14431 19274
rect 11513 19216 11518 19272
rect 11574 19216 14370 19272
rect 14426 19216 14431 19272
rect 11513 19214 14431 19216
rect 11513 19211 11579 19214
rect 14365 19211 14431 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 33777 17642 33843 17645
rect 35249 17642 35315 17645
rect 33777 17640 35315 17642
rect 33777 17584 33782 17640
rect 33838 17584 35254 17640
rect 35310 17584 35315 17640
rect 33777 17582 35315 17584
rect 33777 17579 33843 17582
rect 35249 17579 35315 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4797 16692 4863 16693
rect 4797 16688 4844 16692
rect 4908 16690 4914 16692
rect 4797 16632 4802 16688
rect 4797 16628 4844 16632
rect 4908 16630 4954 16690
rect 4908 16628 4914 16630
rect 4797 16627 4863 16628
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4429 15058 4495 15061
rect 35893 15058 35959 15061
rect 4429 15056 35959 15058
rect 4429 15000 4434 15056
rect 4490 15000 35898 15056
rect 35954 15000 35959 15056
rect 4429 14998 35959 15000
rect 4429 14995 4495 14998
rect 35893 14995 35959 14998
rect 17401 14922 17467 14925
rect 17769 14922 17835 14925
rect 18597 14922 18663 14925
rect 17401 14920 18663 14922
rect 17401 14864 17406 14920
rect 17462 14864 17774 14920
rect 17830 14864 18602 14920
rect 18658 14864 18663 14920
rect 17401 14862 18663 14864
rect 17401 14859 17467 14862
rect 17769 14859 17835 14862
rect 18597 14859 18663 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 3969 13970 4035 13973
rect 34605 13970 34671 13973
rect 3969 13968 34671 13970
rect 3969 13912 3974 13968
rect 4030 13912 34610 13968
rect 34666 13912 34671 13968
rect 3969 13910 34671 13912
rect 3969 13907 4035 13910
rect 34605 13907 34671 13910
rect 9489 13834 9555 13837
rect 30741 13834 30807 13837
rect 9489 13832 30807 13834
rect 9489 13776 9494 13832
rect 9550 13776 30746 13832
rect 30802 13776 30807 13832
rect 9489 13774 30807 13776
rect 9489 13771 9555 13774
rect 30741 13771 30807 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 34513 12882 34579 12885
rect 34646 12882 34652 12884
rect 34513 12880 34652 12882
rect 34513 12824 34518 12880
rect 34574 12824 34652 12880
rect 34513 12822 34652 12824
rect 34513 12819 34579 12822
rect 34646 12820 34652 12822
rect 34716 12820 34722 12884
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 7741 12202 7807 12205
rect 8201 12202 8267 12205
rect 7741 12200 8267 12202
rect 7741 12144 7746 12200
rect 7802 12144 8206 12200
rect 8262 12144 8267 12200
rect 7741 12142 8267 12144
rect 7741 12139 7807 12142
rect 8201 12139 8267 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 8293 11658 8359 11661
rect 33409 11658 33475 11661
rect 8293 11656 33475 11658
rect 8293 11600 8298 11656
rect 8354 11600 33414 11656
rect 33470 11600 33475 11656
rect 8293 11598 33475 11600
rect 8293 11595 8359 11598
rect 33409 11595 33475 11598
rect 24577 11522 24643 11525
rect 28993 11522 29059 11525
rect 24577 11520 29059 11522
rect 24577 11464 24582 11520
rect 24638 11464 28998 11520
rect 29054 11464 29059 11520
rect 24577 11462 29059 11464
rect 24577 11459 24643 11462
rect 28993 11459 29059 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 26049 11114 26115 11117
rect 28349 11114 28415 11117
rect 26049 11112 28415 11114
rect 26049 11056 26054 11112
rect 26110 11056 28354 11112
rect 28410 11056 28415 11112
rect 26049 11054 28415 11056
rect 26049 11051 26115 11054
rect 28349 11051 28415 11054
rect 33961 11114 34027 11117
rect 36353 11114 36419 11117
rect 33961 11112 36419 11114
rect 33961 11056 33966 11112
rect 34022 11056 36358 11112
rect 36414 11056 36419 11112
rect 33961 11054 36419 11056
rect 33961 11051 34027 11054
rect 36353 11051 36419 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 3141 7714 3207 7717
rect 4705 7714 4771 7717
rect 3141 7712 4771 7714
rect 3141 7656 3146 7712
rect 3202 7656 4710 7712
rect 4766 7656 4771 7712
rect 3141 7654 4771 7656
rect 3141 7651 3207 7654
rect 4705 7651 4771 7654
rect 24209 7714 24275 7717
rect 27061 7714 27127 7717
rect 24209 7712 27127 7714
rect 24209 7656 24214 7712
rect 24270 7656 27066 7712
rect 27122 7656 27127 7712
rect 24209 7654 27127 7656
rect 24209 7651 24275 7654
rect 27061 7651 27127 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4153 7306 4219 7309
rect 4797 7306 4863 7309
rect 4153 7304 4863 7306
rect 4153 7248 4158 7304
rect 4214 7248 4802 7304
rect 4858 7248 4863 7304
rect 4153 7246 4863 7248
rect 4153 7243 4219 7246
rect 4797 7243 4863 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 24669 6900 24735 6901
rect 24669 6896 24716 6900
rect 24780 6898 24786 6900
rect 29177 6898 29243 6901
rect 29310 6898 29316 6900
rect 24669 6840 24674 6896
rect 24669 6836 24716 6840
rect 24780 6838 24826 6898
rect 29177 6896 29316 6898
rect 29177 6840 29182 6896
rect 29238 6840 29316 6896
rect 29177 6838 29316 6840
rect 24780 6836 24786 6838
rect 24669 6835 24735 6836
rect 29177 6835 29243 6838
rect 29310 6836 29316 6838
rect 29380 6836 29386 6900
rect 30281 6762 30347 6765
rect 35525 6762 35591 6765
rect 30281 6760 35591 6762
rect 30281 6704 30286 6760
rect 30342 6704 35530 6760
rect 35586 6704 35591 6760
rect 30281 6702 35591 6704
rect 30281 6699 30347 6702
rect 35525 6699 35591 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 30189 6490 30255 6493
rect 37365 6490 37431 6493
rect 30189 6488 37431 6490
rect 30189 6432 30194 6488
rect 30250 6432 37370 6488
rect 37426 6432 37431 6488
rect 30189 6430 37431 6432
rect 30189 6427 30255 6430
rect 37365 6427 37431 6430
rect 11421 6354 11487 6357
rect 17217 6354 17283 6357
rect 18597 6354 18663 6357
rect 11421 6352 18663 6354
rect 11421 6296 11426 6352
rect 11482 6296 17222 6352
rect 17278 6296 18602 6352
rect 18658 6296 18663 6352
rect 11421 6294 18663 6296
rect 11421 6291 11487 6294
rect 17217 6291 17283 6294
rect 18597 6291 18663 6294
rect 30097 6354 30163 6357
rect 30230 6354 30236 6356
rect 30097 6352 30236 6354
rect 30097 6296 30102 6352
rect 30158 6296 30236 6352
rect 30097 6294 30236 6296
rect 30097 6291 30163 6294
rect 30230 6292 30236 6294
rect 30300 6292 30306 6356
rect 3141 6218 3207 6221
rect 4797 6218 4863 6221
rect 3141 6216 4863 6218
rect 3141 6160 3146 6216
rect 3202 6160 4802 6216
rect 4858 6160 4863 6216
rect 3141 6158 4863 6160
rect 3141 6155 3207 6158
rect 4797 6155 4863 6158
rect 7373 6218 7439 6221
rect 19425 6218 19491 6221
rect 7373 6216 19491 6218
rect 7373 6160 7378 6216
rect 7434 6160 19430 6216
rect 19486 6160 19491 6216
rect 7373 6158 19491 6160
rect 7373 6155 7439 6158
rect 19425 6155 19491 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 33409 5810 33475 5813
rect 34237 5810 34303 5813
rect 38285 5810 38351 5813
rect 33409 5808 38351 5810
rect 33409 5752 33414 5808
rect 33470 5752 34242 5808
rect 34298 5752 38290 5808
rect 38346 5752 38351 5808
rect 33409 5750 38351 5752
rect 33409 5747 33475 5750
rect 34237 5747 34303 5750
rect 38285 5747 38351 5750
rect 8661 5674 8727 5677
rect 19609 5674 19675 5677
rect 8661 5672 19675 5674
rect 8661 5616 8666 5672
rect 8722 5616 19614 5672
rect 19670 5616 19675 5672
rect 8661 5614 19675 5616
rect 8661 5611 8727 5614
rect 19609 5611 19675 5614
rect 24485 5674 24551 5677
rect 26182 5674 26188 5676
rect 24485 5672 26188 5674
rect 24485 5616 24490 5672
rect 24546 5616 26188 5672
rect 24485 5614 26188 5616
rect 24485 5611 24551 5614
rect 26182 5612 26188 5614
rect 26252 5612 26258 5676
rect 32213 5674 32279 5677
rect 36353 5674 36419 5677
rect 32213 5672 36419 5674
rect 32213 5616 32218 5672
rect 32274 5616 36358 5672
rect 36414 5616 36419 5672
rect 32213 5614 36419 5616
rect 32213 5611 32279 5614
rect 36353 5611 36419 5614
rect 30465 5538 30531 5541
rect 33869 5538 33935 5541
rect 30465 5536 33935 5538
rect 30465 5480 30470 5536
rect 30526 5480 33874 5536
rect 33930 5480 33935 5536
rect 30465 5478 33935 5480
rect 30465 5475 30531 5478
rect 33869 5475 33935 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 32029 5402 32095 5405
rect 36537 5402 36603 5405
rect 32029 5400 36603 5402
rect 32029 5344 32034 5400
rect 32090 5344 36542 5400
rect 36598 5344 36603 5400
rect 32029 5342 36603 5344
rect 32029 5339 32095 5342
rect 36537 5339 36603 5342
rect 24485 5266 24551 5269
rect 31845 5266 31911 5269
rect 32213 5266 32279 5269
rect 36077 5266 36143 5269
rect 24485 5264 36143 5266
rect 24485 5208 24490 5264
rect 24546 5208 31850 5264
rect 31906 5208 32218 5264
rect 32274 5208 36082 5264
rect 36138 5208 36143 5264
rect 24485 5206 36143 5208
rect 24485 5203 24551 5206
rect 22369 5130 22435 5133
rect 27061 5130 27127 5133
rect 22369 5128 27127 5130
rect 22369 5072 22374 5128
rect 22430 5072 27066 5128
rect 27122 5072 27127 5128
rect 22369 5070 27127 5072
rect 22369 5067 22435 5070
rect 27061 5067 27127 5070
rect 27662 4997 27722 5206
rect 31845 5203 31911 5206
rect 32213 5203 32279 5206
rect 36077 5203 36143 5206
rect 31109 5130 31175 5133
rect 32029 5130 32095 5133
rect 31109 5128 32095 5130
rect 31109 5072 31114 5128
rect 31170 5072 32034 5128
rect 32090 5072 32095 5128
rect 31109 5070 32095 5072
rect 31109 5067 31175 5070
rect 32029 5067 32095 5070
rect 27613 4992 27722 4997
rect 27613 4936 27618 4992
rect 27674 4936 27722 4992
rect 27613 4934 27722 4936
rect 27613 4931 27679 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 30189 4722 30255 4725
rect 33869 4722 33935 4725
rect 30189 4720 33935 4722
rect 30189 4664 30194 4720
rect 30250 4664 33874 4720
rect 33930 4664 33935 4720
rect 30189 4662 33935 4664
rect 30189 4659 30255 4662
rect 33869 4659 33935 4662
rect 34646 4660 34652 4724
rect 34716 4722 34722 4724
rect 34881 4722 34947 4725
rect 34716 4720 34947 4722
rect 34716 4664 34886 4720
rect 34942 4664 34947 4720
rect 34716 4662 34947 4664
rect 34716 4660 34722 4662
rect 34881 4659 34947 4662
rect 11053 4586 11119 4589
rect 16205 4586 16271 4589
rect 11053 4584 16271 4586
rect 11053 4528 11058 4584
rect 11114 4528 16210 4584
rect 16266 4528 16271 4584
rect 11053 4526 16271 4528
rect 11053 4523 11119 4526
rect 16205 4523 16271 4526
rect 29177 4450 29243 4453
rect 33225 4450 33291 4453
rect 37917 4450 37983 4453
rect 29177 4448 37983 4450
rect 29177 4392 29182 4448
rect 29238 4392 33230 4448
rect 33286 4392 37922 4448
rect 37978 4392 37983 4448
rect 29177 4390 37983 4392
rect 29177 4387 29243 4390
rect 33225 4387 33291 4390
rect 37917 4387 37983 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 31477 4178 31543 4181
rect 32673 4178 32739 4181
rect 31477 4176 32739 4178
rect 31477 4120 31482 4176
rect 31538 4120 32678 4176
rect 32734 4120 32739 4176
rect 31477 4118 32739 4120
rect 31477 4115 31543 4118
rect 32673 4115 32739 4118
rect 33593 4178 33659 4181
rect 36905 4178 36971 4181
rect 33593 4176 36971 4178
rect 33593 4120 33598 4176
rect 33654 4120 36910 4176
rect 36966 4120 36971 4176
rect 33593 4118 36971 4120
rect 33593 4115 33659 4118
rect 36905 4115 36971 4118
rect 2865 4042 2931 4045
rect 5073 4042 5139 4045
rect 2865 4040 5139 4042
rect 2865 3984 2870 4040
rect 2926 3984 5078 4040
rect 5134 3984 5139 4040
rect 2865 3982 5139 3984
rect 2865 3979 2931 3982
rect 5073 3979 5139 3982
rect 7833 4042 7899 4045
rect 7966 4042 7972 4044
rect 7833 4040 7972 4042
rect 7833 3984 7838 4040
rect 7894 3984 7972 4040
rect 7833 3982 7972 3984
rect 7833 3979 7899 3982
rect 7966 3980 7972 3982
rect 8036 3980 8042 4044
rect 14825 4042 14891 4045
rect 18597 4042 18663 4045
rect 14825 4040 18663 4042
rect 14825 3984 14830 4040
rect 14886 3984 18602 4040
rect 18658 3984 18663 4040
rect 14825 3982 18663 3984
rect 14825 3979 14891 3982
rect 18597 3979 18663 3982
rect 18965 4044 19031 4045
rect 18965 4040 19012 4044
rect 19076 4042 19082 4044
rect 25681 4042 25747 4045
rect 27429 4042 27495 4045
rect 18965 3984 18970 4040
rect 18965 3980 19012 3984
rect 19076 3982 19122 4042
rect 25681 4040 27495 4042
rect 25681 3984 25686 4040
rect 25742 3984 27434 4040
rect 27490 3984 27495 4040
rect 25681 3982 27495 3984
rect 19076 3980 19082 3982
rect 18965 3979 19031 3980
rect 25681 3979 25747 3982
rect 27429 3979 27495 3982
rect 30097 4042 30163 4045
rect 34421 4042 34487 4045
rect 38837 4042 38903 4045
rect 30097 4040 31770 4042
rect 30097 3984 30102 4040
rect 30158 3984 31770 4040
rect 30097 3982 31770 3984
rect 30097 3979 30163 3982
rect 11237 3906 11303 3909
rect 15009 3906 15075 3909
rect 11237 3904 15075 3906
rect 11237 3848 11242 3904
rect 11298 3848 15014 3904
rect 15070 3848 15075 3904
rect 11237 3846 15075 3848
rect 11237 3843 11303 3846
rect 15009 3843 15075 3846
rect 25589 3906 25655 3909
rect 30189 3906 30255 3909
rect 25589 3904 30255 3906
rect 25589 3848 25594 3904
rect 25650 3848 30194 3904
rect 30250 3848 30255 3904
rect 25589 3846 30255 3848
rect 25589 3843 25655 3846
rect 30189 3843 30255 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 31710 3770 31770 3982
rect 34421 4040 38903 4042
rect 34421 3984 34426 4040
rect 34482 3984 38842 4040
rect 38898 3984 38903 4040
rect 34421 3982 38903 3984
rect 34421 3979 34487 3982
rect 38837 3979 38903 3982
rect 35341 3906 35407 3909
rect 35893 3906 35959 3909
rect 35341 3904 35959 3906
rect 35341 3848 35346 3904
rect 35402 3848 35898 3904
rect 35954 3848 35959 3904
rect 35341 3846 35959 3848
rect 35341 3843 35407 3846
rect 35893 3843 35959 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 31710 3710 34346 3770
rect 2589 3634 2655 3637
rect 2957 3634 3023 3637
rect 2589 3632 3023 3634
rect 2589 3576 2594 3632
rect 2650 3576 2962 3632
rect 3018 3576 3023 3632
rect 2589 3574 3023 3576
rect 2589 3571 2655 3574
rect 2957 3571 3023 3574
rect 3325 3634 3391 3637
rect 4613 3634 4679 3637
rect 32213 3634 32279 3637
rect 3325 3632 32279 3634
rect 3325 3576 3330 3632
rect 3386 3576 4618 3632
rect 4674 3576 32218 3632
rect 32274 3576 32279 3632
rect 3325 3574 32279 3576
rect 34286 3634 34346 3710
rect 36721 3634 36787 3637
rect 34286 3632 36787 3634
rect 34286 3576 36726 3632
rect 36782 3576 36787 3632
rect 34286 3574 36787 3576
rect 3325 3571 3391 3574
rect 4613 3571 4679 3574
rect 32213 3571 32279 3574
rect 36721 3571 36787 3574
rect 2681 3498 2747 3501
rect 4838 3498 4844 3500
rect 2681 3496 4844 3498
rect 2681 3440 2686 3496
rect 2742 3440 4844 3496
rect 2681 3438 4844 3440
rect 2681 3435 2747 3438
rect 4838 3436 4844 3438
rect 4908 3436 4914 3500
rect 14641 3498 14707 3501
rect 23565 3498 23631 3501
rect 14641 3496 23631 3498
rect 14641 3440 14646 3496
rect 14702 3440 23570 3496
rect 23626 3440 23631 3496
rect 14641 3438 23631 3440
rect 14641 3435 14707 3438
rect 23565 3435 23631 3438
rect 23933 3498 23999 3501
rect 26601 3498 26667 3501
rect 23933 3496 26667 3498
rect 23933 3440 23938 3496
rect 23994 3440 26606 3496
rect 26662 3440 26667 3496
rect 23933 3438 26667 3440
rect 23933 3435 23999 3438
rect 26601 3435 26667 3438
rect 30230 3436 30236 3500
rect 30300 3498 30306 3500
rect 37733 3498 37799 3501
rect 30300 3496 37799 3498
rect 30300 3440 37738 3496
rect 37794 3440 37799 3496
rect 30300 3438 37799 3440
rect 30300 3436 30306 3438
rect 37733 3435 37799 3438
rect 2497 3362 2563 3365
rect 5441 3362 5507 3365
rect 14181 3362 14247 3365
rect 2497 3360 14247 3362
rect 2497 3304 2502 3360
rect 2558 3304 5446 3360
rect 5502 3304 14186 3360
rect 14242 3304 14247 3360
rect 2497 3302 14247 3304
rect 2497 3299 2563 3302
rect 5441 3299 5507 3302
rect 14181 3299 14247 3302
rect 32765 3362 32831 3365
rect 37457 3362 37523 3365
rect 32765 3360 37523 3362
rect 32765 3304 32770 3360
rect 32826 3304 37462 3360
rect 37518 3304 37523 3360
rect 32765 3302 37523 3304
rect 32765 3299 32831 3302
rect 37457 3299 37523 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 2957 3226 3023 3229
rect 5165 3226 5231 3229
rect 2957 3224 5231 3226
rect 2957 3168 2962 3224
rect 3018 3168 5170 3224
rect 5226 3168 5231 3224
rect 2957 3166 5231 3168
rect 2957 3163 3023 3166
rect 5165 3163 5231 3166
rect 32305 3226 32371 3229
rect 34053 3226 34119 3229
rect 36353 3226 36419 3229
rect 32305 3224 33058 3226
rect 32305 3168 32310 3224
rect 32366 3168 33058 3224
rect 32305 3166 33058 3168
rect 32305 3163 32371 3166
rect 32998 3090 33058 3166
rect 34053 3224 36419 3226
rect 34053 3168 34058 3224
rect 34114 3168 36358 3224
rect 36414 3168 36419 3224
rect 34053 3166 36419 3168
rect 34053 3163 34119 3166
rect 36353 3163 36419 3166
rect 38561 3090 38627 3093
rect 32998 3088 38627 3090
rect 32998 3032 38566 3088
rect 38622 3032 38627 3088
rect 32998 3030 38627 3032
rect 38561 3027 38627 3030
rect 26182 2892 26188 2956
rect 26252 2892 26258 2956
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 26190 2682 26250 2892
rect 27521 2818 27587 2821
rect 31937 2818 32003 2821
rect 27521 2816 32003 2818
rect 27521 2760 27526 2816
rect 27582 2760 31942 2816
rect 31998 2760 32003 2816
rect 27521 2758 32003 2760
rect 27521 2755 27587 2758
rect 31937 2755 32003 2758
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 26601 2682 26667 2685
rect 26190 2680 26667 2682
rect 26190 2624 26606 2680
rect 26662 2624 26667 2680
rect 26190 2622 26667 2624
rect 26601 2619 26667 2622
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 29316 27704 29380 27708
rect 29316 27648 29330 27704
rect 29330 27648 29380 27704
rect 29316 27644 29380 27648
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 24716 26284 24780 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 7972 22264 8036 22268
rect 7972 22208 8022 22264
rect 8022 22208 8036 22264
rect 7972 22204 8036 22208
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19012 20708 19076 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4844 16688 4908 16692
rect 4844 16632 4858 16688
rect 4858 16632 4908 16688
rect 4844 16628 4908 16632
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 34652 12820 34716 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 24716 6896 24780 6900
rect 24716 6840 24730 6896
rect 24730 6840 24780 6896
rect 24716 6836 24780 6840
rect 29316 6836 29380 6900
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 30236 6292 30300 6356
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 26188 5612 26252 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 34652 4660 34716 4724
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 7972 3980 8036 4044
rect 19012 4040 19076 4044
rect 19012 3984 19026 4040
rect 19026 3984 19076 4040
rect 19012 3980 19076 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4844 3436 4908 3500
rect 30236 3436 30300 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 26188 2892 26252 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 29315 27708 29381 27709
rect 29315 27644 29316 27708
rect 29380 27644 29381 27708
rect 29315 27643 29381 27644
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 24715 26348 24781 26349
rect 24715 26284 24716 26348
rect 24780 26284 24781 26348
rect 24715 26283 24781 26284
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 7971 22268 8037 22269
rect 7971 22204 7972 22268
rect 8036 22204 8037 22268
rect 7971 22203 8037 22204
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4843 16692 4909 16693
rect 4843 16628 4844 16692
rect 4908 16628 4909 16692
rect 4843 16627 4909 16628
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4846 3501 4906 16627
rect 7974 4045 8034 22203
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19011 20772 19077 20773
rect 19011 20708 19012 20772
rect 19076 20708 19077 20772
rect 19011 20707 19077 20708
rect 19014 4045 19074 20707
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 24718 6901 24778 26283
rect 29318 6901 29378 27643
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34651 12884 34717 12885
rect 34651 12820 34652 12884
rect 34716 12820 34717 12884
rect 34651 12819 34717 12820
rect 24715 6900 24781 6901
rect 24715 6836 24716 6900
rect 24780 6836 24781 6900
rect 24715 6835 24781 6836
rect 29315 6900 29381 6901
rect 29315 6836 29316 6900
rect 29380 6836 29381 6900
rect 29315 6835 29381 6836
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 30235 6356 30301 6357
rect 30235 6292 30236 6356
rect 30300 6292 30301 6356
rect 30235 6291 30301 6292
rect 26187 5676 26253 5677
rect 26187 5612 26188 5676
rect 26252 5612 26253 5676
rect 26187 5611 26253 5612
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 7971 4044 8037 4045
rect 7971 3980 7972 4044
rect 8036 3980 8037 4044
rect 7971 3979 8037 3980
rect 19011 4044 19077 4045
rect 19011 3980 19012 4044
rect 19076 3980 19077 4044
rect 19011 3979 19077 3980
rect 4843 3500 4909 3501
rect 4843 3436 4844 3500
rect 4908 3436 4909 3500
rect 4843 3435 4909 3436
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 26190 2957 26250 5611
rect 30238 3501 30298 6291
rect 34654 4725 34714 12819
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34651 4724 34717 4725
rect 34651 4660 34652 4724
rect 34716 4660 34717 4724
rect 34651 4659 34717 4660
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 30235 3500 30301 3501
rect 30235 3436 30236 3500
rect 30300 3436 30301 3500
rect 30235 3435 30301 3436
rect 26187 2956 26253 2957
rect 26187 2892 26188 2956
rect 26252 2892 26253 2956
rect 26187 2891 26253 2892
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _0409_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0410_
timestamp 1688980957
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0411_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 38364 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0412_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0413_
timestamp 1688980957
transform -1 0 29440 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0414_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 32660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0415_
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0416_
timestamp 1688980957
transform 1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0417_
timestamp 1688980957
transform -1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0418_
timestamp 1688980957
transform -1 0 24288 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0419_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14720 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0420_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3220 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0421_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4600 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0422_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0423_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _0424_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4692 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__mux4_1  _0425_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0426_
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0427_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0428_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0429_
timestamp 1688980957
transform -1 0 8832 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0430_
timestamp 1688980957
transform 1 0 3312 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0431_
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0432_
timestamp 1688980957
transform -1 0 5980 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0433_
timestamp 1688980957
transform -1 0 8372 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0434_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0435_
timestamp 1688980957
transform 1 0 5428 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0436_
timestamp 1688980957
transform 1 0 3220 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0437_
timestamp 1688980957
transform -1 0 8832 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0438_
timestamp 1688980957
transform 1 0 3404 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0439_
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0440_
timestamp 1688980957
transform 1 0 7636 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0441_
timestamp 1688980957
transform -1 0 11408 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0442_
timestamp 1688980957
transform 1 0 9476 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0443_
timestamp 1688980957
transform 1 0 10764 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0444_
timestamp 1688980957
transform 1 0 9108 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0445_
timestamp 1688980957
transform 1 0 8188 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0446_
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0447_
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0448_
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0449_
timestamp 1688980957
transform -1 0 13892 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0450_
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0451_
timestamp 1688980957
transform 1 0 13064 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0452_
timestamp 1688980957
transform 1 0 8372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0453_
timestamp 1688980957
transform -1 0 13984 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0454_
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0455_
timestamp 1688980957
transform 1 0 13156 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0456_
timestamp 1688980957
transform 1 0 11592 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0457_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0458_
timestamp 1688980957
transform -1 0 13708 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0459_
timestamp 1688980957
transform -1 0 13800 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0460_
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0461_
timestamp 1688980957
transform -1 0 16008 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0462_
timestamp 1688980957
transform 1 0 13892 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0463_
timestamp 1688980957
transform 1 0 15548 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0464_
timestamp 1688980957
transform 1 0 14536 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0465_
timestamp 1688980957
transform -1 0 18584 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0466_
timestamp 1688980957
transform -1 0 19320 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0467_
timestamp 1688980957
transform 1 0 17296 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0468_
timestamp 1688980957
transform -1 0 15732 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0469_
timestamp 1688980957
transform -1 0 18676 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0470_
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0471_
timestamp 1688980957
transform -1 0 17664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0472_
timestamp 1688980957
transform -1 0 19320 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0473_
timestamp 1688980957
transform -1 0 18952 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0474_
timestamp 1688980957
transform -1 0 18492 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0475_
timestamp 1688980957
transform -1 0 18952 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0476_
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0477_
timestamp 1688980957
transform 1 0 16836 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0478_
timestamp 1688980957
transform 1 0 17112 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0479_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0480_
timestamp 1688980957
transform 1 0 18676 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0481_
timestamp 1688980957
transform 1 0 18584 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0482_
timestamp 1688980957
transform 1 0 18676 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0483_
timestamp 1688980957
transform 1 0 20608 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0484_
timestamp 1688980957
transform 1 0 19780 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0485_
timestamp 1688980957
transform -1 0 23092 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0486_
timestamp 1688980957
transform -1 0 23368 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0487_
timestamp 1688980957
transform -1 0 23092 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0488_
timestamp 1688980957
transform -1 0 24288 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0489_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0490_
timestamp 1688980957
transform -1 0 23000 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0491_
timestamp 1688980957
transform -1 0 24196 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0492_
timestamp 1688980957
transform -1 0 24564 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0493_
timestamp 1688980957
transform 1 0 21988 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0494_
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0495_
timestamp 1688980957
transform -1 0 26036 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0496_
timestamp 1688980957
transform -1 0 25944 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0497_
timestamp 1688980957
transform -1 0 27600 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0498_
timestamp 1688980957
transform -1 0 27416 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0499_
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0500_
timestamp 1688980957
transform -1 0 26772 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0501_
timestamp 1688980957
transform -1 0 24840 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0502_
timestamp 1688980957
transform 1 0 22632 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0503_
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0504_
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0505_
timestamp 1688980957
transform -1 0 28888 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0506_
timestamp 1688980957
transform -1 0 28888 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0507_
timestamp 1688980957
transform 1 0 27784 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0508_
timestamp 1688980957
transform -1 0 28152 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0509_
timestamp 1688980957
transform -1 0 30452 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0510_
timestamp 1688980957
transform 1 0 24840 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0511_
timestamp 1688980957
transform -1 0 28612 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0512_
timestamp 1688980957
transform -1 0 32016 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0513_
timestamp 1688980957
transform -1 0 29072 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0514_
timestamp 1688980957
transform 1 0 27140 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0515_
timestamp 1688980957
transform -1 0 29348 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0516_
timestamp 1688980957
transform 1 0 28980 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0517_
timestamp 1688980957
transform -1 0 31464 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0518_
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1688980957
transform -1 0 30452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0520_
timestamp 1688980957
transform -1 0 34132 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0521_
timestamp 1688980957
transform -1 0 32384 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0522_
timestamp 1688980957
transform -1 0 32660 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1688980957
transform -1 0 32936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0524_
timestamp 1688980957
transform -1 0 35972 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0525_
timestamp 1688980957
transform -1 0 34040 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0526_
timestamp 1688980957
transform -1 0 34040 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0527_
timestamp 1688980957
transform -1 0 33764 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0528_
timestamp 1688980957
transform -1 0 35144 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0529_
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0530_
timestamp 1688980957
transform 1 0 30452 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0531_
timestamp 1688980957
transform -1 0 32936 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0532_
timestamp 1688980957
transform 1 0 34132 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0533_
timestamp 1688980957
transform -1 0 37168 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0534_
timestamp 1688980957
transform -1 0 37076 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0535_
timestamp 1688980957
transform -1 0 37076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0536_
timestamp 1688980957
transform -1 0 38456 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0537_
timestamp 1688980957
transform -1 0 37168 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0538_
timestamp 1688980957
transform -1 0 37720 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1688980957
transform -1 0 37168 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0540_
timestamp 1688980957
transform -1 0 38548 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0541_
timestamp 1688980957
transform -1 0 37168 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0542_
timestamp 1688980957
transform -1 0 37444 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0543_
timestamp 1688980957
transform -1 0 38088 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0544_
timestamp 1688980957
transform -1 0 38456 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0545_
timestamp 1688980957
transform 1 0 35052 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0546_
timestamp 1688980957
transform -1 0 37076 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0547_
timestamp 1688980957
transform -1 0 38088 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0548_
timestamp 1688980957
transform -1 0 38456 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0549_
timestamp 1688980957
transform -1 0 37720 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0550_
timestamp 1688980957
transform 1 0 33580 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp 1688980957
transform -1 0 38088 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0552_
timestamp 1688980957
transform -1 0 38456 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0553_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0554_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0555_
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0556_
timestamp 1688980957
transform -1 0 14444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0557_
timestamp 1688980957
transform -1 0 12420 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1688980957
transform -1 0 15180 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1688980957
transform -1 0 17480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1688980957
transform -1 0 18124 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1688980957
transform 1 0 18768 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1688980957
transform -1 0 23644 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 1688980957
transform 1 0 22172 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1688980957
transform -1 0 27784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0568_
timestamp 1688980957
transform -1 0 24012 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1688980957
transform -1 0 28428 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1688980957
transform 1 0 30452 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1688980957
transform -1 0 29256 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0572_
timestamp 1688980957
transform -1 0 31280 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0573_
timestamp 1688980957
transform 1 0 32384 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1688980957
transform -1 0 32936 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0575_
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1688980957
transform -1 0 36800 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0577_
timestamp 1688980957
transform -1 0 36892 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0578_
timestamp 1688980957
transform -1 0 38088 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 1688980957
transform -1 0 36340 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1688980957
transform -1 0 37168 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0581_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _0582_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0583_
timestamp 1688980957
transform -1 0 7176 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0587_
timestamp 1688980957
transform 1 0 10764 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1688980957
transform 1 0 10120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1688980957
transform 1 0 13892 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1688980957
transform 1 0 12972 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 1688980957
transform -1 0 13340 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1688980957
transform 1 0 15548 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1688980957
transform 1 0 18676 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1688980957
transform -1 0 18952 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1688980957
transform -1 0 18492 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1688980957
transform -1 0 20516 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1688980957
transform -1 0 22448 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1688980957
transform -1 0 23460 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1688980957
transform -1 0 24012 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1688980957
transform -1 0 27784 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1688980957
transform 1 0 24840 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1688980957
transform -1 0 29716 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1688980957
transform -1 0 29992 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0606_
timestamp 1688980957
transform -1 0 31188 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1688980957
transform 1 0 32936 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1688980957
transform -1 0 33856 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1688980957
transform -1 0 33764 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 1688980957
transform 1 0 37628 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0611_
timestamp 1688980957
transform 1 0 37260 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0612_
timestamp 1688980957
transform 1 0 37076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1688980957
transform -1 0 38088 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1688980957
transform -1 0 38088 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_1  _0615_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3036 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0616_
timestamp 1688980957
transform 1 0 3772 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0617_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1688980957
transform 1 0 2760 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1688980957
transform 1 0 3128 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1688980957
transform -1 0 3680 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1688980957
transform 1 0 3220 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1688980957
transform 1 0 10212 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1688980957
transform 1 0 8648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0625_
timestamp 1688980957
transform 1 0 11776 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1688980957
transform 1 0 12144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1688980957
transform 1 0 13156 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1688980957
transform 1 0 17112 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1688980957
transform -1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1688980957
transform 1 0 16928 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1688980957
transform 1 0 18308 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1688980957
transform -1 0 23184 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform 1 0 26036 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform -1 0 26864 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1688980957
transform 1 0 24564 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1688980957
transform -1 0 29256 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1688980957
transform 1 0 25852 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 30636 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0644_
timestamp 1688980957
transform 1 0 30728 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0646_
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0647_
timestamp 1688980957
transform 1 0 35696 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0648_
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 1688980957
transform -1 0 35512 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0650_
timestamp 1688980957
transform 1 0 4232 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0651_
timestamp 1688980957
transform 1 0 2760 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0652_
timestamp 1688980957
transform -1 0 4600 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0653_
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0654_
timestamp 1688980957
transform 1 0 4600 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 1688980957
transform 1 0 10948 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0656_
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0657_
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1688980957
transform 1 0 10856 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0659_
timestamp 1688980957
transform 1 0 10580 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0660_
timestamp 1688980957
transform 1 0 13156 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0661_
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0662_
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0663_
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0664_
timestamp 1688980957
transform 1 0 16744 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0665_
timestamp 1688980957
transform 1 0 18308 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0666_
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1688980957
transform 1 0 20884 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0668_
timestamp 1688980957
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1688980957
transform 1 0 24656 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0670_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0671_
timestamp 1688980957
transform 1 0 26864 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform -1 0 26680 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0673_
timestamp 1688980957
transform 1 0 26036 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0674_
timestamp 1688980957
transform 1 0 25760 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0675_
timestamp 1688980957
transform 1 0 30452 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0676_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1688980957
transform 1 0 29624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1688980957
transform -1 0 34592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1688980957
transform 1 0 34960 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0681_
timestamp 1688980957
transform 1 0 34040 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0682_
timestamp 1688980957
transform 1 0 32752 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0683_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0685_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1688980957
transform -1 0 2208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1688980957
transform 1 0 2944 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1688980957
transform 1 0 9752 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1688980957
transform 1 0 8096 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1688980957
transform -1 0 12420 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1688980957
transform -1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1688980957
transform -1 0 18952 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1688980957
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1688980957
transform -1 0 17940 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1688980957
transform 1 0 19044 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1688980957
transform -1 0 19780 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1688980957
transform -1 0 22724 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1688980957
transform 1 0 23276 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0701_
timestamp 1688980957
transform 1 0 25576 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1688980957
transform -1 0 26680 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1688980957
transform -1 0 24288 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1688980957
transform -1 0 26864 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1688980957
transform -1 0 26680 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1688980957
transform 1 0 27324 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1688980957
transform -1 0 27784 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1688980957
transform -1 0 33488 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1688980957
transform -1 0 33580 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1688980957
transform -1 0 31740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1688980957
transform -1 0 36248 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1688980957
transform -1 0 36800 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1688980957
transform -1 0 36524 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1688980957
transform 1 0 33488 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _0716_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5612 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0717_
timestamp 1688980957
transform 1 0 3956 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1688980957
transform -1 0 4600 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform -1 0 12328 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0722_
timestamp 1688980957
transform -1 0 9752 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1688980957
transform -1 0 12880 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1688980957
transform -1 0 14628 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1688980957
transform 1 0 14444 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1688980957
transform -1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1688980957
transform 1 0 14904 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1688980957
transform -1 0 17756 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1688980957
transform -1 0 19136 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1688980957
transform -1 0 20148 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1688980957
transform -1 0 23552 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0733_
timestamp 1688980957
transform -1 0 23092 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1688980957
transform 1 0 25208 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1688980957
transform -1 0 27784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1688980957
transform -1 0 25392 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1688980957
transform -1 0 30084 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform -1 0 27784 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1688980957
transform -1 0 32936 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform 1 0 34040 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1688980957
transform 1 0 32384 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0745_
timestamp 1688980957
transform 1 0 37720 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform -1 0 36340 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_2  _0749_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0750_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0751_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0752_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0753_
timestamp 1688980957
transform 1 0 3128 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0754_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0755_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4876 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0756_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0757_
timestamp 1688980957
transform -1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0758_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0759_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5888 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0760_
timestamp 1688980957
transform -1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0761_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0762_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3220 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_4  _0763_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1688980957
transform -1 0 4784 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1688980957
transform 1 0 6164 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1688980957
transform -1 0 9016 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 1688980957
transform -1 0 7176 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1688980957
transform 1 0 9476 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1688980957
transform 1 0 7360 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1688980957
transform 1 0 12052 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 1688980957
transform -1 0 18676 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1688980957
transform -1 0 17020 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1688980957
transform -1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1688980957
transform 1 0 18308 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1688980957
transform -1 0 22632 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1688980957
transform -1 0 26404 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1688980957
transform 1 0 22724 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1688980957
transform -1 0 30360 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1688980957
transform -1 0 28520 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1688980957
transform -1 0 30360 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1688980957
transform 1 0 32200 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1688980957
transform 1 0 29808 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1688980957
transform 1 0 34960 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1688980957
transform -1 0 35880 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1688980957
transform -1 0 36156 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0796_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0797_
timestamp 1688980957
transform 1 0 2116 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0798_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0799_
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0800_
timestamp 1688980957
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0801_
timestamp 1688980957
transform -1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0802_
timestamp 1688980957
transform -1 0 4048 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0803_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _0804_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0805_
timestamp 1688980957
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0806_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0807_
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0808_
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0809_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0810_
timestamp 1688980957
transform -1 0 5888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0811_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0812_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1688980957
transform -1 0 5152 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1688980957
transform -1 0 6900 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1688980957
transform 1 0 6992 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1688980957
transform 1 0 11040 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1688980957
transform 1 0 6532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 1688980957
transform 1 0 12972 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 1688980957
transform 1 0 15088 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1688980957
transform 1 0 15364 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1688980957
transform 1 0 18216 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 1688980957
transform 1 0 20884 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform 1 0 20516 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1688980957
transform -1 0 25668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp 1688980957
transform -1 0 24196 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0834_
timestamp 1688980957
transform 1 0 28336 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1688980957
transform 1 0 26864 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 1688980957
transform 1 0 29624 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 1688980957
transform 1 0 31372 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp 1688980957
transform 1 0 30912 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 1688980957
transform -1 0 34592 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp 1688980957
transform -1 0 35236 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1688980957
transform 1 0 34776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0843_
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1688980957
transform 1 0 5428 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1688980957
transform -1 0 6256 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0847_
timestamp 1688980957
transform -1 0 7912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1688980957
transform 1 0 7360 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1688980957
transform 1 0 8464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _0851_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0852_
timestamp 1688980957
transform -1 0 13340 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0853_
timestamp 1688980957
transform -1 0 12512 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0854_
timestamp 1688980957
transform 1 0 13800 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0855_
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0856_
timestamp 1688980957
transform 1 0 16744 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0857_
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0858_
timestamp 1688980957
transform -1 0 18124 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0859_
timestamp 1688980957
transform 1 0 18216 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0860_
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0861_
timestamp 1688980957
transform -1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1688980957
transform 1 0 25392 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1688980957
transform -1 0 25852 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1688980957
transform 1 0 26128 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1688980957
transform -1 0 30084 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1688980957
transform 1 0 28980 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1688980957
transform 1 0 31004 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1688980957
transform 1 0 32384 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1688980957
transform -1 0 31740 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1688980957
transform 1 0 36156 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1688980957
transform -1 0 37904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1688980957
transform 1 0 35604 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1688980957
transform -1 0 36156 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1688980957
transform 1 0 36340 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1688980957
transform -1 0 6256 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1688980957
transform 1 0 6716 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1688980957
transform 1 0 7176 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1688980957
transform 1 0 9568 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1688980957
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1688980957
transform 1 0 12144 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1688980957
transform -1 0 13616 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1688980957
transform -1 0 12880 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1688980957
transform 1 0 17112 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1688980957
transform -1 0 18032 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1688980957
transform -1 0 20700 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1688980957
transform 1 0 21804 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1688980957
transform -1 0 22816 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1688980957
transform -1 0 23368 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1688980957
transform -1 0 29072 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1688980957
transform 1 0 23644 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1688980957
transform -1 0 28888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1688980957
transform -1 0 31004 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1688980957
transform 1 0 27140 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1688980957
transform -1 0 31556 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1688980957
transform 1 0 30452 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1688980957
transform -1 0 32660 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1688980957
transform -1 0 37628 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1688980957
transform 1 0 36800 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1688980957
transform 1 0 36340 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1688980957
transform 1 0 36340 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1688980957
transform 1 0 1932 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1688980957
transform 1 0 2208 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1688980957
transform 1 0 2300 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1688980957
transform 1 0 2208 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1688980957
transform 1 0 8004 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1688980957
transform 1 0 9936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1688980957
transform 1 0 10304 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1688980957
transform 1 0 12420 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1688980957
transform 1 0 16192 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1688980957
transform 1 0 15088 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1688980957
transform 1 0 15732 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1688980957
transform -1 0 18676 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1688980957
transform 1 0 19596 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1688980957
transform -1 0 23368 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1688980957
transform 1 0 24840 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1688980957
transform 1 0 21988 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1688980957
transform 1 0 23368 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1688980957
transform 1 0 25208 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1688980957
transform -1 0 31556 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1688980957
transform 1 0 31096 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1688980957
transform 1 0 29440 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1688980957
transform 1 0 34132 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1688980957
transform -1 0 36708 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1688980957
transform 1 0 33488 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1688980957
transform 1 0 32476 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1688980957
transform -1 0 3496 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1688980957
transform 1 0 2300 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1688980957
transform 1 0 2208 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1688980957
transform 1 0 2208 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1688980957
transform 1 0 8740 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1688980957
transform 1 0 9936 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1688980957
transform -1 0 11960 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1688980957
transform 1 0 13064 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1688980957
transform 1 0 11040 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1688980957
transform -1 0 17112 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1688980957
transform -1 0 16560 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1688980957
transform 1 0 20240 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1688980957
transform -1 0 21712 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1688980957
transform 1 0 21620 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1688980957
transform 1 0 24564 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1688980957
transform 1 0 21804 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1688980957
transform 1 0 26036 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1688980957
transform 1 0 25668 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1688980957
transform 1 0 25024 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1688980957
transform 1 0 29900 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1688980957
transform 1 0 30544 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1688980957
transform 1 0 29256 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1688980957
transform 1 0 33856 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1688980957
transform 1 0 35052 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1688980957
transform -1 0 35696 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1688980957
transform 1 0 33120 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1688980957
transform 1 0 32292 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1688980957
transform 1 0 2208 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1688980957
transform 1 0 2208 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1688980957
transform 1 0 2208 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1688980957
transform 1 0 1932 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1688980957
transform -1 0 10764 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1688980957
transform -1 0 8832 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1688980957
transform -1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1688980957
transform -1 0 13156 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1688980957
transform -1 0 15548 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1688980957
transform -1 0 19136 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1688980957
transform -1 0 13984 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1688980957
transform -1 0 18308 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1688980957
transform -1 0 20700 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1688980957
transform -1 0 23276 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1688980957
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1688980957
transform -1 0 23736 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1688980957
transform 1 0 25392 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1688980957
transform -1 0 23276 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1688980957
transform -1 0 28980 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1688980957
transform -1 0 25852 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1688980957
transform -1 0 33580 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1688980957
transform 1 0 31280 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1688980957
transform -1 0 31372 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1688980957
transform 1 0 35328 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1688980957
transform 1 0 35604 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1688980957
transform 1 0 35512 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1688980957
transform 1 0 35052 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1688980957
transform 1 0 32752 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1688980957
transform -1 0 4876 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1688980957
transform 1 0 1840 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1688980957
transform -1 0 5244 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1688980957
transform -1 0 10948 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1688980957
transform -1 0 8832 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1688980957
transform -1 0 13064 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1688980957
transform -1 0 13524 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1688980957
transform -1 0 15548 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1688980957
transform -1 0 20792 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1688980957
transform -1 0 13984 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1688980957
transform -1 0 18676 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1688980957
transform -1 0 20700 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1688980957
transform -1 0 24840 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1688980957
transform -1 0 28888 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1688980957
transform -1 0 23920 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1688980957
transform 1 0 26496 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1688980957
transform -1 0 28520 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1688980957
transform -1 0 28152 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1688980957
transform -1 0 33028 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1688980957
transform -1 0 34040 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1688980957
transform -1 0 32016 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1688980957
transform 1 0 37076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1688980957
transform -1 0 38180 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1688980957
transform 1 0 36248 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1688980957
transform 1 0 37076 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1688980957
transform -1 0 35236 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1688980957
transform -1 0 4600 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1688980957
transform -1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1688980957
transform -1 0 3680 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1688980957
transform -1 0 7820 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1688980957
transform 1 0 6164 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1688980957
transform -1 0 10120 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1688980957
transform 1 0 8004 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1688980957
transform 1 0 7360 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1688980957
transform 1 0 11592 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1688980957
transform 1 0 9936 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1688980957
transform 1 0 12512 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1688980957
transform 1 0 16652 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1688980957
transform 1 0 17664 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1688980957
transform 1 0 19688 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1688980957
transform -1 0 24104 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1688980957
transform 1 0 25024 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1688980957
transform 1 0 22172 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1688980957
transform 1 0 25944 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1688980957
transform 1 0 27968 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1688980957
transform -1 0 31280 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1688980957
transform 1 0 30452 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1688980957
transform 1 0 30912 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1688980957
transform 1 0 29716 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1688980957
transform 1 0 34408 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1688980957
transform 1 0 35144 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1688980957
transform 1 0 34684 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1688980957
transform 1 0 33120 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1688980957
transform 1 0 35512 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1688980957
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1073_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1074_
timestamp 1688980957
transform 1 0 2576 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1075_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1688980957
transform -1 0 8280 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1077_
timestamp 1688980957
transform 1 0 7176 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1688980957
transform -1 0 7820 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1688980957
transform 1 0 6624 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1688980957
transform 1 0 5612 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1688980957
transform -1 0 8004 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1688980957
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1688980957
transform 1 0 10580 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1688980957
transform 1 0 9936 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1688980957
transform 1 0 14812 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1688980957
transform -1 0 16560 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1688980957
transform 1 0 15088 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1688980957
transform 1 0 15088 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1688980957
transform 1 0 17112 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1688980957
transform 1 0 20240 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1688980957
transform -1 0 21988 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1688980957
transform 1 0 24656 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1688980957
transform 1 0 21896 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1688980957
transform 1 0 25392 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1688980957
transform 1 0 27876 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1688980957
transform 1 0 26220 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1688980957
transform 1 0 27968 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1688980957
transform 1 0 30544 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1688980957
transform 1 0 34960 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1688980957
transform 1 0 33764 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1688980957
transform 1 0 33304 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1688980957
transform 1 0 34040 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1688980957
transform 1 0 4968 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1688980957
transform -1 0 8372 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1688980957
transform 1 0 6440 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1688980957
transform 1 0 6992 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1688980957
transform 1 0 9292 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1688980957
transform -1 0 9384 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0422__B asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__A
timestamp 1688980957
transform -1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0425__S0
timestamp 1688980957
transform 1 0 8004 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0425__S1
timestamp 1688980957
transform 1 0 7728 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0426__S0
timestamp 1688980957
transform 1 0 5888 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0426__S1
timestamp 1688980957
transform 1 0 5704 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__S
timestamp 1688980957
transform 1 0 7360 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__B
timestamp 1688980957
transform -1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0429__S0
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0429__S1
timestamp 1688980957
transform 1 0 10580 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__S0
timestamp 1688980957
transform 1 0 5428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__S1
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0431__S
timestamp 1688980957
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0433__S0
timestamp 1688980957
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0433__S1
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__S0
timestamp 1688980957
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__S1
timestamp 1688980957
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0435__S
timestamp 1688980957
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0437__S0
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0437__S1
timestamp 1688980957
transform 1 0 10304 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__S0
timestamp 1688980957
transform 1 0 5520 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__S1
timestamp 1688980957
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0439__S
timestamp 1688980957
transform 1 0 7820 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0441__S0
timestamp 1688980957
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0441__S1
timestamp 1688980957
transform -1 0 9292 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__S0
timestamp 1688980957
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__S1
timestamp 1688980957
transform 1 0 9292 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__S
timestamp 1688980957
transform 1 0 9108 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__B
timestamp 1688980957
transform -1 0 8004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0445__S0
timestamp 1688980957
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0445__S1
timestamp 1688980957
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__S0
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__S1
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__S
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__S0
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__S1
timestamp 1688980957
transform 1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__S0
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__S1
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__S
timestamp 1688980957
transform -1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__S0
timestamp 1688980957
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__S1
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__S0
timestamp 1688980957
transform 1 0 12052 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__S1
timestamp 1688980957
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__S
timestamp 1688980957
transform 1 0 13800 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0457__S0
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0457__S1
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__S0
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__S1
timestamp 1688980957
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__S
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0461__S0
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0461__S1
timestamp 1688980957
transform 1 0 13432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__S0
timestamp 1688980957
transform 1 0 13524 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__S1
timestamp 1688980957
transform 1 0 13708 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__S
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__B
timestamp 1688980957
transform 1 0 14720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__S0
timestamp 1688980957
transform -1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__S1
timestamp 1688980957
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__S0
timestamp 1688980957
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__S1
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__S
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__S0
timestamp 1688980957
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__S1
timestamp 1688980957
transform 1 0 15824 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__S0
timestamp 1688980957
transform 1 0 11960 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__S1
timestamp 1688980957
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__S
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__S0
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__S1
timestamp 1688980957
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__S0
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__S1
timestamp 1688980957
transform 1 0 18676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__S
timestamp 1688980957
transform 1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__S0
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__S1
timestamp 1688980957
transform 1 0 14904 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__S0
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__S1
timestamp 1688980957
transform 1 0 16928 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__S
timestamp 1688980957
transform -1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__S0
timestamp 1688980957
transform -1 0 17112 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__S1
timestamp 1688980957
transform -1 0 17664 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__S0
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__S1
timestamp 1688980957
transform 1 0 17020 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__S
timestamp 1688980957
transform 1 0 20884 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__B
timestamp 1688980957
transform -1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__S0
timestamp 1688980957
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__S1
timestamp 1688980957
transform 1 0 24104 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__S0
timestamp 1688980957
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__S1
timestamp 1688980957
transform 1 0 23552 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__S
timestamp 1688980957
transform 1 0 24196 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__S0
timestamp 1688980957
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__S1
timestamp 1688980957
transform 1 0 24564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__S0
timestamp 1688980957
transform -1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__S1
timestamp 1688980957
transform -1 0 28152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__S
timestamp 1688980957
transform -1 0 20700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__S0
timestamp 1688980957
transform 1 0 24564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__S1
timestamp 1688980957
transform 1 0 24196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__S0
timestamp 1688980957
transform 1 0 26220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__S1
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__S
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__S0
timestamp 1688980957
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__S1
timestamp 1688980957
transform 1 0 27968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__S0
timestamp 1688980957
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__S1
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__S
timestamp 1688980957
transform 1 0 27508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__S0
timestamp 1688980957
transform 1 0 25852 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__S1
timestamp 1688980957
transform 1 0 24840 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__S0
timestamp 1688980957
transform 1 0 26036 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__S1
timestamp 1688980957
transform 1 0 25576 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__S
timestamp 1688980957
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__S0
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__S1
timestamp 1688980957
transform 1 0 26956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__S0
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__S1
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__S
timestamp 1688980957
transform 1 0 28060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__S0
timestamp 1688980957
transform 1 0 28152 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__S1
timestamp 1688980957
transform 1 0 28336 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__S0
timestamp 1688980957
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__S1
timestamp 1688980957
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__S
timestamp 1688980957
transform 1 0 27600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__S0
timestamp 1688980957
transform 1 0 26772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__S1
timestamp 1688980957
transform 1 0 27140 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__S0
timestamp 1688980957
transform 1 0 26772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__S1
timestamp 1688980957
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__S
timestamp 1688980957
transform -1 0 29348 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__S0
timestamp 1688980957
transform 1 0 29164 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__S1
timestamp 1688980957
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__S0
timestamp 1688980957
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__S1
timestamp 1688980957
transform 1 0 27232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__S
timestamp 1688980957
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__S0
timestamp 1688980957
transform 1 0 29992 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__S1
timestamp 1688980957
transform -1 0 30452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__S0
timestamp 1688980957
transform 1 0 30360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__S1
timestamp 1688980957
transform 1 0 29716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__S
timestamp 1688980957
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__S0
timestamp 1688980957
transform -1 0 31924 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__S1
timestamp 1688980957
transform 1 0 34224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__S0
timestamp 1688980957
transform 1 0 30912 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__S1
timestamp 1688980957
transform 1 0 31464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__S
timestamp 1688980957
transform 1 0 32752 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__B
timestamp 1688980957
transform 1 0 34500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__S0
timestamp 1688980957
transform 1 0 30084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__S1
timestamp 1688980957
transform 1 0 33028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__S0
timestamp 1688980957
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__S1
timestamp 1688980957
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__S
timestamp 1688980957
transform 1 0 32660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__S0
timestamp 1688980957
transform 1 0 33672 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__S1
timestamp 1688980957
transform 1 0 31556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__S0
timestamp 1688980957
transform 1 0 29348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__S1
timestamp 1688980957
transform 1 0 28520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__S
timestamp 1688980957
transform 1 0 29900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__S0
timestamp 1688980957
transform 1 0 34868 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__S1
timestamp 1688980957
transform 1 0 35236 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__S0
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__S1
timestamp 1688980957
transform 1 0 36708 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__S
timestamp 1688980957
transform 1 0 35052 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__B
timestamp 1688980957
transform 1 0 38180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__S0
timestamp 1688980957
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__S1
timestamp 1688980957
transform 1 0 33580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__S0
timestamp 1688980957
transform -1 0 36892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__S1
timestamp 1688980957
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__S
timestamp 1688980957
transform 1 0 37720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__S0
timestamp 1688980957
transform 1 0 32752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__S1
timestamp 1688980957
transform 1 0 33120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__S0
timestamp 1688980957
transform -1 0 36892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__S1
timestamp 1688980957
transform 1 0 32936 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__S
timestamp 1688980957
transform -1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__S0
timestamp 1688980957
transform 1 0 35420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__S1
timestamp 1688980957
transform -1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__S0
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__S1
timestamp 1688980957
transform 1 0 34132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__S
timestamp 1688980957
transform -1 0 13156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__S
timestamp 1688980957
transform 1 0 13524 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__S
timestamp 1688980957
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__S
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__S
timestamp 1688980957
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__S
timestamp 1688980957
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__S
timestamp 1688980957
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__S
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__S
timestamp 1688980957
transform 1 0 20240 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__S
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__S
timestamp 1688980957
transform 1 0 23828 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__S
timestamp 1688980957
transform 1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__S
timestamp 1688980957
transform 1 0 28704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__S
timestamp 1688980957
transform 1 0 23000 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__S
timestamp 1688980957
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__S
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__S
timestamp 1688980957
transform 1 0 29716 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__S
timestamp 1688980957
transform 1 0 30636 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__S
timestamp 1688980957
transform 1 0 33396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__S
timestamp 1688980957
transform 1 0 31096 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__S
timestamp 1688980957
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__S
timestamp 1688980957
transform -1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__S
timestamp 1688980957
transform 1 0 35880 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__S
timestamp 1688980957
transform -1 0 38456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__S
timestamp 1688980957
transform 1 0 33304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__S
timestamp 1688980957
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__S
timestamp 1688980957
transform 1 0 7360 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__S
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__S
timestamp 1688980957
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__S
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__S
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__S
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__S
timestamp 1688980957
transform -1 0 13984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__S
timestamp 1688980957
transform 1 0 13984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__S
timestamp 1688980957
transform 1 0 13524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__S
timestamp 1688980957
transform 1 0 16192 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__S
timestamp 1688980957
transform 1 0 18400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__S
timestamp 1688980957
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__S
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__S
timestamp 1688980957
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1688980957
transform -1 0 19688 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__S
timestamp 1688980957
transform 1 0 22448 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1688980957
transform -1 0 24748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__S
timestamp 1688980957
transform 1 0 24564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1688980957
transform 1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__S
timestamp 1688980957
transform 1 0 24656 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1688980957
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__S
timestamp 1688980957
transform 1 0 28888 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1688980957
transform 1 0 30544 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__S
timestamp 1688980957
transform -1 0 31556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__S
timestamp 1688980957
transform 1 0 33856 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__S
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__S
timestamp 1688980957
transform 1 0 38180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__S
timestamp 1688980957
transform -1 0 38456 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__S
timestamp 1688980957
transform 1 0 38088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__S
timestamp 1688980957
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__S
timestamp 1688980957
transform 1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__S
timestamp 1688980957
transform 1 0 4692 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__S
timestamp 1688980957
transform -1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__S
timestamp 1688980957
transform 1 0 5060 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__S
timestamp 1688980957
transform 1 0 9844 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__S
timestamp 1688980957
transform 1 0 8464 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__S
timestamp 1688980957
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__S
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__S
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__S
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__S
timestamp 1688980957
transform 1 0 16928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__S
timestamp 1688980957
transform 1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__S
timestamp 1688980957
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__S
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__S
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__S
timestamp 1688980957
transform 1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1688980957
transform 1 0 21620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__S
timestamp 1688980957
transform 1 0 24564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__S
timestamp 1688980957
transform 1 0 33028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__S
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__S
timestamp 1688980957
transform 1 0 27324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__S
timestamp 1688980957
transform 1 0 24564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__S
timestamp 1688980957
transform 1 0 28336 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__S
timestamp 1688980957
transform 1 0 25668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__S
timestamp 1688980957
transform 1 0 30452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__S
timestamp 1688980957
transform -1 0 31280 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__S
timestamp 1688980957
transform 1 0 29716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__S
timestamp 1688980957
transform 1 0 28980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__S
timestamp 1688980957
transform -1 0 38456 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__S
timestamp 1688980957
transform 1 0 34040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__S
timestamp 1688980957
transform 1 0 34868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__S
timestamp 1688980957
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__S
timestamp 1688980957
transform 1 0 1840 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__S
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__S
timestamp 1688980957
transform -1 0 1932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__S
timestamp 1688980957
transform 1 0 5704 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__S
timestamp 1688980957
transform 1 0 10948 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__S
timestamp 1688980957
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__S
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__S
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__S
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__S
timestamp 1688980957
transform -1 0 12972 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__S
timestamp 1688980957
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__S
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__S
timestamp 1688980957
transform 1 0 15088 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__S
timestamp 1688980957
transform 1 0 15640 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__S
timestamp 1688980957
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__S
timestamp 1688980957
transform 1 0 21712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__S
timestamp 1688980957
transform -1 0 20148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__S
timestamp 1688980957
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__S
timestamp 1688980957
transform 1 0 29072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__S
timestamp 1688980957
transform -1 0 22448 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__S
timestamp 1688980957
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__S
timestamp 1688980957
transform 1 0 25668 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__S
timestamp 1688980957
transform 1 0 26404 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__S
timestamp 1688980957
transform 1 0 25576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__S
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__S
timestamp 1688980957
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__S
timestamp 1688980957
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__S
timestamp 1688980957
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__S
timestamp 1688980957
transform 1 0 34868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__S
timestamp 1688980957
transform 1 0 34040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__S
timestamp 1688980957
transform -1 0 33304 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__S
timestamp 1688980957
transform 1 0 32568 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__S
timestamp 1688980957
transform -1 0 4876 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__S
timestamp 1688980957
transform 1 0 4876 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__S
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__S
timestamp 1688980957
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__S
timestamp 1688980957
transform 1 0 8832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__S
timestamp 1688980957
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__S
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__S
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__S
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__S
timestamp 1688980957
transform 1 0 14352 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__S
timestamp 1688980957
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__S
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__S
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__S
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__S
timestamp 1688980957
transform -1 0 19044 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__S
timestamp 1688980957
transform 1 0 24564 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__S
timestamp 1688980957
transform -1 0 19872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__S
timestamp 1688980957
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__S
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__S
timestamp 1688980957
transform -1 0 23920 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__S
timestamp 1688980957
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__S
timestamp 1688980957
transform 1 0 27600 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__S
timestamp 1688980957
transform 1 0 27140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__S
timestamp 1688980957
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__S
timestamp 1688980957
transform 1 0 32476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__S
timestamp 1688980957
transform 1 0 34868 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__S
timestamp 1688980957
transform 1 0 30728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__S
timestamp 1688980957
transform 1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__S
timestamp 1688980957
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__S
timestamp 1688980957
transform -1 0 38456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__S
timestamp 1688980957
transform -1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__S
timestamp 1688980957
transform 1 0 32476 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__S
timestamp 1688980957
transform 1 0 4784 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__S
timestamp 1688980957
transform 1 0 4692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__S
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__S
timestamp 1688980957
transform 1 0 4692 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__S
timestamp 1688980957
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__S
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__S
timestamp 1688980957
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__S
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__S
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__S
timestamp 1688980957
transform -1 0 14444 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__S
timestamp 1688980957
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__S
timestamp 1688980957
transform 1 0 15272 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__S
timestamp 1688980957
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__S
timestamp 1688980957
transform 1 0 18584 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__S
timestamp 1688980957
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__S
timestamp 1688980957
transform 1 0 24288 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__S
timestamp 1688980957
transform -1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__S
timestamp 1688980957
transform 1 0 26036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__S
timestamp 1688980957
transform 1 0 29716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__S
timestamp 1688980957
transform -1 0 25760 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S
timestamp 1688980957
transform 1 0 27968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__S
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__S
timestamp 1688980957
transform 1 0 27600 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S
timestamp 1688980957
transform 1 0 31924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__S
timestamp 1688980957
transform 1 0 34224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__S
timestamp 1688980957
transform 1 0 33028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__S
timestamp 1688980957
transform 1 0 28152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__S
timestamp 1688980957
transform -1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S
timestamp 1688980957
transform 1 0 37076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S
timestamp 1688980957
transform -1 0 38456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__S
timestamp 1688980957
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__S
timestamp 1688980957
transform 1 0 4508 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S
timestamp 1688980957
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__S
timestamp 1688980957
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__S
timestamp 1688980957
transform -1 0 10488 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S
timestamp 1688980957
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__S
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S
timestamp 1688980957
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__S
timestamp 1688980957
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__S
timestamp 1688980957
transform -1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__S
timestamp 1688980957
transform 1 0 16652 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__S
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S
timestamp 1688980957
transform 1 0 23368 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__S
timestamp 1688980957
transform -1 0 23368 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__S
timestamp 1688980957
transform 1 0 25300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S
timestamp 1688980957
transform 1 0 28060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S
timestamp 1688980957
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__S
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__S
timestamp 1688980957
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S
timestamp 1688980957
transform -1 0 27508 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S
timestamp 1688980957
transform -1 0 29532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp 1688980957
transform 1 0 32292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__S
timestamp 1688980957
transform 1 0 30728 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S
timestamp 1688980957
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S
timestamp 1688980957
transform 1 0 31188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp 1688980957
transform -1 0 38456 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__S
timestamp 1688980957
transform 1 0 34868 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S
timestamp 1688980957
transform 1 0 35604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S
timestamp 1688980957
transform -1 0 38456 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__D
timestamp 1688980957
transform -1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A1
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A1
timestamp 1688980957
transform -1 0 3680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1688980957
transform -1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A
timestamp 1688980957
transform -1 0 5336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__S
timestamp 1688980957
transform -1 0 4324 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__S
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__S
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__S
timestamp 1688980957
transform 1 0 8004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__S
timestamp 1688980957
transform 1 0 9384 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S
timestamp 1688980957
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S
timestamp 1688980957
transform -1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__S
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__S
timestamp 1688980957
transform 1 0 10488 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S
timestamp 1688980957
transform -1 0 12880 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__S
timestamp 1688980957
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__S
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__S
timestamp 1688980957
transform -1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__S
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__S
timestamp 1688980957
transform 1 0 17296 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__S
timestamp 1688980957
transform 1 0 21988 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__S
timestamp 1688980957
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__S
timestamp 1688980957
transform 1 0 21712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__S
timestamp 1688980957
transform -1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__S
timestamp 1688980957
transform 1 0 21712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__S
timestamp 1688980957
transform 1 0 25944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__S
timestamp 1688980957
transform 1 0 27784 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__S
timestamp 1688980957
transform -1 0 26864 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__S
timestamp 1688980957
transform 1 0 28704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__S
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__S
timestamp 1688980957
transform 1 0 30452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S
timestamp 1688980957
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__S
timestamp 1688980957
transform 1 0 34868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__S
timestamp 1688980957
transform 1 0 34868 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__S
timestamp 1688980957
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__S
timestamp 1688980957
transform 1 0 33672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__S
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__S
timestamp 1688980957
transform 1 0 7268 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__S
timestamp 1688980957
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__S
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__S
timestamp 1688980957
transform 1 0 8372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__S
timestamp 1688980957
transform 1 0 12788 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__S
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1688980957
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1688980957
transform 1 0 14260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1688980957
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1688980957
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1688980957
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1688980957
transform 1 0 24472 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1688980957
transform 1 0 25300 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1688980957
transform 1 0 26404 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1688980957
transform 1 0 30912 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1688980957
transform 1 0 35328 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1688980957
transform 1 0 34960 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1688980957
transform 1 0 29808 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1688980957
transform 1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1688980957
transform 1 0 29532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1688980957
transform 1 0 34316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1688980957
transform 1 0 32292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1688980957
transform 1 0 25300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1688980957
transform 1 0 25668 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1688980957
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1688980957
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform -1 0 24288 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1688980957
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 1688980957
transform 1 0 24656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 1688980957
transform 1 0 4508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 1688980957
transform -1 0 22172 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1688980957
transform -1 0 10212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 1688980957
transform -1 0 23736 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 1688980957
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 1688980957
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 1688980957
transform 1 0 19596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout123_A
timestamp 1688980957
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_A
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp 1688980957
transform 1 0 24932 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout129_A
timestamp 1688980957
transform -1 0 8372 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout130_A
timestamp 1688980957
transform 1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout131_A
timestamp 1688980957
transform 1 0 24564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold561_A
timestamp 1688980957
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold563_A
timestamp 1688980957
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 9660 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 28612 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1688980957
transform 1 0 4232 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1688980957
transform 1 0 11592 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1688980957
transform -1 0 5612 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1688980957
transform 1 0 4416 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1688980957
transform -1 0 13340 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1688980957
transform 1 0 17020 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1688980957
transform -1 0 23920 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1688980957
transform 1 0 23276 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1688980957
transform -1 0 26864 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1688980957
transform 1 0 31096 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1688980957
transform 1 0 35512 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1688980957
transform 1 0 27968 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1688980957
transform 1 0 25024 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1688980957
transform 1 0 30176 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1688980957
transform 1 0 34960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1688980957
transform 1 0 34408 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1688980957
transform -1 0 34132 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1688980957
transform -1 0 27876 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1688980957
transform 1 0 22172 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1688980957
transform 1 0 16008 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1688980957
transform -1 0 16560 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  fanout102 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23184 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout103
timestamp 1688980957
transform 1 0 3772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout104
timestamp 1688980957
transform 1 0 22080 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout105
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout106
timestamp 1688980957
transform 1 0 23276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout107
timestamp 1688980957
transform 1 0 10212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout108
timestamp 1688980957
transform 1 0 24840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout109
timestamp 1688980957
transform -1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout110 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21712 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout111
timestamp 1688980957
transform 1 0 4232 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout112
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout113
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout114
timestamp 1688980957
transform 1 0 23276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout115
timestamp 1688980957
transform 1 0 9108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout116
timestamp 1688980957
transform 1 0 22080 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout117
timestamp 1688980957
transform 1 0 9384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout121
timestamp 1688980957
transform -1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout122
timestamp 1688980957
transform 1 0 23368 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout123 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9292 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout124
timestamp 1688980957
transform 1 0 6808 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout125
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout126
timestamp 1688980957
transform -1 0 24288 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout127 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6440 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout128
timestamp 1688980957
transform -1 0 6256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout129
timestamp 1688980957
transform 1 0 8096 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout130
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout131
timestamp 1688980957
transform -1 0 24380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_116 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_120
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_200
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_204
timestamp 1688980957
transform 1 0 19872 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_406
timestamp 1688980957
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_44
timestamp 1688980957
transform 1 0 5152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_135
timestamp 1688980957
transform 1 0 13524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_175
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_276
timestamp 1688980957
transform 1 0 26496 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_319
timestamp 1688980957
transform 1 0 30452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_343
timestamp 1688980957
transform 1 0 32660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_406
timestamp 1688980957
transform 1 0 38456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_16
timestamp 1688980957
transform 1 0 2576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_20
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_72
timestamp 1688980957
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_96
timestamp 1688980957
transform 1 0 9936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_124
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_136
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_156
timestamp 1688980957
transform 1 0 15456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_304
timestamp 1688980957
transform 1 0 29072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_379
timestamp 1688980957
transform 1 0 35972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_405
timestamp 1688980957
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_13
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_89
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_138
timestamp 1688980957
transform 1 0 13800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_150
timestamp 1688980957
transform 1 0 14904 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_290
timestamp 1688980957
transform 1 0 27784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_345
timestamp 1688980957
transform 1 0 32844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_388
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_20
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_24
timestamp 1688980957
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_32
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_92
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_21
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_32
timestamp 1688980957
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_40 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_46
timestamp 1688980957
transform 1 0 5336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_60
timestamp 1688980957
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_71
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_185
timestamp 1688980957
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_198
timestamp 1688980957
transform 1 0 19320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_228
timestamp 1688980957
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_257
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_306
timestamp 1688980957
transform 1 0 29256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_375
timestamp 1688980957
transform 1 0 35604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_45
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_51
timestamp 1688980957
transform 1 0 5796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_55
timestamp 1688980957
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_74
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_111
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_127
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_131
timestamp 1688980957
transform 1 0 13156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_168
timestamp 1688980957
transform 1 0 16560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_193
timestamp 1688980957
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_203
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_256
timestamp 1688980957
transform 1 0 24656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_270
timestamp 1688980957
transform 1 0 25944 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_318
timestamp 1688980957
transform 1 0 30360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_38
timestamp 1688980957
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_74
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_78
timestamp 1688980957
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_82
timestamp 1688980957
transform 1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_86
timestamp 1688980957
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_91
timestamp 1688980957
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_96
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_100
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_139
timestamp 1688980957
transform 1 0 13892 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_143
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_146
timestamp 1688980957
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_150
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_159
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_188
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_192
timestamp 1688980957
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_204
timestamp 1688980957
transform 1 0 19872 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_209
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_229
timestamp 1688980957
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_238
timestamp 1688980957
transform 1 0 23000 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_252
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_259
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 1688980957
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_294
timestamp 1688980957
transform 1 0 28152 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_301
timestamp 1688980957
transform 1 0 28796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_308
timestamp 1688980957
transform 1 0 29440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_345
timestamp 1688980957
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_406
timestamp 1688980957
transform 1 0 38456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_11
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_32
timestamp 1688980957
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_36
timestamp 1688980957
transform 1 0 4416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_55
timestamp 1688980957
transform 1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_63
timestamp 1688980957
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 1688980957
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_108
timestamp 1688980957
transform 1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_136
timestamp 1688980957
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_149
timestamp 1688980957
transform 1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_159
timestamp 1688980957
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_164
timestamp 1688980957
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_213
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_217
timestamp 1688980957
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_257
timestamp 1688980957
transform 1 0 24748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_261
timestamp 1688980957
transform 1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_291
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_295
timestamp 1688980957
transform 1 0 28244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_299
timestamp 1688980957
transform 1 0 28612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_303
timestamp 1688980957
transform 1 0 28980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_313
timestamp 1688980957
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_330
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_360
timestamp 1688980957
transform 1 0 34224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_405
timestamp 1688980957
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_65
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_91
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_95
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_99
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_107
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_156
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_165
timestamp 1688980957
transform 1 0 16284 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_202
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_214
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1688980957
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_290
timestamp 1688980957
transform 1 0 27784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_298
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_302
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_306
timestamp 1688980957
transform 1 0 29256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_310
timestamp 1688980957
transform 1 0 29624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_314
timestamp 1688980957
transform 1 0 29992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_333
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_345
timestamp 1688980957
transform 1 0 32844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_353
timestamp 1688980957
transform 1 0 33580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_406
timestamp 1688980957
transform 1 0 38456 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 1688980957
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_59
timestamp 1688980957
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_151
timestamp 1688980957
transform 1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_257
timestamp 1688980957
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_304
timestamp 1688980957
transform 1 0 29072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_350
timestamp 1688980957
transform 1 0 33304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_354
timestamp 1688980957
transform 1 0 33672 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_406
timestamp 1688980957
transform 1 0 38456 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_147
timestamp 1688980957
transform 1 0 14628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_151
timestamp 1688980957
transform 1 0 14996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_173
timestamp 1688980957
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_198
timestamp 1688980957
transform 1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_254
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_306
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_333
timestamp 1688980957
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_355
timestamp 1688980957
transform 1 0 33764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_378
timestamp 1688980957
transform 1 0 35880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_396
timestamp 1688980957
transform 1 0 37536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_400
timestamp 1688980957
transform 1 0 37904 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_40
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_102
timestamp 1688980957
transform 1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_110
timestamp 1688980957
transform 1 0 11224 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 1688980957
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_191
timestamp 1688980957
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_257
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_292
timestamp 1688980957
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_296
timestamp 1688980957
transform 1 0 28336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_300
timestamp 1688980957
transform 1 0 28704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_304
timestamp 1688980957
transform 1 0 29072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_359
timestamp 1688980957
transform 1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_369
timestamp 1688980957
transform 1 0 35052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_396
timestamp 1688980957
transform 1 0 37536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_406
timestamp 1688980957
transform 1 0 38456 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_119
timestamp 1688980957
transform 1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_123
timestamp 1688980957
transform 1 0 12420 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_140
timestamp 1688980957
transform 1 0 13984 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_152
timestamp 1688980957
transform 1 0 15088 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_164
timestamp 1688980957
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_196
timestamp 1688980957
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_248
timestamp 1688980957
transform 1 0 23920 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_285
timestamp 1688980957
transform 1 0 27324 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_301
timestamp 1688980957
transform 1 0 28796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_333
timestamp 1688980957
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_347
timestamp 1688980957
transform 1 0 33028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_351
timestamp 1688980957
transform 1 0 33396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_390
timestamp 1688980957
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_401
timestamp 1688980957
transform 1 0 37996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_24
timestamp 1688980957
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_33
timestamp 1688980957
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_49
timestamp 1688980957
transform 1 0 5612 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_61
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_67
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_70
timestamp 1688980957
transform 1 0 7544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_117
timestamp 1688980957
transform 1 0 11868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_120
timestamp 1688980957
transform 1 0 12144 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_152
timestamp 1688980957
transform 1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_156
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_162
timestamp 1688980957
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_185
timestamp 1688980957
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1688980957
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_237
timestamp 1688980957
transform 1 0 22908 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_240
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_279
timestamp 1688980957
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_291
timestamp 1688980957
transform 1 0 27876 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_295
timestamp 1688980957
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_315
timestamp 1688980957
transform 1 0 30084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_319
timestamp 1688980957
transform 1 0 30452 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_324
timestamp 1688980957
transform 1 0 30912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_329
timestamp 1688980957
transform 1 0 31372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_337
timestamp 1688980957
transform 1 0 32108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_341
timestamp 1688980957
transform 1 0 32476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_349
timestamp 1688980957
transform 1 0 33212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_353
timestamp 1688980957
transform 1 0 33580 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_356
timestamp 1688980957
transform 1 0 33856 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_360
timestamp 1688980957
transform 1 0 34224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_381
timestamp 1688980957
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_406
timestamp 1688980957
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_68
timestamp 1688980957
transform 1 0 7360 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_89
timestamp 1688980957
transform 1 0 9292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1688980957
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_197
timestamp 1688980957
transform 1 0 19228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_209
timestamp 1688980957
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1688980957
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_238
timestamp 1688980957
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_253
timestamp 1688980957
transform 1 0 24380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_257
timestamp 1688980957
transform 1 0 24748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_269
timestamp 1688980957
transform 1 0 25852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_307
timestamp 1688980957
transform 1 0 29348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_315
timestamp 1688980957
transform 1 0 30084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_354
timestamp 1688980957
transform 1 0 33672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_385
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_389
timestamp 1688980957
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_405
timestamp 1688980957
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_57
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_101
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_158
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_191
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_201
timestamp 1688980957
transform 1 0 19596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_213
timestamp 1688980957
transform 1 0 20700 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_242
timestamp 1688980957
transform 1 0 23368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_269
timestamp 1688980957
transform 1 0 25852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_302
timestamp 1688980957
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_306
timestamp 1688980957
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_355
timestamp 1688980957
transform 1 0 33764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_404
timestamp 1688980957
transform 1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_12
timestamp 1688980957
transform 1 0 2208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_50
timestamp 1688980957
transform 1 0 5704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_107
timestamp 1688980957
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_208
timestamp 1688980957
transform 1 0 20240 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_214
timestamp 1688980957
transform 1 0 20792 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_311
timestamp 1688980957
transform 1 0 29716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_353
timestamp 1688980957
transform 1 0 33580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_372
timestamp 1688980957
transform 1 0 35328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_390
timestamp 1688980957
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_402
timestamp 1688980957
transform 1 0 38088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_406
timestamp 1688980957
transform 1 0 38456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 1688980957
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_36
timestamp 1688980957
transform 1 0 4416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_48
timestamp 1688980957
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_111
timestamp 1688980957
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_120
timestamp 1688980957
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_135
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_248
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_271
timestamp 1688980957
transform 1 0 26036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_317
timestamp 1688980957
transform 1 0 30268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_360
timestamp 1688980957
transform 1 0 34224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_386
timestamp 1688980957
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_390
timestamp 1688980957
transform 1 0 36984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_393
timestamp 1688980957
transform 1 0 37260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_398
timestamp 1688980957
transform 1 0 37720 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_34
timestamp 1688980957
transform 1 0 4232 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_46
timestamp 1688980957
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_102
timestamp 1688980957
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_117
timestamp 1688980957
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_145
timestamp 1688980957
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_157
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_183
timestamp 1688980957
transform 1 0 17940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_187
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_195
timestamp 1688980957
transform 1 0 19044 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_207
timestamp 1688980957
transform 1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_269
timestamp 1688980957
transform 1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_306
timestamp 1688980957
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_310
timestamp 1688980957
transform 1 0 29624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_330
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_354
timestamp 1688980957
transform 1 0 33672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_362
timestamp 1688980957
transform 1 0 34408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_389
timestamp 1688980957
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_401
timestamp 1688980957
transform 1 0 37996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_19
timestamp 1688980957
transform 1 0 2852 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_73
timestamp 1688980957
transform 1 0 7820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_101
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_134
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_157
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_191
timestamp 1688980957
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 1688980957
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_269
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_273
timestamp 1688980957
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_279
timestamp 1688980957
transform 1 0 26772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_283
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_287
timestamp 1688980957
transform 1 0 27508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_295
timestamp 1688980957
transform 1 0 28244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_299
timestamp 1688980957
transform 1 0 28612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_317
timestamp 1688980957
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_336
timestamp 1688980957
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_340
timestamp 1688980957
transform 1 0 32384 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_343
timestamp 1688980957
transform 1 0 32660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_355
timestamp 1688980957
transform 1 0 33764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_360
timestamp 1688980957
transform 1 0 34224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_404
timestamp 1688980957
transform 1 0 38272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_11
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_14
timestamp 1688980957
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_25
timestamp 1688980957
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_41
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_49
timestamp 1688980957
transform 1 0 5612 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_61
timestamp 1688980957
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_65
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_87
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_91
timestamp 1688980957
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_134
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_144
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_152
timestamp 1688980957
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_201
timestamp 1688980957
transform 1 0 19596 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_221
timestamp 1688980957
transform 1 0 21436 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_257
timestamp 1688980957
transform 1 0 24748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_267
timestamp 1688980957
transform 1 0 25668 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_297
timestamp 1688980957
transform 1 0 28428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_319
timestamp 1688980957
transform 1 0 30452 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_328
timestamp 1688980957
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_341
timestamp 1688980957
transform 1 0 32476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_402
timestamp 1688980957
transform 1 0 38088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_406
timestamp 1688980957
transform 1 0 38456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_54
timestamp 1688980957
transform 1 0 6072 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_71
timestamp 1688980957
transform 1 0 7636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_75
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_89
timestamp 1688980957
transform 1 0 9292 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_154
timestamp 1688980957
transform 1 0 15272 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_214
timestamp 1688980957
transform 1 0 20792 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_226
timestamp 1688980957
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_246
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_261
timestamp 1688980957
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_271
timestamp 1688980957
transform 1 0 26036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_275
timestamp 1688980957
transform 1 0 26404 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_361
timestamp 1688980957
transform 1 0 34316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_400
timestamp 1688980957
transform 1 0 37904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_404
timestamp 1688980957
transform 1 0 38272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_46
timestamp 1688980957
transform 1 0 5336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_94
timestamp 1688980957
transform 1 0 9752 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_108
timestamp 1688980957
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_138
timestamp 1688980957
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_142
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_146
timestamp 1688980957
transform 1 0 14536 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_156
timestamp 1688980957
transform 1 0 15456 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_275
timestamp 1688980957
transform 1 0 26404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_310
timestamp 1688980957
transform 1 0 29624 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_359
timestamp 1688980957
transform 1 0 34132 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_379
timestamp 1688980957
transform 1 0 35972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_383
timestamp 1688980957
transform 1 0 36340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_401
timestamp 1688980957
transform 1 0 37996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_79
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_99
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_107
timestamp 1688980957
transform 1 0 10948 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_203
timestamp 1688980957
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_212
timestamp 1688980957
transform 1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_220
timestamp 1688980957
transform 1 0 21344 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_248
timestamp 1688980957
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_270
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_303
timestamp 1688980957
transform 1 0 28980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_349
timestamp 1688980957
transform 1 0 33212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_353
timestamp 1688980957
transform 1 0 33580 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_373
timestamp 1688980957
transform 1 0 35420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_381
timestamp 1688980957
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_386
timestamp 1688980957
transform 1 0 36616 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_406
timestamp 1688980957
transform 1 0 38456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_29
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_42
timestamp 1688980957
transform 1 0 4968 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_91
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_99
timestamp 1688980957
transform 1 0 10212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_123
timestamp 1688980957
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_135
timestamp 1688980957
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_147
timestamp 1688980957
transform 1 0 14628 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_155
timestamp 1688980957
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_186
timestamp 1688980957
transform 1 0 18216 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_190
timestamp 1688980957
transform 1 0 18584 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_202
timestamp 1688980957
transform 1 0 19688 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_214
timestamp 1688980957
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1688980957
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_258
timestamp 1688980957
transform 1 0 24840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_297
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_370
timestamp 1688980957
transform 1 0 35144 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_388
timestamp 1688980957
transform 1 0 36800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_402
timestamp 1688980957
transform 1 0 38088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_406
timestamp 1688980957
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_38
timestamp 1688980957
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 1688980957
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1688980957
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_257
timestamp 1688980957
transform 1 0 24748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_264
timestamp 1688980957
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_268
timestamp 1688980957
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 1688980957
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_317
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_343
timestamp 1688980957
transform 1 0 32660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_347
timestamp 1688980957
transform 1 0 33028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_381
timestamp 1688980957
transform 1 0 36156 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_34
timestamp 1688980957
transform 1 0 4232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_43
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_61
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_79
timestamp 1688980957
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_83
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_92
timestamp 1688980957
transform 1 0 9568 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_142
timestamp 1688980957
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_198
timestamp 1688980957
transform 1 0 19320 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_210
timestamp 1688980957
transform 1 0 20424 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_214
timestamp 1688980957
transform 1 0 20792 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_253
timestamp 1688980957
transform 1 0 24380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_265
timestamp 1688980957
transform 1 0 25484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_276
timestamp 1688980957
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_297
timestamp 1688980957
transform 1 0 28428 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_303
timestamp 1688980957
transform 1 0 28980 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_308
timestamp 1688980957
transform 1 0 29440 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_316
timestamp 1688980957
transform 1 0 30176 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_319
timestamp 1688980957
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_331
timestamp 1688980957
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_343
timestamp 1688980957
transform 1 0 32660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_346
timestamp 1688980957
transform 1 0 32936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_366
timestamp 1688980957
transform 1 0 34776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_390
timestamp 1688980957
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_402
timestamp 1688980957
transform 1 0 38088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_406
timestamp 1688980957
transform 1 0 38456 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_37
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_45
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_57
timestamp 1688980957
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_74
timestamp 1688980957
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_82
timestamp 1688980957
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1688980957
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_149
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_186
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_190
timestamp 1688980957
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_239
timestamp 1688980957
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_257
timestamp 1688980957
transform 1 0 24748 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_261
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_273
timestamp 1688980957
transform 1 0 26220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_282
timestamp 1688980957
transform 1 0 27048 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_286
timestamp 1688980957
transform 1 0 27416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_290
timestamp 1688980957
transform 1 0 27784 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_294
timestamp 1688980957
transform 1 0 28152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_306
timestamp 1688980957
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_313
timestamp 1688980957
transform 1 0 29900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_325
timestamp 1688980957
transform 1 0 31004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_337
timestamp 1688980957
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_349
timestamp 1688980957
transform 1 0 33212 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_352
timestamp 1688980957
transform 1 0 33488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_391
timestamp 1688980957
transform 1 0 37076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_402
timestamp 1688980957
transform 1 0 38088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_406
timestamp 1688980957
transform 1 0 38456 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_11
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_46
timestamp 1688980957
transform 1 0 5336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_97
timestamp 1688980957
transform 1 0 10028 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_100
timestamp 1688980957
transform 1 0 10304 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_138
timestamp 1688980957
transform 1 0 13800 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_150
timestamp 1688980957
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_173
timestamp 1688980957
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_183
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_207
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_253
timestamp 1688980957
transform 1 0 24380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_257
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_265
timestamp 1688980957
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_277
timestamp 1688980957
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_298
timestamp 1688980957
transform 1 0 28520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_319
timestamp 1688980957
transform 1 0 30452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_323
timestamp 1688980957
transform 1 0 30820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_368
timestamp 1688980957
transform 1 0 34960 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_389
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_402
timestamp 1688980957
transform 1 0 38088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_406
timestamp 1688980957
transform 1 0 38456 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_80
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_105
timestamp 1688980957
transform 1 0 10764 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_114
timestamp 1688980957
transform 1 0 11592 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1688980957
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_175
timestamp 1688980957
transform 1 0 17204 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_184
timestamp 1688980957
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_242
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_246
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1688980957
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_259
timestamp 1688980957
transform 1 0 24932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_302
timestamp 1688980957
transform 1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_327
timestamp 1688980957
transform 1 0 31188 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_331
timestamp 1688980957
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_369
timestamp 1688980957
transform 1 0 35052 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_7
timestamp 1688980957
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_45
timestamp 1688980957
transform 1 0 5244 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_61
timestamp 1688980957
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_101
timestamp 1688980957
transform 1 0 10396 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_109
timestamp 1688980957
transform 1 0 11132 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_130
timestamp 1688980957
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_139
timestamp 1688980957
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_192
timestamp 1688980957
transform 1 0 18768 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_204
timestamp 1688980957
transform 1 0 19872 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_212
timestamp 1688980957
transform 1 0 20608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_257
timestamp 1688980957
transform 1 0 24748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_276
timestamp 1688980957
transform 1 0 26496 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_302
timestamp 1688980957
transform 1 0 28888 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_345
timestamp 1688980957
transform 1 0 32844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_385
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_389
timestamp 1688980957
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_401
timestamp 1688980957
transform 1 0 37996 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_11
timestamp 1688980957
transform 1 0 2116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_79
timestamp 1688980957
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_135
timestamp 1688980957
transform 1 0 13524 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_149
timestamp 1688980957
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_157
timestamp 1688980957
transform 1 0 15548 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_191
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_205
timestamp 1688980957
transform 1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_290
timestamp 1688980957
transform 1 0 27784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_354
timestamp 1688980957
transform 1 0 33672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_397
timestamp 1688980957
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_11
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_43
timestamp 1688980957
transform 1 0 5060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_49
timestamp 1688980957
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_88
timestamp 1688980957
transform 1 0 9200 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_147
timestamp 1688980957
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_151
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_204
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_216
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_250
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_260
timestamp 1688980957
transform 1 0 25024 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_289
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_351
timestamp 1688980957
transform 1 0 33396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_357
timestamp 1688980957
transform 1 0 33948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_366
timestamp 1688980957
transform 1 0 34776 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_370
timestamp 1688980957
transform 1 0 35144 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_374
timestamp 1688980957
transform 1 0 35512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_386
timestamp 1688980957
transform 1 0 36616 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_405
timestamp 1688980957
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_23
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_75
timestamp 1688980957
transform 1 0 8004 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_79
timestamp 1688980957
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_105
timestamp 1688980957
transform 1 0 10764 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_149
timestamp 1688980957
transform 1 0 14812 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_206
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_269
timestamp 1688980957
transform 1 0 25852 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_275
timestamp 1688980957
transform 1 0 26404 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_292
timestamp 1688980957
transform 1 0 27968 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_304
timestamp 1688980957
transform 1 0 29072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_314
timestamp 1688980957
transform 1 0 29992 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_331
timestamp 1688980957
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_343
timestamp 1688980957
transform 1 0 32660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_360
timestamp 1688980957
transform 1 0 34224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_385
timestamp 1688980957
transform 1 0 36524 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_393
timestamp 1688980957
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_397
timestamp 1688980957
transform 1 0 37628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_405
timestamp 1688980957
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_19
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_49
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_75
timestamp 1688980957
transform 1 0 8004 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_87
timestamp 1688980957
transform 1 0 9108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_95
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_136
timestamp 1688980957
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_140
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_152
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_179
timestamp 1688980957
transform 1 0 17572 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_198
timestamp 1688980957
transform 1 0 19320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_202
timestamp 1688980957
transform 1 0 19688 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_248
timestamp 1688980957
transform 1 0 23920 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_252
timestamp 1688980957
transform 1 0 24288 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_256
timestamp 1688980957
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_268
timestamp 1688980957
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_334
timestamp 1688980957
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_341
timestamp 1688980957
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_390
timestamp 1688980957
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_402
timestamp 1688980957
transform 1 0 38088 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_406
timestamp 1688980957
transform 1 0 38456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_11
timestamp 1688980957
transform 1 0 2116 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_45
timestamp 1688980957
transform 1 0 5244 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_50
timestamp 1688980957
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_54
timestamp 1688980957
transform 1 0 6072 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_66
timestamp 1688980957
transform 1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_105
timestamp 1688980957
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_188
timestamp 1688980957
transform 1 0 18400 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_192
timestamp 1688980957
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 1688980957
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_248
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_261
timestamp 1688980957
transform 1 0 25116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_269
timestamp 1688980957
transform 1 0 25852 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_279
timestamp 1688980957
transform 1 0 26772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_291
timestamp 1688980957
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_295
timestamp 1688980957
transform 1 0 28244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_298
timestamp 1688980957
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_361
timestamp 1688980957
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1688980957
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_92
timestamp 1688980957
transform 1 0 9568 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_96
timestamp 1688980957
transform 1 0 9936 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_138
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_142
timestamp 1688980957
transform 1 0 14168 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_154
timestamp 1688980957
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_250
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_254
timestamp 1688980957
transform 1 0 24472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_287
timestamp 1688980957
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_315
timestamp 1688980957
transform 1 0 30084 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_319
timestamp 1688980957
transform 1 0 30452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_331
timestamp 1688980957
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_371
timestamp 1688980957
transform 1 0 35236 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_381
timestamp 1688980957
transform 1 0 36156 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_402
timestamp 1688980957
transform 1 0 38088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_406
timestamp 1688980957
transform 1 0 38456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_11
timestamp 1688980957
transform 1 0 2116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_94
timestamp 1688980957
transform 1 0 9752 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_98
timestamp 1688980957
transform 1 0 10120 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_102
timestamp 1688980957
transform 1 0 10488 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_149
timestamp 1688980957
transform 1 0 14812 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_155
timestamp 1688980957
transform 1 0 15364 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_178
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_201
timestamp 1688980957
transform 1 0 19596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_240
timestamp 1688980957
transform 1 0 23184 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_244
timestamp 1688980957
transform 1 0 23552 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_248
timestamp 1688980957
transform 1 0 23920 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_286
timestamp 1688980957
transform 1 0 27416 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_290
timestamp 1688980957
transform 1 0 27784 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_325
timestamp 1688980957
transform 1 0 31004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_337
timestamp 1688980957
transform 1 0 32108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_351
timestamp 1688980957
transform 1 0 33396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_361
timestamp 1688980957
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_374
timestamp 1688980957
transform 1 0 35512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_406
timestamp 1688980957
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_48
timestamp 1688980957
transform 1 0 5520 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_52
timestamp 1688980957
transform 1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_98
timestamp 1688980957
transform 1 0 10120 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_119
timestamp 1688980957
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_145
timestamp 1688980957
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_209
timestamp 1688980957
transform 1 0 20332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_229
timestamp 1688980957
transform 1 0 22172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_234
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_390
timestamp 1688980957
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_401
timestamp 1688980957
transform 1 0 37996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_405
timestamp 1688980957
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_37
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_45
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_80
timestamp 1688980957
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_94
timestamp 1688980957
transform 1 0 9752 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_106
timestamp 1688980957
transform 1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_149
timestamp 1688980957
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_155
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_192
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_249
timestamp 1688980957
transform 1 0 24012 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_286
timestamp 1688980957
transform 1 0 27416 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_290
timestamp 1688980957
transform 1 0 27784 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_342
timestamp 1688980957
transform 1 0 32568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_354
timestamp 1688980957
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_29
timestamp 1688980957
transform 1 0 3772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_38
timestamp 1688980957
transform 1 0 4600 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_42
timestamp 1688980957
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_54
timestamp 1688980957
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_63
timestamp 1688980957
transform 1 0 6900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_73
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_144
timestamp 1688980957
transform 1 0 14352 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_156
timestamp 1688980957
transform 1 0 15456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_185
timestamp 1688980957
transform 1 0 18124 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_195
timestamp 1688980957
transform 1 0 19044 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_207
timestamp 1688980957
transform 1 0 20148 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_219
timestamp 1688980957
transform 1 0 21252 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_245
timestamp 1688980957
transform 1 0 23644 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_289
timestamp 1688980957
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_292
timestamp 1688980957
transform 1 0 27968 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_330
timestamp 1688980957
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_371
timestamp 1688980957
transform 1 0 35236 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_380
timestamp 1688980957
transform 1 0 36064 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_401
timestamp 1688980957
transform 1 0 37996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_9
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_48
timestamp 1688980957
transform 1 0 5520 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_52
timestamp 1688980957
transform 1 0 5888 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_60
timestamp 1688980957
transform 1 0 6624 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_71
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 1688980957
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_93
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_105
timestamp 1688980957
transform 1 0 10764 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_125
timestamp 1688980957
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_134
timestamp 1688980957
transform 1 0 13432 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_146
timestamp 1688980957
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_158
timestamp 1688980957
transform 1 0 15640 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_174
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_182
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_191
timestamp 1688980957
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_205
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_217
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_229
timestamp 1688980957
transform 1 0 22172 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_249
timestamp 1688980957
transform 1 0 24012 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_257
timestamp 1688980957
transform 1 0 24748 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_276
timestamp 1688980957
transform 1 0 26496 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_288
timestamp 1688980957
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_300
timestamp 1688980957
transform 1 0 28704 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_304
timestamp 1688980957
transform 1 0 29072 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_317
timestamp 1688980957
transform 1 0 30268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_329
timestamp 1688980957
transform 1 0 31372 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_341
timestamp 1688980957
transform 1 0 32476 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_346
timestamp 1688980957
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_358
timestamp 1688980957
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_371
timestamp 1688980957
transform 1 0 35236 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_392
timestamp 1688980957
transform 1 0 37168 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_402
timestamp 1688980957
transform 1 0 38088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_406
timestamp 1688980957
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_49
timestamp 1688980957
transform 1 0 5612 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_53
timestamp 1688980957
transform 1 0 5980 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_66
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_70
timestamp 1688980957
transform 1 0 7544 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_82
timestamp 1688980957
transform 1 0 8648 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_108
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_121
timestamp 1688980957
transform 1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_129
timestamp 1688980957
transform 1 0 12972 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_155
timestamp 1688980957
transform 1 0 15364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_196
timestamp 1688980957
transform 1 0 19136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_215
timestamp 1688980957
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_265
timestamp 1688980957
transform 1 0 25484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_277
timestamp 1688980957
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_294
timestamp 1688980957
transform 1 0 28152 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_298
timestamp 1688980957
transform 1 0 28520 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_310
timestamp 1688980957
transform 1 0 29624 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_322
timestamp 1688980957
transform 1 0 30728 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_332
timestamp 1688980957
transform 1 0 31648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_355
timestamp 1688980957
transform 1 0 33764 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_365
timestamp 1688980957
transform 1 0 34684 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_369
timestamp 1688980957
transform 1 0 35052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_401
timestamp 1688980957
transform 1 0 37996 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_11
timestamp 1688980957
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_50
timestamp 1688980957
transform 1 0 5704 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_54
timestamp 1688980957
transform 1 0 6072 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_66
timestamp 1688980957
transform 1 0 7176 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_70
timestamp 1688980957
transform 1 0 7544 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_74
timestamp 1688980957
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_116
timestamp 1688980957
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_120
timestamp 1688980957
transform 1 0 12144 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_250
timestamp 1688980957
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_269
timestamp 1688980957
transform 1 0 25852 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_273
timestamp 1688980957
transform 1 0 26220 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_281
timestamp 1688980957
transform 1 0 26956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_306
timestamp 1688980957
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_317
timestamp 1688980957
transform 1 0 30268 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_323
timestamp 1688980957
transform 1 0 30820 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_358
timestamp 1688980957
transform 1 0 34040 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_362
timestamp 1688980957
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_9
timestamp 1688980957
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_35
timestamp 1688980957
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_73
timestamp 1688980957
transform 1 0 7820 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_122
timestamp 1688980957
transform 1 0 12328 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_264
timestamp 1688980957
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_268
timestamp 1688980957
transform 1 0 25760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_315
timestamp 1688980957
transform 1 0 30084 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_319
timestamp 1688980957
transform 1 0 30452 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_367
timestamp 1688980957
transform 1 0 34868 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_389
timestamp 1688980957
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_402
timestamp 1688980957
transform 1 0 38088 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_406
timestamp 1688980957
transform 1 0 38456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_7
timestamp 1688980957
transform 1 0 1748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_122
timestamp 1688980957
transform 1 0 12328 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_166
timestamp 1688980957
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_170
timestamp 1688980957
transform 1 0 16744 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_176
timestamp 1688980957
transform 1 0 17296 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_213
timestamp 1688980957
transform 1 0 20700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_217
timestamp 1688980957
transform 1 0 21068 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_262
timestamp 1688980957
transform 1 0 25208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_266
timestamp 1688980957
transform 1 0 25576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_304
timestamp 1688980957
transform 1 0 29072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_317
timestamp 1688980957
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_369
timestamp 1688980957
transform 1 0 35052 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_403
timestamp 1688980957
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_11
timestamp 1688980957
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_29
timestamp 1688980957
transform 1 0 3772 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_73
timestamp 1688980957
transform 1 0 7820 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_77
timestamp 1688980957
transform 1 0 8188 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_83
timestamp 1688980957
transform 1 0 8740 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_121
timestamp 1688980957
transform 1 0 12236 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_162
timestamp 1688980957
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_203
timestamp 1688980957
transform 1 0 19780 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_214
timestamp 1688980957
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_229
timestamp 1688980957
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_264
timestamp 1688980957
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_268
timestamp 1688980957
transform 1 0 25760 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_297
timestamp 1688980957
transform 1 0 28428 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_315
timestamp 1688980957
transform 1 0 30084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_323
timestamp 1688980957
transform 1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_378
timestamp 1688980957
transform 1 0 35880 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_388
timestamp 1688980957
transform 1 0 36800 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_401
timestamp 1688980957
transform 1 0 37996 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_37
timestamp 1688980957
transform 1 0 4508 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_74
timestamp 1688980957
transform 1 0 7912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_82
timestamp 1688980957
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_101
timestamp 1688980957
transform 1 0 10396 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_110
timestamp 1688980957
transform 1 0 11224 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_122
timestamp 1688980957
transform 1 0 12328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_134
timestamp 1688980957
transform 1 0 13432 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1688980957
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_191
timestamp 1688980957
transform 1 0 18676 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_206
timestamp 1688980957
transform 1 0 20056 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_218
timestamp 1688980957
transform 1 0 21160 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_230
timestamp 1688980957
transform 1 0 22264 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_244
timestamp 1688980957
transform 1 0 23552 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_248
timestamp 1688980957
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_261
timestamp 1688980957
transform 1 0 25116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_273
timestamp 1688980957
transform 1 0 26220 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_303
timestamp 1688980957
transform 1 0 28980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 1688980957
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_371
timestamp 1688980957
transform 1 0 35236 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_402
timestamp 1688980957
transform 1 0 38088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_406
timestamp 1688980957
transform 1 0 38456 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_35
timestamp 1688980957
transform 1 0 4324 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_65
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_107
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_139
timestamp 1688980957
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_151
timestamp 1688980957
transform 1 0 14996 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 1688980957
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_175
timestamp 1688980957
transform 1 0 17204 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_203
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_215
timestamp 1688980957
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_243
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_246
timestamp 1688980957
transform 1 0 23736 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_260
timestamp 1688980957
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_272
timestamp 1688980957
transform 1 0 26128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_285
timestamp 1688980957
transform 1 0 27324 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_297
timestamp 1688980957
transform 1 0 28428 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_309
timestamp 1688980957
transform 1 0 29532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_321
timestamp 1688980957
transform 1 0 30636 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_324
timestamp 1688980957
transform 1 0 30912 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_354
timestamp 1688980957
transform 1 0 33672 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_358
timestamp 1688980957
transform 1 0 34040 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_366
timestamp 1688980957
transform 1 0 34776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_369
timestamp 1688980957
transform 1 0 35052 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_373
timestamp 1688980957
transform 1 0 35420 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_377
timestamp 1688980957
transform 1 0 35788 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_389
timestamp 1688980957
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_401
timestamp 1688980957
transform 1 0 37996 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_45
timestamp 1688980957
transform 1 0 5244 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_54
timestamp 1688980957
transform 1 0 6072 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_63
timestamp 1688980957
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_75
timestamp 1688980957
transform 1 0 8004 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_81
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_89
timestamp 1688980957
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_125
timestamp 1688980957
transform 1 0 12604 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_129
timestamp 1688980957
transform 1 0 12972 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_136
timestamp 1688980957
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_206
timestamp 1688980957
transform 1 0 20056 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_210
timestamp 1688980957
transform 1 0 20424 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_222
timestamp 1688980957
transform 1 0 21528 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_234
timestamp 1688980957
transform 1 0 22632 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_267
timestamp 1688980957
transform 1 0 25668 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_271
timestamp 1688980957
transform 1 0 26036 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_281
timestamp 1688980957
transform 1 0 26956 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_299
timestamp 1688980957
transform 1 0 28612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_317
timestamp 1688980957
transform 1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_402
timestamp 1688980957
transform 1 0 38088 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_406
timestamp 1688980957
transform 1 0 38456 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_122
timestamp 1688980957
transform 1 0 12328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_162
timestamp 1688980957
transform 1 0 16008 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_166
timestamp 1688980957
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_219
timestamp 1688980957
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_258
timestamp 1688980957
transform 1 0 24840 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_358
timestamp 1688980957
transform 1 0 34040 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_402
timestamp 1688980957
transform 1 0 38088 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_406
timestamp 1688980957
transform 1 0 38456 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_122
timestamp 1688980957
transform 1 0 12328 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_174
timestamp 1688980957
transform 1 0 17112 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_269
timestamp 1688980957
transform 1 0 25852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_305
timestamp 1688980957
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_318
timestamp 1688980957
transform 1 0 30360 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_322
timestamp 1688980957
transform 1 0 30728 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_400
timestamp 1688980957
transform 1 0 37904 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_406
timestamp 1688980957
transform 1 0 38456 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_108
timestamp 1688980957
transform 1 0 11040 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_162
timestamp 1688980957
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_185
timestamp 1688980957
transform 1 0 18124 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_219
timestamp 1688980957
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_277
timestamp 1688980957
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_322
timestamp 1688980957
transform 1 0 30728 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_330
timestamp 1688980957
transform 1 0 31464 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_369
timestamp 1688980957
transform 1 0 35052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_386
timestamp 1688980957
transform 1 0 36616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_401
timestamp 1688980957
transform 1 0 37996 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_101
timestamp 1688980957
transform 1 0 10396 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_111
timestamp 1688980957
transform 1 0 11316 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_123
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_128
timestamp 1688980957
transform 1 0 12880 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_150
timestamp 1688980957
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_159
timestamp 1688980957
transform 1 0 15732 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_171
timestamp 1688980957
transform 1 0 16836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_183
timestamp 1688980957
transform 1 0 17940 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_187
timestamp 1688980957
transform 1 0 18308 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_210
timestamp 1688980957
transform 1 0 20424 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_222
timestamp 1688980957
transform 1 0 21528 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_234
timestamp 1688980957
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_249
timestamp 1688980957
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_269
timestamp 1688980957
transform 1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_306
timestamp 1688980957
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_313
timestamp 1688980957
transform 1 0 29900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_325
timestamp 1688980957
transform 1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_343
timestamp 1688980957
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_355
timestamp 1688980957
transform 1 0 33764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_403
timestamp 1688980957
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_99
timestamp 1688980957
transform 1 0 10212 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_102
timestamp 1688980957
transform 1 0 10488 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_110
timestamp 1688980957
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_133
timestamp 1688980957
transform 1 0 13340 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_142
timestamp 1688980957
transform 1 0 14168 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_151
timestamp 1688980957
transform 1 0 14996 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_163
timestamp 1688980957
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_265
timestamp 1688980957
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_277
timestamp 1688980957
transform 1 0 26588 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_303
timestamp 1688980957
transform 1 0 28980 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_315
timestamp 1688980957
transform 1 0 30084 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_327
timestamp 1688980957
transform 1 0 31188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_373
timestamp 1688980957
transform 1 0 35420 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_381
timestamp 1688980957
transform 1 0 36156 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1688980957
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_401
timestamp 1688980957
transform 1 0 37996 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1688980957
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1688980957
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_401
timestamp 1688980957
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_401
timestamp 1688980957
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_401
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1688980957
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1688980957
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1688980957
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1688980957
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1688980957
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1688980957
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1688980957
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 1688980957
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 1688980957
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1688980957
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_225
timestamp 1688980957
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_237
timestamp 1688980957
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_249
timestamp 1688980957
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 1688980957
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_293
timestamp 1688980957
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 1688980957
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 1688980957
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 1688980957
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 1688980957
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 1688980957
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_405
timestamp 1688980957
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 37996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 30360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold5
timestamp 1688980957
transform -1 0 28520 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 29348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 32108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 32844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 33304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 28520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 28520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 33396 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 31372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 31740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 33672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 32844 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 33396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold20
timestamp 1688980957
transform 1 0 33856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 33120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold23
timestamp 1688980957
transform -1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 27232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 26864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 24012 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 23828 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform -1 0 35420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 24472 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 23920 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 37996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 37076 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 37168 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 34868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 22264 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 24196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 38272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 27140 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 26220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 20148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 20700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 25116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 22816 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 27968 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 25116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 27600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 24748 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 32292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 34132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 31464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 29900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 29532 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold60
timestamp 1688980957
transform 1 0 37628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 36892 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 37996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 37536 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 34592 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 28520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 34500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 34500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 36432 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 37996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 38548 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 37996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 35972 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 37720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 33856 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 36800 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 35604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 34224 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold81
timestamp 1688980957
transform -1 0 33580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 34224 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 36984 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 36064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 28336 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold86
timestamp 1688980957
transform -1 0 28520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 26864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 28612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 30268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 33672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 15088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold93
timestamp 1688980957
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 19596 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 26588 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold96
timestamp 1688980957
transform -1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 27876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 26864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 29992 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold101 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 38088 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 10764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold104
timestamp 1688980957
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 29256 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 28520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 37996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 25116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 22540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 25116 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 28428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 30268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 8464 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 6624 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 35420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 34040 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 36156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 34592 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 29716 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 38456 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 37996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 32016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 30636 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 33948 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform -1 0 33212 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform -1 0 20792 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 33580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 32844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 29256 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 32016 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 30544 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 29624 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform -1 0 28428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform -1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 33672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold147
timestamp 1688980957
transform -1 0 37720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform -1 0 37996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform -1 0 10856 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 24748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform -1 0 24748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 8832 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 36064 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform -1 0 35236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 35328 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform -1 0 36800 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 38548 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform -1 0 37996 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 36984 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform -1 0 36248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 6624 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform 1 0 6532 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform -1 0 25116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 34868 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 36340 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 38548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform -1 0 38456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 34040 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 33396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 34316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold176
timestamp 1688980957
transform -1 0 30084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform -1 0 27692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform -1 0 32936 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 32200 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 20148 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 20148 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 28520 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 28888 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform -1 0 38456 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform -1 0 38548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform 1 0 8372 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform 1 0 6624 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform -1 0 35420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform -1 0 34592 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 31832 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 29440 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold195
timestamp 1688980957
transform -1 0 24104 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 23368 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold198
timestamp 1688980957
transform -1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform -1 0 21252 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 27232 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 24748 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 21620 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 24012 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 23368 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 36892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold209
timestamp 1688980957
transform 1 0 33764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 34316 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform -1 0 32660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 33672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform -1 0 34684 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 37076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform -1 0 34592 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 27692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform -1 0 25668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform -1 0 31740 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold222
timestamp 1688980957
transform -1 0 29440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 28244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 30728 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 29256 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform -1 0 34776 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform -1 0 30084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 30268 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 34592 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 34592 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 32016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform -1 0 27508 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 26772 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 17664 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold237
timestamp 1688980957
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 14444 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 32660 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform -1 0 31372 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 32016 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 29624 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform -1 0 33672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform -1 0 32016 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform -1 0 24104 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 15640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 15088 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform 1 0 28520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold250
timestamp 1688980957
transform -1 0 28244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 26496 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform -1 0 20056 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform 1 0 20056 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform -1 0 24748 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 24104 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform -1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 32016 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform -1 0 18952 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform -1 0 22632 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform -1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform -1 0 21436 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform -1 0 31832 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform -1 0 32568 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform 1 0 27600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold267
timestamp 1688980957
transform -1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform -1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform -1 0 25116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform -1 0 24288 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform -1 0 28980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform -1 0 28244 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform -1 0 29992 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform -1 0 26864 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform -1 0 32016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform -1 0 31096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform -1 0 35052 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform -1 0 34316 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform -1 0 33672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 31280 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform -1 0 31464 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform -1 0 30268 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform -1 0 30728 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform -1 0 28520 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 24748 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform 1 0 24748 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform 1 0 31648 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold288
timestamp 1688980957
transform -1 0 36616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform -1 0 35972 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform -1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold291
timestamp 1688980957
transform 1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform -1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform -1 0 24564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform 1 0 15640 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform 1 0 26036 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform -1 0 26772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform -1 0 18952 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform -1 0 18400 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform -1 0 13616 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform -1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform -1 0 37444 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 37996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 35144 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold308
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform -1 0 16560 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform -1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform -1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform -1 0 26588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform -1 0 25852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform 1 0 37444 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform 1 0 35052 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform -1 0 4232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform -1 0 3496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform 1 0 34408 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform -1 0 38088 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform -1 0 37996 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform -1 0 37996 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform 1 0 14352 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform -1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform -1 0 8648 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform -1 0 7636 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1688980957
transform -1 0 16468 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform -1 0 15088 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform -1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform 1 0 21252 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform 1 0 29808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform -1 0 29808 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform 1 0 35604 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform 1 0 37352 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform -1 0 25852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform -1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform 1 0 22908 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform -1 0 24656 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform -1 0 13616 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform -1 0 14168 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform -1 0 20240 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform -1 0 19228 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform -1 0 37076 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform -1 0 6256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform -1 0 3680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform 1 0 1472 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1688980957
transform -1 0 18676 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform -1 0 17112 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1688980957
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1688980957
transform -1 0 30268 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1688980957
transform 1 0 26680 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 1688980957
transform -1 0 27416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1688980957
transform 1 0 24656 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold359
timestamp 1688980957
transform -1 0 25116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1688980957
transform -1 0 14352 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold362
timestamp 1688980957
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1688980957
transform -1 0 9752 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1688980957
transform -1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold365
timestamp 1688980957
transform -1 0 12144 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1688980957
transform -1 0 17388 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1688980957
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1688980957
transform -1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 1688980957
transform -1 0 8372 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1688980957
transform -1 0 6440 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1688980957
transform 1 0 1564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1688980957
transform -1 0 13800 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 1688980957
transform -1 0 11592 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 1688980957
transform -1 0 4784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold375
timestamp 1688980957
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold376
timestamp 1688980957
transform -1 0 3128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold377
timestamp 1688980957
transform -1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 1688980957
transform 1 0 6440 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 1688980957
transform -1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 1688980957
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 1688980957
transform -1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold382
timestamp 1688980957
transform 1 0 1472 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold383
timestamp 1688980957
transform -1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 1688980957
transform -1 0 18860 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 1688980957
transform -1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 1688980957
transform 1 0 6532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 1688980957
transform -1 0 6072 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold388
timestamp 1688980957
transform -1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold389
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 1688980957
transform -1 0 13064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 1688980957
transform -1 0 19320 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold392
timestamp 1688980957
transform -1 0 17940 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold393
timestamp 1688980957
transform -1 0 15456 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold394
timestamp 1688980957
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold395
timestamp 1688980957
transform -1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 1688980957
transform -1 0 9936 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold397
timestamp 1688980957
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold399
timestamp 1688980957
transform -1 0 5336 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold400
timestamp 1688980957
transform -1 0 3680 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold401
timestamp 1688980957
transform -1 0 23184 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold402
timestamp 1688980957
transform -1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold403
timestamp 1688980957
transform 1 0 18768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold404
timestamp 1688980957
transform -1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 1688980957
transform -1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold406
timestamp 1688980957
transform -1 0 13616 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold407
timestamp 1688980957
transform -1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold408
timestamp 1688980957
transform -1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold409
timestamp 1688980957
transform -1 0 16008 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 1688980957
transform -1 0 14996 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold411
timestamp 1688980957
transform -1 0 13984 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold412
timestamp 1688980957
transform 1 0 12236 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold413
timestamp 1688980957
transform -1 0 17112 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold414
timestamp 1688980957
transform -1 0 15732 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold415
timestamp 1688980957
transform -1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold416
timestamp 1688980957
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold417
timestamp 1688980957
transform -1 0 14996 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 1688980957
transform -1 0 14168 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 1688980957
transform 1 0 17848 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 1688980957
transform -1 0 19320 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 1688980957
transform -1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 1688980957
transform -1 0 16284 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 1688980957
transform -1 0 12328 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 1688980957
transform -1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 1688980957
transform -1 0 20332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 1688980957
transform -1 0 18768 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 1688980957
transform -1 0 11316 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 1688980957
transform -1 0 3680 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold432
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 1688980957
transform -1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 1688980957
transform 1 0 17572 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 1688980957
transform 1 0 17940 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 1688980957
transform -1 0 6072 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold437
timestamp 1688980957
transform 1 0 7176 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 1688980957
transform -1 0 21252 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 1688980957
transform -1 0 18216 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 1688980957
transform -1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 1688980957
transform -1 0 11776 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 1688980957
transform -1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 1688980957
transform -1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 1688980957
transform -1 0 18308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 1688980957
transform -1 0 12328 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 1688980957
transform -1 0 11040 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 1688980957
transform -1 0 5520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 1688980957
transform -1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 1688980957
transform -1 0 11316 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 1688980957
transform -1 0 9752 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 1688980957
transform -1 0 19044 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 1688980957
transform -1 0 13432 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold456
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold457
timestamp 1688980957
transform -1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold458
timestamp 1688980957
transform -1 0 3220 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold459
timestamp 1688980957
transform -1 0 18032 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold460
timestamp 1688980957
transform -1 0 17204 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 1688980957
transform -1 0 12604 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 1688980957
transform -1 0 10948 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold464
timestamp 1688980957
transform -1 0 3772 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold465
timestamp 1688980957
transform -1 0 5612 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 1688980957
transform 1 0 3864 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 1688980957
transform -1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 1688980957
transform -1 0 11408 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 1688980957
transform 1 0 2024 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold470
timestamp 1688980957
transform 1 0 2300 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 1688980957
transform -1 0 13616 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold473
timestamp 1688980957
transform -1 0 13340 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 1688980957
transform -1 0 11408 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold475
timestamp 1688980957
transform -1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold476
timestamp 1688980957
transform -1 0 19136 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 1688980957
transform -1 0 9568 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 1688980957
transform 1 0 6164 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold481
timestamp 1688980957
transform -1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold482
timestamp 1688980957
transform -1 0 16560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold483
timestamp 1688980957
transform -1 0 6164 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 1688980957
transform -1 0 3588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 1688980957
transform -1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold486
timestamp 1688980957
transform -1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold487
timestamp 1688980957
transform -1 0 14444 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold488
timestamp 1688980957
transform 1 0 12420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 1688980957
transform -1 0 10396 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 1688980957
transform -1 0 9476 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold491
timestamp 1688980957
transform 1 0 9016 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold492
timestamp 1688980957
transform -1 0 8924 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold493
timestamp 1688980957
transform 1 0 4784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold494
timestamp 1688980957
transform -1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold495
timestamp 1688980957
transform -1 0 4784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold496
timestamp 1688980957
transform -1 0 6072 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold497
timestamp 1688980957
transform 1 0 6256 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold498
timestamp 1688980957
transform 1 0 6900 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold499
timestamp 1688980957
transform 1 0 6440 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold500
timestamp 1688980957
transform -1 0 8556 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold501
timestamp 1688980957
transform -1 0 16008 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold502
timestamp 1688980957
transform 1 0 14444 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold503
timestamp 1688980957
transform -1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold504
timestamp 1688980957
transform -1 0 10764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold505
timestamp 1688980957
transform -1 0 8464 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold506
timestamp 1688980957
transform 1 0 8924 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold507
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold508
timestamp 1688980957
transform -1 0 16836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold509
timestamp 1688980957
transform -1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold510
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold511
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold512
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold513
timestamp 1688980957
transform -1 0 12052 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold514
timestamp 1688980957
transform -1 0 11408 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold515
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold516
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold517
timestamp 1688980957
transform -1 0 10488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold518
timestamp 1688980957
transform -1 0 14628 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold519
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold520
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold521
timestamp 1688980957
transform -1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold522
timestamp 1688980957
transform -1 0 17296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold523
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold524
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold525
timestamp 1688980957
transform -1 0 16836 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold526
timestamp 1688980957
transform -1 0 16100 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold527
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold528
timestamp 1688980957
transform -1 0 13800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold529
timestamp 1688980957
transform -1 0 14352 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold530
timestamp 1688980957
transform -1 0 13616 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 1688980957
transform 1 0 14352 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 1688980957
transform -1 0 15732 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold533
timestamp 1688980957
transform -1 0 15456 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold534
timestamp 1688980957
transform -1 0 13892 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold535
timestamp 1688980957
transform -1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold536
timestamp 1688980957
transform -1 0 19688 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold537
timestamp 1688980957
transform -1 0 19320 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold538
timestamp 1688980957
transform -1 0 19136 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold539
timestamp 1688980957
transform -1 0 18400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold540
timestamp 1688980957
transform -1 0 18676 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold541
timestamp 1688980957
transform -1 0 18492 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold542
timestamp 1688980957
transform -1 0 17664 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold543
timestamp 1688980957
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold544
timestamp 1688980957
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold545
timestamp 1688980957
transform -1 0 3680 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold546
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold547
timestamp 1688980957
transform -1 0 3772 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold548 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold549
timestamp 1688980957
transform -1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold550 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3036 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold551
timestamp 1688980957
transform 1 0 4508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold552
timestamp 1688980957
transform -1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold553
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold554
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold555
timestamp 1688980957
transform 1 0 4232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold556
timestamp 1688980957
transform -1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold557
timestamp 1688980957
transform -1 0 3312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold558
timestamp 1688980957
transform -1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold559
timestamp 1688980957
transform -1 0 2208 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold560
timestamp 1688980957
transform 1 0 2668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold561
timestamp 1688980957
transform -1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold562
timestamp 1688980957
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold563
timestamp 1688980957
transform -1 0 8740 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold564
timestamp 1688980957
transform -1 0 24288 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold565
timestamp 1688980957
transform -1 0 36708 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold566
timestamp 1688980957
transform -1 0 29256 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold567
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold568
timestamp 1688980957
transform -1 0 32844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold569
timestamp 1688980957
transform -1 0 21160 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold570
timestamp 1688980957
transform -1 0 33672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold571
timestamp 1688980957
transform 1 0 32384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold572
timestamp 1688980957
transform 1 0 19688 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold573
timestamp 1688980957
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold574
timestamp 1688980957
transform -1 0 18860 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold575
timestamp 1688980957
transform 1 0 27232 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold576
timestamp 1688980957
transform -1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold577
timestamp 1688980957
transform -1 0 34408 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold578
timestamp 1688980957
transform -1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold579
timestamp 1688980957
transform -1 0 18860 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold580
timestamp 1688980957
transform -1 0 36616 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold581
timestamp 1688980957
transform -1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold582
timestamp 1688980957
transform -1 0 11224 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold583
timestamp 1688980957
transform -1 0 28980 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold584
timestamp 1688980957
transform -1 0 38548 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold585
timestamp 1688980957
transform -1 0 6900 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold586
timestamp 1688980957
transform -1 0 13708 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold587
timestamp 1688980957
transform -1 0 11408 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold588
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold589
timestamp 1688980957
transform 1 0 18124 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold590
timestamp 1688980957
transform -1 0 13616 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold591
timestamp 1688980957
transform -1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold592
timestamp 1688980957
transform -1 0 37076 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold593
timestamp 1688980957
transform 1 0 13616 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold594
timestamp 1688980957
transform -1 0 25852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold595
timestamp 1688980957
transform -1 0 29164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 24288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 29440 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 33580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 37536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform -1 0 32292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform -1 0 32016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform -1 0 11040 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform -1 0 14628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform -1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 19320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform -1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform -1 0 26864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 24472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform -1 0 30452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 29624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 28520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform -1 0 29440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform -1 0 33672 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 35880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 34132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform -1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform -1 0 38364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 38272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform -1 0 9016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform -1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 11040 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input68
timestamp 1688980957
transform 1 0 2944 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  max_cap118
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  max_cap119
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  output69 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1472 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform -1 0 5152 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform -1 0 18768 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform -1 0 19136 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform -1 0 23276 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform -1 0 24288 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform -1 0 25852 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform -1 0 26496 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform 1 0 27232 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform -1 0 30176 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform -1 0 32016 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform -1 0 33580 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform -1 0 34224 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1688980957
transform -1 0 36432 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1688980957
transform -1 0 37536 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1688980957
transform -1 0 38548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1688980957
transform -1 0 37168 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1688980957
transform -1 0 34592 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1688980957
transform 1 0 8096 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform 1 0 15088 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire120
timestamp 1688980957
transform -1 0 1932 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 1030 0 1086 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 5 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 6 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 7 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 8 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 9 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 10 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 11 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 12 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 13 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 14 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 15 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 16 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 17 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 18 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 19 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 20 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 21 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 22 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 23 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 24 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 25 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 26 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 27 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 28 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 29 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 30 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 31 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 32 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 33 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 34 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 35 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 36 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 37 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 38 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 40 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 41 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 42 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 43 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 44 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 45 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 46 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 47 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 48 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 49 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 50 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 51 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 52 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 53 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 54 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 55 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 56 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 57 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 58 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 59 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 60 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 61 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 62 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 63 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 64 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 65 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 66 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 67 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 68 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 69 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 70 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 71 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 72 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 73 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 74 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 75 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 76 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 77 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 78 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 79 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 80 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 81 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 82 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 83 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 84 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 85 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 86 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 87 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 88 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 89 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 90 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 91 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 92 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 93 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 94 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 95 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 96 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 97 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 98 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 99 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 100 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 101 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 102 nsew signal input
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 103 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 104 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 105 nsew signal input
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 106 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 wbs_we_i
port 107 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
