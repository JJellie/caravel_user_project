magic
tech sky130A
magscale 1 2
timestamp 1725975754
<< obsli1 >>
rect 1104 2159 58880 27761
<< obsm1 >>
rect 1104 1504 59142 27792
<< metal2 >>
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
<< obsm2 >>
rect 938 856 59136 27781
rect 1050 734 1434 856
rect 1602 734 1986 856
rect 2154 734 2538 856
rect 2706 734 3090 856
rect 3258 734 3642 856
rect 3810 734 4194 856
rect 4362 734 4746 856
rect 4914 734 5298 856
rect 5466 734 5850 856
rect 6018 734 6402 856
rect 6570 734 6954 856
rect 7122 734 7506 856
rect 7674 734 8058 856
rect 8226 734 8610 856
rect 8778 734 9162 856
rect 9330 734 9714 856
rect 9882 734 10266 856
rect 10434 734 10818 856
rect 10986 734 11370 856
rect 11538 734 11922 856
rect 12090 734 12474 856
rect 12642 734 13026 856
rect 13194 734 13578 856
rect 13746 734 14130 856
rect 14298 734 14682 856
rect 14850 734 15234 856
rect 15402 734 15786 856
rect 15954 734 16338 856
rect 16506 734 16890 856
rect 17058 734 17442 856
rect 17610 734 17994 856
rect 18162 734 18546 856
rect 18714 734 19098 856
rect 19266 734 19650 856
rect 19818 734 20202 856
rect 20370 734 20754 856
rect 20922 734 21306 856
rect 21474 734 21858 856
rect 22026 734 22410 856
rect 22578 734 22962 856
rect 23130 734 23514 856
rect 23682 734 24066 856
rect 24234 734 24618 856
rect 24786 734 25170 856
rect 25338 734 25722 856
rect 25890 734 26274 856
rect 26442 734 26826 856
rect 26994 734 27378 856
rect 27546 734 27930 856
rect 28098 734 28482 856
rect 28650 734 29034 856
rect 29202 734 29586 856
rect 29754 734 30138 856
rect 30306 734 30690 856
rect 30858 734 31242 856
rect 31410 734 31794 856
rect 31962 734 32346 856
rect 32514 734 32898 856
rect 33066 734 33450 856
rect 33618 734 34002 856
rect 34170 734 34554 856
rect 34722 734 35106 856
rect 35274 734 35658 856
rect 35826 734 36210 856
rect 36378 734 36762 856
rect 36930 734 37314 856
rect 37482 734 37866 856
rect 38034 734 38418 856
rect 38586 734 38970 856
rect 39138 734 39522 856
rect 39690 734 40074 856
rect 40242 734 40626 856
rect 40794 734 41178 856
rect 41346 734 41730 856
rect 41898 734 42282 856
rect 42450 734 42834 856
rect 43002 734 43386 856
rect 43554 734 43938 856
rect 44106 734 44490 856
rect 44658 734 45042 856
rect 45210 734 45594 856
rect 45762 734 46146 856
rect 46314 734 46698 856
rect 46866 734 47250 856
rect 47418 734 47802 856
rect 47970 734 48354 856
rect 48522 734 48906 856
rect 49074 734 49458 856
rect 49626 734 50010 856
rect 50178 734 50562 856
rect 50730 734 51114 856
rect 51282 734 51666 856
rect 51834 734 52218 856
rect 52386 734 52770 856
rect 52938 734 53322 856
rect 53490 734 53874 856
rect 54042 734 54426 856
rect 54594 734 54978 856
rect 55146 734 55530 856
rect 55698 734 56082 856
rect 56250 734 56634 856
rect 56802 734 57186 856
rect 57354 734 57738 856
rect 57906 734 58290 856
rect 58458 734 58842 856
rect 59010 734 59136 856
<< obsm3 >>
rect 933 2143 59038 27777
<< metal4 >>
rect 8166 2128 8486 27792
rect 15388 2128 15708 27792
rect 22610 2128 22930 27792
rect 29832 2128 30152 27792
rect 37054 2128 37374 27792
rect 44276 2128 44596 27792
rect 51498 2128 51818 27792
rect 58720 2128 59040 27792
<< obsm4 >>
rect 57099 3979 57165 11117
<< labels >>
rlabel metal4 s 8166 2128 8486 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 22610 2128 22930 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 37054 2128 37374 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 51498 2128 51818 27792 6 vccd1
port 1 nsew power bidirectional
rlabel metal4 s 15388 2128 15708 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal4 s 29832 2128 30152 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal4 s 44276 2128 44596 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal4 s 58720 2128 59040 27792 6 vssd1
port 2 nsew ground bidirectional
rlabel metal2 s 938 0 994 800 6 wb_clk_i
port 3 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 4 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_ack_o
port 5 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[0]
port 6 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[10]
port 7 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[11]
port 8 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[12]
port 9 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[13]
port 10 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[14]
port 11 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[15]
port 12 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[16]
port 13 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[17]
port 14 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[18]
port 15 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[19]
port 16 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[1]
port 17 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[20]
port 18 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_adr_i[21]
port 19 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[22]
port 20 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_adr_i[23]
port 21 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_adr_i[24]
port 22 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_adr_i[25]
port 23 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[26]
port 24 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[27]
port 25 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[28]
port 26 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_adr_i[29]
port 27 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[2]
port 28 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_adr_i[30]
port 29 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_adr_i[31]
port 30 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[3]
port 31 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[4]
port 32 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[5]
port 33 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[6]
port 34 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[7]
port 35 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[8]
port 36 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[9]
port 37 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_cyc_i
port 38 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_i[0]
port 39 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[10]
port 40 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[11]
port 41 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[12]
port 42 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[13]
port 43 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[14]
port 44 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[15]
port 45 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[16]
port 46 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[17]
port 47 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[18]
port 48 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[19]
port 49 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[1]
port 50 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[20]
port 51 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[21]
port 52 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[22]
port 53 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[23]
port 54 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_i[24]
port 55 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_i[25]
port 56 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[26]
port 57 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[27]
port 58 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_i[28]
port 59 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_i[29]
port 60 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_i[2]
port 61 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_i[30]
port 62 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_i[31]
port 63 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[3]
port 64 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[4]
port 65 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[5]
port 66 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[6]
port 67 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[7]
port 68 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[8]
port 69 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_i[9]
port 70 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_o[0]
port 71 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[10]
port 72 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[11]
port 73 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[12]
port 74 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[13]
port 75 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[14]
port 76 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[15]
port 77 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[16]
port 78 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[17]
port 79 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[18]
port 80 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[19]
port 81 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_o[1]
port 82 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[20]
port 83 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 wbs_dat_o[21]
port 84 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_o[22]
port 85 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_o[23]
port 86 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_o[24]
port 87 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 wbs_dat_o[25]
port 88 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_o[26]
port 89 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_o[27]
port 90 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[28]
port 91 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_o[29]
port 92 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[2]
port 93 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_o[30]
port 94 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[31]
port 95 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[3]
port 96 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[4]
port 97 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[5]
port 98 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[6]
port 99 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[7]
port 100 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[8]
port 101 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[9]
port 102 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_sel_i[0]
port 103 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_sel_i[1]
port 104 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_sel_i[2]
port 105 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_sel_i[3]
port 106 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_stb_i
port 107 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_we_i
port 108 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3823736
string GDS_FILE /home/jelmer/Documents/stage/efabless/caravel_user_project/openlane/wishbone_nn/runs/24_09_10_15_39/results/signoff/wishbone_nn.magic.gds
string GDS_START 392402
<< end >>

