magic
tech sky130A
magscale 1 2
timestamp 1725975750
<< viali >>
rect 38853 23069 38887 23103
rect 47869 23069 47903 23103
rect 39405 22933 39439 22967
rect 40049 22933 40083 22967
rect 48513 22933 48547 22967
rect 47860 22661 47894 22695
rect 38301 22593 38335 22627
rect 38568 22593 38602 22627
rect 49065 22593 49099 22627
rect 24777 22525 24811 22559
rect 39773 22525 39807 22559
rect 47593 22525 47627 22559
rect 50721 22525 50755 22559
rect 51365 22525 51399 22559
rect 52929 22525 52963 22559
rect 55045 22525 55079 22559
rect 55873 22525 55907 22559
rect 48973 22457 49007 22491
rect 24317 22389 24351 22423
rect 24685 22389 24719 22423
rect 25421 22389 25455 22423
rect 38209 22389 38243 22423
rect 39681 22389 39715 22423
rect 40417 22389 40451 22423
rect 47409 22389 47443 22423
rect 49709 22389 49743 22423
rect 51273 22389 51307 22423
rect 52009 22389 52043 22423
rect 52377 22389 52411 22423
rect 53573 22389 53607 22423
rect 55597 22389 55631 22423
rect 56425 22389 56459 22423
rect 56701 22389 56735 22423
rect 47777 22185 47811 22219
rect 55321 22185 55355 22219
rect 56517 22117 56551 22151
rect 24409 22049 24443 22083
rect 37473 22049 37507 22083
rect 39589 22049 39623 22083
rect 40509 22049 40543 22083
rect 47685 22049 47719 22083
rect 48329 22049 48363 22083
rect 55781 22049 55815 22083
rect 55965 22049 55999 22083
rect 56333 22049 56367 22083
rect 57069 22049 57103 22083
rect 57345 22049 57379 22083
rect 10517 21981 10551 22015
rect 23673 21981 23707 22015
rect 24676 21981 24710 22015
rect 25881 21981 25915 22015
rect 39865 21981 39899 22015
rect 48237 21981 48271 22015
rect 49985 21981 50019 22015
rect 50169 21981 50203 22015
rect 51641 21981 51675 22015
rect 53113 21981 53147 22015
rect 53849 21981 53883 22015
rect 14841 21913 14875 21947
rect 37740 21913 37774 21947
rect 50436 21913 50470 21947
rect 51908 21913 51942 21947
rect 53757 21913 53791 21947
rect 56977 21913 57011 21947
rect 6377 21845 6411 21879
rect 11069 21845 11103 21879
rect 11345 21845 11379 21879
rect 23029 21845 23063 21879
rect 24225 21845 24259 21879
rect 25789 21845 25823 21879
rect 26525 21845 26559 21879
rect 38853 21845 38887 21879
rect 38945 21845 38979 21879
rect 39313 21845 39347 21879
rect 39405 21845 39439 21879
rect 48145 21845 48179 21879
rect 51549 21845 51583 21879
rect 53021 21845 53055 21879
rect 54493 21845 54527 21879
rect 54769 21845 54803 21879
rect 55689 21845 55723 21879
rect 56885 21845 56919 21879
rect 57989 21845 58023 21879
rect 4445 21641 4479 21675
rect 10517 21641 10551 21675
rect 10977 21641 11011 21675
rect 12173 21641 12207 21675
rect 23581 21641 23615 21675
rect 24777 21641 24811 21675
rect 25237 21641 25271 21675
rect 38853 21641 38887 21675
rect 40325 21641 40359 21675
rect 50721 21641 50755 21675
rect 51181 21641 51215 21675
rect 52101 21641 52135 21675
rect 55689 21641 55723 21675
rect 58541 21641 58575 21675
rect 39313 21573 39347 21607
rect 56416 21573 56450 21607
rect 6469 21505 6503 21539
rect 9229 21505 9263 21539
rect 10885 21505 10919 21539
rect 23489 21505 23523 21539
rect 25145 21505 25179 21539
rect 39221 21505 39255 21539
rect 39681 21505 39715 21539
rect 51089 21505 51123 21539
rect 52009 21505 52043 21539
rect 52745 21505 52779 21539
rect 53012 21505 53046 21539
rect 54309 21505 54343 21539
rect 54576 21505 54610 21539
rect 56057 21505 56091 21539
rect 3157 21437 3191 21471
rect 4077 21437 4111 21471
rect 5641 21437 5675 21471
rect 7481 21437 7515 21471
rect 8401 21437 8435 21471
rect 11069 21437 11103 21471
rect 11529 21437 11563 21471
rect 13921 21437 13955 21471
rect 15209 21437 15243 21471
rect 18705 21437 18739 21471
rect 22477 21437 22511 21471
rect 23765 21437 23799 21471
rect 23949 21437 23983 21471
rect 25329 21437 25363 21471
rect 26065 21437 26099 21471
rect 30205 21437 30239 21471
rect 39405 21437 39439 21471
rect 42717 21437 42751 21471
rect 46673 21437 46707 21471
rect 50629 21437 50663 21471
rect 51365 21437 51399 21471
rect 52285 21437 52319 21471
rect 56149 21437 56183 21471
rect 57897 21437 57931 21471
rect 8217 21369 8251 21403
rect 13737 21369 13771 21403
rect 23121 21369 23155 21403
rect 38117 21369 38151 21403
rect 42257 21369 42291 21403
rect 51641 21369 51675 21403
rect 3709 21301 3743 21335
rect 6193 21301 6227 21335
rect 7113 21301 7147 21335
rect 8953 21301 8987 21335
rect 9781 21301 9815 21335
rect 10149 21301 10183 21335
rect 14473 21301 14507 21335
rect 15025 21301 15059 21335
rect 15853 21301 15887 21335
rect 19349 21301 19383 21335
rect 19625 21301 19659 21335
rect 23029 21301 23063 21335
rect 24593 21301 24627 21335
rect 25789 21301 25823 21335
rect 26617 21301 26651 21335
rect 30849 21301 30883 21335
rect 38393 21301 38427 21335
rect 41889 21301 41923 21335
rect 43269 21301 43303 21335
rect 43637 21301 43671 21335
rect 45937 21301 45971 21335
rect 46489 21301 46523 21335
rect 47225 21301 47259 21335
rect 47869 21301 47903 21335
rect 50169 21301 50203 21335
rect 54125 21301 54159 21335
rect 57529 21301 57563 21335
rect 6285 21097 6319 21131
rect 8769 21097 8803 21131
rect 15025 21097 15059 21131
rect 22385 21097 22419 21131
rect 26341 21097 26375 21131
rect 30021 21097 30055 21131
rect 30205 21097 30239 21131
rect 39589 21097 39623 21131
rect 41429 21097 41463 21131
rect 46765 21097 46799 21131
rect 53665 21097 53699 21131
rect 2881 21029 2915 21063
rect 14105 21029 14139 21063
rect 23857 21029 23891 21063
rect 43913 21029 43947 21063
rect 55137 21029 55171 21063
rect 2237 20961 2271 20995
rect 3525 20961 3559 20995
rect 6745 20961 6779 20995
rect 6929 20961 6963 20995
rect 7389 20961 7423 20995
rect 9413 20961 9447 20995
rect 9597 20961 9631 20995
rect 13185 20961 13219 20995
rect 14565 20961 14599 20995
rect 14749 20961 14783 20995
rect 15577 20961 15611 20995
rect 22477 20961 22511 20995
rect 24409 20961 24443 20995
rect 24593 20961 24627 20995
rect 25053 20961 25087 20995
rect 26801 20961 26835 20995
rect 26893 20961 26927 20995
rect 30757 20961 30791 20995
rect 45753 20961 45787 20995
rect 47409 20961 47443 20995
rect 51641 20961 51675 20995
rect 52101 20961 52135 20995
rect 52377 20961 52411 20995
rect 52653 20961 52687 20995
rect 55689 20961 55723 20995
rect 56333 20961 56367 20995
rect 56726 20961 56760 20995
rect 56885 20961 56919 20995
rect 58173 20961 58207 20995
rect 3985 20893 4019 20927
rect 4813 20893 4847 20927
rect 7656 20893 7690 20927
rect 10057 20893 10091 20927
rect 16037 20893 16071 20927
rect 16681 20893 16715 20927
rect 18245 20893 18279 20927
rect 19901 20893 19935 20927
rect 20637 20893 20671 20927
rect 22744 20893 22778 20927
rect 25329 20893 25363 20927
rect 25446 20893 25480 20927
rect 25605 20893 25639 20927
rect 27169 20893 27203 20927
rect 27997 20893 28031 20927
rect 28825 20893 28859 20927
rect 31033 20893 31067 20927
rect 32873 20893 32907 20927
rect 33701 20893 33735 20927
rect 34989 20893 35023 20927
rect 36093 20893 36127 20927
rect 37565 20893 37599 20927
rect 38301 20893 38335 20927
rect 41797 20893 41831 20927
rect 42441 20893 42475 20927
rect 45017 20893 45051 20927
rect 47685 20893 47719 20927
rect 49157 20893 49191 20927
rect 50813 20893 50847 20927
rect 51457 20893 51491 20927
rect 52494 20893 52528 20927
rect 53757 20893 53791 20927
rect 55873 20893 55907 20927
rect 56609 20893 56643 20927
rect 5080 20825 5114 20859
rect 10324 20825 10358 20859
rect 11805 20825 11839 20859
rect 13001 20825 13035 20859
rect 15485 20825 15519 20859
rect 17325 20825 17359 20859
rect 17969 20825 18003 20859
rect 24133 20825 24167 20859
rect 26709 20825 26743 20859
rect 27813 20825 27847 20859
rect 46397 20825 46431 20859
rect 47133 20825 47167 20859
rect 48973 20825 49007 20859
rect 54024 20825 54058 20859
rect 58081 20825 58115 20859
rect 2789 20757 2823 20791
rect 3249 20757 3283 20791
rect 3341 20757 3375 20791
rect 4537 20757 4571 20791
rect 6193 20757 6227 20791
rect 6653 20757 6687 20791
rect 8953 20757 8987 20791
rect 9321 20757 9355 20791
rect 11437 20757 11471 20791
rect 13737 20757 13771 20791
rect 14473 20757 14507 20791
rect 15393 20757 15427 20791
rect 16589 20757 16623 20791
rect 18797 20757 18831 20791
rect 19533 20757 19567 20791
rect 20545 20757 20579 20791
rect 21281 20757 21315 20791
rect 26249 20757 26283 20791
rect 28549 20757 28583 20791
rect 29377 20757 29411 20791
rect 30573 20757 30607 20791
rect 30665 20757 30699 20791
rect 31677 20757 31711 20791
rect 33425 20757 33459 20791
rect 34253 20757 34287 20791
rect 35357 20757 35391 20791
rect 36737 20757 36771 20791
rect 37381 20757 37415 20791
rect 38117 20757 38151 20791
rect 38853 20757 38887 20791
rect 39221 20757 39255 20791
rect 42349 20757 42383 20791
rect 44649 20757 44683 20791
rect 45661 20757 45695 20791
rect 47225 20757 47259 20791
rect 48237 20757 48271 20791
rect 48605 20757 48639 20791
rect 49709 20757 49743 20791
rect 51089 20757 51123 20791
rect 53297 20757 53331 20791
rect 55505 20757 55539 20791
rect 57529 20757 57563 20791
rect 57621 20757 57655 20791
rect 57989 20757 58023 20791
rect 3801 20553 3835 20587
rect 6837 20553 6871 20587
rect 7573 20553 7607 20587
rect 13093 20553 13127 20587
rect 18521 20553 18555 20587
rect 22201 20553 22235 20587
rect 23673 20553 23707 20587
rect 24133 20553 24167 20587
rect 26709 20553 26743 20587
rect 27905 20553 27939 20587
rect 28089 20553 28123 20587
rect 28549 20553 28583 20587
rect 31585 20553 31619 20587
rect 32965 20553 32999 20587
rect 33425 20553 33459 20587
rect 37565 20553 37599 20587
rect 37933 20553 37967 20587
rect 40785 20553 40819 20587
rect 42441 20553 42475 20587
rect 42901 20553 42935 20587
rect 49525 20553 49559 20587
rect 52745 20553 52779 20587
rect 57713 20553 57747 20587
rect 11980 20485 12014 20519
rect 15292 20485 15326 20519
rect 28457 20485 28491 20519
rect 30104 20485 30138 20519
rect 42809 20485 42843 20519
rect 46296 20485 46330 20519
rect 49893 20485 49927 20519
rect 50997 20485 51031 20519
rect 56885 20485 56919 20519
rect 2053 20417 2087 20451
rect 2320 20417 2354 20451
rect 4997 20417 5031 20451
rect 6745 20417 6779 20451
rect 7665 20417 7699 20451
rect 7932 20417 7966 20451
rect 9505 20417 9539 20451
rect 10425 20417 10459 20451
rect 13185 20417 13219 20451
rect 18429 20417 18463 20451
rect 19533 20417 19567 20451
rect 19800 20417 19834 20451
rect 22293 20417 22327 20451
rect 22560 20417 22594 20451
rect 25596 20417 25630 20451
rect 33333 20417 33367 20451
rect 34796 20417 34830 20451
rect 36645 20417 36679 20451
rect 38393 20417 38427 20451
rect 39313 20417 39347 20451
rect 39589 20417 39623 20451
rect 41144 20417 41178 20451
rect 43361 20417 43395 20451
rect 43628 20417 43662 20451
rect 46029 20417 46063 20451
rect 47593 20417 47627 20451
rect 53113 20417 53147 20451
rect 54309 20417 54343 20451
rect 55045 20417 55079 20451
rect 56149 20417 56183 20451
rect 57069 20417 57103 20451
rect 57897 20417 57931 20451
rect 4077 20349 4111 20383
rect 4261 20349 4295 20383
rect 5114 20349 5148 20383
rect 5273 20349 5307 20383
rect 7021 20349 7055 20383
rect 9689 20349 9723 20383
rect 10542 20349 10576 20383
rect 10701 20349 10735 20383
rect 11713 20349 11747 20383
rect 14933 20349 14967 20383
rect 15025 20349 15059 20383
rect 17417 20349 17451 20383
rect 18705 20349 18739 20383
rect 21097 20349 21131 20383
rect 24225 20349 24259 20383
rect 24317 20349 24351 20383
rect 25329 20349 25363 20383
rect 28641 20349 28675 20383
rect 28917 20349 28951 20383
rect 29837 20349 29871 20383
rect 32873 20349 32907 20383
rect 33517 20349 33551 20383
rect 33793 20349 33827 20383
rect 34529 20349 34563 20383
rect 36001 20349 36035 20383
rect 38025 20349 38059 20383
rect 38117 20349 38151 20383
rect 38577 20349 38611 20383
rect 39430 20349 39464 20383
rect 40877 20349 40911 20383
rect 43085 20349 43119 20383
rect 44925 20349 44959 20383
rect 45753 20349 45787 20383
rect 47777 20349 47811 20383
rect 48513 20349 48547 20383
rect 48630 20349 48664 20383
rect 48789 20349 48823 20383
rect 49985 20349 50019 20383
rect 50169 20349 50203 20383
rect 50445 20349 50479 20383
rect 51365 20349 51399 20383
rect 53205 20349 53239 20383
rect 53389 20349 53423 20383
rect 53757 20349 53791 20383
rect 55137 20349 55171 20383
rect 55229 20349 55263 20383
rect 55597 20349 55631 20383
rect 3433 20281 3467 20315
rect 4721 20281 4755 20315
rect 10149 20281 10183 20315
rect 18061 20281 18095 20315
rect 24869 20281 24903 20315
rect 39037 20281 39071 20315
rect 47409 20281 47443 20315
rect 48237 20281 48271 20315
rect 52561 20281 52595 20315
rect 5917 20213 5951 20247
rect 6377 20213 6411 20247
rect 9045 20213 9079 20247
rect 9413 20213 9447 20247
rect 11345 20213 11379 20247
rect 16405 20213 16439 20247
rect 16865 20213 16899 20247
rect 17969 20213 18003 20247
rect 19073 20213 19107 20247
rect 20913 20213 20947 20247
rect 21649 20213 21683 20247
rect 23765 20213 23799 20247
rect 27261 20213 27295 20247
rect 29561 20213 29595 20247
rect 31217 20213 31251 20247
rect 31861 20213 31895 20247
rect 34437 20213 34471 20247
rect 35909 20213 35943 20247
rect 36921 20213 36955 20247
rect 40233 20213 40267 20247
rect 42257 20213 42291 20247
rect 44741 20213 44775 20247
rect 45477 20213 45511 20247
rect 49433 20213 49467 20247
rect 52009 20213 52043 20247
rect 54677 20213 54711 20247
rect 58541 20213 58575 20247
rect 3801 20009 3835 20043
rect 6653 20009 6687 20043
rect 7665 20009 7699 20043
rect 8769 20009 8803 20043
rect 11897 20009 11931 20043
rect 18797 20009 18831 20043
rect 23857 20009 23891 20043
rect 28825 20009 28859 20043
rect 31769 20009 31803 20043
rect 33517 20009 33551 20043
rect 38393 20009 38427 20043
rect 38945 20009 38979 20043
rect 45017 20009 45051 20043
rect 55045 20009 55079 20043
rect 58265 20009 58299 20043
rect 3433 19941 3467 19975
rect 8953 19941 8987 19975
rect 13921 19941 13955 19975
rect 33425 19941 33459 19975
rect 52285 19941 52319 19975
rect 4445 19873 4479 19907
rect 6745 19873 6779 19907
rect 8217 19873 8251 19907
rect 9597 19873 9631 19907
rect 9781 19873 9815 19907
rect 12449 19873 12483 19907
rect 12541 19873 12575 19907
rect 14289 19873 14323 19907
rect 14933 19873 14967 19907
rect 15326 19873 15360 19907
rect 16681 19873 16715 19907
rect 16865 19873 16899 19907
rect 19901 19873 19935 19907
rect 20294 19873 20328 19907
rect 20453 19873 20487 19907
rect 21741 19873 21775 19907
rect 23305 19873 23339 19907
rect 29561 19873 29595 19907
rect 30205 19873 30239 19907
rect 30481 19873 30515 19907
rect 30598 19873 30632 19907
rect 30757 19873 30791 19907
rect 34161 19873 34195 19907
rect 34897 19873 34931 19907
rect 35357 19873 35391 19907
rect 35750 19873 35784 19907
rect 39497 19873 39531 19907
rect 42165 19873 42199 19907
rect 42533 19873 42567 19907
rect 42901 19873 42935 19907
rect 43361 19873 43395 19907
rect 43754 19873 43788 19907
rect 43913 19873 43947 19907
rect 45569 19873 45603 19907
rect 47961 19873 47995 19907
rect 48329 19873 48363 19907
rect 52377 19873 52411 19907
rect 54493 19873 54527 19907
rect 2053 19805 2087 19839
rect 4169 19805 4203 19839
rect 5273 19805 5307 19839
rect 10517 19805 10551 19839
rect 14473 19805 14507 19839
rect 15209 19805 15243 19839
rect 15485 19805 15519 19839
rect 16589 19805 16623 19839
rect 17325 19805 17359 19839
rect 17417 19805 17451 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 20177 19805 20211 19839
rect 21557 19805 21591 19839
rect 22017 19805 22051 19839
rect 27353 19805 27387 19839
rect 27445 19805 27479 19839
rect 29745 19805 29779 19839
rect 31401 19805 31435 19839
rect 32045 19805 32079 19839
rect 32312 19805 32346 19839
rect 34713 19805 34747 19839
rect 35633 19805 35667 19839
rect 35909 19805 35943 19839
rect 37013 19805 37047 19839
rect 38761 19805 38795 19839
rect 39865 19805 39899 19839
rect 42717 19805 42751 19839
rect 43637 19805 43671 19839
rect 45937 19805 45971 19839
rect 47869 19805 47903 19839
rect 48596 19805 48630 19839
rect 50905 19805 50939 19839
rect 51172 19805 51206 19839
rect 56885 19805 56919 19839
rect 57152 19805 57186 19839
rect 2320 19737 2354 19771
rect 5540 19737 5574 19771
rect 7389 19737 7423 19771
rect 9321 19737 9355 19771
rect 10425 19737 10459 19771
rect 10784 19737 10818 19771
rect 12808 19737 12842 19771
rect 17684 19737 17718 19771
rect 27712 19737 27746 19771
rect 36829 19737 36863 19771
rect 37280 19737 37314 19771
rect 39405 19737 39439 19771
rect 40132 19737 40166 19771
rect 46204 19737 46238 19771
rect 4261 19669 4295 19703
rect 5089 19669 5123 19703
rect 9413 19669 9447 19703
rect 16129 19669 16163 19703
rect 16221 19669 16255 19703
rect 21097 19669 21131 19703
rect 21189 19669 21223 19703
rect 21649 19669 21683 19703
rect 22661 19669 22695 19703
rect 24225 19669 24259 19703
rect 29285 19669 29319 19703
rect 33885 19669 33919 19703
rect 33977 19669 34011 19703
rect 36553 19669 36587 19703
rect 39313 19669 39347 19703
rect 41245 19669 41279 19703
rect 41521 19669 41555 19703
rect 41889 19669 41923 19703
rect 41981 19669 42015 19703
rect 44557 19669 44591 19703
rect 45385 19669 45419 19703
rect 45477 19669 45511 19703
rect 47317 19669 47351 19703
rect 47409 19669 47443 19703
rect 47777 19669 47811 19703
rect 49709 19669 49743 19703
rect 53021 19669 53055 19703
rect 54217 19669 54251 19703
rect 4077 19465 4111 19499
rect 4721 19465 4755 19499
rect 7021 19465 7055 19499
rect 7297 19465 7331 19499
rect 11345 19465 11379 19499
rect 16497 19465 16531 19499
rect 18705 19465 18739 19499
rect 21189 19465 21223 19499
rect 28641 19465 28675 19499
rect 29101 19465 29135 19499
rect 31217 19465 31251 19499
rect 33701 19465 33735 19499
rect 35725 19465 35759 19499
rect 35817 19465 35851 19499
rect 36185 19465 36219 19499
rect 36921 19465 36955 19499
rect 40233 19465 40267 19499
rect 44557 19465 44591 19499
rect 44649 19465 44683 19499
rect 46489 19465 46523 19499
rect 51457 19465 51491 19499
rect 51825 19465 51859 19499
rect 56977 19465 57011 19499
rect 57345 19465 57379 19499
rect 11989 19397 12023 19431
rect 13645 19397 13679 19431
rect 15025 19397 15059 19431
rect 17500 19397 17534 19431
rect 20076 19397 20110 19431
rect 43085 19397 43119 19431
rect 43444 19397 43478 19431
rect 48973 19397 49007 19431
rect 3525 19329 3559 19363
rect 6469 19329 6503 19363
rect 11897 19329 11931 19363
rect 13001 19329 13035 19363
rect 13553 19329 13587 19363
rect 14657 19329 14691 19363
rect 15117 19329 15151 19363
rect 15384 19329 15418 19363
rect 17141 19329 17175 19363
rect 17233 19329 17267 19363
rect 19073 19329 19107 19363
rect 19165 19329 19199 19363
rect 19809 19329 19843 19363
rect 27261 19329 27295 19363
rect 27528 19329 27562 19363
rect 29193 19329 29227 19363
rect 29837 19329 29871 19363
rect 30104 19329 30138 19363
rect 31309 19329 31343 19363
rect 32321 19329 32355 19363
rect 32588 19329 32622 19363
rect 34069 19329 34103 19363
rect 34345 19329 34379 19363
rect 34612 19329 34646 19363
rect 38761 19329 38795 19363
rect 40785 19329 40819 19363
rect 41052 19329 41086 19363
rect 42533 19329 42567 19363
rect 43177 19329 43211 19363
rect 45017 19329 45051 19363
rect 46121 19329 46155 19363
rect 47593 19329 47627 19363
rect 48237 19329 48271 19363
rect 48421 19329 48455 19363
rect 51917 19329 51951 19363
rect 58541 19329 58575 19363
rect 10793 19261 10827 19295
rect 12081 19261 12115 19295
rect 12357 19261 12391 19295
rect 13737 19261 13771 19295
rect 14105 19261 14139 19295
rect 19257 19261 19291 19295
rect 29285 19261 29319 19295
rect 36277 19261 36311 19295
rect 36461 19261 36495 19295
rect 39589 19261 39623 19295
rect 45109 19261 45143 19295
rect 45201 19261 45235 19295
rect 45569 19261 45603 19295
rect 50537 19261 50571 19295
rect 52009 19261 52043 19295
rect 54033 19261 54067 19295
rect 57437 19261 57471 19295
rect 57529 19261 57563 19295
rect 57897 19261 57931 19295
rect 11529 19193 11563 19227
rect 18613 19193 18647 19227
rect 37565 19193 37599 19227
rect 42165 19193 42199 19227
rect 6193 19125 6227 19159
rect 9229 19125 9263 19159
rect 9781 19125 9815 19159
rect 13185 19125 13219 19159
rect 21557 19125 21591 19159
rect 28733 19125 28767 19159
rect 31953 19125 31987 19159
rect 38301 19125 38335 19159
rect 39037 19125 39071 19159
rect 47225 19125 47259 19159
rect 50353 19125 50387 19159
rect 51181 19125 51215 19159
rect 54585 19125 54619 19159
rect 56793 19125 56827 19159
rect 12081 18921 12115 18955
rect 12909 18921 12943 18955
rect 13645 18921 13679 18955
rect 14933 18921 14967 18955
rect 16957 18921 16991 18955
rect 18337 18921 18371 18955
rect 19073 18921 19107 18955
rect 19901 18921 19935 18955
rect 28825 18921 28859 18955
rect 31677 18921 31711 18955
rect 33609 18921 33643 18955
rect 36185 18921 36219 18955
rect 41061 18921 41095 18955
rect 41981 18921 42015 18955
rect 42349 18921 42383 18955
rect 43085 18921 43119 18955
rect 44557 18921 44591 18955
rect 48421 18921 48455 18955
rect 50169 18921 50203 18955
rect 54125 18921 54159 18955
rect 57897 18921 57931 18955
rect 12449 18853 12483 18887
rect 27721 18853 27755 18887
rect 30205 18853 30239 18887
rect 34713 18853 34747 18887
rect 38393 18853 38427 18887
rect 45201 18853 45235 18887
rect 13093 18785 13127 18819
rect 14381 18785 14415 18819
rect 16313 18785 16347 18819
rect 18521 18785 18555 18819
rect 20453 18785 20487 18819
rect 25697 18785 25731 18819
rect 26433 18785 26467 18819
rect 28273 18785 28307 18819
rect 30113 18785 30147 18819
rect 30757 18785 30791 18819
rect 31033 18785 31067 18819
rect 33701 18785 33735 18819
rect 34345 18785 34379 18819
rect 35357 18785 35391 18819
rect 35541 18785 35575 18819
rect 36277 18785 36311 18819
rect 37013 18785 37047 18819
rect 39129 18785 39163 18819
rect 40417 18785 40451 18819
rect 41337 18785 41371 18819
rect 49985 18785 50019 18819
rect 50721 18785 50755 18819
rect 54677 18785 54711 18819
rect 55413 18785 55447 18819
rect 3065 18717 3099 18751
rect 4261 18717 4295 18751
rect 8953 18717 8987 18751
rect 20361 18717 20395 18751
rect 22753 18717 22787 18751
rect 23581 18717 23615 18751
rect 26157 18717 26191 18751
rect 26617 18717 26651 18751
rect 30573 18717 30607 18751
rect 47501 18717 47535 18751
rect 50997 18717 51031 18751
rect 52837 18717 52871 18751
rect 56517 18717 56551 18751
rect 35173 18649 35207 18683
rect 36921 18649 36955 18683
rect 37280 18649 37314 18683
rect 50537 18649 50571 18683
rect 51641 18649 51675 18683
rect 54493 18649 54527 18683
rect 55965 18649 55999 18683
rect 56784 18649 56818 18683
rect 3617 18581 3651 18615
rect 4813 18581 4847 18615
rect 5273 18581 5307 18615
rect 6009 18581 6043 18615
rect 9597 18581 9631 18615
rect 9965 18581 9999 18615
rect 19717 18581 19751 18615
rect 20269 18581 20303 18615
rect 23305 18581 23339 18615
rect 24133 18581 24167 18615
rect 25789 18581 25823 18615
rect 26249 18581 26283 18615
rect 27261 18581 27295 18615
rect 28089 18581 28123 18615
rect 29101 18581 29135 18615
rect 30665 18581 30699 18615
rect 35081 18581 35115 18615
rect 38485 18581 38519 18615
rect 38853 18581 38887 18615
rect 38945 18581 38979 18615
rect 48053 18581 48087 18615
rect 50629 18581 50663 18615
rect 53481 18581 53515 18615
rect 54033 18581 54067 18615
rect 54585 18581 54619 18615
rect 3433 18377 3467 18411
rect 4445 18377 4479 18411
rect 8401 18377 8435 18411
rect 19625 18377 19659 18411
rect 22845 18377 22879 18411
rect 23213 18377 23247 18411
rect 24869 18377 24903 18411
rect 38577 18377 38611 18411
rect 39313 18377 39347 18411
rect 48513 18377 48547 18411
rect 54861 18377 54895 18411
rect 57345 18377 57379 18411
rect 58541 18377 58575 18411
rect 4077 18309 4111 18343
rect 25504 18309 25538 18343
rect 49884 18309 49918 18343
rect 53748 18309 53782 18343
rect 55229 18309 55263 18343
rect 3341 18241 3375 18275
rect 4813 18241 4847 18275
rect 4905 18241 4939 18275
rect 5917 18241 5951 18275
rect 8769 18241 8803 18275
rect 8861 18241 8895 18275
rect 9873 18241 9907 18275
rect 23305 18241 23339 18275
rect 25237 18241 25271 18275
rect 29653 18241 29687 18275
rect 38025 18241 38059 18275
rect 38669 18241 38703 18275
rect 53481 18241 53515 18275
rect 55689 18241 55723 18275
rect 56542 18241 56576 18275
rect 2329 18173 2363 18207
rect 3617 18173 3651 18207
rect 5089 18173 5123 18207
rect 5273 18173 5307 18207
rect 6653 18173 6687 18207
rect 7757 18173 7791 18207
rect 9045 18173 9079 18207
rect 9229 18173 9263 18207
rect 11621 18173 11655 18207
rect 14657 18173 14691 18207
rect 20085 18173 20119 18207
rect 23397 18173 23431 18207
rect 23857 18173 23891 18207
rect 26985 18173 27019 18207
rect 28641 18173 28675 18207
rect 29193 18173 29227 18207
rect 29745 18173 29779 18207
rect 29837 18173 29871 18207
rect 30205 18173 30239 18207
rect 33333 18173 33367 18207
rect 33977 18173 34011 18207
rect 47593 18173 47627 18207
rect 49617 18173 49651 18207
rect 52837 18173 52871 18207
rect 55505 18173 55539 18207
rect 56149 18173 56183 18207
rect 56425 18173 56459 18207
rect 56701 18173 56735 18207
rect 57897 18173 57931 18207
rect 2973 18105 3007 18139
rect 26617 18105 26651 18139
rect 46949 18105 46983 18139
rect 2881 18037 2915 18071
rect 7297 18037 7331 18071
rect 8309 18037 8343 18071
rect 10149 18037 10183 18071
rect 12265 18037 12299 18071
rect 12633 18037 12667 18071
rect 13921 18037 13955 18071
rect 15301 18037 15335 18071
rect 20729 18037 20763 18071
rect 22661 18037 22695 18071
rect 24501 18037 24535 18071
rect 27629 18037 27663 18071
rect 29285 18037 29319 18071
rect 30849 18037 30883 18071
rect 33885 18037 33919 18071
rect 34621 18037 34655 18071
rect 34989 18037 35023 18071
rect 35633 18037 35667 18071
rect 41429 18037 41463 18071
rect 47409 18037 47443 18071
rect 48237 18037 48271 18071
rect 50997 18037 51031 18071
rect 52561 18037 52595 18071
rect 53389 18037 53423 18071
rect 3249 17833 3283 17867
rect 8953 17833 8987 17867
rect 26249 17833 26283 17867
rect 26341 17833 26375 17867
rect 30205 17833 30239 17867
rect 57437 17833 57471 17867
rect 57529 17833 57563 17867
rect 8769 17765 8803 17799
rect 19993 17765 20027 17799
rect 23581 17765 23615 17799
rect 47041 17765 47075 17799
rect 3801 17697 3835 17731
rect 4445 17697 4479 17731
rect 9505 17697 9539 17731
rect 10517 17697 10551 17731
rect 12633 17697 12667 17731
rect 20545 17697 20579 17731
rect 20821 17697 20855 17731
rect 24593 17697 24627 17731
rect 25053 17697 25087 17731
rect 25446 17697 25480 17731
rect 26985 17697 27019 17731
rect 28825 17697 28859 17731
rect 30113 17697 30147 17731
rect 30757 17697 30791 17731
rect 33057 17697 33091 17731
rect 33241 17697 33275 17731
rect 34253 17697 34287 17731
rect 40785 17697 40819 17731
rect 43821 17697 43855 17731
rect 44557 17697 44591 17731
rect 46397 17697 46431 17731
rect 47685 17697 47719 17731
rect 48329 17697 48363 17731
rect 48789 17697 48823 17731
rect 49182 17697 49216 17731
rect 49341 17697 49375 17731
rect 50813 17697 50847 17731
rect 51181 17697 51215 17731
rect 58081 17697 58115 17731
rect 1869 17629 1903 17663
rect 3985 17629 4019 17663
rect 4721 17629 4755 17663
rect 4859 17629 4893 17663
rect 4997 17629 5031 17663
rect 5733 17629 5767 17663
rect 7389 17629 7423 17663
rect 9781 17629 9815 17663
rect 10784 17629 10818 17663
rect 12357 17629 12391 17663
rect 12909 17629 12943 17663
rect 14197 17629 14231 17663
rect 15669 17629 15703 17663
rect 17601 17629 17635 17663
rect 20361 17629 20395 17663
rect 22201 17629 22235 17663
rect 22468 17629 22502 17663
rect 24409 17629 24443 17663
rect 25329 17629 25363 17663
rect 25605 17629 25639 17663
rect 26709 17629 26743 17663
rect 27629 17629 27663 17663
rect 30665 17629 30699 17663
rect 31125 17629 31159 17663
rect 32873 17629 32907 17663
rect 34713 17629 34747 17663
rect 38393 17629 38427 17663
rect 40141 17629 40175 17663
rect 41521 17629 41555 17663
rect 44281 17629 44315 17663
rect 45201 17629 45235 17663
rect 48145 17629 48179 17663
rect 49065 17629 49099 17663
rect 50537 17629 50571 17663
rect 51733 17629 51767 17663
rect 56057 17629 56091 17663
rect 57897 17629 57931 17663
rect 2136 17561 2170 17595
rect 6000 17561 6034 17595
rect 7656 17561 7690 17595
rect 9321 17561 9355 17595
rect 10425 17561 10459 17595
rect 12449 17561 12483 17595
rect 14464 17561 14498 17595
rect 16313 17561 16347 17595
rect 26801 17561 26835 17595
rect 30573 17561 30607 17595
rect 31677 17561 31711 17595
rect 39589 17561 39623 17595
rect 49985 17561 50019 17595
rect 50629 17561 50663 17595
rect 52000 17561 52034 17595
rect 53205 17561 53239 17595
rect 55505 17561 55539 17595
rect 56324 17561 56358 17595
rect 5641 17493 5675 17527
rect 7113 17493 7147 17527
rect 9413 17493 9447 17527
rect 11897 17493 11931 17527
rect 11989 17493 12023 17527
rect 13461 17493 13495 17527
rect 13829 17493 13863 17527
rect 15577 17493 15611 17527
rect 18153 17493 18187 17527
rect 19901 17493 19935 17527
rect 20453 17493 20487 17527
rect 21465 17493 21499 17527
rect 22109 17493 22143 17527
rect 24133 17493 24167 17527
rect 27353 17493 27387 17527
rect 28273 17493 28307 17527
rect 29377 17493 29411 17527
rect 32413 17493 32447 17527
rect 32781 17493 32815 17527
rect 33885 17493 33919 17527
rect 35357 17493 35391 17527
rect 37749 17493 37783 17527
rect 38209 17493 38243 17527
rect 38945 17493 38979 17527
rect 40693 17493 40727 17527
rect 41429 17493 41463 17527
rect 42165 17493 42199 17527
rect 43913 17493 43947 17527
rect 44373 17493 44407 17527
rect 45845 17493 45879 17527
rect 46949 17493 46983 17527
rect 47409 17493 47443 17527
rect 47501 17493 47535 17527
rect 50169 17493 50203 17527
rect 53113 17493 53147 17527
rect 54493 17493 54527 17527
rect 57989 17493 58023 17527
rect 3157 17289 3191 17323
rect 5825 17289 5859 17323
rect 6377 17289 6411 17323
rect 6745 17289 6779 17323
rect 9137 17289 9171 17323
rect 11345 17289 11379 17323
rect 11529 17289 11563 17323
rect 13001 17289 13035 17323
rect 13461 17289 13495 17323
rect 14473 17289 14507 17323
rect 14749 17289 14783 17323
rect 15209 17289 15243 17323
rect 17693 17289 17727 17323
rect 23581 17289 23615 17323
rect 24133 17289 24167 17323
rect 25881 17289 25915 17323
rect 29193 17289 29227 17323
rect 31861 17289 31895 17323
rect 33793 17289 33827 17323
rect 34253 17289 34287 17323
rect 41245 17289 41279 17323
rect 41521 17289 41555 17323
rect 44925 17289 44959 17323
rect 47409 17289 47443 17323
rect 47593 17289 47627 17323
rect 47961 17289 47995 17323
rect 49341 17289 49375 17323
rect 52745 17289 52779 17323
rect 53205 17289 53239 17323
rect 55045 17289 55079 17323
rect 56793 17289 56827 17323
rect 3792 17221 3826 17255
rect 5733 17221 5767 17255
rect 8024 17221 8058 17255
rect 13369 17221 13403 17255
rect 15945 17221 15979 17255
rect 18061 17221 18095 17255
rect 19533 17221 19567 17255
rect 21281 17221 21315 17255
rect 24041 17221 24075 17255
rect 28080 17221 28114 17255
rect 32404 17221 32438 17255
rect 37565 17221 37599 17255
rect 40132 17221 40166 17255
rect 52469 17221 52503 17255
rect 1777 17153 1811 17187
rect 2044 17153 2078 17187
rect 3525 17153 3559 17187
rect 7757 17153 7791 17187
rect 10542 17153 10576 17187
rect 11897 17153 11931 17187
rect 13829 17153 13863 17187
rect 15117 17153 15151 17187
rect 18153 17153 18187 17187
rect 19165 17153 19199 17187
rect 19625 17153 19659 17187
rect 19892 17153 19926 17187
rect 22201 17153 22235 17187
rect 22468 17153 22502 17187
rect 24501 17153 24535 17187
rect 24768 17153 24802 17187
rect 25973 17153 26007 17187
rect 29745 17153 29779 17187
rect 31493 17153 31527 17187
rect 32137 17153 32171 17187
rect 34161 17153 34195 17187
rect 35173 17153 35207 17187
rect 36277 17153 36311 17187
rect 38117 17153 38151 17187
rect 39865 17153 39899 17187
rect 41889 17153 41923 17187
rect 43085 17153 43119 17187
rect 43812 17153 43846 17187
rect 45661 17153 45695 17187
rect 46029 17153 46063 17187
rect 46296 17153 46330 17187
rect 48053 17153 48087 17187
rect 49433 17153 49467 17187
rect 51181 17153 51215 17187
rect 53113 17153 53147 17187
rect 53932 17153 53966 17187
rect 55781 17153 55815 17187
rect 56885 17153 56919 17187
rect 58541 17153 58575 17187
rect 5917 17085 5951 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 7389 17085 7423 17119
rect 9505 17085 9539 17119
rect 9689 17085 9723 17119
rect 10425 17085 10459 17119
rect 10701 17085 10735 17119
rect 11989 17085 12023 17119
rect 12081 17085 12115 17119
rect 12909 17085 12943 17119
rect 13645 17085 13679 17119
rect 15393 17085 15427 17119
rect 16221 17085 16255 17119
rect 17601 17085 17635 17119
rect 18245 17085 18279 17119
rect 18613 17085 18647 17119
rect 24317 17085 24351 17119
rect 27813 17085 27847 17119
rect 34345 17085 34379 17119
rect 35265 17085 35299 17119
rect 35449 17085 35483 17119
rect 35633 17085 35667 17119
rect 36369 17085 36403 17119
rect 37933 17085 37967 17119
rect 38577 17085 38611 17119
rect 38853 17085 38887 17119
rect 38991 17085 39025 17119
rect 39129 17085 39163 17119
rect 41981 17085 42015 17119
rect 42073 17085 42107 17119
rect 42441 17085 42475 17119
rect 43545 17085 43579 17119
rect 45017 17085 45051 17119
rect 48145 17085 48179 17119
rect 49525 17085 49559 17119
rect 49801 17085 49835 17119
rect 50537 17085 50571 17119
rect 53297 17085 53331 17119
rect 53665 17085 53699 17119
rect 55137 17085 55171 17119
rect 56977 17085 57011 17119
rect 57897 17085 57931 17119
rect 4905 17017 4939 17051
rect 10149 17017 10183 17051
rect 34805 17017 34839 17051
rect 48605 17017 48639 17051
rect 48973 17017 49007 17051
rect 5365 16949 5399 16983
rect 21005 16949 21039 16983
rect 23673 16949 23707 16983
rect 26617 16949 26651 16983
rect 27261 16949 27295 16983
rect 29561 16949 29595 16983
rect 33517 16949 33551 16983
rect 37013 16949 37047 16983
rect 39773 16949 39807 16983
rect 43453 16949 43487 16983
rect 50445 16949 50479 16983
rect 56333 16949 56367 16983
rect 56425 16949 56459 16983
rect 57437 16949 57471 16983
rect 2789 16745 2823 16779
rect 6101 16745 6135 16779
rect 6929 16745 6963 16779
rect 11897 16745 11931 16779
rect 12173 16745 12207 16779
rect 18337 16745 18371 16779
rect 22201 16745 22235 16779
rect 23765 16745 23799 16779
rect 24133 16745 24167 16779
rect 29377 16745 29411 16779
rect 29837 16745 29871 16779
rect 31677 16745 31711 16779
rect 32965 16745 32999 16779
rect 36461 16745 36495 16779
rect 38945 16745 38979 16779
rect 39865 16745 39899 16779
rect 42165 16745 42199 16779
rect 44557 16745 44591 16779
rect 45017 16745 45051 16779
rect 49801 16745 49835 16779
rect 54217 16745 54251 16779
rect 57069 16745 57103 16779
rect 2881 16677 2915 16711
rect 9321 16677 9355 16711
rect 9689 16677 9723 16711
rect 13737 16677 13771 16711
rect 34529 16677 34563 16711
rect 38025 16677 38059 16711
rect 46029 16677 46063 16711
rect 55965 16677 55999 16711
rect 2237 16609 2271 16643
rect 3341 16609 3375 16643
rect 3525 16609 3559 16643
rect 3893 16609 3927 16643
rect 5825 16609 5859 16643
rect 6377 16609 6411 16643
rect 11345 16609 11379 16643
rect 14105 16609 14139 16643
rect 14289 16609 14323 16643
rect 14749 16609 14783 16643
rect 15025 16609 15059 16643
rect 15301 16609 15335 16643
rect 15945 16609 15979 16643
rect 16497 16609 16531 16643
rect 16589 16609 16623 16643
rect 16957 16609 16991 16643
rect 19257 16609 19291 16643
rect 19441 16609 19475 16643
rect 19901 16609 19935 16643
rect 21097 16609 21131 16643
rect 21649 16609 21683 16643
rect 21833 16609 21867 16643
rect 23213 16609 23247 16643
rect 24869 16609 24903 16643
rect 25513 16609 25547 16643
rect 25697 16609 25731 16643
rect 27353 16609 27387 16643
rect 29929 16609 29963 16643
rect 33149 16609 33183 16643
rect 34713 16609 34747 16643
rect 36645 16609 36679 16643
rect 38669 16609 38703 16643
rect 39589 16609 39623 16643
rect 40417 16609 40451 16643
rect 42717 16609 42751 16643
rect 43361 16609 43395 16643
rect 43754 16609 43788 16643
rect 45477 16609 45511 16643
rect 45661 16609 45695 16643
rect 48421 16609 48455 16643
rect 51733 16609 51767 16643
rect 54677 16609 54711 16643
rect 54769 16609 54803 16643
rect 55413 16609 55447 16643
rect 56425 16609 56459 16643
rect 12357 16541 12391 16575
rect 12624 16541 12658 16575
rect 15142 16541 15176 16575
rect 16405 16541 16439 16575
rect 17224 16541 17258 16575
rect 18521 16541 18555 16575
rect 20177 16541 20211 16575
rect 20294 16541 20328 16575
rect 20453 16541 20487 16575
rect 25421 16541 25455 16575
rect 26709 16541 26743 16575
rect 27620 16541 27654 16575
rect 30196 16541 30230 16575
rect 32137 16541 32171 16575
rect 33416 16541 33450 16575
rect 34980 16541 35014 16575
rect 40785 16541 40819 16575
rect 41052 16541 41086 16575
rect 42901 16541 42935 16575
rect 43637 16541 43671 16575
rect 43913 16541 43947 16575
rect 46489 16541 46523 16575
rect 48688 16541 48722 16575
rect 53205 16541 53239 16575
rect 54585 16541 54619 16575
rect 3249 16473 3283 16507
rect 4445 16473 4479 16507
rect 21557 16473 21591 16507
rect 26249 16473 26283 16507
rect 36912 16473 36946 16507
rect 40233 16473 40267 16507
rect 45385 16473 45419 16507
rect 46756 16473 46790 16507
rect 52000 16473 52034 16507
rect 53849 16473 53883 16507
rect 16037 16405 16071 16439
rect 19073 16405 19107 16439
rect 21189 16405 21223 16439
rect 25053 16405 25087 16439
rect 27261 16405 27295 16439
rect 28733 16405 28767 16439
rect 31309 16405 31343 16439
rect 32689 16405 32723 16439
rect 36093 16405 36127 16439
rect 38117 16405 38151 16439
rect 38485 16405 38519 16439
rect 38577 16405 38611 16439
rect 39313 16405 39347 16439
rect 39405 16405 39439 16439
rect 40325 16405 40359 16439
rect 42533 16405 42567 16439
rect 47869 16405 47903 16439
rect 53113 16405 53147 16439
rect 3709 16201 3743 16235
rect 8217 16201 8251 16235
rect 14013 16201 14047 16235
rect 18337 16201 18371 16235
rect 18797 16201 18831 16235
rect 20913 16201 20947 16235
rect 25605 16201 25639 16235
rect 27445 16201 27479 16235
rect 27629 16201 27663 16235
rect 28089 16201 28123 16235
rect 30757 16201 30791 16235
rect 32229 16201 32263 16235
rect 32689 16201 32723 16235
rect 33333 16201 33367 16235
rect 35725 16201 35759 16235
rect 37013 16201 37047 16235
rect 38669 16201 38703 16235
rect 39037 16201 39071 16235
rect 39681 16201 39715 16235
rect 40601 16201 40635 16235
rect 42257 16201 42291 16235
rect 44925 16201 44959 16235
rect 45937 16201 45971 16235
rect 48329 16201 48363 16235
rect 51089 16201 51123 16235
rect 51457 16201 51491 16235
rect 52745 16201 52779 16235
rect 54585 16201 54619 16235
rect 18889 16133 18923 16167
rect 37556 16133 37590 16167
rect 39589 16133 39623 16167
rect 9045 16065 9079 16099
rect 11069 16065 11103 16099
rect 12348 16065 12382 16099
rect 13921 16065 13955 16099
rect 15025 16065 15059 16099
rect 16957 16065 16991 16099
rect 17224 16065 17258 16099
rect 19800 16065 19834 16099
rect 25053 16065 25087 16099
rect 27997 16065 28031 16099
rect 28457 16065 28491 16099
rect 28641 16065 28675 16099
rect 29653 16065 29687 16099
rect 32597 16065 32631 16099
rect 33425 16065 33459 16099
rect 34345 16065 34379 16099
rect 37289 16065 37323 16099
rect 40877 16065 40911 16099
rect 41144 16065 41178 16099
rect 43085 16065 43119 16099
rect 43812 16065 43846 16099
rect 45661 16065 45695 16099
rect 47777 16065 47811 16099
rect 53113 16065 53147 16099
rect 54217 16065 54251 16099
rect 5457 15997 5491 16031
rect 12081 15997 12115 16031
rect 14197 15997 14231 16031
rect 14473 15997 14507 16031
rect 15117 15997 15151 16031
rect 19073 15997 19107 16031
rect 19533 15997 19567 16031
rect 21005 15997 21039 16031
rect 28181 15997 28215 16031
rect 29377 15997 29411 16031
rect 29515 15997 29549 16031
rect 30297 15997 30331 16031
rect 30849 15997 30883 16031
rect 30941 15997 30975 16031
rect 32873 15997 32907 16031
rect 33609 15997 33643 16031
rect 34462 15997 34496 16031
rect 34621 15997 34655 16031
rect 35265 15997 35299 16031
rect 35817 15997 35851 16031
rect 36001 15997 36035 16031
rect 39865 15997 39899 16031
rect 42441 15997 42475 16031
rect 43545 15997 43579 16031
rect 45017 15997 45051 16031
rect 53205 15997 53239 16031
rect 53389 15997 53423 16031
rect 53573 15997 53607 16031
rect 55689 15997 55723 16031
rect 57897 15997 57931 16031
rect 13461 15929 13495 15963
rect 26801 15929 26835 15963
rect 29101 15929 29135 15963
rect 34069 15929 34103 15963
rect 46765 15929 46799 15963
rect 6009 15861 6043 15895
rect 10333 15861 10367 15895
rect 13553 15861 13587 15895
rect 15761 15861 15795 15895
rect 18429 15861 18463 15895
rect 21649 15861 21683 15895
rect 23581 15861 23615 15895
rect 30389 15861 30423 15895
rect 35357 15861 35391 15895
rect 39221 15861 39255 15895
rect 40325 15861 40359 15895
rect 43453 15861 43487 15895
rect 46397 15861 46431 15895
rect 48881 15861 48915 15895
rect 52561 15861 52595 15895
rect 55229 15861 55263 15895
rect 56241 15861 56275 15895
rect 58541 15861 58575 15895
rect 5549 15657 5583 15691
rect 11161 15657 11195 15691
rect 13645 15657 13679 15691
rect 14381 15657 14415 15691
rect 18521 15657 18555 15691
rect 19533 15657 19567 15691
rect 21373 15657 21407 15691
rect 28089 15657 28123 15691
rect 33609 15657 33643 15691
rect 34897 15657 34931 15691
rect 38209 15657 38243 15691
rect 38945 15657 38979 15691
rect 39681 15657 39715 15691
rect 41429 15657 41463 15691
rect 41521 15657 41555 15691
rect 43913 15657 43947 15691
rect 46305 15657 46339 15691
rect 48605 15657 48639 15691
rect 50445 15657 50479 15691
rect 56333 15657 56367 15691
rect 19901 15589 19935 15623
rect 32873 15589 32907 15623
rect 48329 15589 48363 15623
rect 52009 15589 52043 15623
rect 55321 15589 55355 15623
rect 6101 15521 6135 15555
rect 7941 15521 7975 15555
rect 9781 15521 9815 15555
rect 11989 15521 12023 15555
rect 13093 15521 13127 15555
rect 14749 15521 14783 15555
rect 17969 15521 18003 15555
rect 20545 15521 20579 15555
rect 20729 15521 20763 15555
rect 26709 15521 26743 15555
rect 28641 15521 28675 15555
rect 28825 15521 28859 15555
rect 29745 15521 29779 15555
rect 33057 15521 33091 15555
rect 37657 15521 37691 15555
rect 38393 15521 38427 15555
rect 42073 15521 42107 15555
rect 42441 15521 42475 15555
rect 43821 15521 43855 15555
rect 44557 15521 44591 15555
rect 45017 15521 45051 15555
rect 51365 15521 51399 15555
rect 51549 15521 51583 15555
rect 52561 15521 52595 15555
rect 53849 15521 53883 15555
rect 54585 15521 54619 15555
rect 55873 15521 55907 15555
rect 56793 15521 56827 15555
rect 6469 15453 6503 15487
rect 8125 15453 8159 15487
rect 8953 15453 8987 15487
rect 11253 15453 11287 15487
rect 15016 15453 15050 15487
rect 16221 15453 16255 15487
rect 20361 15453 20395 15487
rect 22845 15453 22879 15487
rect 25513 15453 25547 15487
rect 30205 15453 30239 15487
rect 31493 15453 31527 15487
rect 31760 15453 31794 15487
rect 39037 15453 39071 15487
rect 50721 15453 50755 15487
rect 52285 15453 52319 15487
rect 52402 15453 52436 15487
rect 53665 15453 53699 15487
rect 7665 15385 7699 15419
rect 10048 15385 10082 15419
rect 11897 15385 11931 15419
rect 26976 15385 27010 15419
rect 28549 15385 28583 15419
rect 41889 15385 41923 15419
rect 44281 15385 44315 15419
rect 45661 15385 45695 15419
rect 53205 15385 53239 15419
rect 53757 15385 53791 15419
rect 57060 15385 57094 15419
rect 5917 15317 5951 15351
rect 6009 15317 6043 15351
rect 7021 15317 7055 15351
rect 7297 15317 7331 15351
rect 7757 15317 7791 15351
rect 8769 15317 8803 15351
rect 9597 15317 9631 15351
rect 12633 15317 12667 15351
rect 16129 15317 16163 15351
rect 16865 15317 16899 15351
rect 18889 15317 18923 15351
rect 20269 15317 20303 15351
rect 23397 15317 23431 15351
rect 26065 15317 26099 15351
rect 28181 15317 28215 15351
rect 29285 15317 29319 15351
rect 31309 15317 31343 15351
rect 33977 15317 34011 15351
rect 35357 15317 35391 15351
rect 40141 15317 40175 15351
rect 41981 15317 42015 15351
rect 42993 15317 43027 15351
rect 44373 15317 44407 15351
rect 47409 15317 47443 15351
rect 51273 15317 51307 15351
rect 53297 15317 53331 15351
rect 55137 15317 55171 15351
rect 55689 15317 55723 15351
rect 55781 15317 55815 15351
rect 58173 15317 58207 15351
rect 6193 15113 6227 15147
rect 6561 15113 6595 15147
rect 10057 15113 10091 15147
rect 10241 15113 10275 15147
rect 10701 15113 10735 15147
rect 13461 15113 13495 15147
rect 15117 15113 15151 15147
rect 15485 15113 15519 15147
rect 18337 15113 18371 15147
rect 20361 15113 20395 15147
rect 21189 15113 21223 15147
rect 21557 15113 21591 15147
rect 26709 15113 26743 15147
rect 28273 15113 28307 15147
rect 29009 15113 29043 15147
rect 33149 15113 33183 15147
rect 40417 15113 40451 15147
rect 42717 15113 42751 15147
rect 48973 15113 49007 15147
rect 50721 15113 50755 15147
rect 53113 15113 53147 15147
rect 53849 15113 53883 15147
rect 58541 15113 58575 15147
rect 8944 15045 8978 15079
rect 22284 15045 22318 15079
rect 24225 15045 24259 15079
rect 45477 15045 45511 15079
rect 4813 14977 4847 15011
rect 5080 14977 5114 15011
rect 6929 14977 6963 15011
rect 10609 14977 10643 15011
rect 15577 14977 15611 15011
rect 22017 14977 22051 15011
rect 24317 14977 24351 15011
rect 24584 14977 24618 15011
rect 26433 14977 26467 15011
rect 27721 14977 27755 15011
rect 45569 14977 45603 15011
rect 47317 14977 47351 15011
rect 47860 14977 47894 15011
rect 51089 14977 51123 15011
rect 52193 14977 52227 15011
rect 54208 14977 54242 15011
rect 55873 14977 55907 15011
rect 56885 14977 56919 15011
rect 6745 14909 6779 14943
rect 7665 14909 7699 14943
rect 7782 14909 7816 14943
rect 7941 14909 7975 14943
rect 8677 14909 8711 14943
rect 10793 14909 10827 14943
rect 11253 14909 11287 14943
rect 15669 14909 15703 14943
rect 19165 14909 19199 14943
rect 23673 14909 23707 14943
rect 25881 14909 25915 14943
rect 28365 14909 28399 14943
rect 36553 14909 36587 14943
rect 43545 14909 43579 14943
rect 45661 14909 45695 14943
rect 45937 14909 45971 14943
rect 46765 14909 46799 14943
rect 47593 14909 47627 14943
rect 49065 14909 49099 14943
rect 49801 14909 49835 14943
rect 51181 14909 51215 14943
rect 51365 14909 51399 14943
rect 51641 14909 51675 14943
rect 53941 14909 53975 14943
rect 55689 14909 55723 14943
rect 56609 14909 56643 14943
rect 56726 14909 56760 14943
rect 57897 14909 57931 14943
rect 7389 14841 7423 14875
rect 40141 14841 40175 14875
rect 45109 14841 45143 14875
rect 50445 14841 50479 14875
rect 56333 14841 56367 14875
rect 8585 14773 8619 14807
rect 14933 14773 14967 14807
rect 18889 14773 18923 14807
rect 19717 14773 19751 14807
rect 20085 14773 20119 14807
rect 23397 14773 23431 14807
rect 25697 14773 25731 14807
rect 27445 14773 27479 14807
rect 33517 14773 33551 14807
rect 37105 14773 37139 14807
rect 37473 14773 37507 14807
rect 39681 14773 39715 14807
rect 44189 14773 44223 14807
rect 44925 14773 44959 14807
rect 46581 14773 46615 14807
rect 49709 14773 49743 14807
rect 55321 14773 55355 14807
rect 57529 14773 57563 14807
rect 6101 14569 6135 14603
rect 8125 14569 8159 14603
rect 8953 14569 8987 14603
rect 19257 14569 19291 14603
rect 23213 14569 23247 14603
rect 26065 14569 26099 14603
rect 31033 14569 31067 14603
rect 32413 14569 32447 14603
rect 41705 14569 41739 14603
rect 49249 14569 49283 14603
rect 51549 14569 51583 14603
rect 55137 14569 55171 14603
rect 57529 14569 57563 14603
rect 57621 14569 57655 14603
rect 31861 14501 31895 14535
rect 39865 14501 39899 14535
rect 42717 14501 42751 14535
rect 46397 14501 46431 14535
rect 4721 14433 4755 14467
rect 9413 14433 9447 14467
rect 9505 14433 9539 14467
rect 9873 14433 9907 14467
rect 19809 14433 19843 14467
rect 21741 14433 21775 14467
rect 23765 14433 23799 14467
rect 26525 14433 26559 14467
rect 26617 14433 26651 14467
rect 34805 14433 34839 14467
rect 39129 14433 39163 14467
rect 40417 14433 40451 14467
rect 42441 14433 42475 14467
rect 43361 14433 43395 14467
rect 43545 14433 43579 14467
rect 47133 14433 47167 14467
rect 47409 14433 47443 14467
rect 47685 14433 47719 14467
rect 48973 14433 49007 14467
rect 49709 14433 49743 14467
rect 49801 14433 49835 14467
rect 52285 14433 52319 14467
rect 53757 14433 53791 14467
rect 55781 14433 55815 14467
rect 55873 14433 55907 14467
rect 58173 14433 58207 14467
rect 2237 14365 2271 14399
rect 6745 14365 6779 14399
rect 12357 14365 12391 14399
rect 14289 14365 14323 14399
rect 17601 14365 17635 14399
rect 18245 14365 18279 14399
rect 20085 14365 20119 14399
rect 20821 14365 20855 14399
rect 24593 14365 24627 14399
rect 26893 14365 26927 14399
rect 28089 14365 28123 14399
rect 28825 14365 28859 14399
rect 29929 14365 29963 14399
rect 35909 14365 35943 14399
rect 37381 14365 37415 14399
rect 40693 14365 40727 14399
rect 42257 14365 42291 14399
rect 43085 14365 43119 14399
rect 45017 14365 45051 14399
rect 45284 14365 45318 14399
rect 46489 14365 46523 14399
rect 46673 14365 46707 14399
rect 47526 14365 47560 14399
rect 50169 14365 50203 14399
rect 52469 14365 52503 14399
rect 56149 14365 56183 14399
rect 57989 14365 58023 14399
rect 4988 14297 5022 14331
rect 7012 14297 7046 14331
rect 9321 14297 9355 14331
rect 10425 14297 10459 14331
rect 22008 14297 22042 14331
rect 23581 14297 23615 14331
rect 23673 14297 23707 14331
rect 24860 14297 24894 14331
rect 36176 14297 36210 14331
rect 40233 14297 40267 14331
rect 41337 14297 41371 14331
rect 43177 14297 43211 14331
rect 50436 14297 50470 14331
rect 54024 14297 54058 14331
rect 55689 14297 55723 14331
rect 56416 14297 56450 14331
rect 2881 14229 2915 14263
rect 6653 14229 6687 14263
rect 8769 14229 8803 14263
rect 12909 14229 12943 14263
rect 14933 14229 14967 14263
rect 17325 14229 17359 14263
rect 18153 14229 18187 14263
rect 18889 14229 18923 14263
rect 19625 14229 19659 14263
rect 19717 14229 19751 14263
rect 20729 14229 20763 14263
rect 21465 14229 21499 14263
rect 23121 14229 23155 14263
rect 25973 14229 26007 14263
rect 26433 14229 26467 14263
rect 27537 14229 27571 14263
rect 28641 14229 28675 14263
rect 29377 14229 29411 14263
rect 30573 14229 30607 14263
rect 31401 14229 31435 14263
rect 35357 14229 35391 14263
rect 37289 14229 37323 14263
rect 38025 14229 38059 14263
rect 39681 14229 39715 14263
rect 40325 14229 40359 14263
rect 41889 14229 41923 14263
rect 42349 14229 42383 14263
rect 44189 14229 44223 14263
rect 44741 14229 44775 14263
rect 48329 14229 48363 14263
rect 48421 14229 48455 14263
rect 48789 14229 48823 14263
rect 48881 14229 48915 14263
rect 49617 14229 49651 14263
rect 51641 14229 51675 14263
rect 52009 14229 52043 14263
rect 52101 14229 52135 14263
rect 53113 14229 53147 14263
rect 55321 14229 55355 14263
rect 58081 14229 58115 14263
rect 3249 14025 3283 14059
rect 5917 14025 5951 14059
rect 7849 14025 7883 14059
rect 10241 14025 10275 14059
rect 14105 14025 14139 14059
rect 14565 14025 14599 14059
rect 18061 14025 18095 14059
rect 19993 14025 20027 14059
rect 20085 14025 20119 14059
rect 25789 14025 25823 14059
rect 28181 14025 28215 14059
rect 28641 14025 28675 14059
rect 31677 14025 31711 14059
rect 33977 14025 34011 14059
rect 34989 14025 35023 14059
rect 37289 14025 37323 14059
rect 37749 14025 37783 14059
rect 39865 14025 39899 14059
rect 42257 14025 42291 14059
rect 46305 14025 46339 14059
rect 49709 14025 49743 14059
rect 55413 14025 55447 14059
rect 56149 14025 56183 14059
rect 56885 14025 56919 14059
rect 2136 13957 2170 13991
rect 11796 13957 11830 13991
rect 18880 13957 18914 13991
rect 22293 13957 22327 13991
rect 29828 13957 29862 13991
rect 36921 13957 36955 13991
rect 42708 13957 42742 13991
rect 46213 13957 46247 13991
rect 47317 13957 47351 13991
rect 1869 13889 1903 13923
rect 3341 13889 3375 13923
rect 5825 13889 5859 13923
rect 7021 13889 7055 13923
rect 7297 13889 7331 13923
rect 14473 13889 14507 13923
rect 15117 13889 15151 13923
rect 16948 13889 16982 13923
rect 18613 13889 18647 13923
rect 20453 13889 20487 13923
rect 21557 13889 21591 13923
rect 22845 13889 22879 13923
rect 23673 13889 23707 13923
rect 24547 13889 24581 13923
rect 26433 13889 26467 13923
rect 27353 13889 27387 13923
rect 28549 13889 28583 13923
rect 29561 13889 29595 13923
rect 32597 13889 32631 13923
rect 32864 13889 32898 13923
rect 34713 13889 34747 13923
rect 35532 13889 35566 13923
rect 37657 13889 37691 13923
rect 38485 13889 38519 13923
rect 38752 13889 38786 13923
rect 40417 13889 40451 13923
rect 40601 13889 40635 13923
rect 44640 13889 44674 13923
rect 46765 13889 46799 13923
rect 47860 13889 47894 13923
rect 49065 13889 49099 13923
rect 50261 13889 50295 13923
rect 50528 13889 50562 13923
rect 51733 13889 51767 13923
rect 52377 13889 52411 13923
rect 54861 13889 54895 13923
rect 55597 13889 55631 13923
rect 56977 13889 57011 13923
rect 58541 13889 58575 13923
rect 6009 13821 6043 13855
rect 6469 13821 6503 13855
rect 9229 13821 9263 13855
rect 11529 13821 11563 13855
rect 13093 13821 13127 13855
rect 14013 13821 14047 13855
rect 14749 13821 14783 13855
rect 16681 13821 16715 13855
rect 18521 13821 18555 13855
rect 20545 13821 20579 13855
rect 20637 13821 20671 13855
rect 21005 13821 21039 13855
rect 22937 13821 22971 13855
rect 23121 13821 23155 13855
rect 23489 13821 23523 13855
rect 24409 13821 24443 13855
rect 24685 13821 24719 13855
rect 25881 13821 25915 13855
rect 26065 13821 26099 13855
rect 27445 13821 27479 13855
rect 28733 13821 28767 13855
rect 31033 13821 31067 13855
rect 34069 13821 34103 13855
rect 35265 13821 35299 13855
rect 37841 13821 37875 13855
rect 38301 13821 38335 13855
rect 41337 13821 41371 13855
rect 41454 13821 41488 13855
rect 41613 13821 41647 13855
rect 42441 13821 42475 13855
rect 44373 13821 44407 13855
rect 46397 13821 46431 13855
rect 47593 13821 47627 13855
rect 54585 13821 54619 13855
rect 57069 13821 57103 13855
rect 57529 13821 57563 13855
rect 57897 13821 57931 13855
rect 12909 13753 12943 13787
rect 24133 13753 24167 13787
rect 30941 13753 30975 13787
rect 41061 13753 41095 13787
rect 43821 13753 43855 13787
rect 45753 13753 45787 13787
rect 48973 13753 49007 13787
rect 51641 13753 51675 13787
rect 3985 13685 4019 13719
rect 5457 13685 5491 13719
rect 9873 13685 9907 13719
rect 13645 13685 13679 13719
rect 15761 13685 15795 13719
rect 22477 13685 22511 13719
rect 25329 13685 25363 13719
rect 25421 13685 25455 13719
rect 28089 13685 28123 13719
rect 32413 13685 32447 13719
rect 36645 13685 36679 13719
rect 40233 13685 40267 13719
rect 44097 13685 44131 13719
rect 45845 13685 45879 13719
rect 56517 13685 56551 13719
rect 5917 13481 5951 13515
rect 6285 13481 6319 13515
rect 12633 13481 12667 13515
rect 13645 13481 13679 13515
rect 17969 13481 18003 13515
rect 22937 13481 22971 13515
rect 23673 13481 23707 13515
rect 25789 13481 25823 13515
rect 26065 13481 26099 13515
rect 38117 13481 38151 13515
rect 39681 13481 39715 13515
rect 42073 13481 42107 13515
rect 45937 13481 45971 13515
rect 46305 13481 46339 13515
rect 48789 13481 48823 13515
rect 49157 13481 49191 13515
rect 51549 13481 51583 13515
rect 57161 13481 57195 13515
rect 3617 13413 3651 13447
rect 22201 13413 22235 13447
rect 36645 13413 36679 13447
rect 2237 13345 2271 13379
rect 3801 13345 3835 13379
rect 5365 13345 5399 13379
rect 8953 13345 8987 13379
rect 11161 13345 11195 13379
rect 13093 13345 13127 13379
rect 13277 13345 13311 13379
rect 14105 13345 14139 13379
rect 18429 13345 18463 13379
rect 18613 13345 18647 13379
rect 19257 13345 19291 13379
rect 19901 13345 19935 13379
rect 20294 13345 20328 13379
rect 20453 13345 20487 13379
rect 22385 13345 22419 13379
rect 23121 13345 23155 13379
rect 25237 13345 25271 13379
rect 29561 13345 29595 13379
rect 30205 13345 30239 13379
rect 32045 13345 32079 13379
rect 34897 13345 34931 13379
rect 35357 13345 35391 13379
rect 35633 13345 35667 13379
rect 35771 13345 35805 13379
rect 35907 13345 35941 13379
rect 37197 13345 37231 13379
rect 37473 13345 37507 13379
rect 38301 13345 38335 13379
rect 40417 13345 40451 13379
rect 40693 13345 40727 13379
rect 45385 13345 45419 13379
rect 48237 13345 48271 13379
rect 56517 13345 56551 13379
rect 10425 13277 10459 13311
rect 14372 13277 14406 13311
rect 16497 13277 16531 13311
rect 18337 13277 18371 13311
rect 19441 13277 19475 13311
rect 20177 13277 20211 13311
rect 27445 13277 27479 13311
rect 27712 13277 27746 13311
rect 29745 13277 29779 13311
rect 30481 13277 30515 13311
rect 30598 13277 30632 13311
rect 30757 13277 30791 13311
rect 32505 13277 32539 13311
rect 34161 13277 34195 13311
rect 34713 13277 34747 13311
rect 37105 13277 37139 13311
rect 38568 13277 38602 13311
rect 42165 13277 42199 13311
rect 2504 13209 2538 13243
rect 9220 13209 9254 13243
rect 11428 13209 11462 13243
rect 13001 13209 13035 13243
rect 16764 13209 16798 13243
rect 31401 13209 31435 13243
rect 32772 13209 32806 13243
rect 40960 13209 40994 13243
rect 43913 13209 43947 13243
rect 4445 13141 4479 13175
rect 10333 13141 10367 13175
rect 11069 13141 11103 13175
rect 12541 13141 12575 13175
rect 15485 13141 15519 13175
rect 17877 13141 17911 13175
rect 18981 13141 19015 13175
rect 21097 13141 21131 13175
rect 23949 13141 23983 13175
rect 24593 13141 24627 13175
rect 27261 13141 27295 13175
rect 28825 13141 28859 13175
rect 31493 13141 31527 13175
rect 31861 13141 31895 13175
rect 31953 13141 31987 13175
rect 33885 13141 33919 13175
rect 36553 13141 36587 13175
rect 37013 13141 37047 13175
rect 39865 13141 39899 13175
rect 40233 13141 40267 13175
rect 40325 13141 40359 13175
rect 44189 13141 44223 13175
rect 47409 13141 47443 13175
rect 56333 13141 56367 13175
rect 2145 12937 2179 12971
rect 3341 12937 3375 12971
rect 8769 12937 8803 12971
rect 9229 12937 9263 12971
rect 9597 12937 9631 12971
rect 11345 12937 11379 12971
rect 15209 12937 15243 12971
rect 17601 12937 17635 12971
rect 21005 12937 21039 12971
rect 23305 12937 23339 12971
rect 24777 12937 24811 12971
rect 28733 12937 28767 12971
rect 33977 12937 34011 12971
rect 34437 12937 34471 12971
rect 37105 12937 37139 12971
rect 39957 12937 39991 12971
rect 42073 12937 42107 12971
rect 43085 12937 43119 12971
rect 47869 12937 47903 12971
rect 53297 12937 53331 12971
rect 55689 12937 55723 12971
rect 56977 12937 57011 12971
rect 2513 12869 2547 12903
rect 3709 12869 3743 12903
rect 7849 12869 7883 12903
rect 10333 12869 10367 12903
rect 17049 12869 17083 12903
rect 19892 12869 19926 12903
rect 27528 12869 27562 12903
rect 33609 12869 33643 12903
rect 34345 12869 34379 12903
rect 35081 12869 35115 12903
rect 40785 12869 40819 12903
rect 41337 12869 41371 12903
rect 2329 12801 2363 12835
rect 2605 12801 2639 12835
rect 3433 12801 3467 12835
rect 3617 12801 3651 12835
rect 3801 12801 3835 12835
rect 12081 12801 12115 12835
rect 13737 12801 13771 12835
rect 14013 12801 14047 12835
rect 15117 12801 15151 12835
rect 16221 12801 16255 12835
rect 17509 12801 17543 12835
rect 18613 12801 18647 12835
rect 19165 12801 19199 12835
rect 24869 12801 24903 12835
rect 29101 12801 29135 12835
rect 29193 12801 29227 12835
rect 30205 12801 30239 12835
rect 32137 12801 32171 12835
rect 33517 12801 33551 12835
rect 35725 12801 35759 12835
rect 36553 12801 36587 12835
rect 39405 12801 39439 12835
rect 40233 12801 40267 12835
rect 41521 12801 41555 12835
rect 42441 12801 42475 12835
rect 47409 12801 47443 12835
rect 53205 12801 53239 12835
rect 57069 12801 57103 12835
rect 58541 12801 58575 12835
rect 2789 12733 2823 12767
rect 7021 12733 7055 12767
rect 9689 12733 9723 12767
rect 9873 12733 9907 12767
rect 12173 12733 12207 12767
rect 12265 12733 12299 12767
rect 12817 12733 12851 12767
rect 13001 12733 13035 12767
rect 13854 12733 13888 12767
rect 15301 12733 15335 12767
rect 15577 12733 15611 12767
rect 17693 12733 17727 12767
rect 17969 12733 18003 12767
rect 19533 12733 19567 12767
rect 19625 12733 19659 12767
rect 22385 12733 22419 12767
rect 24961 12733 24995 12767
rect 25329 12733 25363 12767
rect 27261 12733 27295 12767
rect 29285 12733 29319 12767
rect 33793 12733 33827 12767
rect 34621 12733 34655 12767
rect 48237 12733 48271 12767
rect 50997 12733 51031 12767
rect 51733 12733 51767 12767
rect 53481 12733 53515 12767
rect 55965 12733 55999 12767
rect 57161 12733 57195 12767
rect 57897 12733 57931 12767
rect 3985 12665 4019 12699
rect 13461 12665 13495 12699
rect 28641 12665 28675 12699
rect 35357 12665 35391 12699
rect 36369 12665 36403 12699
rect 56609 12665 56643 12699
rect 7573 12597 7607 12631
rect 8309 12597 8343 12631
rect 11713 12597 11747 12631
rect 14657 12597 14691 12631
rect 14749 12597 14783 12631
rect 17141 12597 17175 12631
rect 22937 12597 22971 12631
rect 24225 12597 24259 12631
rect 24409 12597 24443 12631
rect 25973 12597 26007 12631
rect 26709 12597 26743 12631
rect 31493 12597 31527 12631
rect 32781 12597 32815 12631
rect 33149 12597 33183 12631
rect 39129 12597 39163 12631
rect 48881 12597 48915 12631
rect 51549 12597 51583 12631
rect 52377 12597 52411 12631
rect 54125 12597 54159 12631
rect 56517 12597 56551 12631
rect 7021 12393 7055 12427
rect 12265 12393 12299 12427
rect 13001 12393 13035 12427
rect 15485 12393 15519 12427
rect 17601 12393 17635 12427
rect 22201 12393 22235 12427
rect 22385 12393 22419 12427
rect 24225 12393 24259 12427
rect 29377 12393 29411 12427
rect 31401 12393 31435 12427
rect 32137 12393 32171 12427
rect 33609 12393 33643 12427
rect 34437 12393 34471 12427
rect 40141 12393 40175 12427
rect 40509 12393 40543 12427
rect 51825 12393 51859 12427
rect 52193 12393 52227 12427
rect 58449 12393 58483 12427
rect 16773 12325 16807 12359
rect 25053 12325 25087 12359
rect 28549 12325 28583 12359
rect 41705 12325 41739 12359
rect 48421 12325 48455 12359
rect 7665 12257 7699 12291
rect 9505 12257 9539 12291
rect 11713 12257 11747 12291
rect 12357 12257 12391 12291
rect 17049 12257 17083 12291
rect 22937 12257 22971 12291
rect 25513 12257 25547 12291
rect 25605 12257 25639 12291
rect 26157 12257 26191 12291
rect 28825 12257 28859 12291
rect 31493 12257 31527 12291
rect 33057 12257 33091 12291
rect 33885 12257 33919 12291
rect 42717 12257 42751 12291
rect 48145 12257 48179 12291
rect 49065 12257 49099 12291
rect 49249 12257 49283 12291
rect 3065 12189 3099 12223
rect 3433 12189 3467 12223
rect 3801 12189 3835 12223
rect 5549 12189 5583 12223
rect 7389 12189 7423 12223
rect 7941 12189 7975 12223
rect 9321 12189 9355 12223
rect 14105 12189 14139 12223
rect 19901 12189 19935 12223
rect 22753 12189 22787 12223
rect 23305 12189 23339 12223
rect 30021 12189 30055 12223
rect 34713 12189 34747 12223
rect 36001 12189 36035 12223
rect 37013 12189 37047 12223
rect 42533 12189 42567 12223
rect 45293 12189 45327 12223
rect 46029 12189 46063 12223
rect 46857 12189 46891 12223
rect 47961 12189 47995 12223
rect 48789 12189 48823 12223
rect 50445 12189 50479 12223
rect 52285 12189 52319 12223
rect 53757 12189 53791 12223
rect 54493 12189 54527 12223
rect 55321 12189 55355 12223
rect 56425 12189 56459 12223
rect 56692 12189 56726 12223
rect 3249 12121 3283 12155
rect 3341 12121 3375 12155
rect 4068 12121 4102 12155
rect 6929 12121 6963 12155
rect 14372 12121 14406 12155
rect 18061 12121 18095 12155
rect 20361 12121 20395 12155
rect 30288 12121 30322 12155
rect 50712 12121 50746 12155
rect 52552 12121 52586 12155
rect 58357 12121 58391 12155
rect 3617 12053 3651 12087
rect 5181 12053 5215 12087
rect 7481 12053 7515 12087
rect 8493 12053 8527 12087
rect 8953 12053 8987 12087
rect 9413 12053 9447 12087
rect 13277 12053 13311 12087
rect 13921 12053 13955 12087
rect 15853 12053 15887 12087
rect 21833 12053 21867 12087
rect 22845 12053 22879 12087
rect 23857 12053 23891 12087
rect 24869 12053 24903 12087
rect 25421 12053 25455 12087
rect 26801 12053 26835 12087
rect 35357 12053 35391 12087
rect 36645 12053 36679 12087
rect 39037 12053 39071 12087
rect 42073 12053 42107 12087
rect 42165 12053 42199 12087
rect 42625 12053 42659 12087
rect 45937 12053 45971 12087
rect 46673 12053 46707 12087
rect 47409 12053 47443 12087
rect 47593 12053 47627 12087
rect 48053 12053 48087 12087
rect 48881 12053 48915 12087
rect 49893 12053 49927 12087
rect 53665 12053 53699 12087
rect 54401 12053 54435 12087
rect 55137 12053 55171 12087
rect 55965 12053 55999 12087
rect 56333 12053 56367 12087
rect 57805 12053 57839 12087
rect 2697 11849 2731 11883
rect 3433 11849 3467 11883
rect 4261 11849 4295 11883
rect 4997 11849 5031 11883
rect 6193 11849 6227 11883
rect 10425 11849 10459 11883
rect 12541 11849 12575 11883
rect 15209 11849 15243 11883
rect 17601 11849 17635 11883
rect 19349 11849 19383 11883
rect 21189 11849 21223 11883
rect 23213 11849 23247 11883
rect 30021 11849 30055 11883
rect 30389 11849 30423 11883
rect 30481 11849 30515 11883
rect 31493 11849 31527 11883
rect 34345 11849 34379 11883
rect 36001 11849 36035 11883
rect 42441 11849 42475 11883
rect 42809 11849 42843 11883
rect 43913 11849 43947 11883
rect 45017 11849 45051 11883
rect 45201 11849 45235 11883
rect 45661 11849 45695 11883
rect 46397 11849 46431 11883
rect 47133 11849 47167 11883
rect 49341 11849 49375 11883
rect 50629 11849 50663 11883
rect 51089 11849 51123 11883
rect 51549 11849 51583 11883
rect 52745 11849 52779 11883
rect 53113 11849 53147 11883
rect 55321 11849 55355 11883
rect 6736 11781 6770 11815
rect 9873 11781 9907 11815
rect 15577 11781 15611 11815
rect 18061 11781 18095 11815
rect 20269 11781 20303 11815
rect 22100 11781 22134 11815
rect 25145 11781 25179 11815
rect 25504 11781 25538 11815
rect 33425 11781 33459 11815
rect 35725 11781 35759 11815
rect 39681 11781 39715 11815
rect 45569 11781 45603 11815
rect 47860 11781 47894 11815
rect 54208 11781 54242 11815
rect 2881 11713 2915 11747
rect 3065 11713 3099 11747
rect 3157 11713 3191 11747
rect 3249 11713 3283 11747
rect 3433 11713 3467 11747
rect 4353 11713 4387 11747
rect 6469 11713 6503 11747
rect 8217 11713 8251 11747
rect 14657 11713 14691 11747
rect 21833 11713 21867 11747
rect 24501 11713 24535 11747
rect 25237 11713 25271 11747
rect 29837 11713 29871 11747
rect 33517 11713 33551 11747
rect 34253 11713 34287 11747
rect 35357 11713 35391 11747
rect 36369 11713 36403 11747
rect 36461 11713 36495 11747
rect 37933 11713 37967 11747
rect 39589 11713 39623 11747
rect 44005 11713 44039 11747
rect 46489 11713 46523 11747
rect 51457 11713 51491 11747
rect 53205 11713 53239 11747
rect 53757 11713 53791 11747
rect 53941 11713 53975 11747
rect 55965 11713 55999 11747
rect 56701 11713 56735 11747
rect 56818 11713 56852 11747
rect 3709 11645 3743 11679
rect 8033 11645 8067 11679
rect 8953 11645 8987 11679
rect 9091 11645 9125 11679
rect 9229 11645 9263 11679
rect 16681 11645 16715 11679
rect 20361 11645 20395 11679
rect 20453 11645 20487 11679
rect 23305 11645 23339 11679
rect 23489 11645 23523 11679
rect 24225 11645 24259 11679
rect 24342 11645 24376 11679
rect 28365 11645 28399 11679
rect 30573 11645 30607 11679
rect 32413 11645 32447 11679
rect 33701 11645 33735 11679
rect 34437 11645 34471 11679
rect 34713 11645 34747 11679
rect 36645 11645 36679 11679
rect 37289 11645 37323 11679
rect 38577 11645 38611 11679
rect 39773 11645 39807 11679
rect 40049 11645 40083 11679
rect 40785 11645 40819 11679
rect 42901 11645 42935 11679
rect 42993 11645 43027 11679
rect 43361 11645 43395 11679
rect 45753 11645 45787 11679
rect 46673 11645 46707 11679
rect 47593 11645 47627 11679
rect 51733 11645 51767 11679
rect 52009 11645 52043 11679
rect 53389 11645 53423 11679
rect 55781 11645 55815 11679
rect 56977 11645 57011 11679
rect 7849 11577 7883 11611
rect 8677 11577 8711 11611
rect 21557 11577 21591 11611
rect 23949 11577 23983 11611
rect 26617 11577 26651 11611
rect 33057 11577 33091 11611
rect 39221 11577 39255 11611
rect 41429 11577 41463 11611
rect 56425 11577 56459 11611
rect 17325 11509 17359 11543
rect 19901 11509 19935 11543
rect 28917 11509 28951 11543
rect 29285 11509 29319 11543
rect 32965 11509 32999 11543
rect 33885 11509 33919 11543
rect 37013 11509 37047 11543
rect 39129 11509 39163 11543
rect 40693 11509 40727 11543
rect 42257 11509 42291 11543
rect 44649 11509 44683 11543
rect 46029 11509 46063 11543
rect 48973 11509 49007 11543
rect 50905 11509 50939 11543
rect 52561 11509 52595 11543
rect 55597 11509 55631 11543
rect 57621 11509 57655 11543
rect 2881 11305 2915 11339
rect 3065 11305 3099 11339
rect 3985 11305 4019 11339
rect 4537 11305 4571 11339
rect 7665 11305 7699 11339
rect 10333 11305 10367 11339
rect 11989 11305 12023 11339
rect 19073 11305 19107 11339
rect 21649 11305 21683 11339
rect 23121 11305 23155 11339
rect 25789 11305 25823 11339
rect 29745 11305 29779 11339
rect 33793 11305 33827 11339
rect 39681 11305 39715 11339
rect 39865 11305 39899 11339
rect 42809 11305 42843 11339
rect 54401 11305 54435 11339
rect 20729 11237 20763 11271
rect 36645 11237 36679 11271
rect 41613 11237 41647 11271
rect 44281 11237 44315 11271
rect 46397 11237 46431 11271
rect 48421 11237 48455 11271
rect 48513 11237 48547 11271
rect 51549 11237 51583 11271
rect 55321 11237 55355 11271
rect 56885 11237 56919 11271
rect 3249 11169 3283 11203
rect 4077 11169 4111 11203
rect 4813 11169 4847 11203
rect 8401 11169 8435 11203
rect 8953 11169 8987 11203
rect 10425 11169 10459 11203
rect 14933 11169 14967 11203
rect 19349 11169 19383 11203
rect 21741 11169 21775 11203
rect 23765 11169 23799 11203
rect 25881 11169 25915 11203
rect 33885 11169 33919 11203
rect 34897 11169 34931 11203
rect 35357 11169 35391 11203
rect 35750 11169 35784 11203
rect 35909 11169 35943 11203
rect 37105 11169 37139 11203
rect 37197 11169 37231 11203
rect 38301 11169 38335 11203
rect 40325 11169 40359 11203
rect 40417 11169 40451 11203
rect 40969 11169 41003 11203
rect 41889 11169 41923 11203
rect 42901 11169 42935 11203
rect 46581 11169 46615 11203
rect 47225 11169 47259 11203
rect 47618 11169 47652 11203
rect 47777 11169 47811 11203
rect 49065 11169 49099 11203
rect 49341 11169 49375 11203
rect 50169 11169 50203 11203
rect 51641 11169 51675 11203
rect 51825 11169 51859 11203
rect 52285 11169 52319 11203
rect 52561 11169 52595 11203
rect 52837 11169 52871 11203
rect 54953 11169 54987 11203
rect 55873 11169 55907 11203
rect 56149 11169 56183 11203
rect 57437 11169 57471 11203
rect 57897 11169 57931 11203
rect 2789 11101 2823 11135
rect 2973 11101 3007 11135
rect 3341 11101 3375 11135
rect 3433 11101 3467 11135
rect 3525 11101 3559 11135
rect 3985 11101 4019 11135
rect 4445 11101 4479 11135
rect 4537 11101 4571 11135
rect 6285 11101 6319 11135
rect 11437 11101 11471 11135
rect 14197 11101 14231 11135
rect 15945 11101 15979 11135
rect 16212 11101 16246 11135
rect 17509 11101 17543 11135
rect 24409 11101 24443 11135
rect 27813 11101 27847 11135
rect 28549 11101 28583 11135
rect 32413 11101 32447 11135
rect 32680 11101 32714 11135
rect 34713 11101 34747 11135
rect 35633 11101 35667 11135
rect 37473 11101 37507 11135
rect 38568 11101 38602 11135
rect 41153 11101 41187 11135
rect 42006 11101 42040 11135
rect 42165 11101 42199 11135
rect 45017 11101 45051 11135
rect 45284 11101 45318 11135
rect 46765 11101 46799 11135
rect 47501 11101 47535 11135
rect 49985 11101 50019 11135
rect 50436 11101 50470 11135
rect 52678 11101 52712 11135
rect 54217 11101 54251 11135
rect 54769 11101 54803 11135
rect 57253 11101 57287 11135
rect 6552 11033 6586 11067
rect 8125 11033 8159 11067
rect 9220 11033 9254 11067
rect 12449 11033 12483 11067
rect 19616 11033 19650 11067
rect 22008 11033 22042 11067
rect 23673 11033 23707 11067
rect 24676 11033 24710 11067
rect 29101 11033 29135 11067
rect 34529 11033 34563 11067
rect 36553 11033 36587 11067
rect 37013 11033 37047 11067
rect 40233 11033 40267 11067
rect 43168 11033 43202 11067
rect 48973 11033 49007 11067
rect 53481 11033 53515 11067
rect 54861 11033 54895 11067
rect 55689 11033 55723 11067
rect 57345 11033 57379 11067
rect 4353 10965 4387 10999
rect 4629 10965 4663 10999
rect 7757 10965 7791 10999
rect 8217 10965 8251 10999
rect 11069 10965 11103 10999
rect 14841 10965 14875 10999
rect 15577 10965 15611 10999
rect 17325 10965 17359 10999
rect 18061 10965 18095 10999
rect 18429 10965 18463 10999
rect 23213 10965 23247 10999
rect 23581 10965 23615 10999
rect 26525 10965 26559 10999
rect 28365 10965 28399 10999
rect 30205 10965 30239 10999
rect 38117 10965 38151 10999
rect 44741 10965 44775 10999
rect 48881 10965 48915 10999
rect 55781 10965 55815 10999
rect 56793 10965 56827 10999
rect 3617 10761 3651 10795
rect 4537 10761 4571 10795
rect 6929 10761 6963 10795
rect 7849 10761 7883 10795
rect 8585 10761 8619 10795
rect 9505 10761 9539 10795
rect 11989 10761 12023 10795
rect 13829 10761 13863 10795
rect 14197 10761 14231 10795
rect 15761 10761 15795 10795
rect 16681 10761 16715 10795
rect 17141 10761 17175 10795
rect 19717 10761 19751 10795
rect 21097 10761 21131 10795
rect 31585 10761 31619 10795
rect 33885 10761 33919 10795
rect 34713 10761 34747 10795
rect 37013 10761 37047 10795
rect 37289 10761 37323 10795
rect 38853 10761 38887 10795
rect 41061 10761 41095 10795
rect 41521 10761 41555 10795
rect 43821 10761 43855 10795
rect 44557 10761 44591 10795
rect 47041 10761 47075 10795
rect 48973 10761 49007 10795
rect 49709 10761 49743 10795
rect 51733 10761 51767 10795
rect 55689 10761 55723 10795
rect 57713 10761 57747 10795
rect 8861 10693 8895 10727
rect 10517 10693 10551 10727
rect 16221 10693 16255 10727
rect 19809 10693 19843 10727
rect 39037 10693 39071 10727
rect 52101 10693 52135 10727
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 3433 10625 3467 10659
rect 4445 10625 4479 10659
rect 4721 10625 4755 10659
rect 4905 10625 4939 10659
rect 5181 10625 5215 10659
rect 5335 10625 5369 10659
rect 5641 10625 5675 10659
rect 5795 10625 5829 10659
rect 7297 10625 7331 10659
rect 8033 10625 8067 10659
rect 9413 10625 9447 10659
rect 11897 10625 11931 10659
rect 13001 10625 13035 10659
rect 13737 10625 13771 10659
rect 16129 10625 16163 10659
rect 17049 10625 17083 10659
rect 17877 10625 17911 10659
rect 18797 10625 18831 10659
rect 22753 10625 22787 10659
rect 23305 10625 23339 10659
rect 23397 10625 23431 10659
rect 24041 10625 24075 10659
rect 24409 10625 24443 10659
rect 25145 10625 25179 10659
rect 27261 10625 27295 10659
rect 27528 10625 27562 10659
rect 29101 10625 29135 10659
rect 29193 10625 29227 10659
rect 30205 10625 30239 10659
rect 30297 10625 30331 10659
rect 31033 10625 31067 10659
rect 32772 10625 32806 10659
rect 34621 10625 34655 10659
rect 35900 10625 35934 10659
rect 37657 10625 37691 10659
rect 42441 10625 42475 10659
rect 42708 10625 42742 10659
rect 45100 10625 45134 10659
rect 47860 10625 47894 10659
rect 49065 10625 49099 10659
rect 50528 10625 50562 10659
rect 52193 10625 52227 10659
rect 53389 10625 53423 10659
rect 54309 10625 54343 10659
rect 54576 10625 54610 10659
rect 56333 10625 56367 10659
rect 56600 10625 56634 10659
rect 58541 10625 58575 10659
rect 3157 10557 3191 10591
rect 3249 10557 3283 10591
rect 6009 10557 6043 10591
rect 9597 10557 9631 10591
rect 9873 10557 9907 10591
rect 10793 10557 10827 10591
rect 12173 10557 12207 10591
rect 12357 10557 12391 10591
rect 14289 10557 14323 10591
rect 14473 10557 14507 10591
rect 15117 10557 15151 10591
rect 16313 10557 16347 10591
rect 17233 10557 17267 10591
rect 18061 10557 18095 10591
rect 18914 10557 18948 10591
rect 19073 10557 19107 10591
rect 25237 10557 25271 10591
rect 25329 10557 25363 10591
rect 25605 10557 25639 10591
rect 26249 10557 26283 10591
rect 29285 10557 29319 10591
rect 29653 10557 29687 10591
rect 32505 10557 32539 10591
rect 35633 10557 35667 10591
rect 37749 10557 37783 10591
rect 37933 10557 37967 10591
rect 43913 10557 43947 10591
rect 44833 10557 44867 10591
rect 46489 10557 46523 10591
rect 47593 10557 47627 10591
rect 50169 10557 50203 10591
rect 50261 10557 50295 10591
rect 52285 10557 52319 10591
rect 52745 10557 52779 10591
rect 57897 10557 57931 10591
rect 9045 10489 9079 10523
rect 11529 10489 11563 10523
rect 18521 10489 18555 10523
rect 24777 10489 24811 10523
rect 28641 10489 28675 10523
rect 35449 10489 35483 10523
rect 46213 10489 46247 10523
rect 47409 10489 47443 10523
rect 51641 10489 51675 10523
rect 4813 10421 4847 10455
rect 5365 10421 5399 10455
rect 6561 10421 6595 10455
rect 11345 10421 11379 10455
rect 14933 10421 14967 10455
rect 15669 10421 15703 10455
rect 17693 10421 17727 10455
rect 26801 10421 26835 10455
rect 28733 10421 28767 10455
rect 34253 10421 34287 10455
rect 35081 10421 35115 10455
rect 38301 10421 38335 10455
rect 40325 10421 40359 10455
rect 55965 10421 55999 10455
rect 2789 10217 2823 10251
rect 4169 10217 4203 10251
rect 5733 10217 5767 10251
rect 9965 10217 9999 10251
rect 15485 10217 15519 10251
rect 17049 10217 17083 10251
rect 18521 10217 18555 10251
rect 21281 10217 21315 10251
rect 28825 10217 28859 10251
rect 34989 10217 35023 10251
rect 37289 10217 37323 10251
rect 38025 10217 38059 10251
rect 40509 10217 40543 10251
rect 41061 10217 41095 10251
rect 42257 10217 42291 10251
rect 44097 10217 44131 10251
rect 44741 10217 44775 10251
rect 46489 10217 46523 10251
rect 49525 10217 49559 10251
rect 56425 10217 56459 10251
rect 56885 10217 56919 10251
rect 11897 10149 11931 10183
rect 19809 10149 19843 10183
rect 30205 10149 30239 10183
rect 39681 10149 39715 10183
rect 2973 10081 3007 10115
rect 9597 10081 9631 10115
rect 10517 10081 10551 10115
rect 12265 10081 12299 10115
rect 12725 10081 12759 10115
rect 13001 10081 13035 10115
rect 13139 10081 13173 10115
rect 19717 10081 19751 10115
rect 20361 10081 20395 10115
rect 20637 10081 20671 10115
rect 30481 10081 30515 10115
rect 30598 10081 30632 10115
rect 30757 10081 30791 10115
rect 32045 10081 32079 10115
rect 37381 10081 37415 10115
rect 38301 10081 38335 10115
rect 39957 10081 39991 10115
rect 42165 10081 42199 10115
rect 42809 10081 42843 10115
rect 43177 10081 43211 10115
rect 51457 10081 51491 10115
rect 51549 10081 51583 10115
rect 51917 10081 51951 10115
rect 55873 10081 55907 10115
rect 57437 10081 57471 10115
rect 57713 10081 57747 10115
rect 3065 10013 3099 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 6561 10013 6595 10047
rect 7481 10013 7515 10047
rect 8033 10013 8067 10047
rect 8769 10013 8803 10047
rect 9045 10013 9079 10047
rect 12081 10013 12115 10047
rect 13277 10013 13311 10047
rect 14105 10013 14139 10047
rect 15669 10013 15703 10047
rect 15936 10013 15970 10047
rect 17141 10013 17175 10047
rect 18797 10013 18831 10047
rect 21557 10013 21591 10047
rect 27445 10013 27479 10047
rect 27712 10013 27746 10047
rect 29561 10013 29595 10047
rect 29745 10013 29779 10047
rect 32689 10013 32723 10047
rect 33425 10013 33459 10047
rect 35909 10013 35943 10047
rect 38568 10013 38602 10047
rect 49433 10013 49467 10047
rect 2789 9945 2823 9979
rect 3157 9945 3191 9979
rect 6837 9945 6871 9979
rect 10784 9945 10818 9979
rect 14372 9945 14406 9979
rect 17408 9945 17442 9979
rect 20269 9945 20303 9979
rect 24593 9945 24627 9979
rect 31401 9945 31435 9979
rect 31953 9945 31987 9979
rect 36176 9945 36210 9979
rect 42625 9945 42659 9979
rect 43729 9945 43763 9979
rect 51365 9945 51399 9979
rect 52469 9945 52503 9979
rect 57253 9945 57287 9979
rect 58357 9945 58391 9979
rect 10333 9877 10367 9911
rect 13921 9877 13955 9911
rect 20177 9877 20211 9911
rect 22201 9877 22235 9911
rect 23121 9877 23155 9911
rect 27353 9877 27387 9911
rect 29377 9877 29411 9911
rect 31493 9877 31527 9911
rect 31861 9877 31895 9911
rect 33241 9877 33275 9911
rect 33977 9877 34011 9911
rect 34437 9877 34471 9911
rect 35541 9877 35575 9911
rect 42717 9877 42751 9911
rect 48421 9877 48455 9911
rect 50905 9877 50939 9911
rect 50997 9877 51031 9911
rect 56793 9877 56827 9911
rect 57345 9877 57379 9911
rect 3341 9673 3375 9707
rect 7665 9673 7699 9707
rect 13829 9673 13863 9707
rect 14289 9673 14323 9707
rect 17693 9673 17727 9707
rect 20453 9673 20487 9707
rect 28273 9673 28307 9707
rect 30021 9673 30055 9707
rect 31493 9673 31527 9707
rect 32413 9673 32447 9707
rect 32689 9673 32723 9707
rect 51825 9673 51859 9707
rect 54033 9673 54067 9707
rect 6193 9605 6227 9639
rect 9781 9605 9815 9639
rect 10232 9605 10266 9639
rect 14933 9605 14967 9639
rect 15945 9605 15979 9639
rect 33057 9605 33091 9639
rect 35265 9605 35299 9639
rect 39957 9605 39991 9639
rect 40325 9605 40359 9639
rect 43821 9605 43855 9639
rect 44925 9605 44959 9639
rect 46949 9605 46983 9639
rect 51457 9605 51491 9639
rect 52561 9605 52595 9639
rect 52745 9605 52779 9639
rect 58449 9605 58483 9639
rect 2881 9537 2915 9571
rect 3065 9537 3099 9571
rect 3157 9537 3191 9571
rect 3249 9537 3283 9571
rect 5917 9537 5951 9571
rect 6469 9537 6503 9571
rect 7205 9537 7239 9571
rect 7481 9537 7515 9571
rect 7757 9537 7791 9571
rect 9965 9537 9999 9571
rect 11897 9537 11931 9571
rect 11989 9537 12023 9571
rect 12449 9537 12483 9571
rect 12716 9537 12750 9571
rect 14381 9537 14415 9571
rect 15485 9537 15519 9571
rect 17325 9537 17359 9571
rect 18153 9537 18187 9571
rect 18245 9537 18279 9571
rect 19257 9537 19291 9571
rect 19901 9537 19935 9571
rect 27445 9537 27479 9571
rect 27629 9537 27663 9571
rect 28181 9537 28215 9571
rect 28641 9537 28675 9571
rect 28908 9537 28942 9571
rect 30380 9537 30414 9571
rect 33517 9537 33551 9571
rect 34805 9537 34839 9571
rect 39773 9537 39807 9571
rect 43637 9537 43671 9571
rect 46765 9537 46799 9571
rect 50905 9537 50939 9571
rect 5825 9469 5859 9503
rect 8125 9469 8159 9503
rect 8401 9469 8435 9503
rect 12081 9469 12115 9503
rect 14565 9469 14599 9503
rect 15669 9469 15703 9503
rect 16681 9469 16715 9503
rect 18337 9469 18371 9503
rect 18613 9469 18647 9503
rect 20637 9469 20671 9503
rect 21833 9469 21867 9503
rect 24225 9469 24259 9503
rect 26249 9469 26283 9503
rect 28365 9469 28399 9503
rect 30113 9469 30147 9503
rect 33149 9469 33183 9503
rect 33241 9469 33275 9503
rect 34345 9469 34379 9503
rect 36001 9469 36035 9503
rect 40417 9469 40451 9503
rect 41153 9469 41187 9503
rect 42441 9469 42475 9503
rect 44097 9469 44131 9503
rect 45477 9469 45511 9503
rect 48053 9469 48087 9503
rect 48789 9469 48823 9503
rect 49525 9469 49559 9503
rect 54585 9469 54619 9503
rect 56149 9469 56183 9503
rect 2881 9401 2915 9435
rect 6009 9401 6043 9435
rect 11345 9401 11379 9435
rect 35817 9401 35851 9435
rect 3801 9333 3835 9367
rect 6101 9333 6135 9367
rect 7481 9333 7515 9367
rect 11529 9333 11563 9367
rect 13921 9333 13955 9367
rect 17785 9333 17819 9367
rect 21281 9333 21315 9367
rect 22477 9333 22511 9367
rect 22845 9333 22879 9367
rect 23397 9333 23431 9367
rect 24041 9333 24075 9367
rect 24777 9333 24811 9367
rect 25145 9333 25179 9367
rect 26801 9333 26835 9367
rect 27169 9333 27203 9367
rect 27813 9333 27847 9367
rect 31769 9333 31803 9367
rect 36553 9333 36587 9367
rect 36829 9333 36863 9367
rect 37749 9333 37783 9367
rect 41061 9333 41095 9367
rect 41797 9333 41831 9367
rect 43085 9333 43119 9367
rect 44649 9333 44683 9367
rect 46121 9333 46155 9367
rect 46489 9333 46523 9367
rect 48605 9333 48639 9367
rect 49341 9333 49375 9367
rect 50077 9333 50111 9367
rect 55229 9333 55263 9367
rect 56793 9333 56827 9367
rect 57069 9333 57103 9367
rect 57437 9333 57471 9367
rect 58081 9333 58115 9367
rect 2973 9129 3007 9163
rect 3893 9129 3927 9163
rect 6837 9129 6871 9163
rect 8309 9129 8343 9163
rect 11805 9129 11839 9163
rect 12633 9129 12667 9163
rect 14749 9129 14783 9163
rect 18245 9129 18279 9163
rect 20085 9129 20119 9163
rect 24869 9129 24903 9163
rect 26709 9129 26743 9163
rect 29377 9129 29411 9163
rect 39865 9129 39899 9163
rect 48053 9129 48087 9163
rect 56057 9129 56091 9163
rect 56885 9129 56919 9163
rect 11069 9061 11103 9095
rect 13001 9061 13035 9095
rect 19809 9061 19843 9095
rect 23305 9061 23339 9095
rect 26341 9061 26375 9095
rect 29561 9061 29595 9095
rect 41153 9061 41187 9095
rect 43361 9061 43395 9095
rect 46121 9061 46155 9095
rect 2697 8993 2731 9027
rect 3433 8993 3467 9027
rect 10609 8993 10643 9027
rect 11253 8993 11287 9027
rect 12081 8993 12115 9027
rect 13553 8993 13587 9027
rect 14105 8993 14139 9027
rect 17693 8993 17727 9027
rect 20821 8993 20855 9027
rect 24041 8993 24075 9027
rect 24961 8993 24995 9027
rect 26893 8993 26927 9027
rect 30113 8993 30147 9027
rect 30941 8993 30975 9027
rect 31309 8993 31343 9027
rect 40509 8993 40543 9027
rect 41613 8993 41647 9027
rect 41797 8993 41831 9027
rect 41981 8993 42015 9027
rect 43821 8993 43855 9027
rect 44005 8993 44039 9027
rect 44189 8993 44223 9027
rect 45845 8993 45879 9027
rect 46581 8993 46615 9027
rect 46673 8993 46707 9027
rect 46949 8993 46983 9027
rect 48513 8993 48547 9027
rect 48697 8993 48731 9027
rect 54953 8993 54987 9027
rect 55965 8993 55999 9027
rect 56609 8993 56643 9027
rect 57437 8993 57471 9027
rect 57713 8993 57747 9027
rect 2605 8925 2639 8959
rect 3065 8925 3099 8959
rect 3219 8925 3253 8959
rect 3801 8925 3835 8959
rect 3985 8925 4019 8959
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 6929 8925 6963 8959
rect 7185 8925 7219 8959
rect 8953 8925 8987 8959
rect 9781 8925 9815 8959
rect 18521 8925 18555 8959
rect 21088 8925 21122 8959
rect 22385 8925 22419 8959
rect 23857 8925 23891 8959
rect 25228 8925 25262 8959
rect 28641 8925 28675 8959
rect 28825 8925 28859 8959
rect 32505 8925 32539 8959
rect 34897 8925 34931 8959
rect 35449 8925 35483 8959
rect 36553 8925 36587 8959
rect 37657 8925 37691 8959
rect 38853 8925 38887 8959
rect 41521 8925 41555 8959
rect 43269 8925 43303 8959
rect 45017 8925 45051 8959
rect 48881 8925 48915 8959
rect 50169 8925 50203 8959
rect 52837 8925 52871 8959
rect 54677 8925 54711 8959
rect 57253 8925 57287 8959
rect 5365 8857 5399 8891
rect 5457 8857 5491 8891
rect 6193 8857 6227 8891
rect 10885 8857 10919 8891
rect 13369 8857 13403 8891
rect 16221 8857 16255 8891
rect 19993 8857 20027 8891
rect 30021 8857 30055 8891
rect 30757 8857 30791 8891
rect 31861 8857 31895 8891
rect 36277 8857 36311 8891
rect 37381 8857 37415 8891
rect 40325 8857 40359 8891
rect 43729 8857 43763 8891
rect 47869 8857 47903 8891
rect 53104 8857 53138 8891
rect 54769 8857 54803 8891
rect 56517 8857 56551 8891
rect 58357 8857 58391 8891
rect 4813 8789 4847 8823
rect 5089 8789 5123 8823
rect 8677 8789 8711 8823
rect 9597 8789 9631 8823
rect 10333 8789 10367 8823
rect 13461 8789 13495 8823
rect 17417 8789 17451 8823
rect 19073 8789 19107 8823
rect 20729 8789 20763 8823
rect 22201 8789 22235 8823
rect 23029 8789 23063 8823
rect 23489 8789 23523 8823
rect 23949 8789 23983 8823
rect 27537 8789 27571 8823
rect 29929 8789 29963 8823
rect 30389 8789 30423 8823
rect 30849 8789 30883 8823
rect 33977 8789 34011 8823
rect 35265 8789 35299 8823
rect 38301 8789 38335 8823
rect 39405 8789 39439 8823
rect 40233 8789 40267 8823
rect 40969 8789 41003 8823
rect 42625 8789 42659 8823
rect 44833 8789 44867 8823
rect 46489 8789 46523 8823
rect 47593 8789 47627 8823
rect 48421 8789 48455 8823
rect 49525 8789 49559 8823
rect 50813 8789 50847 8823
rect 54217 8789 54251 8823
rect 54309 8789 54343 8823
rect 55505 8789 55539 8823
rect 56425 8789 56459 8823
rect 57345 8789 57379 8823
rect 3617 8585 3651 8619
rect 4169 8585 4203 8619
rect 4451 8585 4485 8619
rect 7665 8585 7699 8619
rect 8585 8585 8619 8619
rect 9045 8585 9079 8619
rect 13553 8585 13587 8619
rect 13921 8585 13955 8619
rect 19717 8585 19751 8619
rect 20085 8585 20119 8619
rect 20545 8585 20579 8619
rect 20913 8585 20947 8619
rect 21281 8585 21315 8619
rect 26985 8585 27019 8619
rect 27445 8585 27479 8619
rect 29193 8585 29227 8619
rect 30297 8585 30331 8619
rect 31033 8585 31067 8619
rect 36737 8585 36771 8619
rect 39221 8585 39255 8619
rect 40693 8585 40727 8619
rect 44465 8585 44499 8619
rect 47317 8585 47351 8619
rect 48973 8585 49007 8619
rect 53481 8585 53515 8619
rect 57345 8585 57379 8619
rect 57713 8585 57747 8619
rect 4721 8517 4755 8551
rect 4921 8517 4955 8551
rect 8125 8517 8159 8551
rect 11989 8517 12023 8551
rect 18245 8517 18279 8551
rect 18582 8517 18616 8551
rect 32404 8517 32438 8551
rect 42984 8517 43018 8551
rect 49608 8517 49642 8551
rect 55873 8517 55907 8551
rect 56232 8517 56266 8551
rect 2973 8449 3007 8483
rect 4353 8449 4387 8483
rect 4537 8449 4571 8483
rect 4629 8449 4663 8483
rect 5365 8449 5399 8483
rect 6745 8449 6779 8483
rect 7757 8449 7791 8483
rect 7941 8449 7975 8483
rect 8033 8449 8067 8483
rect 8217 8449 8251 8483
rect 8953 8449 8987 8483
rect 9413 8449 9447 8483
rect 11897 8449 11931 8483
rect 20453 8449 20487 8483
rect 21373 8449 21407 8483
rect 21833 8449 21867 8483
rect 22100 8449 22134 8483
rect 23305 8449 23339 8483
rect 23572 8449 23606 8483
rect 24777 8449 24811 8483
rect 25814 8449 25848 8483
rect 25973 8449 26007 8483
rect 27353 8449 27387 8483
rect 29101 8449 29135 8483
rect 29653 8449 29687 8483
rect 33609 8449 33643 8483
rect 34897 8449 34931 8483
rect 35357 8449 35391 8483
rect 35624 8449 35658 8483
rect 37565 8449 37599 8483
rect 37841 8449 37875 8483
rect 38108 8449 38142 8483
rect 39313 8449 39347 8483
rect 39580 8449 39614 8483
rect 40877 8449 40911 8483
rect 41144 8449 41178 8483
rect 44557 8449 44591 8483
rect 44824 8449 44858 8483
rect 46029 8449 46063 8483
rect 47593 8449 47627 8483
rect 47860 8449 47894 8483
rect 49341 8449 49375 8483
rect 51457 8449 51491 8483
rect 53389 8449 53423 8483
rect 55965 8449 55999 8483
rect 57897 8449 57931 8483
rect 3065 8381 3099 8415
rect 3709 8381 3743 8415
rect 6009 8381 6043 8415
rect 7297 8381 7331 8415
rect 9137 8381 9171 8415
rect 9781 8381 9815 8415
rect 10793 8381 10827 8415
rect 12173 8381 12207 8415
rect 13001 8381 13035 8415
rect 15853 8381 15887 8415
rect 16773 8381 16807 8415
rect 17693 8381 17727 8415
rect 18337 8381 18371 8415
rect 20729 8381 20763 8415
rect 21465 8381 21499 8415
rect 24961 8381 24995 8415
rect 25697 8381 25731 8415
rect 27537 8381 27571 8415
rect 27997 8381 28031 8415
rect 30389 8381 30423 8415
rect 32137 8381 32171 8415
rect 34437 8381 34471 8415
rect 42717 8381 42751 8415
rect 46857 8381 46891 8415
rect 50813 8381 50847 8415
rect 51549 8381 51583 8415
rect 53573 8381 53607 8415
rect 54033 8381 54067 8415
rect 54217 8381 54251 8415
rect 54953 8381 54987 8415
rect 55070 8381 55104 8415
rect 55229 8381 55263 8415
rect 3985 8313 4019 8347
rect 5089 8313 5123 8347
rect 7481 8313 7515 8347
rect 11529 8313 11563 8347
rect 12817 8313 12851 8347
rect 23213 8313 23247 8347
rect 24685 8313 24719 8347
rect 25421 8313 25455 8347
rect 26617 8313 26651 8347
rect 42257 8313 42291 8347
rect 44097 8313 44131 8347
rect 45937 8313 45971 8347
rect 54677 8313 54711 8347
rect 58541 8313 58575 8347
rect 4905 8245 4939 8279
rect 11345 8245 11379 8279
rect 15485 8245 15519 8279
rect 16497 8245 16531 8279
rect 17417 8245 17451 8279
rect 33517 8245 33551 8279
rect 37013 8245 37047 8279
rect 50721 8245 50755 8279
rect 52193 8245 52227 8279
rect 52469 8245 52503 8279
rect 53021 8245 53055 8279
rect 3157 8041 3191 8075
rect 4353 8041 4387 8075
rect 7297 8041 7331 8075
rect 7941 8041 7975 8075
rect 8217 8041 8251 8075
rect 8677 8041 8711 8075
rect 10333 8041 10367 8075
rect 13001 8041 13035 8075
rect 18337 8041 18371 8075
rect 24225 8041 24259 8075
rect 27537 8041 27571 8075
rect 29745 8041 29779 8075
rect 39405 8041 39439 8075
rect 43821 8041 43855 8075
rect 47225 8041 47259 8075
rect 48881 8041 48915 8075
rect 49249 8041 49283 8075
rect 51549 8041 51583 8075
rect 53849 8041 53883 8075
rect 55505 8041 55539 8075
rect 55965 8041 55999 8075
rect 58541 8041 58575 8075
rect 15577 7973 15611 8007
rect 16405 7973 16439 8007
rect 33793 7973 33827 8007
rect 45661 7973 45695 8007
rect 57805 7973 57839 8007
rect 2881 7905 2915 7939
rect 4997 7905 5031 7939
rect 12357 7905 12391 7939
rect 14933 7905 14967 7939
rect 16037 7905 16071 7939
rect 16129 7905 16163 7939
rect 17049 7905 17083 7939
rect 17509 7905 17543 7939
rect 18797 7905 18831 7939
rect 18981 7905 19015 7939
rect 19901 7905 19935 7939
rect 20269 7905 20303 7939
rect 20913 7905 20947 7939
rect 21306 7905 21340 7939
rect 24961 7905 24995 7939
rect 25881 7905 25915 7939
rect 34897 7905 34931 7939
rect 35357 7905 35391 7939
rect 35633 7905 35667 7939
rect 35750 7905 35784 7939
rect 35909 7905 35943 7939
rect 37197 7905 37231 7939
rect 37749 7905 37783 7939
rect 40049 7905 40083 7939
rect 40509 7905 40543 7939
rect 40785 7905 40819 7939
rect 42257 7905 42291 7939
rect 42441 7905 42475 7939
rect 44557 7905 44591 7939
rect 45017 7905 45051 7939
rect 45201 7905 45235 7939
rect 46054 7905 46088 7939
rect 46213 7905 46247 7939
rect 49709 7905 49743 7939
rect 49801 7905 49835 7939
rect 54585 7905 54619 7939
rect 56425 7905 56459 7939
rect 57897 7905 57931 7939
rect 2973 7837 3007 7871
rect 3066 7837 3100 7871
rect 5181 7837 5215 7871
rect 5917 7837 5951 7871
rect 8953 7837 8987 7871
rect 11253 7837 11287 7871
rect 12081 7837 12115 7871
rect 13277 7837 13311 7871
rect 14197 7837 14231 7871
rect 16773 7837 16807 7871
rect 18705 7837 18739 7871
rect 19625 7837 19659 7871
rect 20453 7837 20487 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 22845 7837 22879 7871
rect 26157 7837 26191 7871
rect 28641 7837 28675 7871
rect 30849 7837 30883 7871
rect 31861 7837 31895 7871
rect 32229 7837 32263 7871
rect 32413 7837 32447 7871
rect 33885 7837 33919 7871
rect 34713 7837 34747 7871
rect 39865 7837 39899 7871
rect 40902 7837 40936 7871
rect 41061 7837 41095 7871
rect 44373 7837 44407 7871
rect 45937 7837 45971 7871
rect 47501 7837 47535 7871
rect 50169 7837 50203 7871
rect 51641 7837 51675 7871
rect 52469 7837 52503 7871
rect 54309 7837 54343 7871
rect 54401 7837 54435 7871
rect 56692 7837 56726 7871
rect 5733 7769 5767 7803
rect 6162 7769 6196 7803
rect 9220 7769 9254 7803
rect 23112 7769 23146 7803
rect 26424 7769 26458 7803
rect 29653 7769 29687 7803
rect 32680 7769 32714 7803
rect 34529 7769 34563 7803
rect 37013 7769 37047 7803
rect 38016 7769 38050 7803
rect 42708 7769 42742 7803
rect 47768 7769 47802 7803
rect 50436 7769 50470 7803
rect 52285 7769 52319 7803
rect 52736 7769 52770 7803
rect 10701 7701 10735 7735
rect 11161 7701 11195 7735
rect 13921 7701 13955 7735
rect 14749 7701 14783 7735
rect 15485 7701 15519 7735
rect 15945 7701 15979 7735
rect 16865 7701 16899 7735
rect 18153 7701 18187 7735
rect 19257 7701 19291 7735
rect 19717 7701 19751 7735
rect 22109 7701 22143 7735
rect 24409 7701 24443 7735
rect 24777 7701 24811 7735
rect 24869 7701 24903 7735
rect 25329 7701 25363 7735
rect 25697 7701 25731 7735
rect 25789 7701 25823 7735
rect 29193 7701 29227 7735
rect 30205 7701 30239 7735
rect 31493 7701 31527 7735
rect 36553 7701 36587 7735
rect 36645 7701 36679 7735
rect 37105 7701 37139 7735
rect 39129 7701 39163 7735
rect 41705 7701 41739 7735
rect 43913 7701 43947 7735
rect 44281 7701 44315 7735
rect 46857 7701 46891 7735
rect 49617 7701 49651 7735
rect 53941 7701 53975 7735
rect 54953 7701 54987 7735
rect 56241 7701 56275 7735
rect 3801 7497 3835 7531
rect 5825 7497 5859 7531
rect 6193 7497 6227 7531
rect 20545 7497 20579 7531
rect 23949 7497 23983 7531
rect 24685 7497 24719 7531
rect 25421 7497 25455 7531
rect 26617 7497 26651 7531
rect 27629 7497 27663 7531
rect 28733 7497 28767 7531
rect 29101 7497 29135 7531
rect 33149 7497 33183 7531
rect 36093 7497 36127 7531
rect 36553 7497 36587 7531
rect 38209 7497 38243 7531
rect 39313 7497 39347 7531
rect 39681 7497 39715 7531
rect 41429 7497 41463 7531
rect 42165 7497 42199 7531
rect 43269 7497 43303 7531
rect 44005 7497 44039 7531
rect 46489 7497 46523 7531
rect 47961 7497 47995 7531
rect 48421 7497 48455 7531
rect 50813 7497 50847 7531
rect 51181 7497 51215 7531
rect 53573 7497 53607 7531
rect 54309 7497 54343 7531
rect 55045 7497 55079 7531
rect 55321 7497 55355 7531
rect 56057 7497 56091 7531
rect 56885 7497 56919 7531
rect 58449 7497 58483 7531
rect 6929 7429 6963 7463
rect 7205 7429 7239 7463
rect 13360 7429 13394 7463
rect 14841 7429 14875 7463
rect 25789 7429 25823 7463
rect 37933 7429 37967 7463
rect 38945 7429 38979 7463
rect 41061 7429 41095 7463
rect 44741 7429 44775 7463
rect 47777 7429 47811 7463
rect 55781 7429 55815 7463
rect 7389 7361 7423 7395
rect 10232 7361 10266 7395
rect 11529 7361 11563 7395
rect 13093 7361 13127 7395
rect 15292 7361 15326 7395
rect 16681 7361 16715 7395
rect 16948 7361 16982 7395
rect 18429 7361 18463 7395
rect 18696 7361 18730 7395
rect 23397 7361 23431 7395
rect 24133 7361 24167 7395
rect 24777 7361 24811 7395
rect 26985 7361 27019 7395
rect 29193 7361 29227 7395
rect 30205 7361 30239 7395
rect 30564 7361 30598 7395
rect 33517 7361 33551 7395
rect 34888 7361 34922 7395
rect 36461 7361 36495 7395
rect 38853 7361 38887 7395
rect 39773 7361 39807 7395
rect 40785 7361 40819 7395
rect 43453 7361 43487 7395
rect 44097 7361 44131 7395
rect 45109 7361 45143 7395
rect 45376 7361 45410 7395
rect 47225 7361 47259 7395
rect 48329 7361 48363 7395
rect 48881 7361 48915 7395
rect 49065 7361 49099 7395
rect 49918 7361 49952 7395
rect 51273 7361 51307 7395
rect 53021 7361 53055 7395
rect 53757 7361 53791 7395
rect 54493 7361 54527 7395
rect 58357 7361 58391 7395
rect 2605 7293 2639 7327
rect 9229 7293 9263 7327
rect 9965 7293 9999 7327
rect 12173 7293 12207 7327
rect 15025 7293 15059 7327
rect 19901 7293 19935 7327
rect 25973 7293 26007 7327
rect 29285 7293 29319 7327
rect 29653 7293 29687 7327
rect 30297 7293 30331 7327
rect 32137 7293 32171 7327
rect 33609 7293 33643 7327
rect 33793 7293 33827 7327
rect 34253 7293 34287 7327
rect 34621 7293 34655 7327
rect 36737 7293 36771 7327
rect 37289 7293 37323 7327
rect 39037 7293 39071 7327
rect 39865 7293 39899 7327
rect 40141 7293 40175 7327
rect 46581 7293 46615 7327
rect 48513 7293 48547 7327
rect 49801 7293 49835 7327
rect 50077 7293 50111 7327
rect 51365 7293 51399 7327
rect 57069 7293 57103 7327
rect 12817 7225 12851 7259
rect 14473 7225 14507 7259
rect 16405 7225 16439 7259
rect 19809 7225 19843 7259
rect 28549 7225 28583 7259
rect 36001 7225 36035 7259
rect 49525 7225 49559 7259
rect 3249 7157 3283 7191
rect 8677 7157 8711 7191
rect 9873 7157 9907 7191
rect 11345 7157 11379 7191
rect 18061 7157 18095 7191
rect 20913 7157 20947 7191
rect 31677 7157 31711 7191
rect 32781 7157 32815 7191
rect 38485 7157 38519 7191
rect 41889 7157 41923 7191
rect 42625 7157 42659 7191
rect 50721 7157 50755 7191
rect 52193 7157 52227 7191
rect 52561 7157 52595 7191
rect 56517 7157 56551 7191
rect 57713 7157 57747 7191
rect 58081 7157 58115 7191
rect 13185 6953 13219 6987
rect 19901 6953 19935 6987
rect 32045 6953 32079 6987
rect 33517 6953 33551 6987
rect 34345 6953 34379 6987
rect 34989 6953 35023 6987
rect 36737 6953 36771 6987
rect 37749 6953 37783 6987
rect 39681 6953 39715 6987
rect 40141 6953 40175 6987
rect 45477 6953 45511 6987
rect 48605 6953 48639 6987
rect 49525 6953 49559 6987
rect 50721 6953 50755 6987
rect 51641 6953 51675 6987
rect 55873 6953 55907 6987
rect 56609 6953 56643 6987
rect 3525 6885 3559 6919
rect 8769 6885 8803 6919
rect 14105 6885 14139 6919
rect 37105 6885 37139 6919
rect 49065 6885 49099 6919
rect 52745 6885 52779 6919
rect 56241 6885 56275 6919
rect 10149 6817 10183 6851
rect 10542 6817 10576 6851
rect 10701 6817 10735 6851
rect 13737 6817 13771 6851
rect 14657 6817 14691 6851
rect 15025 6817 15059 6851
rect 15669 6817 15703 6851
rect 16062 6817 16096 6851
rect 16221 6817 16255 6851
rect 18245 6817 18279 6851
rect 19257 6817 19291 6851
rect 25053 6817 25087 6851
rect 30573 6817 30607 6851
rect 32597 6817 32631 6851
rect 33793 6817 33827 6851
rect 36185 6817 36219 6851
rect 38393 6817 38427 6851
rect 38945 6817 38979 6851
rect 39129 6817 39163 6851
rect 40417 6817 40451 6851
rect 41889 6817 41923 6851
rect 42257 6817 42291 6851
rect 44465 6817 44499 6851
rect 46121 6817 46155 6851
rect 46949 6817 46983 6851
rect 47777 6817 47811 6851
rect 52009 6817 52043 6851
rect 53389 6817 53423 6851
rect 54217 6817 54251 6851
rect 56793 6817 56827 6851
rect 2145 6749 2179 6783
rect 3893 6749 3927 6783
rect 6745 6749 6779 6783
rect 7389 6749 7423 6783
rect 9505 6749 9539 6783
rect 9689 6749 9723 6783
rect 10425 6749 10459 6783
rect 11437 6749 11471 6783
rect 15209 6749 15243 6783
rect 15945 6749 15979 6783
rect 27997 6749 28031 6783
rect 28264 6749 28298 6783
rect 30840 6749 30874 6783
rect 32873 6749 32907 6783
rect 36001 6749 36035 6783
rect 37473 6749 37507 6783
rect 44741 6749 44775 6783
rect 45845 6749 45879 6783
rect 46305 6749 46339 6783
rect 52193 6749 52227 6783
rect 53297 6749 53331 6783
rect 54033 6749 54067 6783
rect 54585 6749 54619 6783
rect 58449 6749 58483 6783
rect 2412 6681 2446 6715
rect 7634 6681 7668 6715
rect 11704 6681 11738 6715
rect 13553 6681 13587 6715
rect 18981 6681 19015 6715
rect 24869 6681 24903 6715
rect 32505 6681 32539 6715
rect 35817 6681 35851 6715
rect 40877 6681 40911 6715
rect 41705 6681 41739 6715
rect 42993 6681 43027 6715
rect 43361 6681 43395 6715
rect 45293 6681 45327 6715
rect 53205 6681 53239 6715
rect 55137 6681 55171 6715
rect 57060 6681 57094 6715
rect 4445 6613 4479 6647
rect 7297 6613 7331 6647
rect 9321 6613 9355 6647
rect 11345 6613 11379 6647
rect 12817 6613 12851 6647
rect 13645 6613 13679 6647
rect 14473 6613 14507 6647
rect 14565 6613 14599 6647
rect 16865 6613 16899 6647
rect 20269 6613 20303 6647
rect 20637 6613 20671 6647
rect 24593 6613 24627 6647
rect 29377 6613 29411 6647
rect 30113 6613 30147 6647
rect 30481 6613 30515 6647
rect 31953 6613 31987 6647
rect 32413 6613 32447 6647
rect 35357 6613 35391 6647
rect 38209 6613 38243 6647
rect 41153 6613 41187 6647
rect 42533 6613 42567 6647
rect 43729 6613 43763 6647
rect 45937 6613 45971 6647
rect 47225 6613 47259 6647
rect 48237 6613 48271 6647
rect 52837 6613 52871 6647
rect 53665 6613 53699 6647
rect 54125 6613 54159 6647
rect 55505 6613 55539 6647
rect 58173 6613 58207 6647
rect 58265 6613 58299 6647
rect 2237 6409 2271 6443
rect 3341 6409 3375 6443
rect 7665 6409 7699 6443
rect 8033 6409 8067 6443
rect 13093 6409 13127 6443
rect 15301 6409 15335 6443
rect 19257 6409 19291 6443
rect 21557 6409 21591 6443
rect 22201 6409 22235 6443
rect 24317 6409 24351 6443
rect 26433 6409 26467 6443
rect 29561 6409 29595 6443
rect 33425 6409 33459 6443
rect 37565 6409 37599 6443
rect 39497 6409 39531 6443
rect 40969 6409 41003 6443
rect 41337 6409 41371 6443
rect 42165 6409 42199 6443
rect 42993 6409 43027 6443
rect 43361 6409 43395 6443
rect 46029 6409 46063 6443
rect 48881 6409 48915 6443
rect 49249 6409 49283 6443
rect 51181 6409 51215 6443
rect 51549 6409 51583 6443
rect 54493 6409 54527 6443
rect 3801 6341 3835 6375
rect 5457 6341 5491 6375
rect 5834 6341 5868 6375
rect 10241 6341 10275 6375
rect 11989 6341 12023 6375
rect 18889 6341 18923 6375
rect 32781 6341 32815 6375
rect 34161 6341 34195 6375
rect 35725 6341 35759 6375
rect 52990 6341 53024 6375
rect 2053 6273 2087 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2513 6273 2547 6307
rect 2605 6273 2639 6307
rect 3617 6273 3651 6307
rect 6101 6273 6135 6307
rect 7573 6273 7607 6307
rect 8677 6273 8711 6307
rect 9781 6273 9815 6307
rect 10057 6273 10091 6307
rect 11897 6273 11931 6307
rect 13185 6273 13219 6307
rect 13452 6273 13486 6307
rect 19165 6273 19199 6307
rect 20729 6273 20763 6307
rect 24593 6273 24627 6307
rect 27813 6273 27847 6307
rect 28080 6273 28114 6307
rect 29929 6273 29963 6307
rect 30849 6273 30883 6307
rect 33977 6273 34011 6307
rect 34897 6273 34931 6307
rect 36185 6273 36219 6307
rect 40877 6273 40911 6307
rect 45937 6273 45971 6307
rect 50077 6273 50111 6307
rect 52377 6273 52411 6307
rect 52745 6273 52779 6307
rect 54953 6273 54987 6307
rect 55806 6273 55840 6307
rect 57069 6273 57103 6307
rect 57713 6273 57747 6307
rect 2697 6205 2731 6239
rect 8125 6205 8159 6239
rect 8217 6205 8251 6239
rect 8861 6205 8895 6239
rect 12173 6205 12207 6239
rect 12449 6205 12483 6239
rect 14657 6205 14691 6239
rect 19625 6205 19659 6239
rect 19809 6205 19843 6239
rect 20545 6205 20579 6239
rect 25053 6205 25087 6239
rect 25421 6205 25455 6239
rect 30113 6205 30147 6239
rect 30966 6205 31000 6239
rect 31125 6205 31159 6239
rect 32137 6205 32171 6239
rect 37841 6205 37875 6239
rect 38577 6205 38611 6239
rect 42625 6205 42659 6239
rect 44189 6205 44223 6239
rect 44925 6205 44959 6239
rect 47133 6205 47167 6239
rect 49617 6205 49651 6239
rect 52101 6205 52135 6239
rect 54769 6205 54803 6239
rect 55689 6205 55723 6239
rect 55965 6205 55999 6239
rect 57161 6205 57195 6239
rect 57253 6205 57287 6239
rect 57897 6205 57931 6239
rect 2329 6137 2363 6171
rect 11529 6137 11563 6171
rect 14565 6137 14599 6171
rect 17785 6137 17819 6171
rect 21189 6137 21223 6171
rect 22845 6137 22879 6171
rect 29193 6137 29227 6171
rect 30573 6137 30607 6171
rect 36553 6137 36587 6171
rect 38209 6137 38243 6171
rect 46857 6137 46891 6171
rect 47869 6137 47903 6171
rect 48237 6137 48271 6171
rect 48605 6137 48639 6171
rect 52561 6137 52595 6171
rect 55413 6137 55447 6171
rect 56701 6137 56735 6171
rect 3985 6069 4019 6103
rect 5825 6069 5859 6103
rect 15577 6069 15611 6103
rect 16865 6069 16899 6103
rect 18521 6069 18555 6103
rect 20453 6069 20487 6103
rect 20913 6069 20947 6103
rect 22477 6069 22511 6103
rect 23397 6069 23431 6103
rect 26065 6069 26099 6103
rect 31769 6069 31803 6103
rect 33057 6069 33091 6103
rect 34437 6069 34471 6103
rect 36921 6069 36955 6103
rect 39129 6069 39163 6103
rect 39865 6069 39899 6103
rect 40233 6069 40267 6103
rect 40601 6069 40635 6103
rect 41705 6069 41739 6103
rect 43729 6069 43763 6103
rect 44465 6069 44499 6103
rect 45477 6069 45511 6103
rect 46489 6069 46523 6103
rect 50353 6069 50387 6103
rect 50721 6069 50755 6103
rect 54125 6069 54159 6103
rect 56609 6069 56643 6103
rect 57529 6069 57563 6103
rect 58541 6069 58575 6103
rect 5273 5865 5307 5899
rect 8493 5865 8527 5899
rect 9597 5865 9631 5899
rect 11345 5865 11379 5899
rect 12357 5865 12391 5899
rect 13093 5865 13127 5899
rect 14749 5865 14783 5899
rect 17785 5865 17819 5899
rect 28273 5865 28307 5899
rect 30849 5865 30883 5899
rect 33333 5865 33367 5899
rect 34529 5865 34563 5899
rect 38117 5865 38151 5899
rect 38761 5865 38795 5899
rect 45017 5865 45051 5899
rect 46857 5865 46891 5899
rect 49617 5865 49651 5899
rect 54033 5865 54067 5899
rect 57345 5865 57379 5899
rect 57437 5865 57471 5899
rect 58265 5865 58299 5899
rect 12633 5797 12667 5831
rect 37289 5797 37323 5831
rect 41153 5797 41187 5831
rect 50169 5797 50203 5831
rect 4353 5729 4387 5763
rect 11713 5729 11747 5763
rect 14105 5729 14139 5763
rect 15485 5729 15519 5763
rect 19809 5729 19843 5763
rect 19901 5729 19935 5763
rect 22569 5729 22603 5763
rect 22661 5729 22695 5763
rect 24409 5729 24443 5763
rect 26433 5729 26467 5763
rect 29009 5729 29043 5763
rect 31401 5729 31435 5763
rect 32689 5729 32723 5763
rect 35909 5729 35943 5763
rect 39221 5729 39255 5763
rect 39405 5729 39439 5763
rect 41613 5729 41647 5763
rect 41797 5729 41831 5763
rect 41981 5729 42015 5763
rect 45661 5729 45695 5763
rect 47225 5729 47259 5763
rect 50721 5729 50755 5763
rect 51733 5729 51767 5763
rect 52653 5729 52687 5763
rect 55965 5729 55999 5763
rect 57989 5729 58023 5763
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 5641 5661 5675 5695
rect 5825 5661 5859 5695
rect 6285 5661 6319 5695
rect 6929 5661 6963 5695
rect 16497 5661 16531 5695
rect 17877 5661 17911 5695
rect 18061 5661 18095 5695
rect 18521 5661 18555 5695
rect 23397 5661 23431 5695
rect 23673 5661 23707 5695
rect 26709 5661 26743 5695
rect 28917 5661 28951 5695
rect 29745 5661 29779 5695
rect 31861 5661 31895 5695
rect 33609 5661 33643 5695
rect 34713 5661 34747 5695
rect 37381 5661 37415 5695
rect 38301 5661 38335 5695
rect 39865 5661 39899 5695
rect 42901 5661 42935 5695
rect 43269 5661 43303 5695
rect 44005 5661 44039 5695
rect 45385 5661 45419 5695
rect 45845 5661 45879 5695
rect 48697 5661 48731 5695
rect 50537 5661 50571 5695
rect 50997 5661 51031 5695
rect 54125 5661 54159 5695
rect 55137 5661 55171 5695
rect 55505 5661 55539 5695
rect 55689 5661 55723 5695
rect 56232 5661 56266 5695
rect 57805 5661 57839 5695
rect 58449 5661 58483 5695
rect 2697 5593 2731 5627
rect 2881 5593 2915 5627
rect 5089 5593 5123 5627
rect 8217 5593 8251 5627
rect 15117 5593 15151 5627
rect 20269 5593 20303 5627
rect 24676 5593 24710 5627
rect 26249 5593 26283 5627
rect 27353 5593 27387 5627
rect 28825 5593 28859 5627
rect 30573 5593 30607 5627
rect 31309 5593 31343 5627
rect 32321 5593 32355 5627
rect 32965 5593 32999 5627
rect 35541 5593 35575 5627
rect 36176 5593 36210 5627
rect 38025 5593 38059 5627
rect 39129 5593 39163 5627
rect 40509 5593 40543 5627
rect 41521 5593 41555 5627
rect 47492 5593 47526 5627
rect 49341 5593 49375 5627
rect 52920 5593 52954 5627
rect 54769 5593 54803 5627
rect 3065 5525 3099 5559
rect 5273 5525 5307 5559
rect 5457 5525 5491 5559
rect 9229 5525 9263 5559
rect 9965 5525 9999 5559
rect 11069 5525 11103 5559
rect 13369 5525 13403 5559
rect 15853 5525 15887 5559
rect 17141 5525 17175 5559
rect 18245 5525 18279 5559
rect 19073 5525 19107 5559
rect 19349 5525 19383 5559
rect 19717 5525 19751 5559
rect 21557 5525 21591 5559
rect 22109 5525 22143 5559
rect 22477 5525 22511 5559
rect 24225 5525 24259 5559
rect 25789 5525 25823 5559
rect 25881 5525 25915 5559
rect 26341 5525 26375 5559
rect 28457 5525 28491 5559
rect 31217 5525 31251 5559
rect 34161 5525 34195 5559
rect 38669 5525 38703 5559
rect 40785 5525 40819 5559
rect 42625 5525 42659 5559
rect 43821 5525 43855 5559
rect 44649 5525 44683 5559
rect 45477 5525 45511 5559
rect 46489 5525 46523 5559
rect 48605 5525 48639 5559
rect 50629 5525 50663 5559
rect 51641 5525 51675 5559
rect 52377 5525 52411 5559
rect 54953 5525 54987 5559
rect 55873 5525 55907 5559
rect 57897 5525 57931 5559
rect 4537 5321 4571 5355
rect 7849 5321 7883 5355
rect 10241 5321 10275 5355
rect 14473 5321 14507 5355
rect 14749 5321 14783 5355
rect 15577 5321 15611 5355
rect 19717 5321 19751 5355
rect 22293 5321 22327 5355
rect 24133 5321 24167 5355
rect 27353 5321 27387 5355
rect 28917 5321 28951 5355
rect 29009 5321 29043 5355
rect 30205 5321 30239 5355
rect 30941 5321 30975 5355
rect 31309 5321 31343 5355
rect 39313 5321 39347 5355
rect 41797 5321 41831 5355
rect 45661 5321 45695 5355
rect 46121 5321 46155 5355
rect 48145 5321 48179 5355
rect 51825 5321 51859 5355
rect 53757 5321 53791 5355
rect 54769 5321 54803 5355
rect 57713 5321 57747 5355
rect 58541 5321 58575 5355
rect 3801 5253 3835 5287
rect 6561 5253 6595 5287
rect 14381 5253 14415 5287
rect 16497 5253 16531 5287
rect 18604 5253 18638 5287
rect 26801 5253 26835 5287
rect 32321 5253 32355 5287
rect 33324 5253 33358 5287
rect 38200 5253 38234 5287
rect 42984 5253 43018 5287
rect 44548 5253 44582 5287
rect 53297 5253 53331 5287
rect 55505 5253 55539 5287
rect 3893 5185 3927 5219
rect 5365 5185 5399 5219
rect 6653 5185 6687 5219
rect 7021 5185 7055 5219
rect 9689 5185 9723 5219
rect 11529 5185 11563 5219
rect 12541 5185 12575 5219
rect 14933 5185 14967 5219
rect 15209 5185 15243 5219
rect 15761 5185 15795 5219
rect 16865 5185 16899 5219
rect 18081 5183 18115 5217
rect 18337 5185 18371 5219
rect 19809 5185 19843 5219
rect 21005 5185 21039 5219
rect 21649 5185 21683 5219
rect 22201 5185 22235 5219
rect 22753 5185 22787 5219
rect 23020 5185 23054 5219
rect 25605 5185 25639 5219
rect 28365 5185 28399 5219
rect 29193 5185 29227 5219
rect 29653 5185 29687 5219
rect 30481 5185 30515 5219
rect 31217 5185 31251 5219
rect 33057 5185 33091 5219
rect 34805 5185 34839 5219
rect 35081 5185 35115 5219
rect 35265 5185 35299 5219
rect 36001 5185 36035 5219
rect 36277 5185 36311 5219
rect 37657 5185 37691 5219
rect 40325 5185 40359 5219
rect 40442 5185 40476 5219
rect 41245 5185 41279 5219
rect 41705 5185 41739 5219
rect 42717 5185 42751 5219
rect 48053 5185 48087 5219
rect 49433 5185 49467 5219
rect 49709 5185 49743 5219
rect 50445 5185 50479 5219
rect 50712 5185 50746 5219
rect 54033 5185 54067 5219
rect 57069 5185 57103 5219
rect 57897 5185 57931 5219
rect 2145 5117 2179 5151
rect 2421 5117 2455 5151
rect 5273 5117 5307 5151
rect 5825 5117 5859 5151
rect 7113 5117 7147 5151
rect 8033 5117 8067 5151
rect 8861 5117 8895 5151
rect 10793 5117 10827 5151
rect 12173 5117 12207 5151
rect 13093 5117 13127 5151
rect 14197 5117 14231 5151
rect 15025 5117 15059 5151
rect 17417 5117 17451 5151
rect 17877 5117 17911 5151
rect 19993 5117 20027 5151
rect 20729 5117 20763 5151
rect 20846 5117 20880 5151
rect 22385 5117 22419 5151
rect 24409 5117 24443 5151
rect 24593 5117 24627 5151
rect 25329 5117 25363 5151
rect 25446 5117 25480 5151
rect 26249 5117 26283 5151
rect 27445 5117 27479 5151
rect 27537 5117 27571 5151
rect 30297 5117 30331 5151
rect 34621 5117 34655 5151
rect 36118 5117 36152 5151
rect 37473 5117 37507 5151
rect 37933 5117 37967 5151
rect 39405 5117 39439 5151
rect 39589 5117 39623 5151
rect 40601 5117 40635 5151
rect 41981 5117 42015 5151
rect 44281 5117 44315 5151
rect 46213 5117 46247 5151
rect 46397 5117 46431 5151
rect 46857 5117 46891 5151
rect 48237 5117 48271 5151
rect 48513 5117 48547 5151
rect 48697 5117 48731 5151
rect 49550 5117 49584 5151
rect 52561 5117 52595 5151
rect 54217 5117 54251 5151
rect 54953 5117 54987 5151
rect 55689 5117 55723 5151
rect 56333 5117 56367 5151
rect 10517 5049 10551 5083
rect 13461 5049 13495 5083
rect 20453 5049 20487 5083
rect 25053 5049 25087 5083
rect 26985 5049 27019 5083
rect 31769 5049 31803 5083
rect 35725 5049 35759 5083
rect 40049 5049 40083 5083
rect 47685 5049 47719 5083
rect 49157 5049 49191 5083
rect 5733 4981 5767 5015
rect 6101 4981 6135 5015
rect 8585 4981 8619 5015
rect 9413 4981 9447 5015
rect 9781 4981 9815 5015
rect 11345 4981 11379 5015
rect 13829 4981 13863 5015
rect 15393 4981 15427 5015
rect 16037 4981 16071 5015
rect 16957 4981 16991 5015
rect 17785 4981 17819 5015
rect 18245 4981 18279 5015
rect 21833 4981 21867 5015
rect 28181 4981 28215 5015
rect 30665 4981 30699 5015
rect 32689 4981 32723 5015
rect 34437 4981 34471 5015
rect 34989 4981 35023 5015
rect 36921 4981 36955 5015
rect 37841 4981 37875 5015
rect 41337 4981 41371 5015
rect 44097 4981 44131 5015
rect 45753 4981 45787 5015
rect 47409 4981 47443 5015
rect 50353 4981 50387 5015
rect 52101 4981 52135 5015
rect 52929 4981 52963 5015
rect 53849 4981 53883 5015
rect 56241 4981 56275 5015
rect 56977 4981 57011 5015
rect 2145 4777 2179 4811
rect 2697 4777 2731 4811
rect 2881 4777 2915 4811
rect 3985 4777 4019 4811
rect 6009 4777 6043 4811
rect 7849 4777 7883 4811
rect 8033 4777 8067 4811
rect 22293 4777 22327 4811
rect 26801 4777 26835 4811
rect 33609 4777 33643 4811
rect 36093 4777 36127 4811
rect 39681 4777 39715 4811
rect 42349 4777 42383 4811
rect 43085 4777 43119 4811
rect 43361 4777 43395 4811
rect 46857 4777 46891 4811
rect 48329 4777 48363 4811
rect 48421 4777 48455 4811
rect 51825 4777 51859 4811
rect 54953 4777 54987 4811
rect 56333 4777 56367 4811
rect 4169 4709 4203 4743
rect 5549 4709 5583 4743
rect 5641 4709 5675 4743
rect 6331 4709 6365 4743
rect 6469 4709 6503 4743
rect 10241 4709 10275 4743
rect 10517 4709 10551 4743
rect 28089 4709 28123 4743
rect 31217 4709 31251 4743
rect 37013 4709 37047 4743
rect 44189 4709 44223 4743
rect 44557 4709 44591 4743
rect 52561 4709 52595 4743
rect 5181 4641 5215 4675
rect 5733 4641 5767 4675
rect 6561 4641 6595 4675
rect 8493 4641 8527 4675
rect 8677 4641 8711 4675
rect 9321 4641 9355 4675
rect 10977 4641 11011 4675
rect 11069 4641 11103 4675
rect 11713 4641 11747 4675
rect 12449 4641 12483 4675
rect 15945 4641 15979 4675
rect 19257 4641 19291 4675
rect 23949 4641 23983 4675
rect 24133 4641 24167 4675
rect 25053 4641 25087 4675
rect 25145 4641 25179 4675
rect 25421 4641 25455 4675
rect 31861 4641 31895 4675
rect 34069 4641 34103 4675
rect 34253 4641 34287 4675
rect 34713 4641 34747 4675
rect 36645 4641 36679 4675
rect 36737 4641 36771 4675
rect 37657 4641 37691 4675
rect 40509 4641 40543 4675
rect 40969 4641 41003 4675
rect 42441 4641 42475 4675
rect 43913 4641 43947 4675
rect 45017 4641 45051 4675
rect 45201 4641 45235 4675
rect 45661 4641 45695 4675
rect 45937 4641 45971 4675
rect 46213 4641 46247 4675
rect 46949 4641 46983 4675
rect 48973 4641 49007 4675
rect 49341 4641 49375 4675
rect 50629 4641 50663 4675
rect 50813 4641 50847 4675
rect 53113 4641 53147 4675
rect 53389 4641 53423 4675
rect 55965 4641 55999 4675
rect 56793 4641 56827 4675
rect 56977 4641 57011 4675
rect 2053 4573 2087 4607
rect 2237 4573 2271 4607
rect 2329 4573 2363 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 6193 4573 6227 4607
rect 7573 4573 7607 4607
rect 9137 4573 9171 4607
rect 10425 4573 10459 4607
rect 11345 4573 11379 4607
rect 13369 4573 13403 4607
rect 14289 4573 14323 4607
rect 15025 4573 15059 4607
rect 16212 4573 16246 4607
rect 17417 4573 17451 4607
rect 18521 4573 18555 4607
rect 20913 4573 20947 4607
rect 22385 4573 22419 4607
rect 23397 4573 23431 4607
rect 27629 4573 27663 4607
rect 28273 4573 28307 4607
rect 28825 4573 28859 4607
rect 29745 4573 29779 4607
rect 30573 4573 30607 4607
rect 32045 4573 32079 4607
rect 32873 4573 32907 4607
rect 36553 4573 36587 4607
rect 37841 4573 37875 4607
rect 38025 4573 38059 4607
rect 38301 4573 38335 4607
rect 40877 4573 40911 4607
rect 43821 4573 43855 4607
rect 44373 4573 44407 4607
rect 44741 4573 44775 4607
rect 46054 4573 46088 4607
rect 47216 4573 47250 4607
rect 48789 4573 48823 4607
rect 51457 4573 51491 4607
rect 54033 4573 54067 4607
rect 54125 4573 54159 4607
rect 55137 4573 55171 4607
rect 55689 4573 55723 4607
rect 56701 4573 56735 4607
rect 57161 4573 57195 4607
rect 2697 4505 2731 4539
rect 3801 4505 3835 4539
rect 4001 4505 4035 4539
rect 8401 4505 8435 4539
rect 10885 4505 10919 4539
rect 19524 4505 19558 4539
rect 21180 4505 21214 4539
rect 23029 4505 23063 4539
rect 23857 4505 23891 4539
rect 25688 4505 25722 4539
rect 31585 4505 31619 4539
rect 33333 4505 33367 4539
rect 34980 4505 35014 4539
rect 38568 4505 38602 4539
rect 40233 4505 40267 4539
rect 41236 4505 41270 4539
rect 43729 4505 43763 4539
rect 50537 4505 50571 4539
rect 52929 4505 52963 4539
rect 53021 4505 53055 4539
rect 54769 4505 54803 4539
rect 58357 4505 58391 4539
rect 2973 4437 3007 4471
rect 3341 4437 3375 4471
rect 4721 4437 4755 4471
rect 5089 4437 5123 4471
rect 6837 4437 6871 4471
rect 13093 4437 13127 4471
rect 13921 4437 13955 4471
rect 14841 4437 14875 4471
rect 15577 4437 15611 4471
rect 17325 4437 17359 4471
rect 18061 4437 18095 4471
rect 19073 4437 19107 4471
rect 20637 4437 20671 4471
rect 23489 4437 23523 4471
rect 24593 4437 24627 4471
rect 24961 4437 24995 4471
rect 27169 4437 27203 4471
rect 27905 4437 27939 4471
rect 28641 4437 28675 4471
rect 29377 4437 29411 4471
rect 30389 4437 30423 4471
rect 31125 4437 31159 4471
rect 31677 4437 31711 4471
rect 33425 4437 33459 4471
rect 33977 4437 34011 4471
rect 36185 4437 36219 4471
rect 37381 4437 37415 4471
rect 37473 4437 37507 4471
rect 38209 4437 38243 4471
rect 39865 4437 39899 4471
rect 40325 4437 40359 4471
rect 40693 4437 40727 4471
rect 48881 4437 48915 4471
rect 49893 4437 49927 4471
rect 50169 4437 50203 4471
rect 51273 4437 51307 4471
rect 52101 4437 52135 4471
rect 55321 4437 55355 4471
rect 55781 4437 55815 4471
rect 7021 4233 7055 4267
rect 8953 4233 8987 4267
rect 14749 4233 14783 4267
rect 15209 4233 15243 4267
rect 16221 4233 16255 4267
rect 17877 4233 17911 4267
rect 19533 4233 19567 4267
rect 23949 4233 23983 4267
rect 26433 4233 26467 4267
rect 29469 4233 29503 4267
rect 31953 4233 31987 4267
rect 34897 4233 34931 4267
rect 36001 4233 36035 4267
rect 38025 4233 38059 4267
rect 39865 4233 39899 4267
rect 40693 4233 40727 4267
rect 43637 4233 43671 4267
rect 45201 4233 45235 4267
rect 45753 4233 45787 4267
rect 48881 4233 48915 4267
rect 49433 4233 49467 4267
rect 56793 4233 56827 4267
rect 3893 4165 3927 4199
rect 6377 4165 6411 4199
rect 15117 4165 15151 4199
rect 27353 4165 27387 4199
rect 41797 4165 41831 4199
rect 42441 4165 42475 4199
rect 43913 4165 43947 4199
rect 46121 4165 46155 4199
rect 47225 4165 47259 4199
rect 49341 4165 49375 4199
rect 51181 4165 51215 4199
rect 2421 4097 2455 4131
rect 3065 4097 3099 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5457 4097 5491 4131
rect 6193 4097 6227 4131
rect 7205 4097 7239 4131
rect 7840 4097 7874 4131
rect 11345 4097 11379 4131
rect 11529 4097 11563 4131
rect 11796 4097 11830 4131
rect 13185 4097 13219 4131
rect 13277 4097 13311 4131
rect 13544 4097 13578 4131
rect 16497 4097 16531 4131
rect 17049 4097 17083 4131
rect 17141 4097 17175 4131
rect 19625 4097 19659 4131
rect 20269 4097 20303 4131
rect 20913 4097 20947 4131
rect 21557 4097 21591 4131
rect 22477 4097 22511 4131
rect 22845 4097 22879 4131
rect 23029 4097 23063 4131
rect 23397 4097 23431 4131
rect 24225 4097 24259 4131
rect 24409 4097 24443 4131
rect 24685 4097 24719 4131
rect 25329 4097 25363 4131
rect 25605 4097 25639 4131
rect 25881 4097 25915 4131
rect 26801 4097 26835 4131
rect 27169 4097 27203 4131
rect 27629 4097 27663 4131
rect 28356 4097 28390 4131
rect 29653 4097 29687 4131
rect 29745 4097 29779 4131
rect 30113 4097 30147 4131
rect 31309 4097 31343 4131
rect 32229 4097 32263 4131
rect 33241 4097 33275 4131
rect 34989 4097 35023 4131
rect 36093 4097 36127 4131
rect 37105 4097 37139 4131
rect 39037 4097 39071 4131
rect 39313 4097 39347 4131
rect 40049 4097 40083 4131
rect 40877 4097 40911 4131
rect 40969 4097 41003 4131
rect 41429 4097 41463 4131
rect 42073 4097 42107 4131
rect 43085 4097 43119 4131
rect 43545 4097 43579 4131
rect 43821 4097 43855 4131
rect 46581 4097 46615 4131
rect 47869 4097 47903 4131
rect 48237 4097 48271 4131
rect 52745 4097 52779 4131
rect 53012 4097 53046 4131
rect 54401 4097 54435 4131
rect 54677 4097 54711 4131
rect 57437 4097 57471 4131
rect 57897 4097 57931 4131
rect 4353 4029 4387 4063
rect 6745 4029 6779 4063
rect 7573 4029 7607 4063
rect 9045 4029 9079 4063
rect 9229 4029 9263 4063
rect 9965 4029 9999 4063
rect 10103 4029 10137 4063
rect 10241 4029 10275 4063
rect 15301 4029 15335 4063
rect 15577 4029 15611 4063
rect 17233 4029 17267 4063
rect 17969 4029 18003 4063
rect 18061 4029 18095 4063
rect 18429 4029 18463 4063
rect 19717 4029 19751 4063
rect 20085 4029 20119 4063
rect 21005 4029 21039 4063
rect 21097 4029 21131 4063
rect 21925 4029 21959 4063
rect 27445 4029 27479 4063
rect 28089 4029 28123 4063
rect 30297 4029 30331 4063
rect 31033 4029 31067 4063
rect 31171 4029 31205 4063
rect 32965 4029 32999 4063
rect 34069 4029 34103 4063
rect 35081 4029 35115 4063
rect 35357 4029 35391 4063
rect 36737 4029 36771 4063
rect 37381 4029 37415 4063
rect 38117 4029 38151 4063
rect 41245 4029 41279 4063
rect 41981 4029 42015 4063
rect 42809 4029 42843 4063
rect 42901 4029 42935 4063
rect 46213 4029 46247 4063
rect 46305 4029 46339 4063
rect 49525 4029 49559 4063
rect 49801 4029 49835 4063
rect 50537 4029 50571 4063
rect 51641 4029 51675 4063
rect 52009 4029 52043 4063
rect 54493 4029 54527 4063
rect 55413 4029 55447 4063
rect 55530 4029 55564 4063
rect 55689 4029 55723 4063
rect 56333 4029 56367 4063
rect 56885 4029 56919 4063
rect 56977 4029 57011 4063
rect 57253 4029 57287 4063
rect 3249 3961 3283 3995
rect 3893 3961 3927 3995
rect 5089 3961 5123 3995
rect 6561 3961 6595 3995
rect 9689 3961 9723 3995
rect 11161 3961 11195 3995
rect 14657 3961 14691 3995
rect 17509 3961 17543 3995
rect 20453 3961 20487 3995
rect 26617 3961 26651 3995
rect 30757 3961 30791 3995
rect 34529 3961 34563 3995
rect 38853 3961 38887 3995
rect 42257 3961 42291 3995
rect 42625 3961 42659 3995
rect 48973 3961 49007 3995
rect 54125 3961 54159 3995
rect 55137 3961 55171 3995
rect 2973 3893 3007 3927
rect 5825 3893 5859 3927
rect 6377 3893 6411 3927
rect 6653 3893 6687 3927
rect 10885 3893 10919 3927
rect 12909 3893 12943 3927
rect 13001 3893 13035 3927
rect 16313 3893 16347 3927
rect 16681 3893 16715 3927
rect 18981 3893 19015 3927
rect 19165 3893 19199 3927
rect 20545 3893 20579 3927
rect 21373 3893 21407 3927
rect 23213 3893 23247 3927
rect 24593 3893 24627 3927
rect 25421 3893 25455 3927
rect 26985 3893 27019 3927
rect 27353 3893 27387 3927
rect 27813 3893 27847 3927
rect 29929 3893 29963 3927
rect 36921 3893 36955 3927
rect 38761 3893 38795 3927
rect 41153 3893 41187 3927
rect 41613 3893 41647 3927
rect 42073 3893 42107 3927
rect 42441 3893 42475 3927
rect 42717 3893 42751 3927
rect 43269 3893 43303 3927
rect 43361 3893 43395 3927
rect 47685 3893 47719 3927
rect 50445 3893 50479 3927
rect 52561 3893 52595 3927
rect 54217 3893 54251 3927
rect 56425 3893 56459 3927
rect 57621 3893 57655 3927
rect 58541 3893 58575 3927
rect 3157 3689 3191 3723
rect 6561 3689 6595 3723
rect 10057 3689 10091 3723
rect 11989 3689 12023 3723
rect 14933 3689 14967 3723
rect 17325 3689 17359 3723
rect 18797 3689 18831 3723
rect 19993 3689 20027 3723
rect 22201 3689 22235 3723
rect 22293 3689 22327 3723
rect 26709 3689 26743 3723
rect 29561 3689 29595 3723
rect 33609 3689 33643 3723
rect 34437 3689 34471 3723
rect 34713 3689 34747 3723
rect 35173 3689 35207 3723
rect 41337 3689 41371 3723
rect 44649 3689 44683 3723
rect 46489 3689 46523 3723
rect 47409 3689 47443 3723
rect 49801 3689 49835 3723
rect 50721 3689 50755 3723
rect 54953 3689 54987 3723
rect 58357 3689 58391 3723
rect 3433 3621 3467 3655
rect 4169 3621 4203 3655
rect 4445 3621 4479 3655
rect 8677 3621 8711 3655
rect 14105 3621 14139 3655
rect 16129 3621 16163 3655
rect 21465 3621 21499 3655
rect 22753 3621 22787 3655
rect 24225 3621 24259 3655
rect 31769 3621 31803 3655
rect 39681 3621 39715 3655
rect 43729 3621 43763 3655
rect 50445 3621 50479 3655
rect 58265 3621 58299 3655
rect 1777 3553 1811 3587
rect 5089 3553 5123 3587
rect 5365 3553 5399 3587
rect 5457 3553 5491 3587
rect 10609 3553 10643 3587
rect 14565 3553 14599 3587
rect 14749 3553 14783 3587
rect 16522 3553 16556 3587
rect 16681 3553 16715 3587
rect 19349 3553 19383 3587
rect 21557 3553 21591 3587
rect 22385 3553 22419 3587
rect 22845 3553 22879 3587
rect 24869 3553 24903 3587
rect 25053 3553 25087 3587
rect 25329 3553 25363 3587
rect 27077 3553 27111 3587
rect 29101 3553 29135 3587
rect 30113 3553 30147 3587
rect 30389 3553 30423 3587
rect 32229 3553 32263 3587
rect 33885 3553 33919 3587
rect 35265 3553 35299 3587
rect 35909 3553 35943 3587
rect 38301 3553 38335 3587
rect 40509 3553 40543 3587
rect 41429 3553 41463 3587
rect 42349 3553 42383 3587
rect 44281 3553 44315 3587
rect 44465 3553 44499 3587
rect 46581 3553 46615 3587
rect 47593 3553 47627 3587
rect 53389 3553 53423 3587
rect 53757 3553 53791 3587
rect 56885 3553 56919 3587
rect 3617 3485 3651 3519
rect 4813 3485 4847 3519
rect 5825 3485 5859 3519
rect 6009 3485 6043 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 7021 3485 7055 3519
rect 7297 3485 7331 3519
rect 8953 3485 8987 3519
rect 10241 3485 10275 3519
rect 12081 3485 12115 3519
rect 13369 3485 13403 3519
rect 15117 3485 15151 3519
rect 15209 3485 15243 3519
rect 15485 3485 15519 3519
rect 15669 3485 15703 3519
rect 16405 3485 16439 3519
rect 17417 3485 17451 3519
rect 20085 3485 20119 3519
rect 22569 3485 22603 3519
rect 26065 3485 26099 3519
rect 26893 3485 26927 3519
rect 30021 3485 30055 3519
rect 32045 3485 32079 3519
rect 34897 3485 34931 3519
rect 34989 3485 35023 3519
rect 35449 3485 35483 3519
rect 37381 3485 37415 3519
rect 40693 3485 40727 3519
rect 44833 3485 44867 3519
rect 45109 3485 45143 3519
rect 47685 3485 47719 3519
rect 48053 3485 48087 3519
rect 48145 3485 48179 3519
rect 48421 3485 48455 3519
rect 50997 3485 51031 3519
rect 51089 3485 51123 3519
rect 51365 3485 51399 3519
rect 54493 3485 54527 3519
rect 54585 3485 54619 3519
rect 54953 3485 54987 3519
rect 55321 3485 55355 3519
rect 57141 3485 57175 3519
rect 58541 3485 58575 3519
rect 2044 3417 2078 3451
rect 3893 3417 3927 3451
rect 5549 3417 5583 3451
rect 6377 3417 6411 3451
rect 7564 3417 7598 3451
rect 9781 3417 9815 3451
rect 10876 3417 10910 3451
rect 12909 3417 12943 3451
rect 13921 3417 13955 3451
rect 14473 3417 14507 3451
rect 14933 3417 14967 3451
rect 17684 3417 17718 3451
rect 20352 3417 20386 3451
rect 22293 3417 22327 3451
rect 23112 3417 23146 3451
rect 24777 3417 24811 3451
rect 25881 3417 25915 3451
rect 26249 3417 26283 3451
rect 26617 3417 26651 3451
rect 27344 3417 27378 3451
rect 30656 3417 30690 3451
rect 32496 3417 32530 3451
rect 34713 3417 34747 3451
rect 36176 3417 36210 3451
rect 38025 3417 38059 3451
rect 38568 3417 38602 3451
rect 40233 3417 40267 3451
rect 40325 3417 40359 3451
rect 42073 3417 42107 3451
rect 42616 3417 42650 3451
rect 45376 3417 45410 3451
rect 47225 3417 47259 3451
rect 47409 3417 47443 3451
rect 48688 3417 48722 3451
rect 50261 3417 50295 3451
rect 51632 3417 51666 3451
rect 53205 3417 53239 3451
rect 54309 3417 54343 3451
rect 55588 3417 55622 3451
rect 4353 3349 4387 3383
rect 4629 3349 4663 3383
rect 4721 3349 4755 3383
rect 4997 3349 5031 3383
rect 7205 3349 7239 3383
rect 15393 3349 15427 3383
rect 24409 3349 24443 3383
rect 28457 3349 28491 3383
rect 28549 3349 28583 3383
rect 28917 3349 28951 3383
rect 29009 3349 29043 3383
rect 29929 3349 29963 3383
rect 31861 3349 31895 3383
rect 35633 3349 35667 3383
rect 37289 3349 37323 3383
rect 39865 3349 39899 3383
rect 43821 3349 43855 3383
rect 44189 3349 44223 3383
rect 47869 3349 47903 3383
rect 48329 3349 48363 3383
rect 51273 3349 51307 3383
rect 52745 3349 52779 3383
rect 52837 3349 52871 3383
rect 53297 3349 53331 3383
rect 55137 3349 55171 3383
rect 56701 3349 56735 3383
rect 2789 3145 2823 3179
rect 4537 3145 4571 3179
rect 6193 3145 6227 3179
rect 7021 3145 7055 3179
rect 7757 3145 7791 3179
rect 8309 3145 8343 3179
rect 9873 3145 9907 3179
rect 10333 3145 10367 3179
rect 11345 3145 11379 3179
rect 11897 3145 11931 3179
rect 14657 3145 14691 3179
rect 16221 3145 16255 3179
rect 17417 3145 17451 3179
rect 18889 3145 18923 3179
rect 21373 3145 21407 3179
rect 21465 3145 21499 3179
rect 22017 3145 22051 3179
rect 22661 3145 22695 3179
rect 23397 3145 23431 3179
rect 24133 3145 24167 3179
rect 26801 3145 26835 3179
rect 28365 3145 28399 3179
rect 29101 3145 29135 3179
rect 30665 3145 30699 3179
rect 30941 3145 30975 3179
rect 31401 3145 31435 3179
rect 32321 3145 32355 3179
rect 35265 3145 35299 3179
rect 36185 3145 36219 3179
rect 38945 3145 38979 3179
rect 40601 3145 40635 3179
rect 43085 3145 43119 3179
rect 43913 3145 43947 3179
rect 46213 3145 46247 3179
rect 48237 3145 48271 3179
rect 56149 3145 56183 3179
rect 58541 3145 58575 3179
rect 10241 3077 10275 3111
rect 11989 3077 12023 3111
rect 13544 3077 13578 3111
rect 21925 3077 21959 3111
rect 26065 3077 26099 3111
rect 32689 3077 32723 3111
rect 33793 3077 33827 3111
rect 36553 3077 36587 3111
rect 46673 3077 46707 3111
rect 2881 3009 2915 3043
rect 3065 3009 3099 3043
rect 3525 3009 3559 3043
rect 3617 3009 3651 3043
rect 4721 3009 4755 3043
rect 5733 3009 5767 3043
rect 6009 3009 6043 3043
rect 8217 3009 8251 3043
rect 9321 3009 9355 3043
rect 9505 3009 9539 3043
rect 9597 3009 9631 3043
rect 13277 3009 13311 3043
rect 14749 3009 14783 3043
rect 16405 3009 16439 3043
rect 16865 3009 16899 3043
rect 17509 3009 17543 3043
rect 18061 3009 18095 3043
rect 19165 3009 19199 3043
rect 19441 3009 19475 3043
rect 20729 3009 20763 3043
rect 21649 3009 21683 3043
rect 23581 3009 23615 3043
rect 24225 3009 24259 3043
rect 25697 3009 25731 3043
rect 25881 3009 25915 3043
rect 27813 3009 27847 3043
rect 29377 3009 29411 3043
rect 30849 3009 30883 3043
rect 31309 3009 31343 3043
rect 31953 3009 31987 3043
rect 33885 3009 33919 3043
rect 34529 3009 34563 3043
rect 34621 3009 34655 3043
rect 36645 3009 36679 3043
rect 37565 3009 37599 3043
rect 39129 3009 39163 3043
rect 39313 3009 39347 3043
rect 40969 3009 41003 3043
rect 43361 3009 43395 3043
rect 44281 3009 44315 3043
rect 46397 3009 46431 3043
rect 46489 3009 46523 3043
rect 46765 3009 46799 3043
rect 46949 3009 46983 3043
rect 47133 3009 47167 3043
rect 47409 3009 47443 3043
rect 48329 3009 48363 3043
rect 48513 3009 48547 3043
rect 48973 3009 49007 3043
rect 49065 3009 49099 3043
rect 51641 3009 51675 3043
rect 52837 3009 52871 3043
rect 53665 3009 53699 3043
rect 53757 3009 53791 3043
rect 53941 3009 53975 3043
rect 54033 3009 54067 3043
rect 55505 3009 55539 3043
rect 56517 3009 56551 3043
rect 2237 2941 2271 2975
rect 3249 2941 3283 2975
rect 3893 2941 3927 2975
rect 4813 2941 4847 2975
rect 5549 2941 5583 2975
rect 6469 2941 6503 2975
rect 7205 2941 7239 2975
rect 8493 2941 8527 2975
rect 8769 2941 8803 2975
rect 10517 2941 10551 2975
rect 10793 2941 10827 2975
rect 12173 2941 12207 2975
rect 12633 2941 12667 2975
rect 15209 2941 15243 2975
rect 17601 2941 17635 2975
rect 18245 2941 18279 2975
rect 19717 2941 19751 2975
rect 22845 2941 22879 2975
rect 24685 2941 24719 2975
rect 26249 2941 26283 2975
rect 27077 2941 27111 2975
rect 28457 2941 28491 2975
rect 29653 2941 29687 2975
rect 31493 2941 31527 2975
rect 32781 2941 32815 2975
rect 32873 2941 32907 2975
rect 33149 2941 33183 2975
rect 35357 2941 35391 2975
rect 36737 2941 36771 2975
rect 37933 2941 37967 2975
rect 39865 2941 39899 2975
rect 39957 2941 39991 2975
rect 41245 2941 41279 2975
rect 42441 2941 42475 2975
rect 44557 2941 44591 2975
rect 45569 2941 45603 2975
rect 47593 2941 47627 2975
rect 48697 2941 48731 2975
rect 49525 2941 49559 2975
rect 50537 2941 50571 2975
rect 51457 2941 51491 2975
rect 51917 2941 51951 2975
rect 53389 2941 53423 2975
rect 54493 2941 54527 2975
rect 57253 2941 57287 2975
rect 57897 2941 57931 2975
rect 7849 2873 7883 2907
rect 11529 2873 11563 2907
rect 16681 2873 16715 2907
rect 17049 2873 17083 2907
rect 18981 2873 19015 2907
rect 27629 2873 27663 2907
rect 48789 2873 48823 2907
rect 5457 2805 5491 2839
rect 5917 2805 5951 2839
rect 9781 2805 9815 2839
rect 13185 2805 13219 2839
rect 17877 2805 17911 2839
rect 31769 2805 31803 2839
rect 36001 2805 36035 2839
rect 47225 2805 47259 2839
rect 51181 2805 51215 2839
rect 51825 2805 51859 2839
rect 52561 2805 52595 2839
rect 4169 2601 4203 2635
rect 4353 2601 4387 2635
rect 6377 2601 6411 2635
rect 7297 2601 7331 2635
rect 9781 2601 9815 2635
rect 13921 2601 13955 2635
rect 15025 2601 15059 2635
rect 17509 2601 17543 2635
rect 20177 2601 20211 2635
rect 22477 2601 22511 2635
rect 24041 2601 24075 2635
rect 24409 2601 24443 2635
rect 25329 2601 25363 2635
rect 27077 2601 27111 2635
rect 27445 2601 27479 2635
rect 29101 2601 29135 2635
rect 32229 2601 32263 2635
rect 34437 2601 34471 2635
rect 36921 2601 36955 2635
rect 39405 2601 39439 2635
rect 39497 2601 39531 2635
rect 42073 2601 42107 2635
rect 44649 2601 44683 2635
rect 45661 2601 45695 2635
rect 47225 2601 47259 2635
rect 49801 2601 49835 2635
rect 50261 2601 50295 2635
rect 52469 2601 52503 2635
rect 54493 2601 54527 2635
rect 58541 2601 58575 2635
rect 1961 2533 1995 2567
rect 3801 2533 3835 2567
rect 14105 2533 14139 2567
rect 19257 2533 19291 2567
rect 54953 2533 54987 2567
rect 2789 2465 2823 2499
rect 5549 2465 5583 2499
rect 6745 2465 6779 2499
rect 7849 2465 7883 2499
rect 10333 2465 10367 2499
rect 11621 2465 11655 2499
rect 12541 2465 12575 2499
rect 15853 2465 15887 2499
rect 18061 2465 18095 2499
rect 20821 2465 20855 2499
rect 23029 2465 23063 2499
rect 25881 2465 25915 2499
rect 27169 2465 27203 2499
rect 27997 2465 28031 2499
rect 30481 2465 30515 2499
rect 31033 2465 31067 2499
rect 32965 2465 32999 2499
rect 37749 2465 37783 2499
rect 38761 2465 38795 2499
rect 40325 2465 40359 2499
rect 42901 2465 42935 2499
rect 44097 2465 44131 2499
rect 46213 2465 46247 2499
rect 48053 2465 48087 2499
rect 51273 2465 51307 2499
rect 53205 2465 53239 2499
rect 56149 2465 56183 2499
rect 57897 2465 57931 2499
rect 2329 2397 2363 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 6561 2397 6595 2431
rect 7389 2397 7423 2431
rect 9229 2397 9263 2431
rect 9873 2397 9907 2431
rect 11805 2397 11839 2431
rect 11989 2397 12023 2431
rect 12081 2397 12115 2431
rect 13553 2397 13587 2431
rect 13737 2397 13771 2431
rect 14289 2397 14323 2431
rect 14473 2397 14507 2431
rect 15209 2397 15243 2431
rect 16957 2397 16991 2431
rect 17785 2397 17819 2431
rect 19441 2397 19475 2431
rect 19625 2397 19659 2431
rect 20269 2397 20303 2431
rect 21925 2397 21959 2431
rect 22569 2397 22603 2431
rect 24225 2397 24259 2431
rect 24593 2397 24627 2431
rect 24777 2397 24811 2431
rect 25421 2397 25455 2431
rect 27261 2397 27295 2431
rect 27721 2397 27755 2431
rect 29285 2397 29319 2431
rect 29745 2397 29779 2431
rect 29929 2397 29963 2431
rect 30665 2397 30699 2431
rect 32413 2397 32447 2431
rect 32597 2397 32631 2431
rect 34161 2397 34195 2431
rect 34897 2397 34931 2431
rect 36185 2397 36219 2431
rect 37105 2397 37139 2431
rect 37289 2397 37323 2431
rect 39681 2397 39715 2431
rect 39957 2397 39991 2431
rect 41337 2397 41371 2431
rect 41981 2397 42015 2431
rect 42257 2397 42291 2431
rect 42533 2397 42567 2431
rect 45017 2397 45051 2431
rect 45937 2397 45971 2431
rect 47409 2397 47443 2431
rect 47777 2397 47811 2431
rect 49065 2397 49099 2431
rect 49985 2397 50019 2431
rect 50445 2397 50479 2431
rect 50905 2397 50939 2431
rect 52285 2397 52319 2431
rect 52745 2397 52779 2431
rect 54769 2397 54803 2431
rect 55413 2397 55447 2431
rect 55873 2397 55907 2431
rect 57161 2397 57195 2431
rect 57345 2397 57379 2431
rect 1685 2329 1719 2363
rect 4169 2329 4203 2363
rect 26985 2329 27019 2363
rect 35633 2329 35667 2363
rect 57529 2329 57563 2363
rect 4537 2261 4571 2295
rect 29561 2261 29595 2295
rect 36829 2261 36863 2295
rect 49709 2261 49743 2295
rect 55597 2261 55631 2295
<< metal1 >>
rect 1104 27770 58880 27792
rect 1104 27718 8172 27770
rect 8224 27718 8236 27770
rect 8288 27718 8300 27770
rect 8352 27718 8364 27770
rect 8416 27718 8428 27770
rect 8480 27718 22616 27770
rect 22668 27718 22680 27770
rect 22732 27718 22744 27770
rect 22796 27718 22808 27770
rect 22860 27718 22872 27770
rect 22924 27718 37060 27770
rect 37112 27718 37124 27770
rect 37176 27718 37188 27770
rect 37240 27718 37252 27770
rect 37304 27718 37316 27770
rect 37368 27718 51504 27770
rect 51556 27718 51568 27770
rect 51620 27718 51632 27770
rect 51684 27718 51696 27770
rect 51748 27718 51760 27770
rect 51812 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 59040 27248
rect 1104 27174 15394 27226
rect 15446 27174 15458 27226
rect 15510 27174 15522 27226
rect 15574 27174 15586 27226
rect 15638 27174 15650 27226
rect 15702 27174 29838 27226
rect 29890 27174 29902 27226
rect 29954 27174 29966 27226
rect 30018 27174 30030 27226
rect 30082 27174 30094 27226
rect 30146 27174 44282 27226
rect 44334 27174 44346 27226
rect 44398 27174 44410 27226
rect 44462 27174 44474 27226
rect 44526 27174 44538 27226
rect 44590 27174 58726 27226
rect 58778 27174 58790 27226
rect 58842 27174 58854 27226
rect 58906 27174 58918 27226
rect 58970 27174 58982 27226
rect 59034 27174 59040 27226
rect 1104 27152 59040 27174
rect 1104 26682 58880 26704
rect 1104 26630 8172 26682
rect 8224 26630 8236 26682
rect 8288 26630 8300 26682
rect 8352 26630 8364 26682
rect 8416 26630 8428 26682
rect 8480 26630 22616 26682
rect 22668 26630 22680 26682
rect 22732 26630 22744 26682
rect 22796 26630 22808 26682
rect 22860 26630 22872 26682
rect 22924 26630 37060 26682
rect 37112 26630 37124 26682
rect 37176 26630 37188 26682
rect 37240 26630 37252 26682
rect 37304 26630 37316 26682
rect 37368 26630 51504 26682
rect 51556 26630 51568 26682
rect 51620 26630 51632 26682
rect 51684 26630 51696 26682
rect 51748 26630 51760 26682
rect 51812 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 59040 26160
rect 1104 26086 15394 26138
rect 15446 26086 15458 26138
rect 15510 26086 15522 26138
rect 15574 26086 15586 26138
rect 15638 26086 15650 26138
rect 15702 26086 29838 26138
rect 29890 26086 29902 26138
rect 29954 26086 29966 26138
rect 30018 26086 30030 26138
rect 30082 26086 30094 26138
rect 30146 26086 44282 26138
rect 44334 26086 44346 26138
rect 44398 26086 44410 26138
rect 44462 26086 44474 26138
rect 44526 26086 44538 26138
rect 44590 26086 58726 26138
rect 58778 26086 58790 26138
rect 58842 26086 58854 26138
rect 58906 26086 58918 26138
rect 58970 26086 58982 26138
rect 59034 26086 59040 26138
rect 1104 26064 59040 26086
rect 1104 25594 58880 25616
rect 1104 25542 8172 25594
rect 8224 25542 8236 25594
rect 8288 25542 8300 25594
rect 8352 25542 8364 25594
rect 8416 25542 8428 25594
rect 8480 25542 22616 25594
rect 22668 25542 22680 25594
rect 22732 25542 22744 25594
rect 22796 25542 22808 25594
rect 22860 25542 22872 25594
rect 22924 25542 37060 25594
rect 37112 25542 37124 25594
rect 37176 25542 37188 25594
rect 37240 25542 37252 25594
rect 37304 25542 37316 25594
rect 37368 25542 51504 25594
rect 51556 25542 51568 25594
rect 51620 25542 51632 25594
rect 51684 25542 51696 25594
rect 51748 25542 51760 25594
rect 51812 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 59040 25072
rect 1104 24998 15394 25050
rect 15446 24998 15458 25050
rect 15510 24998 15522 25050
rect 15574 24998 15586 25050
rect 15638 24998 15650 25050
rect 15702 24998 29838 25050
rect 29890 24998 29902 25050
rect 29954 24998 29966 25050
rect 30018 24998 30030 25050
rect 30082 24998 30094 25050
rect 30146 24998 44282 25050
rect 44334 24998 44346 25050
rect 44398 24998 44410 25050
rect 44462 24998 44474 25050
rect 44526 24998 44538 25050
rect 44590 24998 58726 25050
rect 58778 24998 58790 25050
rect 58842 24998 58854 25050
rect 58906 24998 58918 25050
rect 58970 24998 58982 25050
rect 59034 24998 59040 25050
rect 1104 24976 59040 24998
rect 1104 24506 58880 24528
rect 1104 24454 8172 24506
rect 8224 24454 8236 24506
rect 8288 24454 8300 24506
rect 8352 24454 8364 24506
rect 8416 24454 8428 24506
rect 8480 24454 22616 24506
rect 22668 24454 22680 24506
rect 22732 24454 22744 24506
rect 22796 24454 22808 24506
rect 22860 24454 22872 24506
rect 22924 24454 37060 24506
rect 37112 24454 37124 24506
rect 37176 24454 37188 24506
rect 37240 24454 37252 24506
rect 37304 24454 37316 24506
rect 37368 24454 51504 24506
rect 51556 24454 51568 24506
rect 51620 24454 51632 24506
rect 51684 24454 51696 24506
rect 51748 24454 51760 24506
rect 51812 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 59040 23984
rect 1104 23910 15394 23962
rect 15446 23910 15458 23962
rect 15510 23910 15522 23962
rect 15574 23910 15586 23962
rect 15638 23910 15650 23962
rect 15702 23910 29838 23962
rect 29890 23910 29902 23962
rect 29954 23910 29966 23962
rect 30018 23910 30030 23962
rect 30082 23910 30094 23962
rect 30146 23910 44282 23962
rect 44334 23910 44346 23962
rect 44398 23910 44410 23962
rect 44462 23910 44474 23962
rect 44526 23910 44538 23962
rect 44590 23910 58726 23962
rect 58778 23910 58790 23962
rect 58842 23910 58854 23962
rect 58906 23910 58918 23962
rect 58970 23910 58982 23962
rect 59034 23910 59040 23962
rect 1104 23888 59040 23910
rect 1104 23418 58880 23440
rect 1104 23366 8172 23418
rect 8224 23366 8236 23418
rect 8288 23366 8300 23418
rect 8352 23366 8364 23418
rect 8416 23366 8428 23418
rect 8480 23366 22616 23418
rect 22668 23366 22680 23418
rect 22732 23366 22744 23418
rect 22796 23366 22808 23418
rect 22860 23366 22872 23418
rect 22924 23366 37060 23418
rect 37112 23366 37124 23418
rect 37176 23366 37188 23418
rect 37240 23366 37252 23418
rect 37304 23366 37316 23418
rect 37368 23366 51504 23418
rect 51556 23366 51568 23418
rect 51620 23366 51632 23418
rect 51684 23366 51696 23418
rect 51748 23366 51760 23418
rect 51812 23366 58880 23418
rect 1104 23344 58880 23366
rect 38838 23060 38844 23112
rect 38896 23060 38902 23112
rect 47854 23060 47860 23112
rect 47912 23060 47918 23112
rect 39390 22924 39396 22976
rect 39448 22924 39454 22976
rect 40034 22924 40040 22976
rect 40092 22924 40098 22976
rect 48498 22924 48504 22976
rect 48556 22924 48562 22976
rect 1104 22874 59040 22896
rect 1104 22822 15394 22874
rect 15446 22822 15458 22874
rect 15510 22822 15522 22874
rect 15574 22822 15586 22874
rect 15638 22822 15650 22874
rect 15702 22822 29838 22874
rect 29890 22822 29902 22874
rect 29954 22822 29966 22874
rect 30018 22822 30030 22874
rect 30082 22822 30094 22874
rect 30146 22822 44282 22874
rect 44334 22822 44346 22874
rect 44398 22822 44410 22874
rect 44462 22822 44474 22874
rect 44526 22822 44538 22874
rect 44590 22822 58726 22874
rect 58778 22822 58790 22874
rect 58842 22822 58854 22874
rect 58906 22822 58918 22874
rect 58970 22822 58982 22874
rect 59034 22822 59040 22874
rect 1104 22800 59040 22822
rect 48498 22720 48504 22772
rect 48556 22720 48562 22772
rect 40034 22692 40040 22704
rect 38304 22664 40040 22692
rect 38304 22636 38332 22664
rect 40034 22652 40040 22664
rect 40092 22652 40098 22704
rect 47578 22652 47584 22704
rect 47636 22652 47642 22704
rect 47848 22695 47906 22701
rect 47848 22661 47860 22695
rect 47894 22692 47906 22695
rect 48516 22692 48544 22720
rect 47894 22664 48544 22692
rect 47894 22661 47906 22664
rect 47848 22655 47906 22661
rect 38286 22584 38292 22636
rect 38344 22584 38350 22636
rect 38556 22627 38614 22633
rect 38556 22593 38568 22627
rect 38602 22624 38614 22627
rect 39390 22624 39396 22636
rect 38602 22596 39396 22624
rect 38602 22593 38614 22596
rect 38556 22587 38614 22593
rect 39390 22584 39396 22596
rect 39448 22584 39454 22636
rect 47596 22624 47624 22652
rect 49053 22627 49111 22633
rect 49053 22624 49065 22627
rect 47596 22596 49065 22624
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 39761 22559 39819 22565
rect 39761 22556 39773 22559
rect 39684 22528 39773 22556
rect 24302 22380 24308 22432
rect 24360 22380 24366 22432
rect 24670 22380 24676 22432
rect 24728 22380 24734 22432
rect 25406 22380 25412 22432
rect 25464 22380 25470 22432
rect 37918 22380 37924 22432
rect 37976 22420 37982 22432
rect 38197 22423 38255 22429
rect 38197 22420 38209 22423
rect 37976 22392 38209 22420
rect 37976 22380 37982 22392
rect 38197 22389 38209 22392
rect 38243 22420 38255 22423
rect 38562 22420 38568 22432
rect 38243 22392 38568 22420
rect 38243 22389 38255 22392
rect 38197 22383 38255 22389
rect 38562 22380 38568 22392
rect 38620 22380 38626 22432
rect 38654 22380 38660 22432
rect 38712 22420 38718 22432
rect 39684 22429 39712 22528
rect 39761 22525 39773 22528
rect 39807 22525 39819 22559
rect 39761 22519 39819 22525
rect 47581 22559 47639 22565
rect 47581 22525 47593 22559
rect 47627 22525 47639 22559
rect 47581 22519 47639 22525
rect 39669 22423 39727 22429
rect 39669 22420 39681 22423
rect 38712 22392 39681 22420
rect 38712 22380 38718 22392
rect 39669 22389 39681 22392
rect 39715 22389 39727 22423
rect 39669 22383 39727 22389
rect 40402 22380 40408 22432
rect 40460 22380 40466 22432
rect 47397 22423 47455 22429
rect 47397 22389 47409 22423
rect 47443 22420 47455 22423
rect 47596 22420 47624 22519
rect 48976 22497 49004 22596
rect 49053 22593 49065 22596
rect 49099 22593 49111 22627
rect 49053 22587 49111 22593
rect 50706 22516 50712 22568
rect 50764 22516 50770 22568
rect 51350 22516 51356 22568
rect 51408 22516 51414 22568
rect 52914 22516 52920 22568
rect 52972 22516 52978 22568
rect 55033 22559 55091 22565
rect 55033 22525 55045 22559
rect 55079 22556 55091 22559
rect 55306 22556 55312 22568
rect 55079 22528 55312 22556
rect 55079 22525 55091 22528
rect 55033 22519 55091 22525
rect 55306 22516 55312 22528
rect 55364 22516 55370 22568
rect 55861 22559 55919 22565
rect 55861 22525 55873 22559
rect 55907 22556 55919 22559
rect 55950 22556 55956 22568
rect 55907 22528 55956 22556
rect 55907 22525 55919 22528
rect 55861 22519 55919 22525
rect 55950 22516 55956 22528
rect 56008 22516 56014 22568
rect 48961 22491 49019 22497
rect 48961 22457 48973 22491
rect 49007 22457 49019 22491
rect 48961 22451 49019 22457
rect 48498 22420 48504 22432
rect 47443 22392 48504 22420
rect 47443 22389 47455 22392
rect 47397 22383 47455 22389
rect 48498 22380 48504 22392
rect 48556 22380 48562 22432
rect 49694 22380 49700 22432
rect 49752 22380 49758 22432
rect 50798 22380 50804 22432
rect 50856 22420 50862 22432
rect 51261 22423 51319 22429
rect 51261 22420 51273 22423
rect 50856 22392 51273 22420
rect 50856 22380 50862 22392
rect 51261 22389 51273 22392
rect 51307 22389 51319 22423
rect 51261 22383 51319 22389
rect 51994 22380 52000 22432
rect 52052 22380 52058 22432
rect 52362 22380 52368 22432
rect 52420 22380 52426 22432
rect 53558 22380 53564 22432
rect 53616 22380 53622 22432
rect 54846 22380 54852 22432
rect 54904 22420 54910 22432
rect 55585 22423 55643 22429
rect 55585 22420 55597 22423
rect 54904 22392 55597 22420
rect 54904 22380 54910 22392
rect 55585 22389 55597 22392
rect 55631 22389 55643 22423
rect 55585 22383 55643 22389
rect 55766 22380 55772 22432
rect 55824 22420 55830 22432
rect 56413 22423 56471 22429
rect 56413 22420 56425 22423
rect 55824 22392 56425 22420
rect 55824 22380 55830 22392
rect 56413 22389 56425 22392
rect 56459 22389 56471 22423
rect 56413 22383 56471 22389
rect 56686 22380 56692 22432
rect 56744 22380 56750 22432
rect 1104 22330 58880 22352
rect 1104 22278 8172 22330
rect 8224 22278 8236 22330
rect 8288 22278 8300 22330
rect 8352 22278 8364 22330
rect 8416 22278 8428 22330
rect 8480 22278 22616 22330
rect 22668 22278 22680 22330
rect 22732 22278 22744 22330
rect 22796 22278 22808 22330
rect 22860 22278 22872 22330
rect 22924 22278 37060 22330
rect 37112 22278 37124 22330
rect 37176 22278 37188 22330
rect 37240 22278 37252 22330
rect 37304 22278 37316 22330
rect 37368 22278 51504 22330
rect 51556 22278 51568 22330
rect 51620 22278 51632 22330
rect 51684 22278 51696 22330
rect 51748 22278 51760 22330
rect 51812 22278 58880 22330
rect 1104 22256 58880 22278
rect 47765 22219 47823 22225
rect 47765 22185 47777 22219
rect 47811 22216 47823 22219
rect 47854 22216 47860 22228
rect 47811 22188 47860 22216
rect 47811 22185 47823 22188
rect 47765 22179 47823 22185
rect 47854 22176 47860 22188
rect 47912 22176 47918 22228
rect 55306 22176 55312 22228
rect 55364 22176 55370 22228
rect 38562 22108 38568 22160
rect 38620 22148 38626 22160
rect 40770 22148 40776 22160
rect 38620 22120 40776 22148
rect 38620 22108 38626 22120
rect 24302 22040 24308 22092
rect 24360 22080 24366 22092
rect 39592 22089 39620 22120
rect 40770 22108 40776 22120
rect 40828 22108 40834 22160
rect 48222 22108 48228 22160
rect 48280 22108 48286 22160
rect 56505 22151 56563 22157
rect 56505 22117 56517 22151
rect 56551 22117 56563 22151
rect 56505 22111 56563 22117
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 24360 22052 24409 22080
rect 24360 22040 24366 22052
rect 24397 22049 24409 22052
rect 24443 22049 24455 22083
rect 24397 22043 24455 22049
rect 37461 22083 37519 22089
rect 37461 22049 37473 22083
rect 37507 22049 37519 22083
rect 37461 22043 37519 22049
rect 39577 22083 39635 22089
rect 39577 22049 39589 22083
rect 39623 22080 39635 22083
rect 40497 22083 40555 22089
rect 40497 22080 40509 22083
rect 39623 22052 39657 22080
rect 39776 22052 40509 22080
rect 39623 22049 39635 22052
rect 39577 22043 39635 22049
rect 10502 21972 10508 22024
rect 10560 21972 10566 22024
rect 23658 21972 23664 22024
rect 23716 21972 23722 22024
rect 24664 22015 24722 22021
rect 24664 21981 24676 22015
rect 24710 22012 24722 22015
rect 25406 22012 25412 22024
rect 24710 21984 25412 22012
rect 24710 21981 24722 21984
rect 24664 21975 24722 21981
rect 25406 21972 25412 21984
rect 25464 21972 25470 22024
rect 25869 22015 25927 22021
rect 25869 22012 25881 22015
rect 25792 21984 25881 22012
rect 14826 21944 14832 21956
rect 12406 21916 14832 21944
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 6365 21879 6423 21885
rect 6365 21876 6377 21879
rect 5408 21848 6377 21876
rect 5408 21836 5414 21848
rect 6365 21845 6377 21848
rect 6411 21876 6423 21879
rect 7558 21876 7564 21888
rect 6411 21848 7564 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 11330 21836 11336 21888
rect 11388 21876 11394 21888
rect 12406 21876 12434 21916
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 11388 21848 12434 21876
rect 11388 21836 11394 21848
rect 23014 21836 23020 21888
rect 23072 21836 23078 21888
rect 24210 21836 24216 21888
rect 24268 21836 24274 21888
rect 24394 21836 24400 21888
rect 24452 21876 24458 21888
rect 25792 21885 25820 21984
rect 25869 21981 25881 21984
rect 25915 21981 25927 22015
rect 37476 22012 37504 22043
rect 38286 22012 38292 22024
rect 37476 21984 38292 22012
rect 25869 21975 25927 21981
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 39776 22012 39804 22052
rect 40497 22049 40509 22052
rect 40543 22049 40555 22083
rect 40497 22043 40555 22049
rect 47673 22083 47731 22089
rect 47673 22049 47685 22083
rect 47719 22080 47731 22083
rect 48240 22080 48268 22108
rect 48317 22083 48375 22089
rect 48317 22080 48329 22083
rect 47719 22052 48329 22080
rect 47719 22049 47731 22052
rect 47673 22043 47731 22049
rect 48317 22049 48329 22052
rect 48363 22049 48375 22083
rect 49694 22080 49700 22092
rect 48317 22043 48375 22049
rect 48424 22052 49700 22080
rect 38856 21984 39804 22012
rect 39853 22015 39911 22021
rect 37728 21947 37786 21953
rect 37728 21913 37740 21947
rect 37774 21944 37786 21947
rect 38856 21944 38884 21984
rect 39853 21981 39865 22015
rect 39899 21981 39911 22015
rect 39853 21975 39911 21981
rect 48225 22015 48283 22021
rect 48225 21981 48237 22015
rect 48271 22012 48283 22015
rect 48424 22012 48452 22052
rect 49694 22040 49700 22052
rect 49752 22040 49758 22092
rect 55766 22040 55772 22092
rect 55824 22040 55830 22092
rect 55858 22040 55864 22092
rect 55916 22080 55922 22092
rect 55953 22083 56011 22089
rect 55953 22080 55965 22083
rect 55916 22052 55965 22080
rect 55916 22040 55922 22052
rect 55953 22049 55965 22052
rect 55999 22080 56011 22083
rect 56321 22083 56379 22089
rect 56321 22080 56333 22083
rect 55999 22052 56333 22080
rect 55999 22049 56011 22052
rect 55953 22043 56011 22049
rect 56321 22049 56333 22052
rect 56367 22049 56379 22083
rect 56321 22043 56379 22049
rect 48271 21984 48452 22012
rect 48271 21981 48283 21984
rect 48225 21975 48283 21981
rect 39868 21944 39896 21975
rect 48498 21972 48504 22024
rect 48556 22012 48562 22024
rect 49973 22015 50031 22021
rect 49973 22012 49985 22015
rect 48556 21984 49985 22012
rect 48556 21972 48562 21984
rect 49973 21981 49985 21984
rect 50019 22012 50031 22015
rect 50157 22015 50215 22021
rect 50157 22012 50169 22015
rect 50019 21984 50169 22012
rect 50019 21981 50031 21984
rect 49973 21975 50031 21981
rect 50157 21981 50169 21984
rect 50203 22012 50215 22015
rect 51629 22015 51687 22021
rect 51629 22012 51641 22015
rect 50203 21984 51641 22012
rect 50203 21981 50215 21984
rect 50157 21975 50215 21981
rect 51629 21981 51641 21984
rect 51675 22012 51687 22015
rect 52362 22012 52368 22024
rect 51675 21984 52368 22012
rect 51675 21981 51687 21984
rect 51629 21975 51687 21981
rect 52362 21972 52368 21984
rect 52420 21972 52426 22024
rect 52454 21972 52460 22024
rect 52512 22012 52518 22024
rect 53101 22015 53159 22021
rect 53101 22012 53113 22015
rect 52512 21984 53113 22012
rect 52512 21972 52518 21984
rect 53101 21981 53113 21984
rect 53147 21981 53159 22015
rect 53101 21975 53159 21981
rect 53837 22015 53895 22021
rect 53837 21981 53849 22015
rect 53883 21981 53895 22015
rect 56520 22012 56548 22111
rect 56686 22108 56692 22160
rect 56744 22148 56750 22160
rect 56744 22120 57100 22148
rect 56744 22108 56750 22120
rect 57072 22094 57100 22120
rect 57072 22089 57137 22094
rect 57057 22083 57137 22089
rect 57057 22049 57069 22083
rect 57103 22066 57137 22083
rect 57333 22083 57391 22089
rect 57103 22049 57115 22066
rect 57057 22043 57115 22049
rect 57333 22049 57345 22083
rect 57379 22049 57391 22083
rect 57333 22043 57391 22049
rect 57348 22012 57376 22043
rect 56520 21984 57376 22012
rect 53837 21975 53895 21981
rect 37774 21916 38884 21944
rect 38948 21916 39896 21944
rect 50424 21947 50482 21953
rect 37774 21913 37786 21916
rect 37728 21907 37786 21913
rect 25777 21879 25835 21885
rect 25777 21876 25789 21879
rect 24452 21848 25789 21876
rect 24452 21836 24458 21848
rect 25777 21845 25789 21848
rect 25823 21845 25835 21879
rect 25777 21839 25835 21845
rect 26510 21836 26516 21888
rect 26568 21836 26574 21888
rect 38746 21836 38752 21888
rect 38804 21876 38810 21888
rect 38948 21885 38976 21916
rect 50424 21913 50436 21947
rect 50470 21944 50482 21947
rect 50798 21944 50804 21956
rect 50470 21916 50804 21944
rect 50470 21913 50482 21916
rect 50424 21907 50482 21913
rect 50798 21904 50804 21916
rect 50856 21904 50862 21956
rect 51896 21947 51954 21953
rect 51896 21913 51908 21947
rect 51942 21944 51954 21947
rect 53745 21947 53803 21953
rect 53745 21944 53757 21947
rect 51942 21916 53757 21944
rect 51942 21913 51954 21916
rect 51896 21907 51954 21913
rect 53745 21913 53757 21916
rect 53791 21913 53803 21947
rect 53745 21907 53803 21913
rect 38841 21879 38899 21885
rect 38841 21876 38853 21879
rect 38804 21848 38853 21876
rect 38804 21836 38810 21848
rect 38841 21845 38853 21848
rect 38887 21845 38899 21879
rect 38841 21839 38899 21845
rect 38933 21879 38991 21885
rect 38933 21845 38945 21879
rect 38979 21845 38991 21879
rect 38933 21839 38991 21845
rect 39206 21836 39212 21888
rect 39264 21876 39270 21888
rect 39301 21879 39359 21885
rect 39301 21876 39313 21879
rect 39264 21848 39313 21876
rect 39264 21836 39270 21848
rect 39301 21845 39313 21848
rect 39347 21845 39359 21879
rect 39301 21839 39359 21845
rect 39390 21836 39396 21888
rect 39448 21836 39454 21888
rect 47302 21836 47308 21888
rect 47360 21876 47366 21888
rect 48133 21879 48191 21885
rect 48133 21876 48145 21879
rect 47360 21848 48145 21876
rect 47360 21836 47366 21848
rect 48133 21845 48145 21848
rect 48179 21845 48191 21879
rect 48133 21839 48191 21845
rect 51350 21836 51356 21888
rect 51408 21876 51414 21888
rect 51537 21879 51595 21885
rect 51537 21876 51549 21879
rect 51408 21848 51549 21876
rect 51408 21836 51414 21848
rect 51537 21845 51549 21848
rect 51583 21876 51595 21879
rect 52178 21876 52184 21888
rect 51583 21848 52184 21876
rect 51583 21845 51595 21848
rect 51537 21839 51595 21845
rect 52178 21836 52184 21848
rect 52236 21836 52242 21888
rect 52730 21836 52736 21888
rect 52788 21876 52794 21888
rect 53009 21879 53067 21885
rect 53009 21876 53021 21879
rect 52788 21848 53021 21876
rect 52788 21836 52794 21848
rect 53009 21845 53021 21848
rect 53055 21876 53067 21879
rect 53852 21876 53880 21975
rect 56965 21947 57023 21953
rect 56965 21913 56977 21947
rect 57011 21944 57023 21947
rect 58526 21944 58532 21956
rect 57011 21916 58532 21944
rect 57011 21913 57023 21916
rect 56965 21907 57023 21913
rect 58526 21904 58532 21916
rect 58584 21904 58590 21956
rect 53055 21848 53880 21876
rect 53055 21845 53067 21848
rect 53009 21839 53067 21845
rect 54478 21836 54484 21888
rect 54536 21836 54542 21888
rect 54754 21836 54760 21888
rect 54812 21836 54818 21888
rect 55677 21879 55735 21885
rect 55677 21845 55689 21879
rect 55723 21876 55735 21879
rect 56873 21879 56931 21885
rect 56873 21876 56885 21879
rect 55723 21848 56885 21876
rect 55723 21845 55735 21848
rect 55677 21839 55735 21845
rect 56873 21845 56885 21848
rect 56919 21876 56931 21879
rect 57790 21876 57796 21888
rect 56919 21848 57796 21876
rect 56919 21845 56931 21848
rect 56873 21839 56931 21845
rect 57790 21836 57796 21848
rect 57848 21836 57854 21888
rect 57974 21836 57980 21888
rect 58032 21836 58038 21888
rect 1104 21786 59040 21808
rect 1104 21734 15394 21786
rect 15446 21734 15458 21786
rect 15510 21734 15522 21786
rect 15574 21734 15586 21786
rect 15638 21734 15650 21786
rect 15702 21734 29838 21786
rect 29890 21734 29902 21786
rect 29954 21734 29966 21786
rect 30018 21734 30030 21786
rect 30082 21734 30094 21786
rect 30146 21734 44282 21786
rect 44334 21734 44346 21786
rect 44398 21734 44410 21786
rect 44462 21734 44474 21786
rect 44526 21734 44538 21786
rect 44590 21734 58726 21786
rect 58778 21734 58790 21786
rect 58842 21734 58854 21786
rect 58906 21734 58918 21786
rect 58970 21734 58982 21786
rect 59034 21734 59040 21786
rect 1104 21712 59040 21734
rect 4430 21632 4436 21684
rect 4488 21672 4494 21684
rect 5810 21672 5816 21684
rect 4488 21644 5816 21672
rect 4488 21632 4494 21644
rect 5810 21632 5816 21644
rect 5868 21672 5874 21684
rect 9858 21672 9864 21684
rect 5868 21644 9864 21672
rect 5868 21632 5874 21644
rect 9858 21632 9864 21644
rect 9916 21632 9922 21684
rect 10502 21632 10508 21684
rect 10560 21632 10566 21684
rect 10965 21675 11023 21681
rect 10965 21641 10977 21675
rect 11011 21672 11023 21675
rect 12161 21675 12219 21681
rect 12161 21672 12173 21675
rect 11011 21644 12173 21672
rect 11011 21641 11023 21644
rect 10965 21635 11023 21641
rect 12161 21641 12173 21644
rect 12207 21641 12219 21675
rect 12161 21635 12219 21641
rect 23569 21675 23627 21681
rect 23569 21641 23581 21675
rect 23615 21672 23627 21675
rect 24210 21672 24216 21684
rect 23615 21644 24216 21672
rect 23615 21641 23627 21644
rect 23569 21635 23627 21641
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 24762 21632 24768 21684
rect 24820 21632 24826 21684
rect 25225 21675 25283 21681
rect 25225 21641 25237 21675
rect 25271 21672 25283 21675
rect 26510 21672 26516 21684
rect 25271 21644 26516 21672
rect 25271 21641 25283 21644
rect 25225 21635 25283 21641
rect 26510 21632 26516 21644
rect 26568 21632 26574 21684
rect 38838 21632 38844 21684
rect 38896 21632 38902 21684
rect 39390 21632 39396 21684
rect 39448 21672 39454 21684
rect 40313 21675 40371 21681
rect 40313 21672 40325 21675
rect 39448 21644 40325 21672
rect 39448 21632 39454 21644
rect 40313 21641 40325 21644
rect 40359 21641 40371 21675
rect 40313 21635 40371 21641
rect 40402 21632 40408 21684
rect 40460 21632 40466 21684
rect 50706 21632 50712 21684
rect 50764 21632 50770 21684
rect 51169 21675 51227 21681
rect 51169 21641 51181 21675
rect 51215 21672 51227 21675
rect 51994 21672 52000 21684
rect 51215 21644 52000 21672
rect 51215 21641 51227 21644
rect 51169 21635 51227 21641
rect 51994 21632 52000 21644
rect 52052 21632 52058 21684
rect 52089 21675 52147 21681
rect 52089 21641 52101 21675
rect 52135 21672 52147 21675
rect 54478 21672 54484 21684
rect 52135 21644 54484 21672
rect 52135 21641 52147 21644
rect 52089 21635 52147 21641
rect 54478 21632 54484 21644
rect 54536 21632 54542 21684
rect 54754 21632 54760 21684
rect 54812 21632 54818 21684
rect 55677 21675 55735 21681
rect 55677 21641 55689 21675
rect 55723 21672 55735 21675
rect 55950 21672 55956 21684
rect 55723 21644 55956 21672
rect 55723 21641 55735 21644
rect 55677 21635 55735 21641
rect 55950 21632 55956 21644
rect 56008 21672 56014 21684
rect 56502 21672 56508 21684
rect 56008 21644 56508 21672
rect 56008 21632 56014 21644
rect 56502 21632 56508 21644
rect 56560 21632 56566 21684
rect 57974 21632 57980 21684
rect 58032 21632 58038 21684
rect 58526 21632 58532 21684
rect 58584 21632 58590 21684
rect 11330 21604 11336 21616
rect 7852 21576 11336 21604
rect 6457 21539 6515 21545
rect 6457 21536 6469 21539
rect 5460 21508 6469 21536
rect 5460 21480 5488 21508
rect 6457 21505 6469 21508
rect 6503 21505 6515 21539
rect 6457 21499 6515 21505
rect 7852 21480 7880 21576
rect 8754 21496 8760 21548
rect 8812 21536 8818 21548
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 8812 21508 9229 21536
rect 8812 21496 8818 21508
rect 9217 21505 9229 21508
rect 9263 21536 9275 21539
rect 10410 21536 10416 21548
rect 9263 21508 10416 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 10873 21539 10931 21545
rect 10873 21505 10885 21539
rect 10919 21505 10931 21539
rect 10873 21499 10931 21505
rect 3142 21428 3148 21480
rect 3200 21428 3206 21480
rect 4062 21428 4068 21480
rect 4120 21468 4126 21480
rect 5350 21468 5356 21480
rect 4120 21440 5356 21468
rect 4120 21428 4126 21440
rect 5350 21428 5356 21440
rect 5408 21428 5414 21480
rect 5442 21428 5448 21480
rect 5500 21428 5506 21480
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21468 5687 21471
rect 6270 21468 6276 21480
rect 5675 21440 6276 21468
rect 5675 21437 5687 21440
rect 5629 21431 5687 21437
rect 6270 21428 6276 21440
rect 6328 21428 6334 21480
rect 7469 21471 7527 21477
rect 7469 21437 7481 21471
rect 7515 21468 7527 21471
rect 7834 21468 7840 21480
rect 7515 21440 7840 21468
rect 7515 21437 7527 21440
rect 7469 21431 7527 21437
rect 7834 21428 7840 21440
rect 7892 21428 7898 21480
rect 8389 21471 8447 21477
rect 8389 21437 8401 21471
rect 8435 21468 8447 21471
rect 8662 21468 8668 21480
rect 8435 21440 8668 21468
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 8662 21428 8668 21440
rect 8720 21428 8726 21480
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 10888 21468 10916 21499
rect 9456 21440 10916 21468
rect 9456 21428 9462 21440
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 11072 21477 11100 21576
rect 11330 21564 11336 21576
rect 11388 21564 11394 21616
rect 18966 21564 18972 21616
rect 19024 21604 19030 21616
rect 23014 21604 23020 21616
rect 19024 21576 23020 21604
rect 19024 21564 19030 21576
rect 23014 21564 23020 21576
rect 23072 21604 23078 21616
rect 27890 21604 27896 21616
rect 23072 21576 27896 21604
rect 23072 21564 23078 21576
rect 23477 21539 23535 21545
rect 23477 21505 23489 21539
rect 23523 21505 23535 21539
rect 23477 21499 23535 21505
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 7558 21360 7564 21412
rect 7616 21400 7622 21412
rect 8205 21403 8263 21409
rect 8205 21400 8217 21403
rect 7616 21372 8217 21400
rect 7616 21360 7622 21372
rect 8205 21369 8217 21372
rect 8251 21400 8263 21403
rect 10980 21400 11008 21428
rect 11532 21400 11560 21431
rect 13906 21428 13912 21480
rect 13964 21428 13970 21480
rect 15194 21428 15200 21480
rect 15252 21428 15258 21480
rect 18690 21428 18696 21480
rect 18748 21428 18754 21480
rect 22465 21471 22523 21477
rect 22465 21437 22477 21471
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 13725 21403 13783 21409
rect 13725 21400 13737 21403
rect 8251 21372 9720 21400
rect 10980 21372 11560 21400
rect 12406 21372 13737 21400
rect 8251 21369 8263 21372
rect 8205 21363 8263 21369
rect 9692 21344 9720 21372
rect 3694 21292 3700 21344
rect 3752 21292 3758 21344
rect 6178 21292 6184 21344
rect 6236 21292 6242 21344
rect 7098 21292 7104 21344
rect 7156 21292 7162 21344
rect 8938 21292 8944 21344
rect 8996 21292 9002 21344
rect 9674 21292 9680 21344
rect 9732 21292 9738 21344
rect 9766 21292 9772 21344
rect 9824 21292 9830 21344
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 10137 21335 10195 21341
rect 10137 21332 10149 21335
rect 9916 21304 10149 21332
rect 9916 21292 9922 21304
rect 10137 21301 10149 21304
rect 10183 21332 10195 21335
rect 12406 21332 12434 21372
rect 13725 21369 13737 21372
rect 13771 21400 13783 21403
rect 14734 21400 14740 21412
rect 13771 21372 14740 21400
rect 13771 21369 13783 21372
rect 13725 21363 13783 21369
rect 14734 21360 14740 21372
rect 14792 21360 14798 21412
rect 22480 21400 22508 21431
rect 23109 21403 23167 21409
rect 23109 21400 23121 21403
rect 22480 21372 23121 21400
rect 23109 21369 23121 21372
rect 23155 21369 23167 21403
rect 23109 21363 23167 21369
rect 10183 21304 12434 21332
rect 10183 21301 10195 21304
rect 10137 21295 10195 21301
rect 14458 21292 14464 21344
rect 14516 21292 14522 21344
rect 14642 21292 14648 21344
rect 14700 21332 14706 21344
rect 15013 21335 15071 21341
rect 15013 21332 15025 21335
rect 14700 21304 15025 21332
rect 14700 21292 14706 21304
rect 15013 21301 15025 21304
rect 15059 21301 15071 21335
rect 15013 21295 15071 21301
rect 15838 21292 15844 21344
rect 15896 21292 15902 21344
rect 19334 21292 19340 21344
rect 19392 21292 19398 21344
rect 19610 21292 19616 21344
rect 19668 21292 19674 21344
rect 23014 21292 23020 21344
rect 23072 21292 23078 21344
rect 23492 21332 23520 21499
rect 23753 21471 23811 21477
rect 23753 21437 23765 21471
rect 23799 21468 23811 21471
rect 23860 21468 23888 21576
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 39301 21607 39359 21613
rect 39301 21573 39313 21607
rect 39347 21604 39359 21607
rect 40420 21604 40448 21632
rect 39347 21576 40448 21604
rect 39347 21573 39359 21576
rect 39301 21567 39359 21573
rect 52362 21564 52368 21616
rect 52420 21604 52426 21616
rect 54772 21604 54800 21632
rect 52420 21576 54800 21604
rect 52420 21564 52426 21576
rect 25133 21539 25191 21545
rect 25133 21536 25145 21539
rect 24044 21508 25145 21536
rect 23799 21440 23888 21468
rect 23799 21437 23811 21440
rect 23753 21431 23811 21437
rect 23934 21428 23940 21480
rect 23992 21428 23998 21480
rect 24044 21344 24072 21508
rect 25133 21505 25145 21508
rect 25179 21536 25191 21539
rect 26786 21536 26792 21548
rect 25179 21508 26792 21536
rect 25179 21505 25191 21508
rect 25133 21499 25191 21505
rect 26786 21496 26792 21508
rect 26844 21496 26850 21548
rect 38746 21496 38752 21548
rect 38804 21496 38810 21548
rect 38930 21496 38936 21548
rect 38988 21536 38994 21548
rect 39206 21536 39212 21548
rect 38988 21508 39212 21536
rect 38988 21496 38994 21508
rect 39206 21496 39212 21508
rect 39264 21496 39270 21548
rect 39669 21539 39727 21545
rect 39669 21536 39681 21539
rect 39316 21508 39681 21536
rect 24854 21428 24860 21480
rect 24912 21468 24918 21480
rect 25317 21471 25375 21477
rect 25317 21468 25329 21471
rect 24912 21440 25329 21468
rect 24912 21428 24918 21440
rect 25317 21437 25329 21440
rect 25363 21437 25375 21471
rect 25317 21431 25375 21437
rect 25332 21400 25360 21431
rect 26050 21428 26056 21480
rect 26108 21428 26114 21480
rect 30190 21428 30196 21480
rect 30248 21428 30254 21480
rect 38764 21468 38792 21496
rect 39316 21480 39344 21508
rect 39669 21505 39681 21508
rect 39715 21505 39727 21539
rect 39669 21499 39727 21505
rect 51077 21539 51135 21545
rect 51077 21505 51089 21539
rect 51123 21536 51135 21539
rect 51997 21539 52055 21545
rect 51997 21536 52009 21539
rect 51123 21508 52009 21536
rect 51123 21505 51135 21508
rect 51077 21499 51135 21505
rect 51997 21505 52009 21508
rect 52043 21536 52055 21539
rect 52086 21536 52092 21548
rect 52043 21508 52092 21536
rect 52043 21505 52055 21508
rect 51997 21499 52055 21505
rect 52086 21496 52092 21508
rect 52144 21496 52150 21548
rect 52454 21496 52460 21548
rect 52512 21496 52518 21548
rect 52748 21545 52776 21576
rect 52733 21539 52791 21545
rect 52733 21505 52745 21539
rect 52779 21505 52791 21539
rect 52733 21499 52791 21505
rect 53000 21539 53058 21545
rect 53000 21505 53012 21539
rect 53046 21536 53058 21539
rect 53558 21536 53564 21548
rect 53046 21508 53564 21536
rect 53046 21505 53058 21508
rect 53000 21499 53058 21505
rect 53558 21496 53564 21508
rect 53616 21496 53622 21548
rect 54312 21545 54340 21576
rect 54846 21564 54852 21616
rect 54904 21564 54910 21616
rect 56404 21607 56462 21613
rect 56404 21573 56416 21607
rect 56450 21604 56462 21607
rect 57992 21604 58020 21632
rect 56450 21576 58020 21604
rect 56450 21573 56462 21576
rect 56404 21567 56462 21573
rect 54297 21539 54355 21545
rect 54297 21505 54309 21539
rect 54343 21505 54355 21539
rect 54297 21499 54355 21505
rect 54564 21539 54622 21545
rect 54564 21505 54576 21539
rect 54610 21536 54622 21539
rect 54864 21536 54892 21564
rect 54610 21508 54892 21536
rect 54610 21505 54622 21508
rect 54564 21499 54622 21505
rect 56042 21496 56048 21548
rect 56100 21536 56106 21548
rect 56870 21536 56876 21548
rect 56100 21508 56876 21536
rect 56100 21496 56106 21508
rect 56870 21496 56876 21508
rect 56928 21496 56934 21548
rect 39298 21468 39304 21480
rect 38764 21440 39304 21468
rect 39298 21428 39304 21440
rect 39356 21428 39362 21480
rect 39393 21471 39451 21477
rect 39393 21437 39405 21471
rect 39439 21437 39451 21471
rect 39393 21431 39451 21437
rect 30006 21400 30012 21412
rect 25332 21372 30012 21400
rect 30006 21360 30012 21372
rect 30064 21360 30070 21412
rect 35342 21360 35348 21412
rect 35400 21400 35406 21412
rect 38105 21403 38163 21409
rect 38105 21400 38117 21403
rect 35400 21372 38117 21400
rect 35400 21360 35406 21372
rect 38105 21369 38117 21372
rect 38151 21400 38163 21403
rect 39022 21400 39028 21412
rect 38151 21372 39028 21400
rect 38151 21369 38163 21372
rect 38105 21363 38163 21369
rect 39022 21360 39028 21372
rect 39080 21360 39086 21412
rect 39408 21400 39436 21431
rect 42702 21428 42708 21480
rect 42760 21428 42766 21480
rect 46658 21428 46664 21480
rect 46716 21428 46722 21480
rect 50617 21471 50675 21477
rect 50617 21437 50629 21471
rect 50663 21468 50675 21471
rect 51350 21468 51356 21480
rect 50663 21440 51356 21468
rect 50663 21437 50675 21440
rect 50617 21431 50675 21437
rect 51350 21428 51356 21440
rect 51408 21428 51414 21480
rect 52270 21468 52276 21480
rect 51552 21440 52276 21468
rect 39224 21372 39436 21400
rect 39224 21344 39252 21372
rect 42242 21360 42248 21412
rect 42300 21400 42306 21412
rect 51552 21400 51580 21440
rect 52270 21428 52276 21440
rect 52328 21428 52334 21480
rect 42300 21372 43668 21400
rect 42300 21360 42306 21372
rect 24026 21332 24032 21344
rect 23492 21304 24032 21332
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24578 21292 24584 21344
rect 24636 21292 24642 21344
rect 25774 21292 25780 21344
rect 25832 21292 25838 21344
rect 26602 21292 26608 21344
rect 26660 21292 26666 21344
rect 30834 21292 30840 21344
rect 30892 21292 30898 21344
rect 38378 21292 38384 21344
rect 38436 21292 38442 21344
rect 39206 21292 39212 21344
rect 39264 21292 39270 21344
rect 41874 21292 41880 21344
rect 41932 21292 41938 21344
rect 43254 21292 43260 21344
rect 43312 21292 43318 21344
rect 43640 21341 43668 21372
rect 51046 21372 51580 21400
rect 51629 21403 51687 21409
rect 43625 21335 43683 21341
rect 43625 21301 43637 21335
rect 43671 21332 43683 21335
rect 43898 21332 43904 21344
rect 43671 21304 43904 21332
rect 43671 21301 43683 21304
rect 43625 21295 43683 21301
rect 43898 21292 43904 21304
rect 43956 21292 43962 21344
rect 45925 21335 45983 21341
rect 45925 21301 45937 21335
rect 45971 21332 45983 21335
rect 46106 21332 46112 21344
rect 45971 21304 46112 21332
rect 45971 21301 45983 21304
rect 45925 21295 45983 21301
rect 46106 21292 46112 21304
rect 46164 21292 46170 21344
rect 46474 21292 46480 21344
rect 46532 21292 46538 21344
rect 47210 21292 47216 21344
rect 47268 21292 47274 21344
rect 47854 21292 47860 21344
rect 47912 21292 47918 21344
rect 48222 21292 48228 21344
rect 48280 21332 48286 21344
rect 50157 21335 50215 21341
rect 50157 21332 50169 21335
rect 48280 21304 50169 21332
rect 48280 21292 48286 21304
rect 50157 21301 50169 21304
rect 50203 21332 50215 21335
rect 51046 21332 51074 21372
rect 51629 21369 51641 21403
rect 51675 21400 51687 21403
rect 52472 21400 52500 21496
rect 56137 21471 56195 21477
rect 56137 21437 56149 21471
rect 56183 21437 56195 21471
rect 56137 21431 56195 21437
rect 57885 21471 57943 21477
rect 57885 21437 57897 21471
rect 57931 21437 57943 21471
rect 57885 21431 57943 21437
rect 51675 21372 52500 21400
rect 51675 21369 51687 21372
rect 51629 21363 51687 21369
rect 50203 21304 51074 21332
rect 50203 21301 50215 21304
rect 50157 21295 50215 21301
rect 51258 21292 51264 21344
rect 51316 21332 51322 21344
rect 52638 21332 52644 21344
rect 51316 21304 52644 21332
rect 51316 21292 51322 21304
rect 52638 21292 52644 21304
rect 52696 21292 52702 21344
rect 53742 21292 53748 21344
rect 53800 21332 53806 21344
rect 54113 21335 54171 21341
rect 54113 21332 54125 21335
rect 53800 21304 54125 21332
rect 53800 21292 53806 21304
rect 54113 21301 54125 21304
rect 54159 21301 54171 21335
rect 56152 21332 56180 21431
rect 56502 21332 56508 21344
rect 56152 21304 56508 21332
rect 54113 21295 54171 21301
rect 56502 21292 56508 21304
rect 56560 21292 56566 21344
rect 57514 21292 57520 21344
rect 57572 21332 57578 21344
rect 57900 21332 57928 21431
rect 57572 21304 57928 21332
rect 57572 21292 57578 21304
rect 1104 21242 58880 21264
rect 1104 21190 8172 21242
rect 8224 21190 8236 21242
rect 8288 21190 8300 21242
rect 8352 21190 8364 21242
rect 8416 21190 8428 21242
rect 8480 21190 22616 21242
rect 22668 21190 22680 21242
rect 22732 21190 22744 21242
rect 22796 21190 22808 21242
rect 22860 21190 22872 21242
rect 22924 21190 37060 21242
rect 37112 21190 37124 21242
rect 37176 21190 37188 21242
rect 37240 21190 37252 21242
rect 37304 21190 37316 21242
rect 37368 21190 51504 21242
rect 51556 21190 51568 21242
rect 51620 21190 51632 21242
rect 51684 21190 51696 21242
rect 51748 21190 51760 21242
rect 51812 21190 58880 21242
rect 1104 21168 58880 21190
rect 4430 21088 4436 21140
rect 4488 21088 4494 21140
rect 6178 21088 6184 21140
rect 6236 21088 6242 21140
rect 6270 21088 6276 21140
rect 6328 21088 6334 21140
rect 7098 21088 7104 21140
rect 7156 21088 7162 21140
rect 7558 21128 7564 21140
rect 7392 21100 7564 21128
rect 2869 21063 2927 21069
rect 2869 21060 2881 21063
rect 2746 21032 2881 21060
rect 2225 20995 2283 21001
rect 2225 20961 2237 20995
rect 2271 20992 2283 20995
rect 2746 20992 2774 21032
rect 2869 21029 2881 21032
rect 2915 21029 2927 21063
rect 2869 21023 2927 21029
rect 2271 20964 2774 20992
rect 3513 20995 3571 21001
rect 2271 20961 2283 20964
rect 2225 20955 2283 20961
rect 3513 20961 3525 20995
rect 3559 20992 3571 20995
rect 4448 20992 4476 21088
rect 3559 20964 4476 20992
rect 3559 20961 3571 20964
rect 3513 20955 3571 20961
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 4801 20927 4859 20933
rect 4801 20893 4813 20927
rect 4847 20924 4859 20927
rect 5350 20924 5356 20936
rect 4847 20896 5356 20924
rect 4847 20893 4859 20896
rect 4801 20887 4859 20893
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 5068 20859 5126 20865
rect 4172 20828 5028 20856
rect 4172 20800 4200 20828
rect 2777 20791 2835 20797
rect 2777 20757 2789 20791
rect 2823 20788 2835 20791
rect 2866 20788 2872 20800
rect 2823 20760 2872 20788
rect 2823 20757 2835 20760
rect 2777 20751 2835 20757
rect 2866 20748 2872 20760
rect 2924 20748 2930 20800
rect 3234 20748 3240 20800
rect 3292 20748 3298 20800
rect 3326 20748 3332 20800
rect 3384 20748 3390 20800
rect 4154 20748 4160 20800
rect 4212 20748 4218 20800
rect 4522 20748 4528 20800
rect 4580 20748 4586 20800
rect 5000 20788 5028 20828
rect 5068 20825 5080 20859
rect 5114 20856 5126 20859
rect 6196 20856 6224 21088
rect 7116 21060 7144 21088
rect 6748 21032 7144 21060
rect 6748 21001 6776 21032
rect 7392 21001 7420 21100
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 8754 21088 8760 21140
rect 8812 21088 8818 21140
rect 8938 21088 8944 21140
rect 8996 21088 9002 21140
rect 9766 21128 9772 21140
rect 9416 21100 9772 21128
rect 6733 20995 6791 21001
rect 6733 20961 6745 20995
rect 6779 20961 6791 20995
rect 6733 20955 6791 20961
rect 6917 20995 6975 21001
rect 6917 20961 6929 20995
rect 6963 20992 6975 20995
rect 7377 20995 7435 21001
rect 6963 20964 7328 20992
rect 6963 20961 6975 20964
rect 6917 20955 6975 20961
rect 5114 20828 6224 20856
rect 7300 20856 7328 20964
rect 7377 20961 7389 20995
rect 7423 20961 7435 20995
rect 7377 20955 7435 20961
rect 7644 20927 7702 20933
rect 7644 20893 7656 20927
rect 7690 20924 7702 20927
rect 8956 20924 8984 21088
rect 9416 21001 9444 21100
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 9858 21088 9864 21140
rect 9916 21088 9922 21140
rect 14458 21088 14464 21140
rect 14516 21088 14522 21140
rect 14826 21088 14832 21140
rect 14884 21088 14890 21140
rect 15013 21131 15071 21137
rect 15013 21097 15025 21131
rect 15059 21128 15071 21131
rect 15194 21128 15200 21140
rect 15059 21100 15200 21128
rect 15059 21097 15071 21100
rect 15013 21091 15071 21097
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 22373 21131 22431 21137
rect 22373 21097 22385 21131
rect 22419 21128 22431 21131
rect 24302 21128 24308 21140
rect 22419 21100 24308 21128
rect 22419 21097 22431 21100
rect 22373 21091 22431 21097
rect 9401 20995 9459 21001
rect 9401 20961 9413 20995
rect 9447 20961 9459 20995
rect 9401 20955 9459 20961
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20992 9643 20995
rect 9876 20992 9904 21088
rect 14093 21063 14151 21069
rect 14093 21029 14105 21063
rect 14139 21029 14151 21063
rect 14093 21023 14151 21029
rect 9631 20964 9904 20992
rect 13173 20995 13231 21001
rect 9631 20961 9643 20964
rect 9585 20955 9643 20961
rect 13173 20961 13185 20995
rect 13219 20992 13231 20995
rect 14108 20992 14136 21023
rect 13219 20964 14136 20992
rect 14476 20992 14504 21088
rect 14553 20995 14611 21001
rect 14553 20992 14565 20995
rect 14476 20964 14565 20992
rect 13219 20961 13231 20964
rect 13173 20955 13231 20961
rect 14553 20961 14565 20964
rect 14599 20961 14611 20995
rect 14553 20955 14611 20961
rect 14734 20952 14740 21004
rect 14792 20952 14798 21004
rect 14844 20992 14872 21088
rect 15565 20995 15623 21001
rect 15565 20992 15577 20995
rect 14844 20964 15577 20992
rect 15565 20961 15577 20964
rect 15611 20961 15623 20995
rect 15565 20955 15623 20961
rect 15672 20964 18000 20992
rect 7690 20896 8984 20924
rect 7690 20893 7702 20896
rect 7644 20887 7702 20893
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 10045 20927 10103 20933
rect 10045 20924 10057 20927
rect 9732 20896 10057 20924
rect 9732 20884 9738 20896
rect 10045 20893 10057 20896
rect 10091 20924 10103 20927
rect 14752 20924 14780 20952
rect 15672 20924 15700 20964
rect 10091 20896 11836 20924
rect 14752 20896 15700 20924
rect 16025 20927 16083 20933
rect 10091 20893 10103 20896
rect 10045 20887 10103 20893
rect 7834 20856 7840 20868
rect 7300 20828 7840 20856
rect 5114 20825 5126 20828
rect 5068 20819 5126 20825
rect 7834 20816 7840 20828
rect 7892 20816 7898 20868
rect 8662 20816 8668 20868
rect 8720 20856 8726 20868
rect 10312 20859 10370 20865
rect 8720 20828 8984 20856
rect 8720 20816 8726 20828
rect 5442 20788 5448 20800
rect 5000 20760 5448 20788
rect 5442 20748 5448 20760
rect 5500 20788 5506 20800
rect 6181 20791 6239 20797
rect 6181 20788 6193 20791
rect 5500 20760 6193 20788
rect 5500 20748 5506 20760
rect 6181 20757 6193 20760
rect 6227 20757 6239 20791
rect 6181 20751 6239 20757
rect 6638 20748 6644 20800
rect 6696 20748 6702 20800
rect 8956 20797 8984 20828
rect 10312 20825 10324 20859
rect 10358 20856 10370 20859
rect 11054 20856 11060 20868
rect 10358 20828 11060 20856
rect 10358 20825 10370 20828
rect 10312 20819 10370 20825
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 11808 20865 11836 20896
rect 16025 20893 16037 20927
rect 16071 20924 16083 20927
rect 16482 20924 16488 20936
rect 16071 20896 16488 20924
rect 16071 20893 16083 20896
rect 16025 20887 16083 20893
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 16666 20884 16672 20936
rect 16724 20884 16730 20936
rect 17972 20865 18000 20964
rect 22186 20952 22192 21004
rect 22244 20992 22250 21004
rect 22480 21001 22508 21100
rect 24302 21088 24308 21100
rect 24360 21088 24366 21140
rect 25314 21128 25320 21140
rect 24504 21100 25320 21128
rect 23658 21020 23664 21072
rect 23716 21060 23722 21072
rect 23845 21063 23903 21069
rect 23845 21060 23857 21063
rect 23716 21032 23857 21060
rect 23716 21020 23722 21032
rect 23845 21029 23857 21032
rect 23891 21060 23903 21063
rect 24504 21060 24532 21100
rect 25314 21088 25320 21100
rect 25372 21088 25378 21140
rect 25774 21088 25780 21140
rect 25832 21128 25838 21140
rect 25832 21100 26004 21128
rect 25832 21088 25838 21100
rect 25976 21060 26004 21100
rect 26050 21088 26056 21140
rect 26108 21128 26114 21140
rect 26329 21131 26387 21137
rect 26329 21128 26341 21131
rect 26108 21100 26341 21128
rect 26108 21088 26114 21100
rect 26329 21097 26341 21100
rect 26375 21097 26387 21131
rect 26329 21091 26387 21097
rect 30006 21088 30012 21140
rect 30064 21088 30070 21140
rect 30190 21088 30196 21140
rect 30248 21088 30254 21140
rect 38378 21128 38384 21140
rect 31726 21100 38384 21128
rect 23891 21032 24532 21060
rect 24596 21032 25176 21060
rect 25976 21032 26924 21060
rect 23891 21029 23903 21032
rect 23845 21023 23903 21029
rect 22465 20995 22523 21001
rect 22465 20992 22477 20995
rect 22244 20964 22477 20992
rect 22244 20952 22250 20964
rect 22465 20961 22477 20964
rect 22511 20961 22523 20995
rect 22465 20955 22523 20961
rect 24394 20952 24400 21004
rect 24452 20952 24458 21004
rect 24596 21001 24624 21032
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20961 24639 20995
rect 24581 20955 24639 20961
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 25004 20964 25053 20992
rect 25004 20952 25010 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25148 20992 25176 21032
rect 26694 20992 26700 21004
rect 25148 20964 26700 20992
rect 25041 20955 25099 20961
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 26786 20952 26792 21004
rect 26844 20952 26850 21004
rect 26896 21001 26924 21032
rect 26881 20995 26939 21001
rect 26881 20961 26893 20995
rect 26927 20961 26939 20995
rect 30024 20992 30052 21088
rect 31726 21072 31754 21100
rect 38378 21088 38384 21100
rect 38436 21128 38442 21140
rect 39482 21128 39488 21140
rect 38436 21100 39488 21128
rect 38436 21088 38442 21100
rect 39482 21088 39488 21100
rect 39540 21088 39546 21140
rect 39577 21131 39635 21137
rect 39577 21097 39589 21131
rect 39623 21128 39635 21131
rect 39942 21128 39948 21140
rect 39623 21100 39948 21128
rect 39623 21097 39635 21100
rect 39577 21091 39635 21097
rect 39942 21088 39948 21100
rect 40000 21088 40006 21140
rect 41414 21088 41420 21140
rect 41472 21128 41478 21140
rect 42242 21128 42248 21140
rect 41472 21100 42248 21128
rect 41472 21088 41478 21100
rect 42242 21088 42248 21100
rect 42300 21088 42306 21140
rect 46658 21088 46664 21140
rect 46716 21128 46722 21140
rect 46753 21131 46811 21137
rect 46753 21128 46765 21131
rect 46716 21100 46765 21128
rect 46716 21088 46722 21100
rect 46753 21097 46765 21100
rect 46799 21097 46811 21131
rect 53653 21131 53711 21137
rect 46753 21091 46811 21097
rect 51644 21100 53052 21128
rect 31662 21020 31668 21072
rect 31720 21032 31754 21072
rect 31720 21020 31726 21032
rect 43898 21020 43904 21072
rect 43956 21060 43962 21072
rect 46106 21060 46112 21072
rect 43956 21032 46112 21060
rect 43956 21020 43962 21032
rect 46106 21020 46112 21032
rect 46164 21020 46170 21072
rect 51074 21020 51080 21072
rect 51132 21060 51138 21072
rect 51132 21032 51580 21060
rect 51132 21020 51138 21032
rect 30745 20995 30803 21001
rect 30745 20992 30757 20995
rect 30024 20964 30757 20992
rect 26881 20955 26939 20961
rect 30745 20961 30757 20964
rect 30791 20961 30803 20995
rect 45741 20995 45799 21001
rect 45741 20992 45753 20995
rect 30745 20955 30803 20961
rect 44744 20964 45753 20992
rect 18230 20884 18236 20936
rect 18288 20884 18294 20936
rect 19886 20884 19892 20936
rect 19944 20884 19950 20936
rect 20622 20884 20628 20936
rect 20680 20884 20686 20936
rect 22732 20927 22790 20933
rect 22732 20893 22744 20927
rect 22778 20924 22790 20927
rect 23014 20924 23020 20936
rect 22778 20896 23020 20924
rect 22778 20893 22790 20896
rect 22732 20887 22790 20893
rect 23014 20884 23020 20896
rect 23072 20884 23078 20936
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 23992 20896 24624 20924
rect 23992 20884 23998 20896
rect 11793 20859 11851 20865
rect 11793 20825 11805 20859
rect 11839 20856 11851 20859
rect 12989 20859 13047 20865
rect 12989 20856 13001 20859
rect 11839 20828 13001 20856
rect 11839 20825 11851 20828
rect 11793 20819 11851 20825
rect 12989 20825 13001 20828
rect 13035 20856 13047 20859
rect 15473 20859 15531 20865
rect 13035 20828 13860 20856
rect 13035 20825 13047 20828
rect 12989 20819 13047 20825
rect 13832 20800 13860 20828
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 17313 20859 17371 20865
rect 17313 20856 17325 20859
rect 15519 20828 17325 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 17313 20825 17325 20828
rect 17359 20825 17371 20859
rect 17313 20819 17371 20825
rect 17957 20859 18015 20865
rect 17957 20825 17969 20859
rect 18003 20856 18015 20859
rect 24121 20859 24179 20865
rect 24121 20856 24133 20859
rect 18003 20828 19012 20856
rect 18003 20825 18015 20828
rect 17957 20819 18015 20825
rect 18984 20800 19012 20828
rect 20456 20828 24133 20856
rect 20456 20800 20484 20828
rect 24121 20825 24133 20828
rect 24167 20856 24179 20859
rect 24302 20856 24308 20868
rect 24167 20828 24308 20856
rect 24167 20825 24179 20828
rect 24121 20819 24179 20825
rect 24302 20816 24308 20828
rect 24360 20816 24366 20868
rect 8941 20791 8999 20797
rect 8941 20757 8953 20791
rect 8987 20757 8999 20791
rect 8941 20751 8999 20757
rect 9309 20791 9367 20797
rect 9309 20757 9321 20791
rect 9355 20788 9367 20791
rect 9398 20788 9404 20800
rect 9355 20760 9404 20788
rect 9355 20757 9367 20760
rect 9309 20751 9367 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 9858 20748 9864 20800
rect 9916 20788 9922 20800
rect 10962 20788 10968 20800
rect 9916 20760 10968 20788
rect 9916 20748 9922 20760
rect 10962 20748 10968 20760
rect 11020 20788 11026 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 11020 20760 11437 20788
rect 11020 20748 11026 20760
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 13722 20748 13728 20800
rect 13780 20748 13786 20800
rect 13814 20748 13820 20800
rect 13872 20748 13878 20800
rect 14461 20791 14519 20797
rect 14461 20757 14473 20791
rect 14507 20788 14519 20791
rect 14918 20788 14924 20800
rect 14507 20760 14924 20788
rect 14507 20757 14519 20760
rect 14461 20751 14519 20757
rect 14918 20748 14924 20760
rect 14976 20788 14982 20800
rect 15381 20791 15439 20797
rect 15381 20788 15393 20791
rect 14976 20760 15393 20788
rect 14976 20748 14982 20760
rect 15381 20757 15393 20760
rect 15427 20757 15439 20791
rect 15381 20751 15439 20757
rect 16574 20748 16580 20800
rect 16632 20748 16638 20800
rect 18782 20748 18788 20800
rect 18840 20748 18846 20800
rect 18966 20748 18972 20800
rect 19024 20748 19030 20800
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20788 19579 20791
rect 19794 20788 19800 20800
rect 19567 20760 19800 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 20438 20748 20444 20800
rect 20496 20748 20502 20800
rect 20530 20748 20536 20800
rect 20588 20748 20594 20800
rect 21266 20748 21272 20800
rect 21324 20748 21330 20800
rect 24596 20788 24624 20896
rect 25314 20884 25320 20936
rect 25372 20884 25378 20936
rect 25406 20884 25412 20936
rect 25464 20933 25470 20936
rect 25464 20927 25492 20933
rect 25480 20893 25492 20927
rect 25464 20887 25492 20893
rect 25464 20884 25470 20887
rect 25590 20884 25596 20936
rect 25648 20884 25654 20936
rect 26712 20924 26740 20952
rect 44744 20936 44772 20964
rect 45741 20961 45753 20964
rect 45787 20961 45799 20995
rect 45741 20955 45799 20961
rect 46474 20952 46480 21004
rect 46532 20992 46538 21004
rect 47397 20995 47455 21001
rect 47397 20992 47409 20995
rect 46532 20964 47409 20992
rect 46532 20952 46538 20964
rect 47397 20961 47409 20964
rect 47443 20992 47455 20995
rect 51350 20992 51356 21004
rect 47443 20964 51356 20992
rect 47443 20961 47455 20964
rect 47397 20955 47455 20961
rect 51350 20952 51356 20964
rect 51408 20952 51414 21004
rect 27157 20927 27215 20933
rect 27157 20924 27169 20927
rect 26712 20896 27169 20924
rect 27157 20893 27169 20896
rect 27203 20893 27215 20927
rect 27157 20887 27215 20893
rect 27982 20884 27988 20936
rect 28040 20884 28046 20936
rect 28810 20884 28816 20936
rect 28868 20884 28874 20936
rect 31018 20884 31024 20936
rect 31076 20884 31082 20936
rect 32858 20884 32864 20936
rect 32916 20884 32922 20936
rect 33686 20884 33692 20936
rect 33744 20884 33750 20936
rect 34977 20927 35035 20933
rect 34977 20893 34989 20927
rect 35023 20924 35035 20927
rect 35342 20924 35348 20936
rect 35023 20896 35348 20924
rect 35023 20893 35035 20896
rect 34977 20887 35035 20893
rect 35342 20884 35348 20896
rect 35400 20884 35406 20936
rect 35894 20884 35900 20936
rect 35952 20924 35958 20936
rect 36081 20927 36139 20933
rect 36081 20924 36093 20927
rect 35952 20896 36093 20924
rect 35952 20884 35958 20896
rect 36081 20893 36093 20896
rect 36127 20893 36139 20927
rect 36081 20887 36139 20893
rect 37550 20884 37556 20936
rect 37608 20884 37614 20936
rect 38286 20884 38292 20936
rect 38344 20884 38350 20936
rect 41782 20884 41788 20936
rect 41840 20884 41846 20936
rect 41874 20884 41880 20936
rect 41932 20924 41938 20936
rect 42429 20927 42487 20933
rect 42429 20924 42441 20927
rect 41932 20896 42441 20924
rect 41932 20884 41938 20896
rect 42429 20893 42441 20896
rect 42475 20893 42487 20927
rect 42429 20887 42487 20893
rect 44726 20884 44732 20936
rect 44784 20884 44790 20936
rect 45002 20884 45008 20936
rect 45060 20884 45066 20936
rect 47670 20884 47676 20936
rect 47728 20884 47734 20936
rect 49145 20927 49203 20933
rect 49145 20893 49157 20927
rect 49191 20924 49203 20927
rect 49510 20924 49516 20936
rect 49191 20896 49516 20924
rect 49191 20893 49203 20896
rect 49145 20887 49203 20893
rect 49510 20884 49516 20896
rect 49568 20884 49574 20936
rect 50801 20927 50859 20933
rect 50801 20893 50813 20927
rect 50847 20924 50859 20927
rect 51258 20924 51264 20936
rect 50847 20896 51264 20924
rect 50847 20893 50859 20896
rect 50801 20887 50859 20893
rect 51258 20884 51264 20896
rect 51316 20884 51322 20936
rect 51445 20927 51503 20933
rect 51445 20893 51457 20927
rect 51491 20893 51503 20927
rect 51552 20924 51580 21032
rect 51644 21001 51672 21100
rect 53024 21060 53052 21100
rect 53653 21097 53665 21131
rect 53699 21128 53711 21131
rect 54754 21128 54760 21140
rect 53699 21100 54760 21128
rect 53699 21097 53711 21100
rect 53653 21091 53711 21097
rect 54754 21088 54760 21100
rect 54812 21088 54818 21140
rect 57514 21128 57520 21140
rect 55692 21100 57520 21128
rect 53742 21060 53748 21072
rect 53024 21032 53748 21060
rect 53742 21020 53748 21032
rect 53800 21020 53806 21072
rect 55125 21063 55183 21069
rect 55125 21029 55137 21063
rect 55171 21060 55183 21063
rect 55171 21032 55628 21060
rect 55171 21029 55183 21032
rect 55125 21023 55183 21029
rect 55600 21004 55628 21032
rect 51629 20995 51687 21001
rect 51629 20961 51641 20995
rect 51675 20961 51687 20995
rect 51994 20992 52000 21004
rect 51629 20955 51687 20961
rect 51828 20964 52000 20992
rect 51828 20924 51856 20964
rect 51994 20952 52000 20964
rect 52052 20992 52058 21004
rect 52089 20995 52147 21001
rect 52089 20992 52101 20995
rect 52052 20964 52101 20992
rect 52052 20952 52058 20964
rect 52089 20961 52101 20964
rect 52135 20961 52147 20995
rect 52089 20955 52147 20961
rect 52178 20952 52184 21004
rect 52236 20992 52242 21004
rect 52365 20995 52423 21001
rect 52365 20992 52377 20995
rect 52236 20964 52377 20992
rect 52236 20952 52242 20964
rect 52365 20961 52377 20964
rect 52411 20961 52423 20995
rect 52365 20955 52423 20961
rect 52638 20952 52644 21004
rect 52696 20992 52702 21004
rect 52696 20964 53880 20992
rect 52696 20952 52702 20964
rect 51552 20896 51856 20924
rect 51445 20887 51503 20893
rect 26697 20859 26755 20865
rect 26697 20825 26709 20859
rect 26743 20856 26755 20859
rect 27801 20859 27859 20865
rect 27801 20856 27813 20859
rect 26743 20828 27813 20856
rect 26743 20825 26755 20828
rect 26697 20819 26755 20825
rect 27801 20825 27813 20828
rect 27847 20825 27859 20859
rect 27801 20819 27859 20825
rect 45370 20816 45376 20868
rect 45428 20856 45434 20868
rect 46385 20859 46443 20865
rect 46385 20856 46397 20859
rect 45428 20828 46397 20856
rect 45428 20816 45434 20828
rect 46385 20825 46397 20828
rect 46431 20825 46443 20859
rect 46385 20819 46443 20825
rect 47121 20859 47179 20865
rect 47121 20825 47133 20859
rect 47167 20856 47179 20859
rect 47302 20856 47308 20868
rect 47167 20828 47308 20856
rect 47167 20825 47179 20828
rect 47121 20819 47179 20825
rect 47302 20816 47308 20828
rect 47360 20816 47366 20868
rect 48682 20816 48688 20868
rect 48740 20856 48746 20868
rect 48961 20859 49019 20865
rect 48961 20856 48973 20859
rect 48740 20828 48973 20856
rect 48740 20816 48746 20828
rect 48961 20825 48973 20828
rect 49007 20856 49019 20859
rect 49007 20828 50200 20856
rect 49007 20825 49019 20828
rect 48961 20819 49019 20825
rect 50172 20800 50200 20828
rect 25406 20788 25412 20800
rect 24596 20760 25412 20788
rect 25406 20748 25412 20760
rect 25464 20748 25470 20800
rect 26142 20748 26148 20800
rect 26200 20788 26206 20800
rect 26237 20791 26295 20797
rect 26237 20788 26249 20791
rect 26200 20760 26249 20788
rect 26200 20748 26206 20760
rect 26237 20757 26249 20760
rect 26283 20757 26295 20791
rect 26237 20751 26295 20757
rect 28534 20748 28540 20800
rect 28592 20748 28598 20800
rect 28902 20748 28908 20800
rect 28960 20788 28966 20800
rect 29365 20791 29423 20797
rect 29365 20788 29377 20791
rect 28960 20760 29377 20788
rect 28960 20748 28966 20760
rect 29365 20757 29377 20760
rect 29411 20757 29423 20791
rect 29365 20751 29423 20757
rect 30558 20748 30564 20800
rect 30616 20748 30622 20800
rect 30653 20791 30711 20797
rect 30653 20757 30665 20791
rect 30699 20788 30711 20791
rect 31665 20791 31723 20797
rect 31665 20788 31677 20791
rect 30699 20760 31677 20788
rect 30699 20757 30711 20760
rect 30653 20751 30711 20757
rect 31665 20757 31677 20760
rect 31711 20757 31723 20791
rect 31665 20751 31723 20757
rect 33410 20748 33416 20800
rect 33468 20748 33474 20800
rect 34238 20748 34244 20800
rect 34296 20748 34302 20800
rect 35345 20791 35403 20797
rect 35345 20757 35357 20791
rect 35391 20788 35403 20791
rect 35802 20788 35808 20800
rect 35391 20760 35808 20788
rect 35391 20757 35403 20760
rect 35345 20751 35403 20757
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 36722 20748 36728 20800
rect 36780 20748 36786 20800
rect 37369 20791 37427 20797
rect 37369 20757 37381 20791
rect 37415 20788 37427 20791
rect 37458 20788 37464 20800
rect 37415 20760 37464 20788
rect 37415 20757 37427 20760
rect 37369 20751 37427 20757
rect 37458 20748 37464 20760
rect 37516 20748 37522 20800
rect 38102 20748 38108 20800
rect 38160 20748 38166 20800
rect 38838 20748 38844 20800
rect 38896 20748 38902 20800
rect 39206 20748 39212 20800
rect 39264 20748 39270 20800
rect 42334 20748 42340 20800
rect 42392 20748 42398 20800
rect 44634 20748 44640 20800
rect 44692 20748 44698 20800
rect 45646 20748 45652 20800
rect 45704 20748 45710 20800
rect 47213 20791 47271 20797
rect 47213 20757 47225 20791
rect 47259 20788 47271 20791
rect 48225 20791 48283 20797
rect 48225 20788 48237 20791
rect 47259 20760 48237 20788
rect 47259 20757 47271 20760
rect 47213 20751 47271 20757
rect 48225 20757 48237 20760
rect 48271 20757 48283 20791
rect 48225 20751 48283 20757
rect 48593 20791 48651 20797
rect 48593 20757 48605 20791
rect 48639 20788 48651 20791
rect 48774 20788 48780 20800
rect 48639 20760 48780 20788
rect 48639 20757 48651 20760
rect 48593 20751 48651 20757
rect 48774 20748 48780 20760
rect 48832 20748 48838 20800
rect 49694 20748 49700 20800
rect 49752 20748 49758 20800
rect 50154 20748 50160 20800
rect 50212 20748 50218 20800
rect 51074 20748 51080 20800
rect 51132 20748 51138 20800
rect 51460 20788 51488 20887
rect 52454 20884 52460 20936
rect 52512 20933 52518 20936
rect 52512 20927 52540 20933
rect 52528 20893 52540 20927
rect 52512 20887 52540 20893
rect 52512 20884 52518 20887
rect 53558 20884 53564 20936
rect 53616 20924 53622 20936
rect 53745 20927 53803 20933
rect 53745 20924 53757 20927
rect 53616 20896 53757 20924
rect 53616 20884 53622 20896
rect 53745 20893 53757 20896
rect 53791 20893 53803 20927
rect 53852 20924 53880 20964
rect 55582 20952 55588 21004
rect 55640 20952 55646 21004
rect 55692 21001 55720 21100
rect 57514 21088 57520 21100
rect 57572 21088 57578 21140
rect 55677 20995 55735 21001
rect 55677 20961 55689 20995
rect 55723 20961 55735 20995
rect 56042 20992 56048 21004
rect 55677 20955 55735 20961
rect 55784 20964 56048 20992
rect 55784 20924 55812 20964
rect 56042 20952 56048 20964
rect 56100 20952 56106 21004
rect 56226 20952 56232 21004
rect 56284 20992 56290 21004
rect 56321 20995 56379 21001
rect 56321 20992 56333 20995
rect 56284 20964 56333 20992
rect 56284 20952 56290 20964
rect 56321 20961 56333 20964
rect 56367 20961 56379 20995
rect 56321 20955 56379 20961
rect 56410 20952 56416 21004
rect 56468 20992 56474 21004
rect 56714 20995 56772 21001
rect 56714 20992 56726 20995
rect 56468 20964 56726 20992
rect 56468 20952 56474 20964
rect 56714 20961 56726 20964
rect 56760 20961 56772 20995
rect 56714 20955 56772 20961
rect 56870 20952 56876 21004
rect 56928 20952 56934 21004
rect 58158 20952 58164 21004
rect 58216 20952 58222 21004
rect 53852 20896 55812 20924
rect 55861 20927 55919 20933
rect 53745 20887 53803 20893
rect 55861 20893 55873 20927
rect 55907 20893 55919 20927
rect 55861 20887 55919 20893
rect 53190 20816 53196 20868
rect 53248 20856 53254 20868
rect 54012 20859 54070 20865
rect 53248 20828 53420 20856
rect 53248 20816 53254 20828
rect 52730 20788 52736 20800
rect 51460 20760 52736 20788
rect 52730 20748 52736 20760
rect 52788 20748 52794 20800
rect 53282 20748 53288 20800
rect 53340 20748 53346 20800
rect 53392 20788 53420 20828
rect 54012 20825 54024 20859
rect 54058 20856 54070 20859
rect 55030 20856 55036 20868
rect 54058 20828 55036 20856
rect 54058 20825 54070 20828
rect 54012 20819 54070 20825
rect 55030 20816 55036 20828
rect 55088 20816 55094 20868
rect 55493 20791 55551 20797
rect 55493 20788 55505 20791
rect 53392 20760 55505 20788
rect 55493 20757 55505 20760
rect 55539 20788 55551 20791
rect 55766 20788 55772 20800
rect 55539 20760 55772 20788
rect 55539 20757 55551 20760
rect 55493 20751 55551 20757
rect 55766 20748 55772 20760
rect 55824 20748 55830 20800
rect 55876 20788 55904 20887
rect 56594 20884 56600 20936
rect 56652 20884 56658 20936
rect 57790 20816 57796 20868
rect 57848 20856 57854 20868
rect 58069 20859 58127 20865
rect 58069 20856 58081 20859
rect 57848 20828 58081 20856
rect 57848 20816 57854 20828
rect 58069 20825 58081 20828
rect 58115 20825 58127 20859
rect 58069 20819 58127 20825
rect 56962 20788 56968 20800
rect 55876 20760 56968 20788
rect 56962 20748 56968 20760
rect 57020 20748 57026 20800
rect 57514 20748 57520 20800
rect 57572 20748 57578 20800
rect 57606 20748 57612 20800
rect 57664 20748 57670 20800
rect 57698 20748 57704 20800
rect 57756 20788 57762 20800
rect 57977 20791 58035 20797
rect 57977 20788 57989 20791
rect 57756 20760 57989 20788
rect 57756 20748 57762 20760
rect 57977 20757 57989 20760
rect 58023 20757 58035 20791
rect 57977 20751 58035 20757
rect 1104 20698 59040 20720
rect 1104 20646 15394 20698
rect 15446 20646 15458 20698
rect 15510 20646 15522 20698
rect 15574 20646 15586 20698
rect 15638 20646 15650 20698
rect 15702 20646 29838 20698
rect 29890 20646 29902 20698
rect 29954 20646 29966 20698
rect 30018 20646 30030 20698
rect 30082 20646 30094 20698
rect 30146 20646 44282 20698
rect 44334 20646 44346 20698
rect 44398 20646 44410 20698
rect 44462 20646 44474 20698
rect 44526 20646 44538 20698
rect 44590 20646 58726 20698
rect 58778 20646 58790 20698
rect 58842 20646 58854 20698
rect 58906 20646 58918 20698
rect 58970 20646 58982 20698
rect 59034 20646 59040 20698
rect 1104 20624 59040 20646
rect 3789 20587 3847 20593
rect 3789 20584 3801 20587
rect 2746 20556 3801 20584
rect 2746 20528 2774 20556
rect 3789 20553 3801 20556
rect 3835 20584 3847 20587
rect 4062 20584 4068 20596
rect 3835 20556 4068 20584
rect 3835 20553 3847 20556
rect 3789 20547 3847 20553
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 4430 20544 4436 20596
rect 4488 20584 4494 20596
rect 6638 20584 6644 20596
rect 4488 20556 6644 20584
rect 4488 20544 4494 20556
rect 6638 20544 6644 20556
rect 6696 20584 6702 20596
rect 6825 20587 6883 20593
rect 6825 20584 6837 20587
rect 6696 20556 6837 20584
rect 6696 20544 6702 20556
rect 6825 20553 6837 20556
rect 6871 20553 6883 20587
rect 6825 20547 6883 20553
rect 7558 20544 7564 20596
rect 7616 20544 7622 20596
rect 13081 20587 13139 20593
rect 13081 20553 13093 20587
rect 13127 20584 13139 20587
rect 13906 20584 13912 20596
rect 13127 20556 13912 20584
rect 13127 20553 13139 20556
rect 13081 20547 13139 20553
rect 13906 20544 13912 20556
rect 13964 20584 13970 20596
rect 18509 20587 18567 20593
rect 13964 20556 15148 20584
rect 13964 20544 13970 20556
rect 2746 20516 2780 20528
rect 2056 20488 2780 20516
rect 2056 20457 2084 20488
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20417 2099 20451
rect 2041 20411 2099 20417
rect 2308 20451 2366 20457
rect 2308 20417 2320 20451
rect 2354 20448 2366 20451
rect 3694 20448 3700 20460
rect 2354 20420 3700 20448
rect 2354 20417 2366 20420
rect 2308 20411 2366 20417
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 3970 20408 3976 20460
rect 4028 20448 4034 20460
rect 4028 20420 4384 20448
rect 4028 20408 4034 20420
rect 3421 20315 3479 20321
rect 3421 20281 3433 20315
rect 3467 20312 3479 20315
rect 3988 20312 4016 20408
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 4154 20380 4160 20392
rect 4111 20352 4160 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20349 4307 20383
rect 4356 20380 4384 20420
rect 4982 20408 4988 20460
rect 5040 20408 5046 20460
rect 6730 20408 6736 20460
rect 6788 20408 6794 20460
rect 7576 20448 7604 20544
rect 11968 20519 12026 20525
rect 11968 20485 11980 20519
rect 12014 20516 12026 20519
rect 13722 20516 13728 20528
rect 12014 20488 13728 20516
rect 12014 20485 12026 20488
rect 11968 20479 12026 20485
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 15120 20460 15148 20556
rect 18509 20553 18521 20587
rect 18555 20584 18567 20587
rect 19334 20584 19340 20596
rect 18555 20556 19340 20584
rect 18555 20553 18567 20556
rect 18509 20547 18567 20553
rect 19334 20544 19340 20556
rect 19392 20544 19398 20596
rect 19518 20584 19524 20596
rect 19444 20556 19524 20584
rect 15280 20519 15338 20525
rect 15280 20485 15292 20519
rect 15326 20516 15338 20519
rect 15838 20516 15844 20528
rect 15326 20488 15844 20516
rect 15326 20485 15338 20488
rect 15280 20479 15338 20485
rect 15838 20476 15844 20488
rect 15896 20476 15902 20528
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 7576 20420 7665 20448
rect 7653 20417 7665 20420
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 7920 20451 7978 20457
rect 7920 20417 7932 20451
rect 7966 20448 7978 20451
rect 8754 20448 8760 20460
rect 7966 20420 8760 20448
rect 7966 20417 7978 20420
rect 7920 20411 7978 20417
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 9493 20451 9551 20457
rect 9493 20417 9505 20451
rect 9539 20448 9551 20451
rect 9858 20448 9864 20460
rect 9539 20420 9864 20448
rect 9539 20417 9551 20420
rect 9493 20411 9551 20417
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 10410 20408 10416 20460
rect 10468 20408 10474 20460
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 14642 20448 14648 20460
rect 13228 20420 14648 20448
rect 13228 20408 13234 20420
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15102 20408 15108 20460
rect 15160 20408 15166 20460
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20448 18475 20451
rect 19150 20448 19156 20460
rect 18463 20420 19156 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 5102 20383 5160 20389
rect 5102 20380 5114 20383
rect 4356 20352 5114 20380
rect 4249 20343 4307 20349
rect 5102 20349 5114 20352
rect 5148 20349 5160 20383
rect 5102 20343 5160 20349
rect 3467 20284 4016 20312
rect 3467 20281 3479 20284
rect 3421 20275 3479 20281
rect 4264 20244 4292 20343
rect 5258 20340 5264 20392
rect 5316 20340 5322 20392
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7282 20380 7288 20392
rect 7055 20352 7288 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7282 20340 7288 20352
rect 7340 20340 7346 20392
rect 9674 20340 9680 20392
rect 9732 20340 9738 20392
rect 10530 20383 10588 20389
rect 10530 20380 10542 20383
rect 9784 20352 10542 20380
rect 4430 20272 4436 20324
rect 4488 20312 4494 20324
rect 4709 20315 4767 20321
rect 4709 20312 4721 20315
rect 4488 20284 4721 20312
rect 4488 20272 4494 20284
rect 4709 20281 4721 20284
rect 4755 20281 4767 20315
rect 6638 20312 6644 20324
rect 4709 20275 4767 20281
rect 5828 20284 6644 20312
rect 5828 20244 5856 20284
rect 6638 20272 6644 20284
rect 6696 20272 6702 20324
rect 9784 20312 9812 20352
rect 10530 20349 10542 20352
rect 10576 20349 10588 20383
rect 10530 20343 10588 20349
rect 10689 20383 10747 20389
rect 10689 20349 10701 20383
rect 10735 20380 10747 20383
rect 11514 20380 11520 20392
rect 10735 20352 11520 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 9048 20284 9812 20312
rect 9048 20256 9076 20284
rect 9858 20272 9864 20324
rect 9916 20312 9922 20324
rect 10137 20315 10195 20321
rect 10137 20312 10149 20315
rect 9916 20284 10149 20312
rect 9916 20272 9922 20284
rect 10137 20281 10149 20284
rect 10183 20281 10195 20315
rect 10137 20275 10195 20281
rect 4264 20216 5856 20244
rect 5902 20204 5908 20256
rect 5960 20204 5966 20256
rect 6362 20204 6368 20256
rect 6420 20204 6426 20256
rect 9030 20204 9036 20256
rect 9088 20204 9094 20256
rect 9401 20247 9459 20253
rect 9401 20213 9413 20247
rect 9447 20244 9459 20247
rect 11072 20244 11100 20352
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 11701 20383 11759 20389
rect 11701 20349 11713 20383
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 9447 20216 11100 20244
rect 11333 20247 11391 20253
rect 9447 20213 9459 20216
rect 9401 20207 9459 20213
rect 11333 20213 11345 20247
rect 11379 20244 11391 20247
rect 11514 20244 11520 20256
rect 11379 20216 11520 20244
rect 11379 20213 11391 20216
rect 11333 20207 11391 20213
rect 11514 20204 11520 20216
rect 11572 20204 11578 20256
rect 11716 20244 11744 20343
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 13872 20352 14933 20380
rect 13872 20340 13878 20352
rect 14921 20349 14933 20352
rect 14967 20380 14979 20383
rect 15010 20380 15016 20392
rect 14967 20352 15016 20380
rect 14967 20349 14979 20352
rect 14921 20343 14979 20349
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 17405 20383 17463 20389
rect 17405 20349 17417 20383
rect 17451 20349 17463 20383
rect 17405 20343 17463 20349
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 18966 20380 18972 20392
rect 18739 20352 18972 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 17420 20312 17448 20343
rect 18966 20340 18972 20352
rect 19024 20340 19030 20392
rect 19444 20380 19472 20556
rect 19518 20544 19524 20556
rect 19576 20584 19582 20596
rect 20438 20584 20444 20596
rect 19576 20556 20444 20584
rect 19576 20544 19582 20556
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 22186 20544 22192 20596
rect 22244 20544 22250 20596
rect 23661 20587 23719 20593
rect 23661 20553 23673 20587
rect 23707 20584 23719 20587
rect 23934 20584 23940 20596
rect 23707 20556 23940 20584
rect 23707 20553 23719 20556
rect 23661 20547 23719 20553
rect 23934 20544 23940 20556
rect 23992 20544 23998 20596
rect 24121 20587 24179 20593
rect 24121 20553 24133 20587
rect 24167 20584 24179 20587
rect 24578 20584 24584 20596
rect 24167 20556 24584 20584
rect 24167 20553 24179 20556
rect 24121 20547 24179 20553
rect 24578 20544 24584 20556
rect 24636 20544 24642 20596
rect 26694 20544 26700 20596
rect 26752 20544 26758 20596
rect 27890 20544 27896 20596
rect 27948 20544 27954 20596
rect 27982 20544 27988 20596
rect 28040 20584 28046 20596
rect 28077 20587 28135 20593
rect 28077 20584 28089 20587
rect 28040 20556 28089 20584
rect 28040 20544 28046 20556
rect 28077 20553 28089 20556
rect 28123 20553 28135 20587
rect 28077 20547 28135 20553
rect 28537 20587 28595 20593
rect 28537 20553 28549 20587
rect 28583 20584 28595 20587
rect 28902 20584 28908 20596
rect 28583 20556 28908 20584
rect 28583 20553 28595 20556
rect 28537 20547 28595 20553
rect 28902 20544 28908 20556
rect 28960 20544 28966 20596
rect 30558 20584 30564 20596
rect 29472 20556 30564 20584
rect 19610 20516 19616 20528
rect 19536 20488 19616 20516
rect 19536 20457 19564 20488
rect 19610 20476 19616 20488
rect 19668 20516 19674 20528
rect 22204 20516 22232 20544
rect 19668 20488 22232 20516
rect 19668 20476 19674 20488
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 19788 20451 19846 20457
rect 19788 20417 19800 20451
rect 19834 20448 19846 20451
rect 20530 20448 20536 20460
rect 19834 20420 20536 20448
rect 19834 20417 19846 20420
rect 19788 20411 19846 20417
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 22204 20448 22232 20488
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 22204 20420 22293 20448
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22548 20451 22606 20457
rect 22548 20417 22560 20451
rect 22594 20448 22606 20451
rect 23842 20448 23848 20460
rect 22594 20420 23848 20448
rect 22594 20417 22606 20420
rect 22548 20411 22606 20417
rect 23842 20408 23848 20420
rect 23900 20408 23906 20460
rect 25584 20451 25642 20457
rect 25584 20417 25596 20451
rect 25630 20448 25642 20451
rect 26602 20448 26608 20460
rect 25630 20420 26608 20448
rect 25630 20417 25642 20420
rect 25584 20411 25642 20417
rect 26602 20408 26608 20420
rect 26660 20408 26666 20460
rect 19076 20352 19472 20380
rect 21085 20383 21143 20389
rect 18049 20315 18107 20321
rect 18049 20312 18061 20315
rect 17420 20284 18061 20312
rect 18049 20281 18061 20284
rect 18095 20281 18107 20315
rect 18049 20275 18107 20281
rect 18138 20272 18144 20324
rect 18196 20272 18202 20324
rect 12066 20244 12072 20256
rect 11716 20216 12072 20244
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 16393 20247 16451 20253
rect 16393 20244 16405 20247
rect 14332 20216 16405 20244
rect 14332 20204 14338 20216
rect 16393 20213 16405 20216
rect 16439 20244 16451 20247
rect 16666 20244 16672 20256
rect 16439 20216 16672 20244
rect 16439 20213 16451 20216
rect 16393 20207 16451 20213
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 16850 20204 16856 20256
rect 16908 20204 16914 20256
rect 17954 20204 17960 20256
rect 18012 20204 18018 20256
rect 18156 20244 18184 20272
rect 19076 20253 19104 20352
rect 21085 20349 21097 20383
rect 21131 20380 21143 20383
rect 21131 20352 21220 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 21192 20256 21220 20352
rect 24026 20340 24032 20392
rect 24084 20380 24090 20392
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 24084 20352 24225 20380
rect 24084 20340 24090 20352
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 24305 20383 24363 20389
rect 24305 20349 24317 20383
rect 24351 20349 24363 20383
rect 24305 20343 24363 20349
rect 25317 20383 25375 20389
rect 25317 20349 25329 20383
rect 25363 20349 25375 20383
rect 27908 20380 27936 20544
rect 29472 20528 29500 20556
rect 30558 20544 30564 20556
rect 30616 20544 30622 20596
rect 30742 20544 30748 20596
rect 30800 20584 30806 20596
rect 31573 20587 31631 20593
rect 31573 20584 31585 20587
rect 30800 20556 31585 20584
rect 30800 20544 30806 20556
rect 31573 20553 31585 20556
rect 31619 20584 31631 20587
rect 31662 20584 31668 20596
rect 31619 20556 31668 20584
rect 31619 20553 31631 20556
rect 31573 20547 31631 20553
rect 31662 20544 31668 20556
rect 31720 20544 31726 20596
rect 32858 20544 32864 20596
rect 32916 20584 32922 20596
rect 32953 20587 33011 20593
rect 32953 20584 32965 20587
rect 32916 20556 32965 20584
rect 32916 20544 32922 20556
rect 32953 20553 32965 20556
rect 32999 20553 33011 20587
rect 32953 20547 33011 20553
rect 33413 20587 33471 20593
rect 33413 20553 33425 20587
rect 33459 20584 33471 20587
rect 34238 20584 34244 20596
rect 33459 20556 34244 20584
rect 33459 20553 33471 20556
rect 33413 20547 33471 20553
rect 34238 20544 34244 20556
rect 34296 20544 34302 20596
rect 37550 20544 37556 20596
rect 37608 20544 37614 20596
rect 37921 20587 37979 20593
rect 37921 20553 37933 20587
rect 37967 20584 37979 20587
rect 38838 20584 38844 20596
rect 37967 20556 38844 20584
rect 37967 20553 37979 20556
rect 37921 20547 37979 20553
rect 38838 20544 38844 20556
rect 38896 20544 38902 20596
rect 40770 20544 40776 20596
rect 40828 20544 40834 20596
rect 41782 20544 41788 20596
rect 41840 20584 41846 20596
rect 42429 20587 42487 20593
rect 42429 20584 42441 20587
rect 41840 20556 42441 20584
rect 41840 20544 41846 20556
rect 42429 20553 42441 20556
rect 42475 20553 42487 20587
rect 42429 20547 42487 20553
rect 42889 20587 42947 20593
rect 42889 20553 42901 20587
rect 42935 20584 42947 20587
rect 43254 20584 43260 20596
rect 42935 20556 43260 20584
rect 42935 20553 42947 20556
rect 42889 20547 42947 20553
rect 43254 20544 43260 20556
rect 43312 20544 43318 20596
rect 48222 20584 48228 20596
rect 45756 20556 48228 20584
rect 28445 20519 28503 20525
rect 28445 20485 28457 20519
rect 28491 20516 28503 20519
rect 29454 20516 29460 20528
rect 28491 20488 29460 20516
rect 28491 20485 28503 20488
rect 28445 20479 28503 20485
rect 29454 20476 29460 20488
rect 29512 20476 29518 20528
rect 30092 20519 30150 20525
rect 30092 20485 30104 20519
rect 30138 20516 30150 20519
rect 30834 20516 30840 20528
rect 30138 20488 30840 20516
rect 30138 20485 30150 20488
rect 30092 20479 30150 20485
rect 30834 20476 30840 20488
rect 30892 20476 30898 20528
rect 34146 20516 34152 20528
rect 33244 20488 34152 20516
rect 30558 20448 30564 20460
rect 28920 20420 30564 20448
rect 28920 20389 28948 20420
rect 30558 20408 30564 20420
rect 30616 20408 30622 20460
rect 28629 20383 28687 20389
rect 28629 20380 28641 20383
rect 27908 20352 28641 20380
rect 25317 20343 25375 20349
rect 28629 20349 28641 20352
rect 28675 20349 28687 20383
rect 28629 20343 28687 20349
rect 28905 20383 28963 20389
rect 28905 20349 28917 20383
rect 28951 20349 28963 20383
rect 28905 20343 28963 20349
rect 24320 20312 24348 20343
rect 24228 20284 24348 20312
rect 24228 20256 24256 20284
rect 24854 20272 24860 20324
rect 24912 20272 24918 20324
rect 25332 20256 25360 20343
rect 28920 20312 28948 20343
rect 29730 20340 29736 20392
rect 29788 20380 29794 20392
rect 29825 20383 29883 20389
rect 29825 20380 29837 20383
rect 29788 20352 29837 20380
rect 29788 20340 29794 20352
rect 29825 20349 29837 20352
rect 29871 20349 29883 20383
rect 29825 20343 29883 20349
rect 32861 20383 32919 20389
rect 32861 20349 32873 20383
rect 32907 20380 32919 20383
rect 33244 20380 33272 20488
rect 34146 20476 34152 20488
rect 34204 20516 34210 20528
rect 37826 20516 37832 20528
rect 34204 20488 37832 20516
rect 34204 20476 34210 20488
rect 37826 20476 37832 20488
rect 37884 20476 37890 20528
rect 41414 20516 41420 20528
rect 40880 20488 41420 20516
rect 33321 20451 33379 20457
rect 33321 20417 33333 20451
rect 33367 20448 33379 20451
rect 33962 20448 33968 20460
rect 33367 20420 33968 20448
rect 33367 20417 33379 20420
rect 33321 20411 33379 20417
rect 33962 20408 33968 20420
rect 34020 20408 34026 20460
rect 34784 20451 34842 20457
rect 34784 20417 34796 20451
rect 34830 20448 34842 20451
rect 36633 20451 36691 20457
rect 36633 20448 36645 20451
rect 34830 20420 36645 20448
rect 34830 20417 34842 20420
rect 34784 20411 34842 20417
rect 36633 20417 36645 20420
rect 36679 20417 36691 20451
rect 38381 20451 38439 20457
rect 36633 20411 36691 20417
rect 37476 20420 38148 20448
rect 37476 20392 37504 20420
rect 33505 20383 33563 20389
rect 33505 20380 33517 20383
rect 32907 20352 33517 20380
rect 32907 20349 32919 20352
rect 32861 20343 32919 20349
rect 33505 20349 33517 20352
rect 33551 20349 33563 20383
rect 33505 20343 33563 20349
rect 33778 20340 33784 20392
rect 33836 20340 33842 20392
rect 34517 20383 34575 20389
rect 34517 20349 34529 20383
rect 34563 20349 34575 20383
rect 34517 20343 34575 20349
rect 26620 20284 27292 20312
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 18156 20216 19073 20244
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 20622 20244 20628 20256
rect 19392 20216 20628 20244
rect 19392 20204 19398 20216
rect 20622 20204 20628 20216
rect 20680 20244 20686 20256
rect 20901 20247 20959 20253
rect 20901 20244 20913 20247
rect 20680 20216 20913 20244
rect 20680 20204 20686 20216
rect 20901 20213 20913 20216
rect 20947 20213 20959 20247
rect 20901 20207 20959 20213
rect 21174 20204 21180 20256
rect 21232 20204 21238 20256
rect 21634 20204 21640 20256
rect 21692 20204 21698 20256
rect 23750 20204 23756 20256
rect 23808 20204 23814 20256
rect 24210 20204 24216 20256
rect 24268 20204 24274 20256
rect 25314 20204 25320 20256
rect 25372 20244 25378 20256
rect 26620 20244 26648 20284
rect 27264 20253 27292 20284
rect 28644 20284 28948 20312
rect 28644 20256 28672 20284
rect 34330 20272 34336 20324
rect 34388 20312 34394 20324
rect 34532 20312 34560 20343
rect 35986 20340 35992 20392
rect 36044 20340 36050 20392
rect 37458 20340 37464 20392
rect 37516 20340 37522 20392
rect 38120 20389 38148 20420
rect 38381 20417 38393 20451
rect 38427 20448 38439 20451
rect 38427 20420 38700 20448
rect 38427 20417 38439 20420
rect 38381 20411 38439 20417
rect 38672 20392 38700 20420
rect 39298 20408 39304 20460
rect 39356 20408 39362 20460
rect 39574 20408 39580 20460
rect 39632 20408 39638 20460
rect 38013 20383 38071 20389
rect 38013 20349 38025 20383
rect 38059 20349 38071 20383
rect 38013 20343 38071 20349
rect 38105 20383 38163 20389
rect 38105 20349 38117 20383
rect 38151 20380 38163 20383
rect 38194 20380 38200 20392
rect 38151 20352 38200 20380
rect 38151 20349 38163 20352
rect 38105 20343 38163 20349
rect 34388 20284 34560 20312
rect 34388 20272 34394 20284
rect 25372 20216 26648 20244
rect 27249 20247 27307 20253
rect 25372 20204 25378 20216
rect 27249 20213 27261 20247
rect 27295 20244 27307 20247
rect 27338 20244 27344 20256
rect 27295 20216 27344 20244
rect 27295 20213 27307 20216
rect 27249 20207 27307 20213
rect 27338 20204 27344 20216
rect 27396 20204 27402 20256
rect 28626 20204 28632 20256
rect 28684 20204 28690 20256
rect 29546 20204 29552 20256
rect 29604 20204 29610 20256
rect 30098 20204 30104 20256
rect 30156 20244 30162 20256
rect 31018 20244 31024 20256
rect 30156 20216 31024 20244
rect 30156 20204 30162 20216
rect 31018 20204 31024 20216
rect 31076 20244 31082 20256
rect 31205 20247 31263 20253
rect 31205 20244 31217 20247
rect 31076 20216 31217 20244
rect 31076 20204 31082 20216
rect 31205 20213 31217 20216
rect 31251 20213 31263 20247
rect 31205 20207 31263 20213
rect 31846 20204 31852 20256
rect 31904 20204 31910 20256
rect 33318 20204 33324 20256
rect 33376 20244 33382 20256
rect 34425 20247 34483 20253
rect 34425 20244 34437 20247
rect 33376 20216 34437 20244
rect 33376 20204 33382 20216
rect 34425 20213 34437 20216
rect 34471 20213 34483 20247
rect 34532 20244 34560 20284
rect 35452 20284 36952 20312
rect 35452 20244 35480 20284
rect 36924 20256 36952 20284
rect 34532 20216 35480 20244
rect 34425 20207 34483 20213
rect 35894 20204 35900 20256
rect 35952 20204 35958 20256
rect 36906 20204 36912 20256
rect 36964 20204 36970 20256
rect 38028 20244 38056 20343
rect 38194 20340 38200 20352
rect 38252 20340 38258 20392
rect 38286 20340 38292 20392
rect 38344 20340 38350 20392
rect 38562 20340 38568 20392
rect 38620 20340 38626 20392
rect 38654 20340 38660 20392
rect 38712 20340 38718 20392
rect 39418 20383 39476 20389
rect 39418 20380 39430 20383
rect 38764 20352 39430 20380
rect 38304 20312 38332 20340
rect 38764 20312 38792 20352
rect 39418 20349 39430 20352
rect 39464 20349 39476 20383
rect 39418 20343 39476 20349
rect 39942 20340 39948 20392
rect 40000 20380 40006 20392
rect 40880 20389 40908 20488
rect 41414 20476 41420 20488
rect 41472 20476 41478 20528
rect 42058 20476 42064 20528
rect 42116 20516 42122 20528
rect 42797 20519 42855 20525
rect 42797 20516 42809 20519
rect 42116 20488 42809 20516
rect 42116 20476 42122 20488
rect 42797 20485 42809 20488
rect 42843 20485 42855 20519
rect 43898 20516 43904 20528
rect 42797 20479 42855 20485
rect 43364 20488 43904 20516
rect 41132 20451 41190 20457
rect 41132 20417 41144 20451
rect 41178 20448 41190 20451
rect 42334 20448 42340 20460
rect 41178 20420 42340 20448
rect 41178 20417 41190 20420
rect 41132 20411 41190 20417
rect 42334 20408 42340 20420
rect 42392 20408 42398 20460
rect 43162 20408 43168 20460
rect 43220 20448 43226 20460
rect 43364 20457 43392 20488
rect 43898 20476 43904 20488
rect 43956 20476 43962 20528
rect 45646 20476 45652 20528
rect 45704 20476 45710 20528
rect 43349 20451 43407 20457
rect 43349 20448 43361 20451
rect 43220 20420 43361 20448
rect 43220 20408 43226 20420
rect 43349 20417 43361 20420
rect 43395 20417 43407 20451
rect 43349 20411 43407 20417
rect 43616 20451 43674 20457
rect 43616 20417 43628 20451
rect 43662 20448 43674 20451
rect 45664 20448 45692 20476
rect 43662 20420 45692 20448
rect 43662 20417 43674 20420
rect 43616 20411 43674 20417
rect 40865 20383 40923 20389
rect 40865 20380 40877 20383
rect 40000 20352 40877 20380
rect 40000 20340 40006 20352
rect 40865 20349 40877 20352
rect 40911 20349 40923 20383
rect 40865 20343 40923 20349
rect 43070 20340 43076 20392
rect 43128 20340 43134 20392
rect 44910 20340 44916 20392
rect 44968 20340 44974 20392
rect 45462 20340 45468 20392
rect 45520 20380 45526 20392
rect 45756 20389 45784 20556
rect 48222 20544 48228 20556
rect 48280 20544 48286 20596
rect 49510 20544 49516 20596
rect 49568 20544 49574 20596
rect 52733 20587 52791 20593
rect 52733 20553 52745 20587
rect 52779 20584 52791 20587
rect 52914 20584 52920 20596
rect 52779 20556 52920 20584
rect 52779 20553 52791 20556
rect 52733 20547 52791 20553
rect 52914 20544 52920 20556
rect 52972 20544 52978 20596
rect 57698 20544 57704 20596
rect 57756 20544 57762 20596
rect 58158 20544 58164 20596
rect 58216 20544 58222 20596
rect 46284 20519 46342 20525
rect 46284 20485 46296 20519
rect 46330 20516 46342 20519
rect 47210 20516 47216 20528
rect 46330 20488 47216 20516
rect 46330 20485 46342 20488
rect 46284 20479 46342 20485
rect 47210 20476 47216 20488
rect 47268 20476 47274 20528
rect 49881 20519 49939 20525
rect 49881 20485 49893 20519
rect 49927 20516 49939 20519
rect 50985 20519 51043 20525
rect 50985 20516 50997 20519
rect 49927 20488 50997 20516
rect 49927 20485 49939 20488
rect 49881 20479 49939 20485
rect 50985 20485 50997 20488
rect 51031 20485 51043 20519
rect 50985 20479 51043 20485
rect 56873 20519 56931 20525
rect 56873 20485 56885 20519
rect 56919 20516 56931 20519
rect 58176 20516 58204 20544
rect 56919 20488 58204 20516
rect 56919 20485 56931 20488
rect 56873 20479 56931 20485
rect 46017 20451 46075 20457
rect 46017 20417 46029 20451
rect 46063 20448 46075 20451
rect 46106 20448 46112 20460
rect 46063 20420 46112 20448
rect 46063 20417 46075 20420
rect 46017 20411 46075 20417
rect 46106 20408 46112 20420
rect 46164 20408 46170 20460
rect 47578 20408 47584 20460
rect 47636 20408 47642 20460
rect 47670 20408 47676 20460
rect 47728 20448 47734 20460
rect 53101 20451 53159 20457
rect 47728 20420 47900 20448
rect 47728 20408 47734 20420
rect 45741 20383 45799 20389
rect 45741 20380 45753 20383
rect 45520 20352 45753 20380
rect 45520 20340 45526 20352
rect 45741 20349 45753 20352
rect 45787 20349 45799 20383
rect 45741 20343 45799 20349
rect 38304 20284 38792 20312
rect 39022 20272 39028 20324
rect 39080 20272 39086 20324
rect 43088 20312 43116 20340
rect 42168 20284 43116 20312
rect 47397 20315 47455 20321
rect 38838 20244 38844 20256
rect 38028 20216 38844 20244
rect 38838 20204 38844 20216
rect 38896 20204 38902 20256
rect 40218 20204 40224 20256
rect 40276 20204 40282 20256
rect 40770 20204 40776 20256
rect 40828 20244 40834 20256
rect 42168 20244 42196 20284
rect 47397 20281 47409 20315
rect 47443 20312 47455 20315
rect 47688 20312 47716 20408
rect 47765 20383 47823 20389
rect 47765 20349 47777 20383
rect 47811 20349 47823 20383
rect 47872 20380 47900 20420
rect 53101 20417 53113 20451
rect 53147 20448 53159 20451
rect 54297 20451 54355 20457
rect 54297 20448 54309 20451
rect 53147 20420 54309 20448
rect 53147 20417 53159 20420
rect 53101 20411 53159 20417
rect 54297 20417 54309 20420
rect 54343 20417 54355 20451
rect 54297 20411 54355 20417
rect 55033 20451 55091 20457
rect 55033 20417 55045 20451
rect 55079 20448 55091 20451
rect 56137 20451 56195 20457
rect 56137 20448 56149 20451
rect 55079 20420 56149 20448
rect 55079 20417 55091 20420
rect 55033 20411 55091 20417
rect 56137 20417 56149 20420
rect 56183 20417 56195 20451
rect 56137 20411 56195 20417
rect 56410 20408 56416 20460
rect 56468 20408 56474 20460
rect 48501 20383 48559 20389
rect 48501 20380 48513 20383
rect 47872 20352 48513 20380
rect 47765 20343 47823 20349
rect 48501 20349 48513 20352
rect 48547 20349 48559 20383
rect 48501 20343 48559 20349
rect 47443 20284 47716 20312
rect 47443 20281 47455 20284
rect 47397 20275 47455 20281
rect 40828 20216 42196 20244
rect 42245 20247 42303 20253
rect 40828 20204 40834 20216
rect 42245 20213 42257 20247
rect 42291 20244 42303 20247
rect 42702 20244 42708 20256
rect 42291 20216 42708 20244
rect 42291 20213 42303 20216
rect 42245 20207 42303 20213
rect 42702 20204 42708 20216
rect 42760 20244 42766 20256
rect 43622 20244 43628 20256
rect 42760 20216 43628 20244
rect 42760 20204 42766 20216
rect 43622 20204 43628 20216
rect 43680 20204 43686 20256
rect 44726 20204 44732 20256
rect 44784 20204 44790 20256
rect 45094 20204 45100 20256
rect 45152 20244 45158 20256
rect 45465 20247 45523 20253
rect 45465 20244 45477 20247
rect 45152 20216 45477 20244
rect 45152 20204 45158 20216
rect 45465 20213 45477 20216
rect 45511 20213 45523 20247
rect 47780 20244 47808 20343
rect 48590 20340 48596 20392
rect 48648 20389 48654 20392
rect 48648 20383 48676 20389
rect 48664 20349 48676 20383
rect 48648 20343 48676 20349
rect 48648 20340 48654 20343
rect 48774 20340 48780 20392
rect 48832 20340 48838 20392
rect 49970 20340 49976 20392
rect 50028 20340 50034 20392
rect 50154 20340 50160 20392
rect 50212 20380 50218 20392
rect 50212 20352 50292 20380
rect 50212 20340 50218 20352
rect 47854 20272 47860 20324
rect 47912 20312 47918 20324
rect 48225 20315 48283 20321
rect 48225 20312 48237 20315
rect 47912 20284 48237 20312
rect 47912 20272 47918 20284
rect 48225 20281 48237 20284
rect 48271 20312 48283 20315
rect 48314 20312 48320 20324
rect 48271 20284 48320 20312
rect 48271 20281 48283 20284
rect 48225 20275 48283 20281
rect 48314 20272 48320 20284
rect 48372 20272 48378 20324
rect 50264 20312 50292 20352
rect 50430 20340 50436 20392
rect 50488 20340 50494 20392
rect 51258 20340 51264 20392
rect 51316 20380 51322 20392
rect 51353 20383 51411 20389
rect 51353 20380 51365 20383
rect 51316 20352 51365 20380
rect 51316 20340 51322 20352
rect 51353 20349 51365 20352
rect 51399 20349 51411 20383
rect 51353 20343 51411 20349
rect 53190 20340 53196 20392
rect 53248 20340 53254 20392
rect 53377 20383 53435 20389
rect 53377 20349 53389 20383
rect 53423 20349 53435 20383
rect 53377 20343 53435 20349
rect 52549 20315 52607 20321
rect 52549 20312 52561 20315
rect 50264 20284 52561 20312
rect 52549 20281 52561 20284
rect 52595 20312 52607 20315
rect 53392 20312 53420 20343
rect 53742 20340 53748 20392
rect 53800 20340 53806 20392
rect 54846 20340 54852 20392
rect 54904 20380 54910 20392
rect 55125 20383 55183 20389
rect 55125 20380 55137 20383
rect 54904 20352 55137 20380
rect 54904 20340 54910 20352
rect 55125 20349 55137 20352
rect 55171 20349 55183 20383
rect 55125 20343 55183 20349
rect 55214 20340 55220 20392
rect 55272 20340 55278 20392
rect 55582 20340 55588 20392
rect 55640 20380 55646 20392
rect 56428 20380 56456 20408
rect 55640 20352 56456 20380
rect 55640 20340 55646 20352
rect 56888 20312 56916 20479
rect 56962 20408 56968 20460
rect 57020 20448 57026 20460
rect 57057 20451 57115 20457
rect 57057 20448 57069 20451
rect 57020 20420 57069 20448
rect 57020 20408 57026 20420
rect 57057 20417 57069 20420
rect 57103 20417 57115 20451
rect 57057 20411 57115 20417
rect 57606 20408 57612 20460
rect 57664 20448 57670 20460
rect 57885 20451 57943 20457
rect 57885 20448 57897 20451
rect 57664 20420 57897 20448
rect 57664 20408 57670 20420
rect 57885 20417 57897 20420
rect 57931 20417 57943 20451
rect 57885 20411 57943 20417
rect 52595 20284 56916 20312
rect 52595 20281 52607 20284
rect 52549 20275 52607 20281
rect 49326 20244 49332 20256
rect 47780 20216 49332 20244
rect 45465 20207 45523 20213
rect 49326 20204 49332 20216
rect 49384 20204 49390 20256
rect 49421 20247 49479 20253
rect 49421 20213 49433 20247
rect 49467 20244 49479 20247
rect 50062 20244 50068 20256
rect 49467 20216 50068 20244
rect 49467 20213 49479 20216
rect 49421 20207 49479 20213
rect 50062 20204 50068 20216
rect 50120 20204 50126 20256
rect 51994 20204 52000 20256
rect 52052 20204 52058 20256
rect 54662 20204 54668 20256
rect 54720 20204 54726 20256
rect 58529 20247 58587 20253
rect 58529 20213 58541 20247
rect 58575 20244 58587 20247
rect 58575 20216 58940 20244
rect 58575 20213 58587 20216
rect 58529 20207 58587 20213
rect 1104 20154 58880 20176
rect 1104 20102 8172 20154
rect 8224 20102 8236 20154
rect 8288 20102 8300 20154
rect 8352 20102 8364 20154
rect 8416 20102 8428 20154
rect 8480 20102 22616 20154
rect 22668 20102 22680 20154
rect 22732 20102 22744 20154
rect 22796 20102 22808 20154
rect 22860 20102 22872 20154
rect 22924 20102 37060 20154
rect 37112 20102 37124 20154
rect 37176 20102 37188 20154
rect 37240 20102 37252 20154
rect 37304 20102 37316 20154
rect 37368 20102 51504 20154
rect 51556 20102 51568 20154
rect 51620 20102 51632 20154
rect 51684 20102 51696 20154
rect 51748 20102 51760 20154
rect 51812 20102 58880 20154
rect 1104 20080 58880 20102
rect 3142 20000 3148 20052
rect 3200 20040 3206 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3200 20012 3801 20040
rect 3200 20000 3206 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 4982 20000 4988 20052
rect 5040 20000 5046 20052
rect 6362 20000 6368 20052
rect 6420 20000 6426 20052
rect 6638 20000 6644 20052
rect 6696 20000 6702 20052
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 7653 20043 7711 20049
rect 7653 20040 7665 20043
rect 7616 20012 7665 20040
rect 7616 20000 7622 20012
rect 7653 20009 7665 20012
rect 7699 20009 7711 20043
rect 7653 20003 7711 20009
rect 8754 20000 8760 20052
rect 8812 20000 8818 20052
rect 9030 20000 9036 20052
rect 9088 20000 9094 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 9732 20012 11897 20040
rect 9732 20000 9738 20012
rect 11885 20009 11897 20012
rect 11931 20040 11943 20043
rect 12342 20040 12348 20052
rect 11931 20012 12348 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 13814 20040 13820 20052
rect 12544 20012 13820 20040
rect 3421 19975 3479 19981
rect 3421 19941 3433 19975
rect 3467 19972 3479 19975
rect 3510 19972 3516 19984
rect 3467 19944 3516 19972
rect 3467 19941 3479 19944
rect 3421 19935 3479 19941
rect 3510 19932 3516 19944
rect 3568 19972 3574 19984
rect 5000 19972 5028 20000
rect 3568 19944 5028 19972
rect 3568 19932 3574 19944
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 6380 19904 6408 20000
rect 8941 19975 8999 19981
rect 8941 19972 8953 19975
rect 8220 19944 8953 19972
rect 8220 19913 8248 19944
rect 8941 19941 8953 19944
rect 8987 19941 8999 19975
rect 9048 19972 9076 20000
rect 9048 19944 9812 19972
rect 8941 19935 8999 19941
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 4479 19876 4752 19904
rect 6380 19876 6745 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19836 2099 19839
rect 2774 19836 2780 19848
rect 2087 19808 2780 19836
rect 2087 19805 2099 19808
rect 2041 19799 2099 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4522 19836 4528 19848
rect 4203 19808 4528 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4724 19780 4752 19876
rect 6733 19873 6745 19876
rect 6779 19873 6791 19907
rect 6733 19867 6791 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 9585 19907 9643 19913
rect 9585 19873 9597 19907
rect 9631 19904 9643 19907
rect 9674 19904 9680 19916
rect 9631 19876 9680 19904
rect 9631 19873 9643 19876
rect 9585 19867 9643 19873
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 5350 19836 5356 19848
rect 5307 19808 5356 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 6086 19836 6092 19848
rect 5460 19808 6092 19836
rect 2308 19771 2366 19777
rect 2308 19737 2320 19771
rect 2354 19768 2366 19771
rect 2866 19768 2872 19780
rect 2354 19740 2872 19768
rect 2354 19737 2366 19740
rect 2308 19731 2366 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 4706 19728 4712 19780
rect 4764 19768 4770 19780
rect 5460 19768 5488 19808
rect 6086 19796 6092 19808
rect 6144 19836 6150 19848
rect 9600 19836 9628 19867
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 9784 19913 9812 19944
rect 9769 19907 9827 19913
rect 9769 19873 9781 19907
rect 9815 19873 9827 19907
rect 9769 19867 9827 19873
rect 12066 19864 12072 19916
rect 12124 19904 12130 19916
rect 12544 19913 12572 20012
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14918 20000 14924 20052
rect 14976 20040 14982 20052
rect 14976 20012 16712 20040
rect 14976 20000 14982 20012
rect 13909 19975 13967 19981
rect 13909 19941 13921 19975
rect 13955 19972 13967 19975
rect 14090 19972 14096 19984
rect 13955 19944 14096 19972
rect 13955 19941 13967 19944
rect 13909 19935 13967 19941
rect 14090 19932 14096 19944
rect 14148 19972 14154 19984
rect 14148 19944 15056 19972
rect 14148 19932 14154 19944
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 12124 19876 12449 19904
rect 12124 19864 12130 19876
rect 12437 19873 12449 19876
rect 12483 19904 12495 19907
rect 12529 19907 12587 19913
rect 12529 19904 12541 19907
rect 12483 19876 12541 19904
rect 12483 19873 12495 19876
rect 12437 19867 12495 19873
rect 12529 19873 12541 19876
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 14274 19864 14280 19916
rect 14332 19864 14338 19916
rect 14921 19907 14979 19913
rect 14921 19904 14933 19907
rect 14384 19876 14933 19904
rect 6144 19808 9628 19836
rect 10505 19839 10563 19845
rect 6144 19796 6150 19808
rect 10505 19805 10517 19839
rect 10551 19836 10563 19839
rect 12084 19836 12112 19864
rect 10551 19808 12112 19836
rect 10551 19805 10563 19808
rect 10505 19799 10563 19805
rect 4764 19740 5488 19768
rect 5528 19771 5586 19777
rect 4764 19728 4770 19740
rect 5528 19737 5540 19771
rect 5574 19768 5586 19771
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 5574 19740 7389 19768
rect 5574 19737 5586 19740
rect 5528 19731 5586 19737
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7377 19731 7435 19737
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 10413 19771 10471 19777
rect 10413 19768 10425 19771
rect 9355 19740 10425 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 10413 19737 10425 19740
rect 10459 19737 10471 19771
rect 10413 19731 10471 19737
rect 10772 19771 10830 19777
rect 10772 19737 10784 19771
rect 10818 19768 10830 19771
rect 11330 19768 11336 19780
rect 10818 19740 11336 19768
rect 10818 19737 10830 19740
rect 10772 19731 10830 19737
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 12796 19771 12854 19777
rect 12796 19737 12808 19771
rect 12842 19768 12854 19771
rect 13630 19768 13636 19780
rect 12842 19740 13636 19768
rect 12842 19737 12854 19740
rect 12796 19731 12854 19737
rect 13630 19728 13636 19740
rect 13688 19728 13694 19780
rect 4249 19703 4307 19709
rect 4249 19669 4261 19703
rect 4295 19700 4307 19703
rect 4338 19700 4344 19712
rect 4295 19672 4344 19700
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 4982 19660 4988 19712
rect 5040 19700 5046 19712
rect 5077 19703 5135 19709
rect 5077 19700 5089 19703
rect 5040 19672 5089 19700
rect 5040 19660 5046 19672
rect 5077 19669 5089 19672
rect 5123 19700 5135 19703
rect 5258 19700 5264 19712
rect 5123 19672 5264 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 8754 19660 8760 19712
rect 8812 19700 8818 19712
rect 9398 19700 9404 19712
rect 8812 19672 9404 19700
rect 8812 19660 8818 19672
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14384 19700 14412 19876
rect 14921 19873 14933 19876
rect 14967 19873 14979 19907
rect 15028 19904 15056 19944
rect 16684 19913 16712 20012
rect 18690 20000 18696 20052
rect 18748 20040 18754 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 18748 20012 18797 20040
rect 18748 20000 18754 20012
rect 18785 20009 18797 20012
rect 18831 20040 18843 20043
rect 20162 20040 20168 20052
rect 18831 20012 20168 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 21634 20040 21640 20052
rect 21560 20012 21640 20040
rect 18598 19932 18604 19984
rect 18656 19972 18662 19984
rect 18656 19944 20024 19972
rect 18656 19932 18662 19944
rect 15314 19907 15372 19913
rect 15314 19904 15326 19907
rect 15028 19876 15326 19904
rect 14921 19867 14979 19873
rect 15314 19873 15326 19876
rect 15360 19873 15372 19907
rect 15314 19867 15372 19873
rect 16669 19907 16727 19913
rect 16669 19873 16681 19907
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 16850 19864 16856 19916
rect 16908 19864 16914 19916
rect 18432 19876 19656 19904
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 13872 19672 14412 19700
rect 14476 19700 14504 19799
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15470 19796 15476 19848
rect 15528 19796 15534 19848
rect 16574 19796 16580 19848
rect 16632 19796 16638 19848
rect 17310 19796 17316 19848
rect 17368 19836 17374 19848
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 17368 19808 17417 19836
rect 17368 19796 17374 19808
rect 17405 19805 17417 19808
rect 17451 19836 17463 19839
rect 18432 19836 18460 19876
rect 19628 19848 19656 19876
rect 19794 19864 19800 19916
rect 19852 19904 19858 19916
rect 19889 19907 19947 19913
rect 19889 19904 19901 19907
rect 19852 19876 19901 19904
rect 19852 19864 19858 19876
rect 19889 19873 19901 19876
rect 19935 19873 19947 19907
rect 19996 19904 20024 19944
rect 20282 19907 20340 19913
rect 20282 19904 20294 19907
rect 19996 19876 20294 19904
rect 19889 19867 19947 19873
rect 20282 19873 20294 19876
rect 20328 19873 20340 19907
rect 20282 19867 20340 19873
rect 20438 19864 20444 19916
rect 20496 19864 20502 19916
rect 17451 19808 18460 19836
rect 19245 19839 19303 19845
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 19245 19805 19257 19839
rect 19291 19836 19303 19839
rect 19334 19836 19340 19848
rect 19291 19808 19340 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 16482 19768 16488 19780
rect 15948 19740 16488 19768
rect 15948 19700 15976 19740
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 17672 19771 17730 19777
rect 17672 19737 17684 19771
rect 17718 19768 17730 19771
rect 17954 19768 17960 19780
rect 17718 19740 17960 19768
rect 17718 19737 17730 19740
rect 17672 19731 17730 19737
rect 17954 19728 17960 19740
rect 18012 19728 18018 19780
rect 14476 19672 15976 19700
rect 13872 19660 13878 19672
rect 16114 19660 16120 19712
rect 16172 19660 16178 19712
rect 16206 19660 16212 19712
rect 16264 19660 16270 19712
rect 19444 19700 19472 19799
rect 19610 19796 19616 19848
rect 19668 19796 19674 19848
rect 20162 19796 20168 19848
rect 20220 19796 20226 19848
rect 21174 19836 21180 19848
rect 21008 19808 21180 19836
rect 21008 19700 21036 19808
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21560 19845 21588 20012
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 23750 20000 23756 20052
rect 23808 20000 23814 20052
rect 23842 20000 23848 20052
rect 23900 20000 23906 20052
rect 28810 20000 28816 20052
rect 28868 20040 28874 20052
rect 31757 20043 31815 20049
rect 28868 20012 30328 20040
rect 28868 20000 28874 20012
rect 21634 19864 21640 19916
rect 21692 19904 21698 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 21692 19876 21741 19904
rect 21692 19864 21698 19876
rect 21729 19873 21741 19876
rect 21775 19904 21787 19907
rect 23293 19907 23351 19913
rect 21775 19876 23244 19904
rect 21775 19873 21787 19876
rect 21729 19867 21787 19873
rect 21545 19839 21603 19845
rect 21545 19805 21557 19839
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19805 22063 19839
rect 23216 19836 23244 19876
rect 23293 19873 23305 19907
rect 23339 19904 23351 19907
rect 23768 19904 23796 20000
rect 29730 19972 29736 19984
rect 23339 19876 23796 19904
rect 28460 19944 29736 19972
rect 23339 19873 23351 19876
rect 23293 19867 23351 19873
rect 25774 19836 25780 19848
rect 23216 19808 25780 19836
rect 22005 19799 22063 19805
rect 22020 19768 22048 19799
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 27338 19796 27344 19848
rect 27396 19836 27402 19848
rect 27433 19839 27491 19845
rect 27433 19836 27445 19839
rect 27396 19808 27445 19836
rect 27396 19796 27402 19808
rect 27433 19805 27445 19808
rect 27479 19836 27491 19839
rect 28460 19836 28488 19944
rect 29730 19932 29736 19944
rect 29788 19932 29794 19984
rect 29549 19907 29607 19913
rect 29549 19873 29561 19907
rect 29595 19904 29607 19907
rect 30098 19904 30104 19916
rect 29595 19876 30104 19904
rect 29595 19873 29607 19876
rect 29549 19867 29607 19873
rect 30098 19864 30104 19876
rect 30156 19864 30162 19916
rect 30190 19864 30196 19916
rect 30248 19864 30254 19916
rect 30300 19904 30328 20012
rect 31757 20009 31769 20043
rect 31803 20040 31815 20043
rect 31846 20040 31852 20052
rect 31803 20012 31852 20040
rect 31803 20009 31815 20012
rect 31757 20003 31815 20009
rect 31846 20000 31852 20012
rect 31904 20000 31910 20052
rect 33318 20000 33324 20052
rect 33376 20000 33382 20052
rect 33505 20043 33563 20049
rect 33505 20009 33517 20043
rect 33551 20040 33563 20043
rect 33778 20040 33784 20052
rect 33551 20012 33784 20040
rect 33551 20009 33563 20012
rect 33505 20003 33563 20009
rect 33778 20000 33784 20012
rect 33836 20000 33842 20052
rect 35894 20040 35900 20052
rect 34900 20012 35900 20040
rect 30469 19907 30527 19913
rect 30469 19904 30481 19907
rect 30300 19876 30481 19904
rect 30469 19873 30481 19876
rect 30515 19873 30527 19907
rect 30469 19867 30527 19873
rect 30558 19864 30564 19916
rect 30616 19913 30622 19916
rect 30616 19907 30644 19913
rect 30632 19873 30644 19907
rect 30616 19867 30644 19873
rect 30616 19864 30622 19867
rect 30742 19864 30748 19916
rect 30800 19864 30806 19916
rect 30926 19864 30932 19916
rect 30984 19904 30990 19916
rect 30984 19876 31432 19904
rect 30984 19864 30990 19876
rect 27479 19808 28488 19836
rect 27479 19805 27491 19808
rect 27433 19799 27491 19805
rect 28534 19796 28540 19848
rect 28592 19796 28598 19848
rect 31404 19845 31432 19876
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 31389 19839 31447 19845
rect 31389 19805 31401 19839
rect 31435 19805 31447 19839
rect 31389 19799 31447 19805
rect 32033 19839 32091 19845
rect 32033 19805 32045 19839
rect 32079 19805 32091 19839
rect 32033 19799 32091 19805
rect 32300 19839 32358 19845
rect 32300 19805 32312 19839
rect 32346 19836 32358 19839
rect 33336 19836 33364 20000
rect 33413 19975 33471 19981
rect 33413 19941 33425 19975
rect 33459 19972 33471 19975
rect 33594 19972 33600 19984
rect 33459 19944 33600 19972
rect 33459 19941 33471 19944
rect 33413 19935 33471 19941
rect 33594 19932 33600 19944
rect 33652 19972 33658 19984
rect 33652 19944 34836 19972
rect 33652 19932 33658 19944
rect 34146 19864 34152 19916
rect 34204 19904 34210 19916
rect 34204 19876 34652 19904
rect 34204 19864 34210 19876
rect 32346 19808 33364 19836
rect 32346 19805 32358 19808
rect 32300 19799 32358 19805
rect 21192 19740 22048 19768
rect 27700 19771 27758 19777
rect 19444 19672 21036 19700
rect 21082 19660 21088 19712
rect 21140 19660 21146 19712
rect 21192 19709 21220 19740
rect 27700 19737 27712 19771
rect 27746 19768 27758 19771
rect 28552 19768 28580 19796
rect 27746 19740 28580 19768
rect 27746 19737 27758 19740
rect 27700 19731 27758 19737
rect 21177 19703 21235 19709
rect 21177 19669 21189 19703
rect 21223 19669 21235 19703
rect 21177 19663 21235 19669
rect 21634 19660 21640 19712
rect 21692 19660 21698 19712
rect 22646 19660 22652 19712
rect 22704 19660 22710 19712
rect 24210 19660 24216 19712
rect 24268 19660 24274 19712
rect 28994 19660 29000 19712
rect 29052 19700 29058 19712
rect 29273 19703 29331 19709
rect 29273 19700 29285 19703
rect 29052 19672 29285 19700
rect 29052 19660 29058 19672
rect 29273 19669 29285 19672
rect 29319 19669 29331 19703
rect 29748 19700 29776 19799
rect 32048 19768 32076 19799
rect 34330 19768 34336 19780
rect 32048 19740 34336 19768
rect 34330 19728 34336 19740
rect 34388 19728 34394 19780
rect 31202 19700 31208 19712
rect 29748 19672 31208 19700
rect 29273 19663 29331 19669
rect 31202 19660 31208 19672
rect 31260 19660 31266 19712
rect 33870 19660 33876 19712
rect 33928 19660 33934 19712
rect 33962 19660 33968 19712
rect 34020 19700 34026 19712
rect 34422 19700 34428 19712
rect 34020 19672 34428 19700
rect 34020 19660 34026 19672
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 34624 19700 34652 19876
rect 34698 19796 34704 19848
rect 34756 19796 34762 19848
rect 34808 19836 34836 19944
rect 34900 19913 34928 20012
rect 35894 20000 35900 20012
rect 35952 20000 35958 20052
rect 38286 20000 38292 20052
rect 38344 20040 38350 20052
rect 38381 20043 38439 20049
rect 38381 20040 38393 20043
rect 38344 20012 38393 20040
rect 38344 20000 38350 20012
rect 38381 20009 38393 20012
rect 38427 20009 38439 20043
rect 38381 20003 38439 20009
rect 38933 20043 38991 20049
rect 38933 20009 38945 20043
rect 38979 20040 38991 20043
rect 40034 20040 40040 20052
rect 38979 20012 40040 20040
rect 38979 20009 38991 20012
rect 38933 20003 38991 20009
rect 40034 20000 40040 20012
rect 40092 20000 40098 20052
rect 44726 20040 44732 20052
rect 42904 20012 44732 20040
rect 34992 19944 35480 19972
rect 34885 19907 34943 19913
rect 34885 19873 34897 19907
rect 34931 19873 34943 19907
rect 34885 19867 34943 19873
rect 34992 19836 35020 19944
rect 35342 19864 35348 19916
rect 35400 19864 35406 19916
rect 35452 19904 35480 19944
rect 38212 19944 39620 19972
rect 38212 19916 38240 19944
rect 35738 19907 35796 19913
rect 35738 19904 35750 19907
rect 35452 19876 35750 19904
rect 35738 19873 35750 19876
rect 35784 19873 35796 19907
rect 35738 19867 35796 19873
rect 38194 19864 38200 19916
rect 38252 19864 38258 19916
rect 39022 19864 39028 19916
rect 39080 19904 39086 19916
rect 39485 19907 39543 19913
rect 39485 19904 39497 19907
rect 39080 19876 39497 19904
rect 39080 19864 39086 19876
rect 39485 19873 39497 19876
rect 39531 19873 39543 19907
rect 39592 19904 39620 19944
rect 42153 19907 42211 19913
rect 42153 19904 42165 19907
rect 39592 19876 39988 19904
rect 39485 19867 39543 19873
rect 34808 19808 35020 19836
rect 35618 19796 35624 19848
rect 35676 19796 35682 19848
rect 35894 19796 35900 19848
rect 35952 19796 35958 19848
rect 36906 19796 36912 19848
rect 36964 19836 36970 19848
rect 37001 19839 37059 19845
rect 37001 19836 37013 19839
rect 36964 19808 37013 19836
rect 36964 19796 36970 19808
rect 37001 19805 37013 19808
rect 37047 19836 37059 19839
rect 38749 19839 38807 19845
rect 38749 19836 38761 19839
rect 37047 19808 38761 19836
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 38749 19805 38761 19808
rect 38795 19836 38807 19839
rect 39853 19839 39911 19845
rect 39853 19836 39865 19839
rect 38795 19808 39865 19836
rect 38795 19805 38807 19808
rect 38749 19799 38807 19805
rect 39853 19805 39865 19808
rect 39899 19805 39911 19839
rect 39960 19836 39988 19876
rect 41386 19876 42165 19904
rect 41386 19836 41414 19876
rect 42153 19873 42165 19876
rect 42199 19904 42211 19907
rect 42521 19907 42579 19913
rect 42521 19904 42533 19907
rect 42199 19876 42533 19904
rect 42199 19873 42211 19876
rect 42153 19867 42211 19873
rect 42521 19873 42533 19876
rect 42567 19873 42579 19907
rect 42521 19867 42579 19873
rect 42610 19864 42616 19916
rect 42668 19904 42674 19916
rect 42904 19913 42932 20012
rect 44726 20000 44732 20012
rect 44784 20000 44790 20052
rect 44910 20000 44916 20052
rect 44968 20040 44974 20052
rect 45005 20043 45063 20049
rect 45005 20040 45017 20043
rect 44968 20012 45017 20040
rect 44968 20000 44974 20012
rect 45005 20009 45017 20012
rect 45051 20009 45063 20043
rect 48498 20040 48504 20052
rect 45005 20003 45063 20009
rect 48332 20012 48504 20040
rect 42996 19944 43484 19972
rect 42889 19907 42947 19913
rect 42668 19876 42840 19904
rect 42668 19864 42674 19876
rect 39960 19808 41414 19836
rect 42705 19839 42763 19845
rect 39853 19799 39911 19805
rect 42705 19805 42717 19839
rect 42751 19805 42763 19839
rect 42812 19836 42840 19876
rect 42889 19873 42901 19907
rect 42935 19873 42947 19907
rect 42889 19867 42947 19873
rect 42996 19836 43024 19944
rect 43254 19864 43260 19916
rect 43312 19904 43318 19916
rect 43349 19907 43407 19913
rect 43349 19904 43361 19907
rect 43312 19876 43361 19904
rect 43312 19864 43318 19876
rect 43349 19873 43361 19876
rect 43395 19873 43407 19907
rect 43456 19904 43484 19944
rect 43742 19907 43800 19913
rect 43742 19904 43754 19907
rect 43456 19876 43754 19904
rect 43349 19867 43407 19873
rect 43742 19873 43754 19876
rect 43788 19873 43800 19907
rect 43742 19867 43800 19873
rect 43901 19907 43959 19913
rect 43901 19873 43913 19907
rect 43947 19904 43959 19907
rect 44082 19904 44088 19916
rect 43947 19876 44088 19904
rect 43947 19873 43959 19876
rect 43901 19867 43959 19873
rect 44082 19864 44088 19876
rect 44140 19904 44146 19916
rect 44634 19904 44640 19916
rect 44140 19876 44640 19904
rect 44140 19864 44146 19876
rect 44634 19864 44640 19876
rect 44692 19864 44698 19916
rect 45462 19864 45468 19916
rect 45520 19904 45526 19916
rect 45557 19907 45615 19913
rect 45557 19904 45569 19907
rect 45520 19876 45569 19904
rect 45520 19864 45526 19876
rect 45557 19873 45569 19876
rect 45603 19873 45615 19907
rect 45557 19867 45615 19873
rect 46934 19864 46940 19916
rect 46992 19904 46998 19916
rect 48332 19913 48360 20012
rect 48498 20000 48504 20012
rect 48556 20000 48562 20052
rect 49694 20000 49700 20052
rect 49752 20000 49758 20052
rect 51994 20000 52000 20052
rect 52052 20000 52058 20052
rect 54662 20000 54668 20052
rect 54720 20000 54726 20052
rect 55030 20000 55036 20052
rect 55088 20000 55094 20052
rect 57054 20000 57060 20052
rect 57112 20040 57118 20052
rect 58253 20043 58311 20049
rect 58253 20040 58265 20043
rect 57112 20012 58265 20040
rect 57112 20000 57118 20012
rect 58253 20009 58265 20012
rect 58299 20009 58311 20043
rect 58253 20003 58311 20009
rect 47949 19907 48007 19913
rect 47949 19904 47961 19907
rect 46992 19876 47961 19904
rect 46992 19864 46998 19876
rect 47949 19873 47961 19876
rect 47995 19873 48007 19907
rect 47949 19867 48007 19873
rect 48317 19907 48375 19913
rect 48317 19873 48329 19907
rect 48363 19873 48375 19907
rect 49712 19904 49740 20000
rect 48317 19867 48375 19873
rect 49344 19876 49740 19904
rect 42812 19808 43024 19836
rect 42705 19799 42763 19805
rect 36817 19771 36875 19777
rect 36817 19768 36829 19771
rect 36464 19740 36829 19768
rect 36464 19700 36492 19740
rect 36817 19737 36829 19740
rect 36863 19737 36875 19771
rect 36817 19731 36875 19737
rect 37268 19771 37326 19777
rect 37268 19737 37280 19771
rect 37314 19768 37326 19771
rect 38102 19768 38108 19780
rect 37314 19740 38108 19768
rect 37314 19737 37326 19740
rect 37268 19731 37326 19737
rect 34624 19672 36492 19700
rect 36538 19660 36544 19712
rect 36596 19660 36602 19712
rect 36832 19700 36860 19731
rect 38102 19728 38108 19740
rect 38160 19728 38166 19780
rect 39393 19771 39451 19777
rect 39393 19768 39405 19771
rect 38856 19740 39405 19768
rect 38856 19712 38884 19740
rect 39393 19737 39405 19740
rect 39439 19737 39451 19771
rect 39868 19768 39896 19799
rect 39942 19768 39948 19780
rect 39868 19740 39948 19768
rect 39393 19731 39451 19737
rect 39942 19728 39948 19740
rect 40000 19728 40006 19780
rect 40120 19771 40178 19777
rect 40120 19737 40132 19771
rect 40166 19768 40178 19771
rect 41046 19768 41052 19780
rect 40166 19740 41052 19768
rect 40166 19737 40178 19740
rect 40120 19731 40178 19737
rect 41046 19728 41052 19740
rect 41104 19728 41110 19780
rect 37458 19700 37464 19712
rect 36832 19672 37464 19700
rect 37458 19660 37464 19672
rect 37516 19660 37522 19712
rect 38838 19660 38844 19712
rect 38896 19660 38902 19712
rect 39298 19660 39304 19712
rect 39356 19660 39362 19712
rect 39574 19660 39580 19712
rect 39632 19700 39638 19712
rect 41233 19703 41291 19709
rect 41233 19700 41245 19703
rect 39632 19672 41245 19700
rect 39632 19660 39638 19672
rect 41233 19669 41245 19672
rect 41279 19669 41291 19703
rect 41233 19663 41291 19669
rect 41506 19660 41512 19712
rect 41564 19660 41570 19712
rect 41782 19660 41788 19712
rect 41840 19700 41846 19712
rect 41877 19703 41935 19709
rect 41877 19700 41889 19703
rect 41840 19672 41889 19700
rect 41840 19660 41846 19672
rect 41877 19669 41889 19672
rect 41923 19669 41935 19703
rect 41877 19663 41935 19669
rect 41969 19703 42027 19709
rect 41969 19669 41981 19703
rect 42015 19700 42027 19703
rect 42058 19700 42064 19712
rect 42015 19672 42064 19700
rect 42015 19669 42027 19672
rect 41969 19663 42027 19669
rect 42058 19660 42064 19672
rect 42116 19660 42122 19712
rect 42720 19700 42748 19799
rect 43622 19796 43628 19848
rect 43680 19796 43686 19848
rect 45925 19839 45983 19845
rect 45925 19805 45937 19839
rect 45971 19836 45983 19839
rect 45971 19808 46152 19836
rect 45971 19805 45983 19808
rect 45925 19799 45983 19805
rect 46124 19712 46152 19808
rect 47302 19796 47308 19848
rect 47360 19836 47366 19848
rect 47857 19839 47915 19845
rect 47857 19836 47869 19839
rect 47360 19808 47869 19836
rect 47360 19796 47366 19808
rect 47857 19805 47869 19808
rect 47903 19805 47915 19839
rect 47857 19799 47915 19805
rect 48584 19839 48642 19845
rect 48584 19805 48596 19839
rect 48630 19836 48642 19839
rect 49344 19836 49372 19876
rect 48630 19808 49372 19836
rect 48630 19805 48642 19808
rect 48584 19799 48642 19805
rect 49602 19796 49608 19848
rect 49660 19836 49666 19848
rect 50893 19839 50951 19845
rect 50893 19836 50905 19839
rect 49660 19808 50905 19836
rect 49660 19796 49666 19808
rect 50893 19805 50905 19808
rect 50939 19836 50951 19839
rect 51160 19839 51218 19845
rect 50939 19808 51074 19836
rect 50939 19805 50951 19808
rect 50893 19799 50951 19805
rect 46192 19771 46250 19777
rect 46192 19737 46204 19771
rect 46238 19768 46250 19771
rect 47210 19768 47216 19780
rect 46238 19740 47216 19768
rect 46238 19737 46250 19740
rect 46192 19731 46250 19737
rect 47210 19728 47216 19740
rect 47268 19728 47274 19780
rect 47320 19740 48636 19768
rect 43990 19700 43996 19712
rect 42720 19672 43996 19700
rect 43990 19660 43996 19672
rect 44048 19660 44054 19712
rect 44174 19660 44180 19712
rect 44232 19700 44238 19712
rect 44545 19703 44603 19709
rect 44545 19700 44557 19703
rect 44232 19672 44557 19700
rect 44232 19660 44238 19672
rect 44545 19669 44557 19672
rect 44591 19669 44603 19703
rect 44545 19663 44603 19669
rect 44910 19660 44916 19712
rect 44968 19700 44974 19712
rect 45373 19703 45431 19709
rect 45373 19700 45385 19703
rect 44968 19672 45385 19700
rect 44968 19660 44974 19672
rect 45373 19669 45385 19672
rect 45419 19669 45431 19703
rect 45373 19663 45431 19669
rect 45462 19660 45468 19712
rect 45520 19660 45526 19712
rect 46106 19660 46112 19712
rect 46164 19660 46170 19712
rect 47320 19709 47348 19740
rect 48608 19712 48636 19740
rect 49326 19728 49332 19780
rect 49384 19768 49390 19780
rect 50430 19768 50436 19780
rect 49384 19740 50436 19768
rect 49384 19728 49390 19740
rect 47305 19703 47363 19709
rect 47305 19669 47317 19703
rect 47351 19669 47363 19703
rect 47305 19663 47363 19669
rect 47394 19660 47400 19712
rect 47452 19660 47458 19712
rect 47762 19660 47768 19712
rect 47820 19660 47826 19712
rect 48590 19660 48596 19712
rect 48648 19660 48654 19712
rect 49712 19709 49740 19740
rect 50430 19728 50436 19740
rect 50488 19728 50494 19780
rect 49697 19703 49755 19709
rect 49697 19669 49709 19703
rect 49743 19669 49755 19703
rect 51046 19700 51074 19808
rect 51160 19805 51172 19839
rect 51206 19836 51218 19839
rect 52012 19836 52040 20000
rect 52273 19975 52331 19981
rect 52273 19941 52285 19975
rect 52319 19972 52331 19975
rect 52319 19944 52408 19972
rect 52319 19941 52331 19944
rect 52273 19935 52331 19941
rect 52380 19913 52408 19944
rect 52365 19907 52423 19913
rect 52365 19873 52377 19907
rect 52411 19904 52423 19907
rect 52454 19904 52460 19916
rect 52411 19876 52460 19904
rect 52411 19873 52423 19876
rect 52365 19867 52423 19873
rect 52454 19864 52460 19876
rect 52512 19864 52518 19916
rect 54481 19907 54539 19913
rect 54481 19873 54493 19907
rect 54527 19904 54539 19907
rect 54680 19904 54708 20000
rect 54527 19876 54708 19904
rect 54527 19873 54539 19876
rect 54481 19867 54539 19873
rect 51206 19808 52040 19836
rect 51206 19805 51218 19808
rect 51160 19799 51218 19805
rect 56502 19796 56508 19848
rect 56560 19836 56566 19848
rect 56873 19839 56931 19845
rect 56873 19836 56885 19839
rect 56560 19808 56885 19836
rect 56560 19796 56566 19808
rect 56873 19805 56885 19808
rect 56919 19805 56931 19839
rect 56873 19799 56931 19805
rect 57140 19839 57198 19845
rect 57140 19805 57152 19839
rect 57186 19836 57198 19839
rect 58912 19836 58940 20216
rect 57186 19808 58940 19836
rect 57186 19805 57198 19808
rect 57140 19799 57198 19805
rect 51350 19700 51356 19712
rect 51046 19672 51356 19700
rect 49697 19663 49755 19669
rect 51350 19660 51356 19672
rect 51408 19660 51414 19712
rect 53006 19660 53012 19712
rect 53064 19660 53070 19712
rect 53926 19660 53932 19712
rect 53984 19700 53990 19712
rect 54205 19703 54263 19709
rect 54205 19700 54217 19703
rect 53984 19672 54217 19700
rect 53984 19660 53990 19672
rect 54205 19669 54217 19672
rect 54251 19700 54263 19703
rect 55122 19700 55128 19712
rect 54251 19672 55128 19700
rect 54251 19669 54263 19672
rect 54205 19663 54263 19669
rect 55122 19660 55128 19672
rect 55180 19660 55186 19712
rect 1104 19610 59040 19632
rect 1104 19558 15394 19610
rect 15446 19558 15458 19610
rect 15510 19558 15522 19610
rect 15574 19558 15586 19610
rect 15638 19558 15650 19610
rect 15702 19558 29838 19610
rect 29890 19558 29902 19610
rect 29954 19558 29966 19610
rect 30018 19558 30030 19610
rect 30082 19558 30094 19610
rect 30146 19558 44282 19610
rect 44334 19558 44346 19610
rect 44398 19558 44410 19610
rect 44462 19558 44474 19610
rect 44526 19558 44538 19610
rect 44590 19558 58726 19610
rect 58778 19558 58790 19610
rect 58842 19558 58854 19610
rect 58906 19558 58918 19610
rect 58970 19558 58982 19610
rect 59034 19558 59040 19610
rect 1104 19536 59040 19558
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 4065 19499 4123 19505
rect 4065 19496 4077 19499
rect 3384 19468 4077 19496
rect 3384 19456 3390 19468
rect 4065 19465 4077 19468
rect 4111 19465 4123 19499
rect 4065 19459 4123 19465
rect 4706 19456 4712 19508
rect 4764 19456 4770 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 6788 19468 7021 19496
rect 6788 19456 6794 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 7282 19456 7288 19508
rect 7340 19456 7346 19508
rect 11330 19456 11336 19508
rect 11388 19456 11394 19508
rect 16482 19456 16488 19508
rect 16540 19456 16546 19508
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 18693 19499 18751 19505
rect 18693 19496 18705 19499
rect 18288 19468 18705 19496
rect 18288 19456 18294 19468
rect 18693 19465 18705 19468
rect 18739 19465 18751 19499
rect 18693 19459 18751 19465
rect 21174 19456 21180 19508
rect 21232 19456 21238 19508
rect 22646 19456 22652 19508
rect 22704 19456 22710 19508
rect 27338 19456 27344 19508
rect 27396 19456 27402 19508
rect 28626 19456 28632 19508
rect 28684 19456 28690 19508
rect 28994 19456 29000 19508
rect 29052 19456 29058 19508
rect 29089 19499 29147 19505
rect 29089 19465 29101 19499
rect 29135 19496 29147 19499
rect 29546 19496 29552 19508
rect 29135 19468 29552 19496
rect 29135 19465 29147 19468
rect 29089 19459 29147 19465
rect 29546 19456 29552 19468
rect 29604 19456 29610 19508
rect 31202 19456 31208 19508
rect 31260 19456 31266 19508
rect 33686 19456 33692 19508
rect 33744 19496 33750 19508
rect 33744 19468 34652 19496
rect 33744 19456 33750 19468
rect 3510 19320 3516 19372
rect 3568 19320 3574 19372
rect 6457 19363 6515 19369
rect 6457 19329 6469 19363
rect 6503 19360 6515 19363
rect 6638 19360 6644 19372
rect 6503 19332 6644 19360
rect 6503 19329 6515 19332
rect 6457 19323 6515 19329
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 7300 19292 7328 19456
rect 11977 19431 12035 19437
rect 11977 19428 11989 19431
rect 11808 19400 11989 19428
rect 11808 19372 11836 19400
rect 11977 19397 11989 19400
rect 12023 19397 12035 19431
rect 11977 19391 12035 19397
rect 13633 19431 13691 19437
rect 13633 19397 13645 19431
rect 13679 19428 13691 19431
rect 13722 19428 13728 19440
rect 13679 19400 13728 19428
rect 13679 19397 13691 19400
rect 13633 19391 13691 19397
rect 13722 19388 13728 19400
rect 13780 19428 13786 19440
rect 14918 19428 14924 19440
rect 13780 19400 14924 19428
rect 13780 19388 13786 19400
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 15010 19388 15016 19440
rect 15068 19428 15074 19440
rect 17488 19431 17546 19437
rect 15068 19400 17172 19428
rect 15068 19388 15074 19400
rect 10704 19332 10916 19360
rect 10704 19292 10732 19332
rect 7300 19264 10732 19292
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19261 10839 19295
rect 10888 19292 10916 19332
rect 11790 19320 11796 19372
rect 11848 19320 11854 19372
rect 15120 19369 15148 19400
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 11931 19332 13001 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19360 13599 19363
rect 14645 19363 14703 19369
rect 14645 19360 14657 19363
rect 13587 19332 14657 19360
rect 13587 19329 13599 19332
rect 13541 19323 13599 19329
rect 14645 19329 14657 19332
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15372 19363 15430 19369
rect 15372 19329 15384 19363
rect 15418 19360 15430 19363
rect 16942 19360 16948 19372
rect 15418 19332 16948 19360
rect 15418 19329 15430 19332
rect 15372 19323 15430 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 17144 19369 17172 19400
rect 17488 19397 17500 19431
rect 17534 19428 17546 19431
rect 18782 19428 18788 19440
rect 17534 19400 18788 19428
rect 17534 19397 17546 19400
rect 17488 19391 17546 19397
rect 18782 19388 18788 19400
rect 18840 19388 18846 19440
rect 20064 19431 20122 19437
rect 20064 19397 20076 19431
rect 20110 19428 20122 19431
rect 22664 19428 22692 19456
rect 20110 19400 22692 19428
rect 20110 19397 20122 19400
rect 20064 19391 20122 19397
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19360 17187 19363
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17175 19332 17233 19360
rect 17175 19329 17187 19332
rect 17129 19323 17187 19329
rect 17221 19329 17233 19332
rect 17267 19360 17279 19363
rect 17310 19360 17316 19372
rect 17267 19332 17316 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 19058 19320 19064 19372
rect 19116 19320 19122 19372
rect 19150 19320 19156 19372
rect 19208 19360 19214 19372
rect 19208 19332 19380 19360
rect 19208 19320 19214 19332
rect 19352 19304 19380 19332
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 19668 19332 19809 19360
rect 19668 19320 19674 19332
rect 19797 19329 19809 19332
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 27249 19363 27307 19369
rect 27249 19329 27261 19363
rect 27295 19360 27307 19363
rect 27356 19360 27384 19456
rect 29012 19428 29040 19456
rect 30190 19428 30196 19440
rect 29012 19400 30196 19428
rect 30190 19388 30196 19400
rect 30248 19388 30254 19440
rect 27295 19332 27384 19360
rect 27516 19363 27574 19369
rect 27295 19329 27307 19332
rect 27249 19323 27307 19329
rect 27516 19329 27528 19363
rect 27562 19360 27574 19363
rect 28810 19360 28816 19372
rect 27562 19332 28816 19360
rect 27562 19329 27574 19332
rect 27516 19323 27574 19329
rect 28810 19320 28816 19332
rect 28868 19320 28874 19372
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19360 29239 19363
rect 29227 19332 29500 19360
rect 29227 19329 29239 19332
rect 29181 19323 29239 19329
rect 29472 19304 29500 19332
rect 29730 19320 29736 19372
rect 29788 19360 29794 19372
rect 29825 19363 29883 19369
rect 29825 19360 29837 19363
rect 29788 19332 29837 19360
rect 29788 19320 29794 19332
rect 29825 19329 29837 19332
rect 29871 19329 29883 19363
rect 29825 19323 29883 19329
rect 30092 19363 30150 19369
rect 30092 19329 30104 19363
rect 30138 19360 30150 19363
rect 30834 19360 30840 19372
rect 30138 19332 30840 19360
rect 30138 19329 30150 19332
rect 30092 19323 30150 19329
rect 30834 19320 30840 19332
rect 30892 19320 30898 19372
rect 31220 19360 31248 19456
rect 34624 19428 34652 19468
rect 34698 19456 34704 19508
rect 34756 19496 34762 19508
rect 35713 19499 35771 19505
rect 35713 19496 35725 19499
rect 34756 19468 35725 19496
rect 34756 19456 34762 19468
rect 35713 19465 35725 19468
rect 35759 19465 35771 19499
rect 35713 19459 35771 19465
rect 35805 19499 35863 19505
rect 35805 19465 35817 19499
rect 35851 19496 35863 19499
rect 35986 19496 35992 19508
rect 35851 19468 35992 19496
rect 35851 19465 35863 19468
rect 35805 19459 35863 19465
rect 35618 19428 35624 19440
rect 32508 19400 34100 19428
rect 34624 19400 35624 19428
rect 31297 19363 31355 19369
rect 31297 19360 31309 19363
rect 31220 19332 31309 19360
rect 31297 19329 31309 19332
rect 31343 19329 31355 19363
rect 31297 19323 31355 19329
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19360 32367 19363
rect 32508 19360 32536 19400
rect 32355 19332 32536 19360
rect 32576 19363 32634 19369
rect 32355 19329 32367 19332
rect 32309 19323 32367 19329
rect 32576 19329 32588 19363
rect 32622 19360 32634 19363
rect 33410 19360 33416 19372
rect 32622 19332 33416 19360
rect 32622 19329 32634 19332
rect 32576 19323 32634 19329
rect 33410 19320 33416 19332
rect 33468 19320 33474 19372
rect 34072 19369 34100 19400
rect 35618 19388 35624 19400
rect 35676 19388 35682 19440
rect 35728 19428 35756 19459
rect 35986 19456 35992 19468
rect 36044 19456 36050 19508
rect 36173 19499 36231 19505
rect 36173 19465 36185 19499
rect 36219 19496 36231 19499
rect 36722 19496 36728 19508
rect 36219 19468 36728 19496
rect 36219 19465 36231 19468
rect 36173 19459 36231 19465
rect 36722 19456 36728 19468
rect 36780 19456 36786 19508
rect 36906 19456 36912 19508
rect 36964 19456 36970 19508
rect 39298 19456 39304 19508
rect 39356 19496 39362 19508
rect 40221 19499 40279 19505
rect 40221 19496 40233 19499
rect 39356 19468 40233 19496
rect 39356 19456 39362 19468
rect 40221 19465 40233 19468
rect 40267 19465 40279 19499
rect 40221 19459 40279 19465
rect 41782 19456 41788 19508
rect 41840 19456 41846 19508
rect 42058 19456 42064 19508
rect 42116 19496 42122 19508
rect 42116 19468 43392 19496
rect 42116 19456 42122 19468
rect 36262 19428 36268 19440
rect 35728 19400 36268 19428
rect 36262 19388 36268 19400
rect 36320 19388 36326 19440
rect 41800 19428 41828 19456
rect 43073 19431 43131 19437
rect 43073 19428 43085 19431
rect 41800 19400 43085 19428
rect 43073 19397 43085 19400
rect 43119 19397 43131 19431
rect 43073 19391 43131 19397
rect 34057 19363 34115 19369
rect 34057 19329 34069 19363
rect 34103 19360 34115 19363
rect 34330 19360 34336 19372
rect 34103 19332 34336 19360
rect 34103 19329 34115 19332
rect 34057 19323 34115 19329
rect 34330 19320 34336 19332
rect 34388 19320 34394 19372
rect 34600 19363 34658 19369
rect 34600 19329 34612 19363
rect 34646 19360 34658 19363
rect 36170 19360 36176 19372
rect 34646 19332 36176 19360
rect 34646 19329 34658 19332
rect 34600 19323 34658 19329
rect 36170 19320 36176 19332
rect 36228 19320 36234 19372
rect 38654 19320 38660 19372
rect 38712 19320 38718 19372
rect 38749 19363 38807 19369
rect 38749 19329 38761 19363
rect 38795 19360 38807 19363
rect 39942 19360 39948 19372
rect 38795 19332 39948 19360
rect 38795 19329 38807 19332
rect 38749 19323 38807 19329
rect 39942 19320 39948 19332
rect 40000 19360 40006 19372
rect 40773 19363 40831 19369
rect 40773 19360 40785 19363
rect 40000 19332 40785 19360
rect 40000 19320 40006 19332
rect 40773 19329 40785 19332
rect 40819 19329 40831 19363
rect 40773 19323 40831 19329
rect 41040 19363 41098 19369
rect 41040 19329 41052 19363
rect 41086 19360 41098 19363
rect 41966 19360 41972 19372
rect 41086 19332 41972 19360
rect 41086 19329 41098 19332
rect 41040 19323 41098 19329
rect 41966 19320 41972 19332
rect 42024 19320 42030 19372
rect 42521 19363 42579 19369
rect 42521 19329 42533 19363
rect 42567 19360 42579 19363
rect 42610 19360 42616 19372
rect 42567 19332 42616 19360
rect 42567 19329 42579 19332
rect 42521 19323 42579 19329
rect 11146 19292 11152 19304
rect 10888 19264 11152 19292
rect 10781 19255 10839 19261
rect 9858 19224 9864 19236
rect 9508 19196 9864 19224
rect 9508 19168 9536 19196
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 10796 19224 10824 19255
rect 11146 19252 11152 19264
rect 11204 19292 11210 19304
rect 12069 19295 12127 19301
rect 12069 19292 12081 19295
rect 11204 19264 12081 19292
rect 11204 19252 11210 19264
rect 12069 19261 12081 19264
rect 12115 19292 12127 19295
rect 12158 19292 12164 19304
rect 12115 19264 12164 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12342 19252 12348 19304
rect 12400 19252 12406 19304
rect 13725 19295 13783 19301
rect 13725 19261 13737 19295
rect 13771 19261 13783 19295
rect 13725 19255 13783 19261
rect 11517 19227 11575 19233
rect 11517 19224 11529 19227
rect 10796 19196 11529 19224
rect 11517 19193 11529 19196
rect 11563 19193 11575 19227
rect 12894 19224 12900 19236
rect 11517 19187 11575 19193
rect 12406 19196 12900 19224
rect 6178 19116 6184 19168
rect 6236 19116 6242 19168
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19156 9275 19159
rect 9490 19156 9496 19168
rect 9263 19128 9496 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9732 19128 9781 19156
rect 9732 19116 9738 19128
rect 9769 19125 9781 19128
rect 9815 19156 9827 19159
rect 12406 19156 12434 19196
rect 12894 19184 12900 19196
rect 12952 19224 12958 19236
rect 13740 19224 13768 19255
rect 14090 19252 14096 19304
rect 14148 19252 14154 19304
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 12952 19196 13768 19224
rect 12952 19184 12958 19196
rect 9815 19128 12434 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 13173 19159 13231 19165
rect 13173 19156 13185 19159
rect 13136 19128 13185 19156
rect 13136 19116 13142 19128
rect 13173 19125 13185 19128
rect 13219 19125 13231 19159
rect 13740 19156 13768 19196
rect 18598 19184 18604 19236
rect 18656 19184 18662 19236
rect 17402 19156 17408 19168
rect 13740 19128 17408 19156
rect 13173 19119 13231 19125
rect 17402 19116 17408 19128
rect 17460 19156 17466 19168
rect 18690 19156 18696 19168
rect 17460 19128 18696 19156
rect 17460 19116 17466 19128
rect 18690 19116 18696 19128
rect 18748 19156 18754 19168
rect 19260 19156 19288 19255
rect 19334 19252 19340 19304
rect 19392 19252 19398 19304
rect 23474 19252 23480 19304
rect 23532 19252 23538 19304
rect 29270 19252 29276 19304
rect 29328 19252 29334 19304
rect 29454 19252 29460 19304
rect 29512 19252 29518 19304
rect 36265 19295 36323 19301
rect 36265 19261 36277 19295
rect 36311 19261 36323 19295
rect 36265 19255 36323 19261
rect 36449 19295 36507 19301
rect 36449 19261 36461 19295
rect 36495 19261 36507 19295
rect 38672 19292 38700 19320
rect 39574 19292 39580 19304
rect 38672 19264 39580 19292
rect 36449 19255 36507 19261
rect 23492 19224 23520 19252
rect 20732 19196 23520 19224
rect 20732 19156 20760 19196
rect 18748 19128 20760 19156
rect 18748 19116 18754 19128
rect 21542 19116 21548 19168
rect 21600 19116 21606 19168
rect 28718 19116 28724 19168
rect 28776 19116 28782 19168
rect 31938 19116 31944 19168
rect 31996 19116 32002 19168
rect 34514 19116 34520 19168
rect 34572 19156 34578 19168
rect 36280 19156 36308 19255
rect 36464 19224 36492 19255
rect 39574 19252 39580 19264
rect 39632 19252 39638 19304
rect 37553 19227 37611 19233
rect 37553 19224 37565 19227
rect 36464 19196 37565 19224
rect 37553 19193 37565 19196
rect 37599 19224 37611 19227
rect 42153 19227 42211 19233
rect 37599 19196 38424 19224
rect 37599 19193 37611 19196
rect 37553 19187 37611 19193
rect 38396 19168 38424 19196
rect 42153 19193 42165 19227
rect 42199 19224 42211 19227
rect 42536 19224 42564 19323
rect 42610 19320 42616 19332
rect 42668 19320 42674 19372
rect 43162 19320 43168 19372
rect 43220 19320 43226 19372
rect 43364 19360 43392 19468
rect 43990 19456 43996 19508
rect 44048 19496 44054 19508
rect 44542 19496 44548 19508
rect 44048 19468 44548 19496
rect 44048 19456 44054 19468
rect 44542 19456 44548 19468
rect 44600 19456 44606 19508
rect 44637 19499 44695 19505
rect 44637 19465 44649 19499
rect 44683 19496 44695 19499
rect 45002 19496 45008 19508
rect 44683 19468 45008 19496
rect 44683 19465 44695 19468
rect 44637 19459 44695 19465
rect 45002 19456 45008 19468
rect 45060 19456 45066 19508
rect 45094 19456 45100 19508
rect 45152 19456 45158 19508
rect 45370 19456 45376 19508
rect 45428 19456 45434 19508
rect 45462 19456 45468 19508
rect 45520 19456 45526 19508
rect 46106 19456 46112 19508
rect 46164 19496 46170 19508
rect 46477 19499 46535 19505
rect 46477 19496 46489 19499
rect 46164 19468 46489 19496
rect 46164 19456 46170 19468
rect 46477 19465 46489 19468
rect 46523 19496 46535 19499
rect 48498 19496 48504 19508
rect 46523 19468 48504 19496
rect 46523 19465 46535 19468
rect 46477 19459 46535 19465
rect 48498 19456 48504 19468
rect 48556 19456 48562 19508
rect 51258 19456 51264 19508
rect 51316 19496 51322 19508
rect 51445 19499 51503 19505
rect 51445 19496 51457 19499
rect 51316 19468 51457 19496
rect 51316 19456 51322 19468
rect 51445 19465 51457 19468
rect 51491 19465 51503 19499
rect 51445 19459 51503 19465
rect 51813 19499 51871 19505
rect 51813 19465 51825 19499
rect 51859 19496 51871 19499
rect 53006 19496 53012 19508
rect 51859 19468 53012 19496
rect 51859 19465 51871 19468
rect 51813 19459 51871 19465
rect 53006 19456 53012 19468
rect 53064 19456 53070 19508
rect 56594 19456 56600 19508
rect 56652 19496 56658 19508
rect 56965 19499 57023 19505
rect 56965 19496 56977 19499
rect 56652 19468 56977 19496
rect 56652 19456 56658 19468
rect 56965 19465 56977 19468
rect 57011 19465 57023 19499
rect 56965 19459 57023 19465
rect 57333 19499 57391 19505
rect 57333 19465 57345 19499
rect 57379 19496 57391 19499
rect 57514 19496 57520 19508
rect 57379 19468 57520 19496
rect 57379 19465 57391 19468
rect 57333 19459 57391 19465
rect 57514 19456 57520 19468
rect 57572 19456 57578 19508
rect 43432 19431 43490 19437
rect 43432 19397 43444 19431
rect 43478 19428 43490 19431
rect 45112 19428 45140 19456
rect 43478 19400 45140 19428
rect 43478 19397 43490 19400
rect 43432 19391 43490 19397
rect 44910 19360 44916 19372
rect 43364 19332 44916 19360
rect 44910 19320 44916 19332
rect 44968 19320 44974 19372
rect 45005 19363 45063 19369
rect 45005 19329 45017 19363
rect 45051 19360 45063 19363
rect 45388 19360 45416 19456
rect 45051 19332 45416 19360
rect 45480 19360 45508 19456
rect 47210 19388 47216 19440
rect 47268 19428 47274 19440
rect 47268 19400 47716 19428
rect 47268 19388 47274 19400
rect 46109 19363 46167 19369
rect 46109 19360 46121 19363
rect 45480 19332 46121 19360
rect 45051 19329 45063 19332
rect 45005 19323 45063 19329
rect 46109 19329 46121 19332
rect 46155 19329 46167 19363
rect 46109 19323 46167 19329
rect 47394 19320 47400 19372
rect 47452 19360 47458 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 47452 19332 47593 19360
rect 47452 19320 47458 19332
rect 47581 19329 47593 19332
rect 47627 19329 47639 19363
rect 47688 19360 47716 19400
rect 47762 19388 47768 19440
rect 47820 19428 47826 19440
rect 48961 19431 49019 19437
rect 48961 19428 48973 19431
rect 47820 19400 48973 19428
rect 47820 19388 47826 19400
rect 48961 19397 48973 19400
rect 49007 19397 49019 19431
rect 48961 19391 49019 19397
rect 48225 19363 48283 19369
rect 48225 19360 48237 19363
rect 47688 19332 48237 19360
rect 47581 19323 47639 19329
rect 48225 19329 48237 19332
rect 48271 19329 48283 19363
rect 48225 19323 48283 19329
rect 48409 19363 48467 19369
rect 48409 19329 48421 19363
rect 48455 19360 48467 19363
rect 48590 19360 48596 19372
rect 48455 19332 48596 19360
rect 48455 19329 48467 19332
rect 48409 19323 48467 19329
rect 48590 19320 48596 19332
rect 48648 19320 48654 19372
rect 48682 19320 48688 19372
rect 48740 19320 48746 19372
rect 51905 19363 51963 19369
rect 51905 19329 51917 19363
rect 51951 19360 51963 19363
rect 52086 19360 52092 19372
rect 51951 19332 52092 19360
rect 51951 19329 51963 19332
rect 51905 19323 51963 19329
rect 52086 19320 52092 19332
rect 52144 19360 52150 19372
rect 53006 19360 53012 19372
rect 52144 19332 53012 19360
rect 52144 19320 52150 19332
rect 53006 19320 53012 19332
rect 53064 19360 53070 19372
rect 53190 19360 53196 19372
rect 53064 19332 53196 19360
rect 53064 19320 53070 19332
rect 53190 19320 53196 19332
rect 53248 19320 53254 19372
rect 58158 19320 58164 19372
rect 58216 19360 58222 19372
rect 58529 19363 58587 19369
rect 58529 19360 58541 19363
rect 58216 19332 58541 19360
rect 58216 19320 58222 19332
rect 58529 19329 58541 19332
rect 58575 19329 58587 19363
rect 58529 19323 58587 19329
rect 44542 19252 44548 19304
rect 44600 19252 44606 19304
rect 44928 19292 44956 19320
rect 45097 19295 45155 19301
rect 45097 19292 45109 19295
rect 44928 19264 45109 19292
rect 45097 19261 45109 19264
rect 45143 19261 45155 19295
rect 45097 19255 45155 19261
rect 45186 19252 45192 19304
rect 45244 19252 45250 19304
rect 45557 19295 45615 19301
rect 45557 19261 45569 19295
rect 45603 19261 45615 19295
rect 45557 19255 45615 19261
rect 42199 19196 42564 19224
rect 44560 19224 44588 19252
rect 45572 19224 45600 19255
rect 48406 19224 48412 19236
rect 44560 19196 45600 19224
rect 45848 19196 48412 19224
rect 42199 19193 42211 19196
rect 42153 19187 42211 19193
rect 34572 19128 36308 19156
rect 34572 19116 34578 19128
rect 38286 19116 38292 19168
rect 38344 19116 38350 19168
rect 38378 19116 38384 19168
rect 38436 19156 38442 19168
rect 39022 19156 39028 19168
rect 38436 19128 39028 19156
rect 38436 19116 38442 19128
rect 39022 19116 39028 19128
rect 39080 19116 39086 19168
rect 45186 19116 45192 19168
rect 45244 19156 45250 19168
rect 45848 19156 45876 19196
rect 48406 19184 48412 19196
rect 48464 19224 48470 19236
rect 48700 19224 48728 19320
rect 50522 19252 50528 19304
rect 50580 19252 50586 19304
rect 51997 19295 52055 19301
rect 51997 19292 52009 19295
rect 51046 19264 52009 19292
rect 48464 19196 48728 19224
rect 48464 19184 48470 19196
rect 45244 19128 45876 19156
rect 45244 19116 45250 19128
rect 46934 19116 46940 19168
rect 46992 19156 46998 19168
rect 47213 19159 47271 19165
rect 47213 19156 47225 19159
rect 46992 19128 47225 19156
rect 46992 19116 46998 19128
rect 47213 19125 47225 19128
rect 47259 19156 47271 19159
rect 50341 19159 50399 19165
rect 50341 19156 50353 19159
rect 47259 19128 50353 19156
rect 47259 19125 47271 19128
rect 47213 19119 47271 19125
rect 50341 19125 50353 19128
rect 50387 19156 50399 19159
rect 51046 19156 51074 19264
rect 51997 19261 52009 19264
rect 52043 19292 52055 19295
rect 53926 19292 53932 19304
rect 52043 19264 53932 19292
rect 52043 19261 52055 19264
rect 51997 19255 52055 19261
rect 53926 19252 53932 19264
rect 53984 19252 53990 19304
rect 54018 19252 54024 19304
rect 54076 19252 54082 19304
rect 57422 19252 57428 19304
rect 57480 19252 57486 19304
rect 57517 19295 57575 19301
rect 57517 19261 57529 19295
rect 57563 19261 57575 19295
rect 57517 19255 57575 19261
rect 57885 19295 57943 19301
rect 57885 19261 57897 19295
rect 57931 19261 57943 19295
rect 57885 19255 57943 19261
rect 57532 19224 57560 19255
rect 56796 19196 57560 19224
rect 56796 19168 56824 19196
rect 57900 19168 57928 19255
rect 50387 19128 51074 19156
rect 50387 19125 50399 19128
rect 50341 19119 50399 19125
rect 51166 19116 51172 19168
rect 51224 19116 51230 19168
rect 54570 19116 54576 19168
rect 54628 19116 54634 19168
rect 56778 19116 56784 19168
rect 56836 19116 56842 19168
rect 57882 19116 57888 19168
rect 57940 19116 57946 19168
rect 1104 19066 58880 19088
rect 1104 19014 8172 19066
rect 8224 19014 8236 19066
rect 8288 19014 8300 19066
rect 8352 19014 8364 19066
rect 8416 19014 8428 19066
rect 8480 19014 22616 19066
rect 22668 19014 22680 19066
rect 22732 19014 22744 19066
rect 22796 19014 22808 19066
rect 22860 19014 22872 19066
rect 22924 19014 37060 19066
rect 37112 19014 37124 19066
rect 37176 19014 37188 19066
rect 37240 19014 37252 19066
rect 37304 19014 37316 19066
rect 37368 19014 51504 19066
rect 51556 19014 51568 19066
rect 51620 19014 51632 19066
rect 51684 19014 51696 19066
rect 51748 19014 51760 19066
rect 51812 19014 58880 19066
rect 1104 18992 58880 19014
rect 12066 18912 12072 18964
rect 12124 18912 12130 18964
rect 12894 18912 12900 18964
rect 12952 18912 12958 18964
rect 13630 18912 13636 18964
rect 13688 18912 13694 18964
rect 14921 18955 14979 18961
rect 14921 18921 14933 18955
rect 14967 18952 14979 18955
rect 15010 18952 15016 18964
rect 14967 18924 15016 18952
rect 14967 18921 14979 18924
rect 14921 18915 14979 18921
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 16850 18912 16856 18964
rect 16908 18912 16914 18964
rect 16942 18912 16948 18964
rect 17000 18912 17006 18964
rect 18325 18955 18383 18961
rect 18325 18921 18337 18955
rect 18371 18952 18383 18955
rect 18690 18952 18696 18964
rect 18371 18924 18696 18952
rect 18371 18921 18383 18924
rect 18325 18915 18383 18921
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 19058 18912 19064 18964
rect 19116 18912 19122 18964
rect 19886 18912 19892 18964
rect 19944 18912 19950 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 24210 18952 24216 18964
rect 23532 18924 24216 18952
rect 23532 18912 23538 18924
rect 24210 18912 24216 18924
rect 24268 18952 24274 18964
rect 24268 18924 26234 18952
rect 24268 18912 24274 18924
rect 12158 18844 12164 18896
rect 12216 18884 12222 18896
rect 12437 18887 12495 18893
rect 12437 18884 12449 18887
rect 12216 18856 12449 18884
rect 12216 18844 12222 18856
rect 12437 18853 12449 18856
rect 12483 18884 12495 18887
rect 16868 18884 16896 18912
rect 24762 18884 24768 18896
rect 12483 18856 16896 18884
rect 20456 18856 24768 18884
rect 12483 18853 12495 18856
rect 12437 18847 12495 18853
rect 13078 18776 13084 18828
rect 13136 18776 13142 18828
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18816 14427 18819
rect 15286 18816 15292 18828
rect 14415 18788 15292 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 16206 18776 16212 18828
rect 16264 18816 16270 18828
rect 20456 18825 20484 18856
rect 24762 18844 24768 18856
rect 24820 18844 24826 18896
rect 26206 18884 26234 18924
rect 28810 18912 28816 18964
rect 28868 18912 28874 18964
rect 29270 18912 29276 18964
rect 29328 18912 29334 18964
rect 30834 18912 30840 18964
rect 30892 18952 30898 18964
rect 31665 18955 31723 18961
rect 31665 18952 31677 18955
rect 30892 18924 31677 18952
rect 30892 18912 30898 18924
rect 31665 18921 31677 18924
rect 31711 18921 31723 18955
rect 31665 18915 31723 18921
rect 33597 18955 33655 18961
rect 33597 18921 33609 18955
rect 33643 18952 33655 18955
rect 34330 18952 34336 18964
rect 33643 18924 34336 18952
rect 33643 18921 33655 18924
rect 33597 18915 33655 18921
rect 34330 18912 34336 18924
rect 34388 18912 34394 18964
rect 36170 18912 36176 18964
rect 36228 18912 36234 18964
rect 41046 18912 41052 18964
rect 41104 18912 41110 18964
rect 41966 18912 41972 18964
rect 42024 18912 42030 18964
rect 42337 18955 42395 18961
rect 42337 18921 42349 18955
rect 42383 18952 42395 18955
rect 43073 18955 43131 18961
rect 43073 18952 43085 18955
rect 42383 18924 43085 18952
rect 42383 18921 42395 18924
rect 42337 18915 42395 18921
rect 43073 18921 43085 18924
rect 43119 18952 43131 18955
rect 43162 18952 43168 18964
rect 43119 18924 43168 18952
rect 43119 18921 43131 18924
rect 43073 18915 43131 18921
rect 43162 18912 43168 18924
rect 43220 18912 43226 18964
rect 44545 18955 44603 18961
rect 44545 18921 44557 18955
rect 44591 18952 44603 18955
rect 45094 18952 45100 18964
rect 44591 18924 45100 18952
rect 44591 18921 44603 18924
rect 44545 18915 44603 18921
rect 45094 18912 45100 18924
rect 45152 18912 45158 18964
rect 48409 18955 48467 18961
rect 48409 18921 48421 18955
rect 48455 18952 48467 18955
rect 48498 18952 48504 18964
rect 48455 18924 48504 18952
rect 48455 18921 48467 18924
rect 48409 18915 48467 18921
rect 48498 18912 48504 18924
rect 48556 18912 48562 18964
rect 50157 18955 50215 18961
rect 50157 18921 50169 18955
rect 50203 18952 50215 18955
rect 50522 18952 50528 18964
rect 50203 18924 50528 18952
rect 50203 18921 50215 18924
rect 50157 18915 50215 18921
rect 50522 18912 50528 18924
rect 50580 18912 50586 18964
rect 54018 18912 54024 18964
rect 54076 18952 54082 18964
rect 54113 18955 54171 18961
rect 54113 18952 54125 18955
rect 54076 18924 54125 18952
rect 54076 18912 54082 18924
rect 54113 18921 54125 18924
rect 54159 18921 54171 18955
rect 57882 18952 57888 18964
rect 54113 18915 54171 18921
rect 55692 18924 57888 18952
rect 27709 18887 27767 18893
rect 27709 18884 27721 18887
rect 26206 18856 27721 18884
rect 27709 18853 27721 18856
rect 27755 18884 27767 18887
rect 29288 18884 29316 18912
rect 55692 18896 55720 18924
rect 57882 18912 57888 18924
rect 57940 18912 57946 18964
rect 27755 18856 29316 18884
rect 30193 18887 30251 18893
rect 27755 18853 27767 18856
rect 27709 18847 27767 18853
rect 30193 18853 30205 18887
rect 30239 18884 30251 18887
rect 30239 18856 31064 18884
rect 30239 18853 30251 18856
rect 30193 18847 30251 18853
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 16264 18788 16313 18816
rect 16264 18776 16270 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 18509 18819 18567 18825
rect 18509 18785 18521 18819
rect 18555 18785 18567 18819
rect 20441 18819 20499 18825
rect 20441 18816 20453 18819
rect 18509 18779 18567 18785
rect 19720 18788 20453 18816
rect 3050 18708 3056 18760
rect 3108 18708 3114 18760
rect 4246 18708 4252 18760
rect 4304 18708 4310 18760
rect 8938 18708 8944 18760
rect 8996 18708 9002 18760
rect 18524 18748 18552 18779
rect 18598 18748 18604 18760
rect 18524 18720 18604 18748
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 9030 18640 9036 18692
rect 9088 18680 9094 18692
rect 9088 18652 9996 18680
rect 9088 18640 9094 18652
rect 3602 18572 3608 18624
rect 3660 18572 3666 18624
rect 4798 18572 4804 18624
rect 4856 18572 4862 18624
rect 5074 18572 5080 18624
rect 5132 18612 5138 18624
rect 5261 18615 5319 18621
rect 5261 18612 5273 18615
rect 5132 18584 5273 18612
rect 5132 18572 5138 18584
rect 5261 18581 5273 18584
rect 5307 18581 5319 18615
rect 5261 18575 5319 18581
rect 5997 18615 6055 18621
rect 5997 18581 6009 18615
rect 6043 18612 6055 18615
rect 6178 18612 6184 18624
rect 6043 18584 6184 18612
rect 6043 18581 6055 18584
rect 5997 18575 6055 18581
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 8018 18572 8024 18624
rect 8076 18612 8082 18624
rect 9968 18621 9996 18652
rect 9585 18615 9643 18621
rect 9585 18612 9597 18615
rect 8076 18584 9597 18612
rect 8076 18572 8082 18584
rect 9585 18581 9597 18584
rect 9631 18581 9643 18615
rect 9585 18575 9643 18581
rect 9953 18615 10011 18621
rect 9953 18581 9965 18615
rect 9999 18612 10011 18615
rect 12710 18612 12716 18624
rect 9999 18584 12716 18612
rect 9999 18581 10011 18584
rect 9953 18575 10011 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 19720 18621 19748 18788
rect 20441 18785 20453 18788
rect 20487 18785 20499 18819
rect 20441 18779 20499 18785
rect 21266 18776 21272 18828
rect 21324 18776 21330 18828
rect 25685 18819 25743 18825
rect 25685 18785 25697 18819
rect 25731 18816 25743 18819
rect 26421 18819 26479 18825
rect 26421 18816 26433 18819
rect 25731 18788 26433 18816
rect 25731 18785 25743 18788
rect 25685 18779 25743 18785
rect 26421 18785 26433 18788
rect 26467 18816 26479 18819
rect 27062 18816 27068 18828
rect 26467 18788 27068 18816
rect 26467 18785 26479 18788
rect 26421 18779 26479 18785
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 28261 18819 28319 18825
rect 28261 18785 28273 18819
rect 28307 18816 28319 18819
rect 28718 18816 28724 18828
rect 28307 18788 28724 18816
rect 28307 18785 28319 18788
rect 28261 18779 28319 18785
rect 28718 18776 28724 18788
rect 28776 18776 28782 18828
rect 30101 18819 30159 18825
rect 30101 18785 30113 18819
rect 30147 18816 30159 18819
rect 30650 18816 30656 18828
rect 30147 18788 30656 18816
rect 30147 18785 30159 18788
rect 30101 18779 30159 18785
rect 30650 18776 30656 18788
rect 30708 18816 30714 18828
rect 31036 18825 31064 18856
rect 33870 18844 33876 18896
rect 33928 18844 33934 18896
rect 34701 18887 34759 18893
rect 34701 18853 34713 18887
rect 34747 18884 34759 18887
rect 38381 18887 38439 18893
rect 34747 18856 35572 18884
rect 34747 18853 34759 18856
rect 34701 18847 34759 18853
rect 30745 18819 30803 18825
rect 30745 18816 30757 18819
rect 30708 18788 30757 18816
rect 30708 18776 30714 18788
rect 30745 18785 30757 18788
rect 30791 18785 30803 18819
rect 30745 18779 30803 18785
rect 31021 18819 31079 18825
rect 31021 18785 31033 18819
rect 31067 18785 31079 18819
rect 31021 18779 31079 18785
rect 33594 18776 33600 18828
rect 33652 18816 33658 18828
rect 33689 18819 33747 18825
rect 33689 18816 33701 18819
rect 33652 18788 33701 18816
rect 33652 18776 33658 18788
rect 33689 18785 33701 18788
rect 33735 18785 33747 18819
rect 33888 18816 33916 18844
rect 35544 18825 35572 18856
rect 38381 18853 38393 18887
rect 38427 18884 38439 18887
rect 38654 18884 38660 18896
rect 38427 18856 38660 18884
rect 38427 18853 38439 18856
rect 38381 18847 38439 18853
rect 38654 18844 38660 18856
rect 38712 18844 38718 18896
rect 43254 18844 43260 18896
rect 43312 18884 43318 18896
rect 45189 18887 45247 18893
rect 45189 18884 45201 18887
rect 43312 18856 45201 18884
rect 43312 18844 43318 18856
rect 45189 18853 45201 18856
rect 45235 18884 45247 18887
rect 45922 18884 45928 18896
rect 45235 18856 45928 18884
rect 45235 18853 45247 18856
rect 45189 18847 45247 18853
rect 45922 18844 45928 18856
rect 45980 18844 45986 18896
rect 55674 18844 55680 18896
rect 55732 18844 55738 18896
rect 34333 18819 34391 18825
rect 34333 18816 34345 18819
rect 33888 18788 34345 18816
rect 33689 18779 33747 18785
rect 34333 18785 34345 18788
rect 34379 18785 34391 18819
rect 34333 18779 34391 18785
rect 35345 18819 35403 18825
rect 35345 18785 35357 18819
rect 35391 18785 35403 18819
rect 35345 18779 35403 18785
rect 35529 18819 35587 18825
rect 35529 18785 35541 18819
rect 35575 18785 35587 18819
rect 35529 18779 35587 18785
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18748 20407 18751
rect 21284 18748 21312 18776
rect 20395 18720 21312 18748
rect 20395 18717 20407 18720
rect 20349 18711 20407 18717
rect 22738 18708 22744 18760
rect 22796 18708 22802 18760
rect 23566 18708 23572 18760
rect 23624 18708 23630 18760
rect 26142 18708 26148 18760
rect 26200 18708 26206 18760
rect 26602 18708 26608 18760
rect 26660 18708 26666 18760
rect 30561 18751 30619 18757
rect 30561 18717 30573 18751
rect 30607 18748 30619 18751
rect 31938 18748 31944 18760
rect 30607 18720 31944 18748
rect 30607 18717 30619 18720
rect 30561 18711 30619 18717
rect 31938 18708 31944 18720
rect 31996 18708 32002 18760
rect 35360 18748 35388 18779
rect 35894 18776 35900 18828
rect 35952 18776 35958 18828
rect 36262 18776 36268 18828
rect 36320 18776 36326 18828
rect 36906 18776 36912 18828
rect 36964 18816 36970 18828
rect 37001 18819 37059 18825
rect 37001 18816 37013 18819
rect 36964 18788 37013 18816
rect 36964 18776 36970 18788
rect 37001 18785 37013 18788
rect 37047 18785 37059 18819
rect 37001 18779 37059 18785
rect 38286 18776 38292 18828
rect 38344 18816 38350 18828
rect 39117 18819 39175 18825
rect 39117 18816 39129 18819
rect 38344 18788 39129 18816
rect 38344 18776 38350 18788
rect 39117 18785 39129 18788
rect 39163 18816 39175 18819
rect 39163 18788 39252 18816
rect 39163 18785 39175 18788
rect 39117 18779 39175 18785
rect 35912 18748 35940 18776
rect 35360 18720 35940 18748
rect 35161 18683 35219 18689
rect 35161 18649 35173 18683
rect 35207 18680 35219 18683
rect 36909 18683 36967 18689
rect 36909 18680 36921 18683
rect 35207 18652 36921 18680
rect 35207 18649 35219 18652
rect 35161 18643 35219 18649
rect 36909 18649 36921 18652
rect 36955 18649 36967 18683
rect 36909 18643 36967 18649
rect 37268 18683 37326 18689
rect 37268 18649 37280 18683
rect 37314 18680 37326 18683
rect 38562 18680 38568 18692
rect 37314 18652 38568 18680
rect 37314 18649 37326 18652
rect 37268 18643 37326 18649
rect 38562 18640 38568 18652
rect 38620 18640 38626 18692
rect 19705 18615 19763 18621
rect 19705 18612 19717 18615
rect 19484 18584 19717 18612
rect 19484 18572 19490 18584
rect 19705 18581 19717 18584
rect 19751 18581 19763 18615
rect 19705 18575 19763 18581
rect 20257 18615 20315 18621
rect 20257 18581 20269 18615
rect 20303 18612 20315 18615
rect 20346 18612 20352 18624
rect 20303 18584 20352 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20346 18572 20352 18584
rect 20404 18612 20410 18624
rect 21634 18612 21640 18624
rect 20404 18584 21640 18612
rect 20404 18572 20410 18584
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 23290 18572 23296 18624
rect 23348 18572 23354 18624
rect 24118 18572 24124 18624
rect 24176 18572 24182 18624
rect 25777 18615 25835 18621
rect 25777 18581 25789 18615
rect 25823 18612 25835 18615
rect 26050 18612 26056 18624
rect 25823 18584 26056 18612
rect 25823 18581 25835 18584
rect 25777 18575 25835 18581
rect 26050 18572 26056 18584
rect 26108 18572 26114 18624
rect 26234 18572 26240 18624
rect 26292 18572 26298 18624
rect 27246 18572 27252 18624
rect 27304 18572 27310 18624
rect 28074 18572 28080 18624
rect 28132 18572 28138 18624
rect 29086 18572 29092 18624
rect 29144 18572 29150 18624
rect 30374 18572 30380 18624
rect 30432 18612 30438 18624
rect 30653 18615 30711 18621
rect 30653 18612 30665 18615
rect 30432 18584 30665 18612
rect 30432 18572 30438 18584
rect 30653 18581 30665 18584
rect 30699 18581 30711 18615
rect 30653 18575 30711 18581
rect 34422 18572 34428 18624
rect 34480 18612 34486 18624
rect 34882 18612 34888 18624
rect 34480 18584 34888 18612
rect 34480 18572 34486 18584
rect 34882 18572 34888 18584
rect 34940 18612 34946 18624
rect 35069 18615 35127 18621
rect 35069 18612 35081 18615
rect 34940 18584 35081 18612
rect 34940 18572 34946 18584
rect 35069 18581 35081 18584
rect 35115 18581 35127 18615
rect 35069 18575 35127 18581
rect 38470 18572 38476 18624
rect 38528 18572 38534 18624
rect 38838 18572 38844 18624
rect 38896 18572 38902 18624
rect 38930 18572 38936 18624
rect 38988 18572 38994 18624
rect 39224 18612 39252 18788
rect 40034 18776 40040 18828
rect 40092 18816 40098 18828
rect 40405 18819 40463 18825
rect 40405 18816 40417 18819
rect 40092 18788 40417 18816
rect 40092 18776 40098 18788
rect 40405 18785 40417 18788
rect 40451 18785 40463 18819
rect 40405 18779 40463 18785
rect 41325 18819 41383 18825
rect 41325 18785 41337 18819
rect 41371 18816 41383 18819
rect 41506 18816 41512 18828
rect 41371 18788 41512 18816
rect 41371 18785 41383 18788
rect 41325 18779 41383 18785
rect 41506 18776 41512 18788
rect 41564 18776 41570 18828
rect 49973 18819 50031 18825
rect 49973 18785 49985 18819
rect 50019 18816 50031 18819
rect 50706 18816 50712 18828
rect 50019 18788 50712 18816
rect 50019 18785 50031 18788
rect 49973 18779 50031 18785
rect 50706 18776 50712 18788
rect 50764 18776 50770 18828
rect 54665 18819 54723 18825
rect 54665 18816 54677 18819
rect 54036 18788 54677 18816
rect 47486 18708 47492 18760
rect 47544 18708 47550 18760
rect 50982 18708 50988 18760
rect 51040 18708 51046 18760
rect 52822 18708 52828 18760
rect 52880 18708 52886 18760
rect 50525 18683 50583 18689
rect 50525 18649 50537 18683
rect 50571 18680 50583 18683
rect 51629 18683 51687 18689
rect 51629 18680 51641 18683
rect 50571 18652 51641 18680
rect 50571 18649 50583 18652
rect 50525 18643 50583 18649
rect 51629 18649 51641 18652
rect 51675 18649 51687 18683
rect 51629 18643 51687 18649
rect 54036 18624 54064 18788
rect 54665 18785 54677 18788
rect 54711 18785 54723 18819
rect 54665 18779 54723 18785
rect 55401 18819 55459 18825
rect 55401 18785 55413 18819
rect 55447 18816 55459 18819
rect 55447 18788 56640 18816
rect 55447 18785 55459 18788
rect 55401 18779 55459 18785
rect 56042 18708 56048 18760
rect 56100 18748 56106 18760
rect 56502 18748 56508 18760
rect 56100 18720 56508 18748
rect 56100 18708 56106 18720
rect 56502 18708 56508 18720
rect 56560 18708 56566 18760
rect 54481 18683 54539 18689
rect 54481 18649 54493 18683
rect 54527 18680 54539 18683
rect 55953 18683 56011 18689
rect 55953 18680 55965 18683
rect 54527 18652 55965 18680
rect 54527 18649 54539 18652
rect 54481 18643 54539 18649
rect 55953 18649 55965 18652
rect 55999 18649 56011 18683
rect 56612 18680 56640 18788
rect 55953 18643 56011 18649
rect 56520 18652 56640 18680
rect 56772 18683 56830 18689
rect 56520 18624 56548 18652
rect 56772 18649 56784 18683
rect 56818 18680 56830 18683
rect 58526 18680 58532 18692
rect 56818 18652 58532 18680
rect 56818 18649 56830 18652
rect 56772 18643 56830 18649
rect 58526 18640 58532 18652
rect 58584 18640 58590 18692
rect 41230 18612 41236 18624
rect 39224 18584 41236 18612
rect 41230 18572 41236 18584
rect 41288 18572 41294 18624
rect 47118 18572 47124 18624
rect 47176 18612 47182 18624
rect 48041 18615 48099 18621
rect 48041 18612 48053 18615
rect 47176 18584 48053 18612
rect 47176 18572 47182 18584
rect 48041 18581 48053 18584
rect 48087 18581 48099 18615
rect 48041 18575 48099 18581
rect 49970 18572 49976 18624
rect 50028 18612 50034 18624
rect 50617 18615 50675 18621
rect 50617 18612 50629 18615
rect 50028 18584 50629 18612
rect 50028 18572 50034 18584
rect 50617 18581 50629 18584
rect 50663 18581 50675 18615
rect 50617 18575 50675 18581
rect 53466 18572 53472 18624
rect 53524 18572 53530 18624
rect 54018 18572 54024 18624
rect 54076 18572 54082 18624
rect 54573 18615 54631 18621
rect 54573 18581 54585 18615
rect 54619 18612 54631 18615
rect 54846 18612 54852 18624
rect 54619 18584 54852 18612
rect 54619 18581 54631 18584
rect 54573 18575 54631 18581
rect 54846 18572 54852 18584
rect 54904 18572 54910 18624
rect 56502 18572 56508 18624
rect 56560 18572 56566 18624
rect 1104 18522 59040 18544
rect 1104 18470 15394 18522
rect 15446 18470 15458 18522
rect 15510 18470 15522 18522
rect 15574 18470 15586 18522
rect 15638 18470 15650 18522
rect 15702 18470 29838 18522
rect 29890 18470 29902 18522
rect 29954 18470 29966 18522
rect 30018 18470 30030 18522
rect 30082 18470 30094 18522
rect 30146 18470 44282 18522
rect 44334 18470 44346 18522
rect 44398 18470 44410 18522
rect 44462 18470 44474 18522
rect 44526 18470 44538 18522
rect 44590 18470 58726 18522
rect 58778 18470 58790 18522
rect 58842 18470 58854 18522
rect 58906 18470 58918 18522
rect 58970 18470 58982 18522
rect 59034 18470 59040 18522
rect 1104 18448 59040 18470
rect 3421 18411 3479 18417
rect 3421 18377 3433 18411
rect 3467 18408 3479 18411
rect 3602 18408 3608 18420
rect 3467 18380 3608 18408
rect 3467 18377 3479 18380
rect 3421 18371 3479 18377
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 4433 18411 4491 18417
rect 4433 18408 4445 18411
rect 4304 18380 4445 18408
rect 4304 18368 4310 18380
rect 4433 18377 4445 18380
rect 4479 18377 4491 18411
rect 4433 18371 4491 18377
rect 8389 18411 8447 18417
rect 8389 18377 8401 18411
rect 8435 18408 8447 18411
rect 8938 18408 8944 18420
rect 8435 18380 8944 18408
rect 8435 18377 8447 18380
rect 8389 18371 8447 18377
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 19610 18368 19616 18420
rect 19668 18368 19674 18420
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 22833 18411 22891 18417
rect 22833 18408 22845 18411
rect 22796 18380 22845 18408
rect 22796 18368 22802 18380
rect 22833 18377 22845 18380
rect 22879 18377 22891 18411
rect 22833 18371 22891 18377
rect 23201 18411 23259 18417
rect 23201 18377 23213 18411
rect 23247 18408 23259 18411
rect 24118 18408 24124 18420
rect 23247 18380 24124 18408
rect 23247 18377 23259 18380
rect 23201 18371 23259 18377
rect 24118 18368 24124 18380
rect 24176 18368 24182 18420
rect 24854 18368 24860 18420
rect 24912 18408 24918 18420
rect 25038 18408 25044 18420
rect 24912 18380 25044 18408
rect 24912 18368 24918 18380
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 27246 18408 27252 18420
rect 26206 18380 27252 18408
rect 4065 18343 4123 18349
rect 4065 18340 4077 18343
rect 3988 18312 4077 18340
rect 3326 18232 3332 18284
rect 3384 18232 3390 18284
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18204 2375 18207
rect 2363 18176 2774 18204
rect 2363 18173 2375 18176
rect 2317 18167 2375 18173
rect 2746 18136 2774 18176
rect 2961 18139 3019 18145
rect 2961 18136 2973 18139
rect 2746 18108 2973 18136
rect 2961 18105 2973 18108
rect 3007 18105 3019 18139
rect 3344 18136 3372 18232
rect 3605 18207 3663 18213
rect 3605 18173 3617 18207
rect 3651 18204 3663 18207
rect 3988 18204 4016 18312
rect 4065 18309 4077 18312
rect 4111 18340 4123 18343
rect 7650 18340 7656 18352
rect 4111 18312 7656 18340
rect 4111 18309 4123 18312
rect 4065 18303 4123 18309
rect 7650 18300 7656 18312
rect 7708 18340 7714 18352
rect 25492 18343 25550 18349
rect 7708 18312 8708 18340
rect 7708 18300 7714 18312
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 3651 18176 4016 18204
rect 4724 18244 4813 18272
rect 3651 18173 3663 18176
rect 3605 18167 3663 18173
rect 4338 18136 4344 18148
rect 3344 18108 4344 18136
rect 2961 18099 3019 18105
rect 4338 18096 4344 18108
rect 4396 18136 4402 18148
rect 4724 18136 4752 18244
rect 4801 18241 4813 18244
rect 4847 18241 4859 18275
rect 4801 18235 4859 18241
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 5905 18275 5963 18281
rect 5905 18272 5917 18275
rect 4939 18244 5917 18272
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 5905 18241 5917 18244
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 5074 18164 5080 18216
rect 5132 18164 5138 18216
rect 5258 18164 5264 18216
rect 5316 18164 5322 18216
rect 6638 18164 6644 18216
rect 6696 18164 6702 18216
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18204 7803 18207
rect 8570 18204 8576 18216
rect 7791 18176 8576 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 8680 18204 8708 18312
rect 25492 18309 25504 18343
rect 25538 18340 25550 18343
rect 26206 18340 26234 18380
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 38470 18368 38476 18420
rect 38528 18368 38534 18420
rect 38562 18368 38568 18420
rect 38620 18368 38626 18420
rect 38930 18368 38936 18420
rect 38988 18408 38994 18420
rect 39301 18411 39359 18417
rect 39301 18408 39313 18411
rect 38988 18380 39313 18408
rect 38988 18368 38994 18380
rect 39301 18377 39313 18380
rect 39347 18377 39359 18411
rect 39301 18371 39359 18377
rect 48314 18368 48320 18420
rect 48372 18408 48378 18420
rect 48501 18411 48559 18417
rect 48501 18408 48513 18411
rect 48372 18380 48513 18408
rect 48372 18368 48378 18380
rect 48501 18377 48513 18380
rect 48547 18408 48559 18411
rect 48682 18408 48688 18420
rect 48547 18380 48688 18408
rect 48547 18377 48559 18380
rect 48501 18371 48559 18377
rect 48682 18368 48688 18380
rect 48740 18408 48746 18420
rect 54849 18411 54907 18417
rect 48740 18380 54800 18408
rect 48740 18368 48746 18380
rect 25538 18312 26234 18340
rect 25538 18309 25550 18312
rect 25492 18303 25550 18309
rect 8754 18232 8760 18284
rect 8812 18232 8818 18284
rect 8849 18275 8907 18281
rect 8849 18241 8861 18275
rect 8895 18272 8907 18275
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 8895 18244 9873 18272
rect 8895 18241 8907 18244
rect 8849 18235 8907 18241
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 25225 18275 25283 18281
rect 23339 18244 24072 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 24044 18216 24072 18244
rect 25225 18241 25237 18275
rect 25271 18272 25283 18275
rect 25314 18272 25320 18284
rect 25271 18244 25320 18272
rect 25271 18241 25283 18244
rect 25225 18235 25283 18241
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 29454 18232 29460 18284
rect 29512 18272 29518 18284
rect 29641 18275 29699 18281
rect 29641 18272 29653 18275
rect 29512 18244 29653 18272
rect 29512 18232 29518 18244
rect 29641 18241 29653 18244
rect 29687 18272 29699 18275
rect 30374 18272 30380 18284
rect 29687 18244 30380 18272
rect 29687 18241 29699 18244
rect 29641 18235 29699 18241
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 38013 18275 38071 18281
rect 38013 18241 38025 18275
rect 38059 18272 38071 18275
rect 38488 18272 38516 18368
rect 47578 18300 47584 18352
rect 47636 18340 47642 18352
rect 48774 18340 48780 18352
rect 47636 18312 48780 18340
rect 47636 18300 47642 18312
rect 48774 18300 48780 18312
rect 48832 18340 48838 18352
rect 49326 18340 49332 18352
rect 48832 18312 49332 18340
rect 48832 18300 48838 18312
rect 49326 18300 49332 18312
rect 49384 18300 49390 18352
rect 49872 18343 49930 18349
rect 49872 18309 49884 18343
rect 49918 18340 49930 18343
rect 51166 18340 51172 18352
rect 49918 18312 51172 18340
rect 49918 18309 49930 18312
rect 49872 18303 49930 18309
rect 51166 18300 51172 18312
rect 51224 18300 51230 18352
rect 53736 18343 53794 18349
rect 53736 18309 53748 18343
rect 53782 18340 53794 18343
rect 54570 18340 54576 18352
rect 53782 18312 54576 18340
rect 53782 18309 53794 18312
rect 53736 18303 53794 18309
rect 54570 18300 54576 18312
rect 54628 18300 54634 18352
rect 54772 18340 54800 18380
rect 54849 18377 54861 18411
rect 54895 18408 54907 18411
rect 56502 18408 56508 18420
rect 54895 18380 56508 18408
rect 54895 18377 54907 18380
rect 54849 18371 54907 18377
rect 56502 18368 56508 18380
rect 56560 18368 56566 18420
rect 57333 18411 57391 18417
rect 57333 18377 57345 18411
rect 57379 18408 57391 18411
rect 57422 18408 57428 18420
rect 57379 18380 57428 18408
rect 57379 18377 57391 18380
rect 57333 18371 57391 18377
rect 57422 18368 57428 18380
rect 57480 18368 57486 18420
rect 58526 18368 58532 18420
rect 58584 18368 58590 18420
rect 55217 18343 55275 18349
rect 55217 18340 55229 18343
rect 54772 18312 55229 18340
rect 55217 18309 55229 18312
rect 55263 18340 55275 18343
rect 55263 18312 55628 18340
rect 55263 18309 55275 18312
rect 55217 18303 55275 18309
rect 38059 18244 38516 18272
rect 38059 18241 38071 18244
rect 38013 18235 38071 18241
rect 38654 18232 38660 18284
rect 38712 18232 38718 18284
rect 53469 18275 53527 18281
rect 53469 18241 53481 18275
rect 53515 18272 53527 18275
rect 53558 18272 53564 18284
rect 53515 18244 53564 18272
rect 53515 18241 53527 18244
rect 53469 18235 53527 18241
rect 53558 18232 53564 18244
rect 53616 18232 53622 18284
rect 9030 18204 9036 18216
rect 8680 18176 9036 18204
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 9214 18164 9220 18216
rect 9272 18164 9278 18216
rect 11606 18164 11612 18216
rect 11664 18164 11670 18216
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 14240 18176 14657 18204
rect 14240 18164 14246 18176
rect 14645 18173 14657 18176
rect 14691 18173 14703 18207
rect 14645 18167 14703 18173
rect 19794 18164 19800 18216
rect 19852 18204 19858 18216
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 19852 18176 20085 18204
rect 19852 18164 19858 18176
rect 20073 18173 20085 18176
rect 20119 18173 20131 18207
rect 20073 18167 20131 18173
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 4396 18108 4752 18136
rect 5092 18136 5120 18164
rect 9950 18136 9956 18148
rect 5092 18108 9956 18136
rect 4396 18096 4402 18108
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 23400 18136 23428 18167
rect 23842 18164 23848 18216
rect 23900 18164 23906 18216
rect 24026 18164 24032 18216
rect 24084 18164 24090 18216
rect 26973 18207 27031 18213
rect 26973 18204 26985 18207
rect 26620 18176 26985 18204
rect 22664 18108 23428 18136
rect 23860 18136 23888 18164
rect 25130 18136 25136 18148
rect 23860 18108 25136 18136
rect 2498 18028 2504 18080
rect 2556 18068 2562 18080
rect 2869 18071 2927 18077
rect 2869 18068 2881 18071
rect 2556 18040 2881 18068
rect 2556 18028 2562 18040
rect 2869 18037 2881 18040
rect 2915 18037 2927 18071
rect 2869 18031 2927 18037
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 6178 18068 6184 18080
rect 4488 18040 6184 18068
rect 4488 18028 4494 18040
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 7282 18028 7288 18080
rect 7340 18028 7346 18080
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8297 18071 8355 18077
rect 8297 18068 8309 18071
rect 7984 18040 8309 18068
rect 7984 18028 7990 18040
rect 8297 18037 8309 18040
rect 8343 18037 8355 18071
rect 8297 18031 8355 18037
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 10137 18071 10195 18077
rect 10137 18068 10149 18071
rect 9456 18040 10149 18068
rect 9456 18028 9462 18040
rect 10137 18037 10149 18040
rect 10183 18037 10195 18071
rect 10137 18031 10195 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 12253 18071 12311 18077
rect 12253 18068 12265 18071
rect 10836 18040 12265 18068
rect 10836 18028 10842 18040
rect 12253 18037 12265 18040
rect 12299 18037 12311 18071
rect 12253 18031 12311 18037
rect 12621 18071 12679 18077
rect 12621 18037 12633 18071
rect 12667 18068 12679 18071
rect 12894 18068 12900 18080
rect 12667 18040 12900 18068
rect 12667 18037 12679 18040
rect 12621 18031 12679 18037
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 13909 18071 13967 18077
rect 13909 18068 13921 18071
rect 13872 18040 13921 18068
rect 13872 18028 13878 18040
rect 13909 18037 13921 18040
rect 13955 18037 13967 18071
rect 13909 18031 13967 18037
rect 15286 18028 15292 18080
rect 15344 18028 15350 18080
rect 20714 18028 20720 18080
rect 20772 18028 20778 18080
rect 22462 18028 22468 18080
rect 22520 18068 22526 18080
rect 22664 18077 22692 18108
rect 25130 18096 25136 18108
rect 25188 18096 25194 18148
rect 26620 18145 26648 18176
rect 26973 18173 26985 18176
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 28626 18164 28632 18216
rect 28684 18164 28690 18216
rect 29086 18164 29092 18216
rect 29144 18164 29150 18216
rect 29181 18207 29239 18213
rect 29181 18173 29193 18207
rect 29227 18204 29239 18207
rect 29733 18207 29791 18213
rect 29733 18204 29745 18207
rect 29227 18176 29745 18204
rect 29227 18173 29239 18176
rect 29181 18167 29239 18173
rect 29733 18173 29745 18176
rect 29779 18173 29791 18207
rect 29733 18167 29791 18173
rect 29825 18207 29883 18213
rect 29825 18173 29837 18207
rect 29871 18173 29883 18207
rect 29825 18167 29883 18173
rect 26605 18139 26663 18145
rect 26605 18136 26617 18139
rect 26206 18108 26617 18136
rect 22649 18071 22707 18077
rect 22649 18068 22661 18071
rect 22520 18040 22661 18068
rect 22520 18028 22526 18040
rect 22649 18037 22661 18040
rect 22695 18037 22707 18071
rect 22649 18031 22707 18037
rect 24486 18028 24492 18080
rect 24544 18028 24550 18080
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 26206 18068 26234 18108
rect 26605 18105 26617 18108
rect 26651 18105 26663 18139
rect 29104 18136 29132 18164
rect 29840 18136 29868 18167
rect 30190 18164 30196 18216
rect 30248 18164 30254 18216
rect 33321 18207 33379 18213
rect 33321 18173 33333 18207
rect 33367 18204 33379 18207
rect 33502 18204 33508 18216
rect 33367 18176 33508 18204
rect 33367 18173 33379 18176
rect 33321 18167 33379 18173
rect 33502 18164 33508 18176
rect 33560 18164 33566 18216
rect 33962 18164 33968 18216
rect 34020 18164 34026 18216
rect 47394 18164 47400 18216
rect 47452 18204 47458 18216
rect 47581 18207 47639 18213
rect 47581 18204 47593 18207
rect 47452 18176 47593 18204
rect 47452 18164 47458 18176
rect 47581 18173 47593 18176
rect 47627 18173 47639 18207
rect 47581 18167 47639 18173
rect 48314 18164 48320 18216
rect 48372 18204 48378 18216
rect 49602 18204 49608 18216
rect 48372 18176 49608 18204
rect 48372 18164 48378 18176
rect 49602 18164 49608 18176
rect 49660 18164 49666 18216
rect 52825 18207 52883 18213
rect 52825 18173 52837 18207
rect 52871 18204 52883 18207
rect 53098 18204 53104 18216
rect 52871 18176 53104 18204
rect 52871 18173 52883 18176
rect 52825 18167 52883 18173
rect 53098 18164 53104 18176
rect 53156 18164 53162 18216
rect 55493 18207 55551 18213
rect 55493 18173 55505 18207
rect 55539 18173 55551 18207
rect 55600 18204 55628 18312
rect 55674 18232 55680 18284
rect 55732 18232 55738 18284
rect 56502 18232 56508 18284
rect 56560 18281 56566 18284
rect 56560 18275 56588 18281
rect 56576 18241 56588 18275
rect 56560 18235 56588 18241
rect 56560 18232 56566 18235
rect 56134 18204 56140 18216
rect 55600 18176 56140 18204
rect 55493 18167 55551 18173
rect 29104 18108 29868 18136
rect 26605 18099 26663 18105
rect 41322 18096 41328 18148
rect 41380 18136 41386 18148
rect 41506 18136 41512 18148
rect 41380 18108 41512 18136
rect 41380 18096 41386 18108
rect 41506 18096 41512 18108
rect 41564 18096 41570 18148
rect 46937 18139 46995 18145
rect 46937 18105 46949 18139
rect 46983 18136 46995 18139
rect 46983 18108 47716 18136
rect 46983 18105 46995 18108
rect 46937 18099 46995 18105
rect 47688 18080 47716 18108
rect 25004 18040 26234 18068
rect 25004 18028 25010 18040
rect 27614 18028 27620 18080
rect 27672 18028 27678 18080
rect 29270 18028 29276 18080
rect 29328 18028 29334 18080
rect 30466 18028 30472 18080
rect 30524 18068 30530 18080
rect 30837 18071 30895 18077
rect 30837 18068 30849 18071
rect 30524 18040 30849 18068
rect 30524 18028 30530 18040
rect 30837 18037 30849 18040
rect 30883 18037 30895 18071
rect 30837 18031 30895 18037
rect 33134 18028 33140 18080
rect 33192 18068 33198 18080
rect 33873 18071 33931 18077
rect 33873 18068 33885 18071
rect 33192 18040 33885 18068
rect 33192 18028 33198 18040
rect 33873 18037 33885 18040
rect 33919 18037 33931 18071
rect 33873 18031 33931 18037
rect 34606 18028 34612 18080
rect 34664 18028 34670 18080
rect 34977 18071 35035 18077
rect 34977 18037 34989 18071
rect 35023 18068 35035 18071
rect 35434 18068 35440 18080
rect 35023 18040 35440 18068
rect 35023 18037 35035 18040
rect 34977 18031 35035 18037
rect 35434 18028 35440 18040
rect 35492 18028 35498 18080
rect 35621 18071 35679 18077
rect 35621 18037 35633 18071
rect 35667 18068 35679 18071
rect 35894 18068 35900 18080
rect 35667 18040 35900 18068
rect 35667 18037 35679 18040
rect 35621 18031 35679 18037
rect 35894 18028 35900 18040
rect 35952 18068 35958 18080
rect 36906 18068 36912 18080
rect 35952 18040 36912 18068
rect 35952 18028 35958 18040
rect 36906 18028 36912 18040
rect 36964 18068 36970 18080
rect 39942 18068 39948 18080
rect 36964 18040 39948 18068
rect 36964 18028 36970 18040
rect 39942 18028 39948 18040
rect 40000 18028 40006 18080
rect 41417 18071 41475 18077
rect 41417 18037 41429 18071
rect 41463 18068 41475 18071
rect 42058 18068 42064 18080
rect 41463 18040 42064 18068
rect 41463 18037 41475 18040
rect 41417 18031 41475 18037
rect 42058 18028 42064 18040
rect 42116 18028 42122 18080
rect 47397 18071 47455 18077
rect 47397 18037 47409 18071
rect 47443 18068 47455 18071
rect 47578 18068 47584 18080
rect 47443 18040 47584 18068
rect 47443 18037 47455 18040
rect 47397 18031 47455 18037
rect 47578 18028 47584 18040
rect 47636 18028 47642 18080
rect 47670 18028 47676 18080
rect 47728 18028 47734 18080
rect 48222 18028 48228 18080
rect 48280 18028 48286 18080
rect 48498 18028 48504 18080
rect 48556 18068 48562 18080
rect 50982 18068 50988 18080
rect 48556 18040 50988 18068
rect 48556 18028 48562 18040
rect 50982 18028 50988 18040
rect 51040 18028 51046 18080
rect 52549 18071 52607 18077
rect 52549 18037 52561 18071
rect 52595 18068 52607 18071
rect 52730 18068 52736 18080
rect 52595 18040 52736 18068
rect 52595 18037 52607 18040
rect 52549 18031 52607 18037
rect 52730 18028 52736 18040
rect 52788 18028 52794 18080
rect 53374 18028 53380 18080
rect 53432 18028 53438 18080
rect 55508 18068 55536 18167
rect 56134 18164 56140 18176
rect 56192 18164 56198 18216
rect 56410 18164 56416 18216
rect 56468 18164 56474 18216
rect 56686 18164 56692 18216
rect 56744 18164 56750 18216
rect 57882 18164 57888 18216
rect 57940 18164 57946 18216
rect 57422 18068 57428 18080
rect 55508 18040 57428 18068
rect 57422 18028 57428 18040
rect 57480 18028 57486 18080
rect 1104 17978 58880 18000
rect 1104 17926 8172 17978
rect 8224 17926 8236 17978
rect 8288 17926 8300 17978
rect 8352 17926 8364 17978
rect 8416 17926 8428 17978
rect 8480 17926 22616 17978
rect 22668 17926 22680 17978
rect 22732 17926 22744 17978
rect 22796 17926 22808 17978
rect 22860 17926 22872 17978
rect 22924 17926 37060 17978
rect 37112 17926 37124 17978
rect 37176 17926 37188 17978
rect 37240 17926 37252 17978
rect 37304 17926 37316 17978
rect 37368 17926 51504 17978
rect 51556 17926 51568 17978
rect 51620 17926 51632 17978
rect 51684 17926 51696 17978
rect 51748 17926 51760 17978
rect 51812 17926 58880 17978
rect 1104 17904 58880 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3237 17867 3295 17873
rect 3237 17864 3249 17867
rect 3108 17836 3249 17864
rect 3108 17824 3114 17836
rect 3237 17833 3249 17836
rect 3283 17864 3295 17867
rect 4706 17864 4712 17876
rect 3283 17836 4712 17864
rect 3283 17833 3295 17836
rect 3237 17827 3295 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 8570 17824 8576 17876
rect 8628 17864 8634 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 8628 17836 8953 17864
rect 8628 17824 8634 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 8941 17827 8999 17833
rect 9306 17824 9312 17876
rect 9364 17864 9370 17876
rect 20438 17864 20444 17876
rect 9364 17836 12940 17864
rect 9364 17824 9370 17836
rect 8757 17799 8815 17805
rect 3804 17768 4568 17796
rect 3804 17737 3832 17768
rect 3789 17731 3847 17737
rect 3789 17697 3801 17731
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 4430 17688 4436 17740
rect 4488 17688 4494 17740
rect 4540 17728 4568 17768
rect 8757 17765 8769 17799
rect 8803 17796 8815 17799
rect 8803 17768 9812 17796
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 5166 17728 5172 17740
rect 4540 17700 5172 17728
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 9398 17728 9404 17740
rect 8628 17700 9404 17728
rect 8628 17688 8634 17700
rect 9398 17688 9404 17700
rect 9456 17728 9462 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9456 17700 9505 17728
rect 9456 17688 9462 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 3973 17663 4031 17669
rect 1903 17632 2774 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 2746 17604 2774 17632
rect 3973 17629 3985 17663
rect 4019 17660 4031 17663
rect 4154 17660 4160 17672
rect 4019 17632 4160 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 4890 17669 4896 17672
rect 4847 17663 4896 17669
rect 4847 17629 4859 17663
rect 4893 17629 4896 17663
rect 4847 17623 4896 17629
rect 4890 17620 4896 17623
rect 4948 17620 4954 17672
rect 4982 17620 4988 17672
rect 5040 17620 5046 17672
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 5552 17632 5733 17660
rect 2124 17595 2182 17601
rect 2124 17561 2136 17595
rect 2170 17592 2182 17595
rect 2498 17592 2504 17604
rect 2170 17564 2504 17592
rect 2170 17561 2182 17564
rect 2124 17555 2182 17561
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 2746 17564 2780 17604
rect 2774 17552 2780 17564
rect 2832 17552 2838 17604
rect 2792 17524 2820 17552
rect 5552 17536 5580 17632
rect 5721 17629 5733 17632
rect 5767 17660 5779 17663
rect 6822 17660 6828 17672
rect 5767 17632 6828 17660
rect 5767 17629 5779 17632
rect 5721 17623 5779 17629
rect 6822 17620 6828 17632
rect 6880 17660 6886 17672
rect 9784 17669 9812 17768
rect 12636 17737 12664 17836
rect 12912 17808 12940 17836
rect 19536 17836 20444 17864
rect 19536 17808 19564 17836
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 25406 17864 25412 17876
rect 25056 17836 25412 17864
rect 12894 17756 12900 17808
rect 12952 17756 12958 17808
rect 19518 17756 19524 17808
rect 19576 17756 19582 17808
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 20027 17768 20852 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 12621 17731 12679 17737
rect 10551 17700 10640 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 6880 17632 7389 17660
rect 6880 17620 6886 17632
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 9815 17632 10548 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 10520 17604 10548 17632
rect 5988 17595 6046 17601
rect 5988 17561 6000 17595
rect 6034 17592 6046 17595
rect 7282 17592 7288 17604
rect 6034 17564 7288 17592
rect 6034 17561 6046 17564
rect 5988 17555 6046 17561
rect 7282 17552 7288 17564
rect 7340 17552 7346 17604
rect 7644 17595 7702 17601
rect 7644 17561 7656 17595
rect 7690 17592 7702 17595
rect 7926 17592 7932 17604
rect 7690 17564 7932 17592
rect 7690 17561 7702 17564
rect 7644 17555 7702 17561
rect 7926 17552 7932 17564
rect 7984 17552 7990 17604
rect 9309 17595 9367 17601
rect 9309 17561 9321 17595
rect 9355 17592 9367 17595
rect 10413 17595 10471 17601
rect 10413 17592 10425 17595
rect 9355 17564 10425 17592
rect 9355 17561 9367 17564
rect 9309 17555 9367 17561
rect 10413 17561 10425 17564
rect 10459 17561 10471 17595
rect 10413 17555 10471 17561
rect 10502 17552 10508 17604
rect 10560 17552 10566 17604
rect 10612 17592 10640 17700
rect 12621 17697 12633 17731
rect 12667 17697 12679 17731
rect 20530 17728 20536 17740
rect 12621 17691 12679 17697
rect 20088 17700 20536 17728
rect 10778 17669 10784 17672
rect 10772 17660 10784 17669
rect 10739 17632 10784 17660
rect 10772 17623 10784 17632
rect 10778 17620 10784 17623
rect 10836 17620 10842 17672
rect 11054 17620 11060 17672
rect 11112 17620 11118 17672
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 11572 17632 12357 17660
rect 11572 17620 11578 17632
rect 12345 17629 12357 17632
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12894 17620 12900 17672
rect 12952 17620 12958 17672
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 14148 17632 14197 17660
rect 14148 17620 14154 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 14792 17632 15669 17660
rect 14792 17620 14798 17632
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 17586 17620 17592 17672
rect 17644 17620 17650 17672
rect 11072 17592 11100 17620
rect 10612 17564 11100 17592
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 12437 17595 12495 17601
rect 12437 17592 12449 17595
rect 11388 17564 12449 17592
rect 11388 17552 11394 17564
rect 12437 17561 12449 17564
rect 12483 17561 12495 17595
rect 12437 17555 12495 17561
rect 14452 17595 14510 17601
rect 14452 17561 14464 17595
rect 14498 17592 14510 17595
rect 16301 17595 16359 17601
rect 16301 17592 16313 17595
rect 14498 17564 16313 17592
rect 14498 17561 14510 17564
rect 14452 17555 14510 17561
rect 16301 17561 16313 17564
rect 16347 17561 16359 17595
rect 16301 17555 16359 17561
rect 20088 17536 20116 17700
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 20824 17737 20852 17768
rect 23566 17756 23572 17808
rect 23624 17796 23630 17808
rect 25056 17796 25084 17836
rect 25406 17824 25412 17836
rect 25464 17824 25470 17876
rect 26234 17824 26240 17876
rect 26292 17824 26298 17876
rect 26329 17867 26387 17873
rect 26329 17833 26341 17867
rect 26375 17864 26387 17867
rect 26602 17864 26608 17876
rect 26375 17836 26608 17864
rect 26375 17833 26387 17836
rect 26329 17827 26387 17833
rect 26602 17824 26608 17836
rect 26660 17824 26666 17876
rect 30190 17824 30196 17876
rect 30248 17824 30254 17876
rect 38286 17824 38292 17876
rect 38344 17824 38350 17876
rect 47394 17824 47400 17876
rect 47452 17864 47458 17876
rect 52454 17864 52460 17876
rect 47452 17836 48912 17864
rect 47452 17824 47458 17836
rect 23624 17768 25084 17796
rect 23624 17756 23630 17768
rect 26142 17756 26148 17808
rect 26200 17796 26206 17808
rect 27614 17796 27620 17808
rect 26200 17768 26648 17796
rect 26200 17756 26206 17768
rect 20809 17731 20867 17737
rect 20809 17697 20821 17731
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24946 17728 24952 17740
rect 24627 17700 24952 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25130 17688 25136 17740
rect 25188 17728 25194 17740
rect 25188 17700 25360 17728
rect 25188 17688 25194 17700
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17660 20407 17663
rect 20714 17660 20720 17672
rect 20395 17632 20720 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22456 17663 22514 17669
rect 22456 17629 22468 17663
rect 22502 17660 22514 17663
rect 23290 17660 23296 17672
rect 22502 17632 23296 17660
rect 22502 17629 22514 17632
rect 22456 17623 22514 17629
rect 22204 17536 22232 17623
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 24397 17663 24455 17669
rect 24397 17629 24409 17663
rect 24443 17660 24455 17663
rect 24762 17660 24768 17672
rect 24443 17632 24768 17660
rect 24443 17629 24455 17632
rect 24397 17623 24455 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25332 17669 25360 17700
rect 25406 17688 25412 17740
rect 25464 17737 25470 17740
rect 25464 17731 25492 17737
rect 25480 17697 25492 17731
rect 26326 17728 26332 17740
rect 25464 17691 25492 17697
rect 25608 17700 26332 17728
rect 25464 17688 25470 17691
rect 25608 17672 25636 17700
rect 26326 17688 26332 17700
rect 26384 17688 26390 17740
rect 25317 17663 25375 17669
rect 25317 17629 25329 17663
rect 25363 17629 25375 17663
rect 25317 17623 25375 17629
rect 25590 17620 25596 17672
rect 25648 17620 25654 17672
rect 26620 17592 26648 17768
rect 26712 17768 27620 17796
rect 26712 17669 26740 17768
rect 27614 17756 27620 17768
rect 27672 17756 27678 17808
rect 38304 17796 38332 17824
rect 47029 17799 47087 17805
rect 47029 17796 47041 17799
rect 28092 17768 30144 17796
rect 26970 17688 26976 17740
rect 27028 17728 27034 17740
rect 28092 17728 28120 17768
rect 27028 17700 28120 17728
rect 28813 17731 28871 17737
rect 27028 17688 27034 17700
rect 28813 17697 28825 17731
rect 28859 17728 28871 17731
rect 29270 17728 29276 17740
rect 28859 17700 29276 17728
rect 28859 17697 28871 17700
rect 28813 17691 28871 17697
rect 29270 17688 29276 17700
rect 29328 17688 29334 17740
rect 30116 17737 30144 17768
rect 33060 17768 34008 17796
rect 33060 17737 33088 17768
rect 30101 17731 30159 17737
rect 30101 17697 30113 17731
rect 30147 17728 30159 17731
rect 30745 17731 30803 17737
rect 30745 17728 30757 17731
rect 30147 17700 30757 17728
rect 30147 17697 30159 17700
rect 30101 17691 30159 17697
rect 30745 17697 30757 17700
rect 30791 17697 30803 17731
rect 30745 17691 30803 17697
rect 33045 17731 33103 17737
rect 33045 17697 33057 17731
rect 33091 17697 33103 17731
rect 33045 17691 33103 17697
rect 33134 17688 33140 17740
rect 33192 17688 33198 17740
rect 33229 17731 33287 17737
rect 33229 17697 33241 17731
rect 33275 17697 33287 17731
rect 33980 17728 34008 17768
rect 36096 17768 38332 17796
rect 46400 17768 47041 17796
rect 34238 17728 34244 17740
rect 33980 17700 34244 17728
rect 33229 17691 33287 17697
rect 26697 17663 26755 17669
rect 26697 17629 26709 17663
rect 26743 17629 26755 17663
rect 26697 17623 26755 17629
rect 27614 17620 27620 17672
rect 27672 17620 27678 17672
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 30653 17663 30711 17669
rect 30653 17660 30665 17663
rect 30432 17632 30665 17660
rect 30432 17620 30438 17632
rect 30653 17629 30665 17632
rect 30699 17629 30711 17663
rect 30653 17623 30711 17629
rect 31110 17620 31116 17672
rect 31168 17620 31174 17672
rect 32861 17663 32919 17669
rect 32861 17629 32873 17663
rect 32907 17660 32919 17663
rect 33152 17660 33180 17688
rect 32907 17632 33180 17660
rect 32907 17629 32919 17632
rect 32861 17623 32919 17629
rect 26789 17595 26847 17601
rect 26789 17592 26801 17595
rect 26620 17564 26801 17592
rect 26789 17561 26801 17564
rect 26835 17592 26847 17595
rect 30561 17595 30619 17601
rect 26835 17564 27476 17592
rect 26835 17561 26847 17564
rect 26789 17555 26847 17561
rect 5534 17524 5540 17536
rect 2792 17496 5540 17524
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 5626 17484 5632 17536
rect 5684 17484 5690 17536
rect 7098 17484 7104 17536
rect 7156 17484 7162 17536
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 9401 17527 9459 17533
rect 9401 17524 9413 17527
rect 8812 17496 9413 17524
rect 8812 17484 8818 17496
rect 9401 17493 9413 17496
rect 9447 17524 9459 17527
rect 10870 17524 10876 17536
rect 9447 17496 10876 17524
rect 9447 17493 9459 17496
rect 9401 17487 9459 17493
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 11885 17527 11943 17533
rect 11885 17524 11897 17527
rect 11480 17496 11897 17524
rect 11480 17484 11486 17496
rect 11885 17493 11897 17496
rect 11931 17493 11943 17527
rect 11885 17487 11943 17493
rect 11974 17484 11980 17536
rect 12032 17484 12038 17536
rect 13446 17484 13452 17536
rect 13504 17484 13510 17536
rect 13814 17484 13820 17536
rect 13872 17484 13878 17536
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 15565 17527 15623 17533
rect 15565 17524 15577 17527
rect 14240 17496 15577 17524
rect 14240 17484 14246 17496
rect 15565 17493 15577 17496
rect 15611 17493 15623 17527
rect 15565 17487 15623 17493
rect 18138 17484 18144 17536
rect 18196 17484 18202 17536
rect 19889 17527 19947 17533
rect 19889 17493 19901 17527
rect 19935 17524 19947 17527
rect 20070 17524 20076 17536
rect 19935 17496 20076 17524
rect 19935 17493 19947 17496
rect 19889 17487 19947 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 20346 17484 20352 17536
rect 20404 17524 20410 17536
rect 20441 17527 20499 17533
rect 20441 17524 20453 17527
rect 20404 17496 20453 17524
rect 20404 17484 20410 17496
rect 20441 17493 20453 17496
rect 20487 17493 20499 17527
rect 20441 17487 20499 17493
rect 21450 17484 21456 17536
rect 21508 17484 21514 17536
rect 22097 17527 22155 17533
rect 22097 17493 22109 17527
rect 22143 17524 22155 17527
rect 22186 17524 22192 17536
rect 22143 17496 22192 17524
rect 22143 17493 22155 17496
rect 22097 17487 22155 17493
rect 22186 17484 22192 17496
rect 22244 17524 22250 17536
rect 23934 17524 23940 17536
rect 22244 17496 23940 17524
rect 22244 17484 22250 17496
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 24118 17484 24124 17536
rect 24176 17484 24182 17536
rect 24302 17484 24308 17536
rect 24360 17524 24366 17536
rect 25590 17524 25596 17536
rect 24360 17496 25596 17524
rect 24360 17484 24366 17496
rect 25590 17484 25596 17496
rect 25648 17484 25654 17536
rect 27338 17484 27344 17536
rect 27396 17484 27402 17536
rect 27448 17524 27476 17564
rect 30561 17561 30573 17595
rect 30607 17592 30619 17595
rect 31665 17595 31723 17601
rect 31665 17592 31677 17595
rect 30607 17564 31677 17592
rect 30607 17561 30619 17564
rect 30561 17555 30619 17561
rect 31665 17561 31677 17564
rect 31711 17561 31723 17595
rect 33244 17592 33272 17691
rect 34238 17688 34244 17700
rect 34296 17728 34302 17740
rect 36096 17728 36124 17768
rect 40770 17728 40776 17740
rect 34296 17700 36124 17728
rect 38120 17700 40776 17728
rect 34296 17688 34302 17700
rect 38120 17672 38148 17700
rect 40770 17688 40776 17700
rect 40828 17688 40834 17740
rect 43346 17688 43352 17740
rect 43404 17728 43410 17740
rect 46400 17737 46428 17768
rect 47029 17765 47041 17768
rect 47075 17765 47087 17799
rect 47029 17759 47087 17765
rect 43809 17731 43867 17737
rect 43809 17728 43821 17731
rect 43404 17700 43821 17728
rect 43404 17688 43410 17700
rect 43809 17697 43821 17700
rect 43855 17728 43867 17731
rect 44545 17731 44603 17737
rect 44545 17728 44557 17731
rect 43855 17700 44557 17728
rect 43855 17697 43867 17700
rect 43809 17691 43867 17697
rect 44545 17697 44557 17700
rect 44591 17728 44603 17731
rect 46385 17731 46443 17737
rect 44591 17700 46336 17728
rect 44591 17697 44603 17700
rect 44545 17691 44603 17697
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 34572 17632 34713 17660
rect 34572 17620 34578 17632
rect 34701 17629 34713 17632
rect 34747 17629 34759 17663
rect 34701 17623 34759 17629
rect 38102 17620 38108 17672
rect 38160 17620 38166 17672
rect 38381 17663 38439 17669
rect 38381 17629 38393 17663
rect 38427 17660 38439 17663
rect 38930 17660 38936 17672
rect 38427 17632 38936 17660
rect 38427 17629 38439 17632
rect 38381 17623 38439 17629
rect 38930 17620 38936 17632
rect 38988 17620 38994 17672
rect 40126 17620 40132 17672
rect 40184 17620 40190 17672
rect 41506 17620 41512 17672
rect 41564 17620 41570 17672
rect 44174 17620 44180 17672
rect 44232 17660 44238 17672
rect 44269 17663 44327 17669
rect 44269 17660 44281 17663
rect 44232 17632 44281 17660
rect 44232 17620 44238 17632
rect 44269 17629 44281 17632
rect 44315 17629 44327 17663
rect 45189 17663 45247 17669
rect 45189 17660 45201 17663
rect 44269 17623 44327 17629
rect 44928 17632 45201 17660
rect 39577 17595 39635 17601
rect 39577 17592 39589 17595
rect 31665 17555 31723 17561
rect 32416 17564 33272 17592
rect 36648 17564 39589 17592
rect 27706 17524 27712 17536
rect 27448 17496 27712 17524
rect 27706 17484 27712 17496
rect 27764 17484 27770 17536
rect 27890 17484 27896 17536
rect 27948 17524 27954 17536
rect 28261 17527 28319 17533
rect 28261 17524 28273 17527
rect 27948 17496 28273 17524
rect 27948 17484 27954 17496
rect 28261 17493 28273 17496
rect 28307 17493 28319 17527
rect 28261 17487 28319 17493
rect 29362 17484 29368 17536
rect 29420 17484 29426 17536
rect 32416 17533 32444 17564
rect 36648 17536 36676 17564
rect 39577 17561 39589 17564
rect 39623 17561 39635 17595
rect 39577 17555 39635 17561
rect 32401 17527 32459 17533
rect 32401 17493 32413 17527
rect 32447 17493 32459 17527
rect 32401 17487 32459 17493
rect 32766 17484 32772 17536
rect 32824 17484 32830 17536
rect 33134 17484 33140 17536
rect 33192 17524 33198 17536
rect 33873 17527 33931 17533
rect 33873 17524 33885 17527
rect 33192 17496 33885 17524
rect 33192 17484 33198 17496
rect 33873 17493 33885 17496
rect 33919 17493 33931 17527
rect 33873 17487 33931 17493
rect 35342 17484 35348 17536
rect 35400 17484 35406 17536
rect 36630 17484 36636 17536
rect 36688 17484 36694 17536
rect 36722 17484 36728 17536
rect 36780 17524 36786 17536
rect 37737 17527 37795 17533
rect 37737 17524 37749 17527
rect 36780 17496 37749 17524
rect 36780 17484 36786 17496
rect 37737 17493 37749 17496
rect 37783 17493 37795 17527
rect 37737 17487 37795 17493
rect 38194 17484 38200 17536
rect 38252 17484 38258 17536
rect 38746 17484 38752 17536
rect 38804 17524 38810 17536
rect 38933 17527 38991 17533
rect 38933 17524 38945 17527
rect 38804 17496 38945 17524
rect 38804 17484 38810 17496
rect 38933 17493 38945 17496
rect 38979 17493 38991 17527
rect 39592 17524 39620 17555
rect 44928 17536 44956 17632
rect 45189 17629 45201 17632
rect 45235 17629 45247 17663
rect 46308 17660 46336 17700
rect 46385 17697 46397 17731
rect 46431 17697 46443 17731
rect 46385 17691 46443 17697
rect 47670 17688 47676 17740
rect 47728 17688 47734 17740
rect 48317 17731 48375 17737
rect 48317 17697 48329 17731
rect 48363 17728 48375 17731
rect 48498 17728 48504 17740
rect 48363 17700 48504 17728
rect 48363 17697 48375 17700
rect 48317 17691 48375 17697
rect 48498 17688 48504 17700
rect 48556 17688 48562 17740
rect 48682 17688 48688 17740
rect 48740 17728 48746 17740
rect 48777 17731 48835 17737
rect 48777 17728 48789 17731
rect 48740 17700 48789 17728
rect 48740 17688 48746 17700
rect 48777 17697 48789 17700
rect 48823 17697 48835 17731
rect 48884 17728 48912 17836
rect 51184 17836 52460 17864
rect 49170 17731 49228 17737
rect 49170 17728 49182 17731
rect 48884 17700 49182 17728
rect 48777 17691 48835 17697
rect 49170 17697 49182 17700
rect 49216 17697 49228 17731
rect 49170 17691 49228 17697
rect 49326 17688 49332 17740
rect 49384 17688 49390 17740
rect 51184 17737 51212 17836
rect 52454 17824 52460 17836
rect 52512 17824 52518 17876
rect 57422 17824 57428 17876
rect 57480 17824 57486 17876
rect 57517 17867 57575 17873
rect 57517 17833 57529 17867
rect 57563 17864 57575 17867
rect 57882 17864 57888 17876
rect 57563 17836 57888 17864
rect 57563 17833 57575 17836
rect 57517 17827 57575 17833
rect 57882 17824 57888 17836
rect 57940 17824 57946 17876
rect 50801 17731 50859 17737
rect 50801 17728 50813 17731
rect 49896 17700 50813 17728
rect 46308 17632 48084 17660
rect 45189 17623 45247 17629
rect 48056 17536 48084 17632
rect 48130 17620 48136 17672
rect 48188 17620 48194 17672
rect 49050 17620 49056 17672
rect 49108 17620 49114 17672
rect 40034 17524 40040 17536
rect 39592 17496 40040 17524
rect 38933 17487 38991 17493
rect 40034 17484 40040 17496
rect 40092 17484 40098 17536
rect 40678 17484 40684 17536
rect 40736 17484 40742 17536
rect 41414 17484 41420 17536
rect 41472 17484 41478 17536
rect 42150 17484 42156 17536
rect 42208 17484 42214 17536
rect 43898 17484 43904 17536
rect 43956 17484 43962 17536
rect 44361 17527 44419 17533
rect 44361 17493 44373 17527
rect 44407 17524 44419 17527
rect 44634 17524 44640 17536
rect 44407 17496 44640 17524
rect 44407 17493 44419 17496
rect 44361 17487 44419 17493
rect 44634 17484 44640 17496
rect 44692 17484 44698 17536
rect 44910 17484 44916 17536
rect 44968 17484 44974 17536
rect 45462 17484 45468 17536
rect 45520 17524 45526 17536
rect 45833 17527 45891 17533
rect 45833 17524 45845 17527
rect 45520 17496 45845 17524
rect 45520 17484 45526 17496
rect 45833 17493 45845 17496
rect 45879 17493 45891 17527
rect 45833 17487 45891 17493
rect 46934 17484 46940 17536
rect 46992 17484 46998 17536
rect 47302 17484 47308 17536
rect 47360 17524 47366 17536
rect 47397 17527 47455 17533
rect 47397 17524 47409 17527
rect 47360 17496 47409 17524
rect 47360 17484 47366 17496
rect 47397 17493 47409 17496
rect 47443 17493 47455 17527
rect 47397 17487 47455 17493
rect 47489 17527 47547 17533
rect 47489 17493 47501 17527
rect 47535 17524 47547 17527
rect 47946 17524 47952 17536
rect 47535 17496 47952 17524
rect 47535 17493 47547 17496
rect 47489 17487 47547 17493
rect 47946 17484 47952 17496
rect 48004 17484 48010 17536
rect 48038 17484 48044 17536
rect 48096 17524 48102 17536
rect 49896 17524 49924 17700
rect 50801 17697 50813 17700
rect 50847 17728 50859 17731
rect 51169 17731 51227 17737
rect 51169 17728 51181 17731
rect 50847 17700 51181 17728
rect 50847 17697 50859 17700
rect 50801 17691 50859 17697
rect 51169 17697 51181 17700
rect 51215 17697 51227 17731
rect 51169 17691 51227 17697
rect 57514 17688 57520 17740
rect 57572 17728 57578 17740
rect 58069 17731 58127 17737
rect 58069 17728 58081 17731
rect 57572 17700 58081 17728
rect 57572 17688 57578 17700
rect 58069 17697 58081 17700
rect 58115 17697 58127 17731
rect 58069 17691 58127 17697
rect 50062 17620 50068 17672
rect 50120 17660 50126 17672
rect 50525 17663 50583 17669
rect 50525 17660 50537 17663
rect 50120 17632 50537 17660
rect 50120 17620 50126 17632
rect 50525 17629 50537 17632
rect 50571 17629 50583 17663
rect 50525 17623 50583 17629
rect 51350 17620 51356 17672
rect 51408 17660 51414 17672
rect 51721 17663 51779 17669
rect 51721 17660 51733 17663
rect 51408 17632 51733 17660
rect 51408 17620 51414 17632
rect 51721 17629 51733 17632
rect 51767 17660 51779 17663
rect 53466 17660 53472 17672
rect 51767 17632 51948 17660
rect 51767 17629 51779 17632
rect 51721 17623 51779 17629
rect 49973 17595 50031 17601
rect 49973 17561 49985 17595
rect 50019 17592 50031 17595
rect 50617 17595 50675 17601
rect 50617 17592 50629 17595
rect 50019 17564 50629 17592
rect 50019 17561 50031 17564
rect 49973 17555 50031 17561
rect 50617 17561 50629 17564
rect 50663 17561 50675 17595
rect 50617 17555 50675 17561
rect 51920 17536 51948 17632
rect 52196 17632 53472 17660
rect 51988 17595 52046 17601
rect 51988 17561 52000 17595
rect 52034 17592 52046 17595
rect 52196 17592 52224 17632
rect 53466 17620 53472 17632
rect 53524 17620 53530 17672
rect 56042 17660 56048 17672
rect 54496 17632 56048 17660
rect 52034 17564 52224 17592
rect 52034 17561 52046 17564
rect 51988 17555 52046 17561
rect 52730 17552 52736 17604
rect 52788 17592 52794 17604
rect 53193 17595 53251 17601
rect 53193 17592 53205 17595
rect 52788 17564 53205 17592
rect 52788 17552 52794 17564
rect 53193 17561 53205 17564
rect 53239 17561 53251 17595
rect 53193 17555 53251 17561
rect 48096 17496 49924 17524
rect 48096 17484 48102 17496
rect 50154 17484 50160 17536
rect 50212 17484 50218 17536
rect 51902 17484 51908 17536
rect 51960 17484 51966 17536
rect 53098 17484 53104 17536
rect 53156 17484 53162 17536
rect 53558 17484 53564 17536
rect 53616 17524 53622 17536
rect 54496 17533 54524 17632
rect 56042 17620 56048 17632
rect 56100 17620 56106 17672
rect 56686 17660 56692 17672
rect 56244 17632 56692 17660
rect 55490 17552 55496 17604
rect 55548 17592 55554 17604
rect 56244 17592 56272 17632
rect 56686 17620 56692 17632
rect 56744 17660 56750 17672
rect 56870 17660 56876 17672
rect 56744 17632 56876 17660
rect 56744 17620 56750 17632
rect 56870 17620 56876 17632
rect 56928 17620 56934 17672
rect 57885 17663 57943 17669
rect 57885 17629 57897 17663
rect 57931 17660 57943 17663
rect 58158 17660 58164 17672
rect 57931 17632 58164 17660
rect 57931 17629 57943 17632
rect 57885 17623 57943 17629
rect 58158 17620 58164 17632
rect 58216 17620 58222 17672
rect 55548 17564 56272 17592
rect 56312 17595 56370 17601
rect 55548 17552 55554 17564
rect 56312 17561 56324 17595
rect 56358 17592 56370 17595
rect 57054 17592 57060 17604
rect 56358 17564 57060 17592
rect 56358 17561 56370 17564
rect 56312 17555 56370 17561
rect 57054 17552 57060 17564
rect 57112 17552 57118 17604
rect 54481 17527 54539 17533
rect 54481 17524 54493 17527
rect 53616 17496 54493 17524
rect 53616 17484 53622 17496
rect 54481 17493 54493 17496
rect 54527 17493 54539 17527
rect 54481 17487 54539 17493
rect 57790 17484 57796 17536
rect 57848 17524 57854 17536
rect 57977 17527 58035 17533
rect 57977 17524 57989 17527
rect 57848 17496 57989 17524
rect 57848 17484 57854 17496
rect 57977 17493 57989 17496
rect 58023 17524 58035 17527
rect 58434 17524 58440 17536
rect 58023 17496 58440 17524
rect 58023 17493 58035 17496
rect 57977 17487 58035 17493
rect 58434 17484 58440 17496
rect 58492 17484 58498 17536
rect 1104 17434 59040 17456
rect 1104 17382 15394 17434
rect 15446 17382 15458 17434
rect 15510 17382 15522 17434
rect 15574 17382 15586 17434
rect 15638 17382 15650 17434
rect 15702 17382 29838 17434
rect 29890 17382 29902 17434
rect 29954 17382 29966 17434
rect 30018 17382 30030 17434
rect 30082 17382 30094 17434
rect 30146 17382 44282 17434
rect 44334 17382 44346 17434
rect 44398 17382 44410 17434
rect 44462 17382 44474 17434
rect 44526 17382 44538 17434
rect 44590 17382 58726 17434
rect 58778 17382 58790 17434
rect 58842 17382 58854 17434
rect 58906 17382 58918 17434
rect 58970 17382 58982 17434
rect 59034 17382 59040 17434
rect 1104 17360 59040 17382
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 3191 17292 4936 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 4908 17264 4936 17292
rect 5626 17280 5632 17332
rect 5684 17320 5690 17332
rect 5813 17323 5871 17329
rect 5813 17320 5825 17323
rect 5684 17292 5825 17320
rect 5684 17280 5690 17292
rect 5813 17289 5825 17292
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 5902 17280 5908 17332
rect 5960 17280 5966 17332
rect 6365 17323 6423 17329
rect 6365 17289 6377 17323
rect 6411 17320 6423 17323
rect 6638 17320 6644 17332
rect 6411 17292 6644 17320
rect 6411 17289 6423 17292
rect 6365 17283 6423 17289
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 6914 17320 6920 17332
rect 6779 17292 6920 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9214 17320 9220 17332
rect 9171 17292 9220 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9692 17292 11284 17320
rect 2774 17252 2780 17264
rect 1780 17224 2780 17252
rect 1780 17193 1808 17224
rect 2774 17212 2780 17224
rect 2832 17252 2838 17264
rect 3780 17255 3838 17261
rect 2832 17224 3556 17252
rect 2832 17212 2838 17224
rect 3528 17193 3556 17224
rect 3780 17221 3792 17255
rect 3826 17252 3838 17255
rect 4798 17252 4804 17264
rect 3826 17224 4804 17252
rect 3826 17221 3838 17224
rect 3780 17215 3838 17221
rect 4798 17212 4804 17224
rect 4856 17212 4862 17264
rect 4890 17212 4896 17264
rect 4948 17212 4954 17264
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 5920 17252 5948 17280
rect 5767 17224 5948 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 8018 17261 8024 17264
rect 8012 17252 8024 17261
rect 6880 17224 7788 17252
rect 7979 17224 8024 17252
rect 6880 17212 6886 17224
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 2032 17187 2090 17193
rect 2032 17153 2044 17187
rect 2078 17184 2090 17187
rect 3513 17187 3571 17193
rect 2078 17156 2820 17184
rect 2078 17153 2090 17156
rect 2032 17147 2090 17153
rect 2792 17128 2820 17156
rect 3513 17153 3525 17187
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 6362 17184 6368 17196
rect 4212 17156 6368 17184
rect 4212 17144 4218 17156
rect 6362 17144 6368 17156
rect 6420 17184 6426 17196
rect 7098 17184 7104 17196
rect 6420 17156 7104 17184
rect 6420 17144 6426 17156
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7760 17193 7788 17224
rect 8012 17215 8024 17224
rect 8018 17212 8024 17215
rect 8076 17212 8082 17264
rect 9692 17252 9720 17292
rect 9048 17224 9720 17252
rect 11256 17252 11284 17292
rect 11330 17280 11336 17332
rect 11388 17280 11394 17332
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17320 11575 17323
rect 11606 17320 11612 17332
rect 11563 17292 11612 17320
rect 11563 17289 11575 17292
rect 11517 17283 11575 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 12894 17280 12900 17332
rect 12952 17320 12958 17332
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 12952 17292 13001 17320
rect 12952 17280 12958 17292
rect 12989 17289 13001 17292
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 13449 17323 13507 17329
rect 13449 17289 13461 17323
rect 13495 17320 13507 17323
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 13495 17292 14473 17320
rect 13495 17289 13507 17292
rect 13449 17283 13507 17289
rect 14461 17289 14473 17292
rect 14507 17289 14519 17323
rect 14461 17283 14519 17289
rect 14734 17280 14740 17332
rect 14792 17280 14798 17332
rect 15197 17323 15255 17329
rect 15197 17289 15209 17323
rect 15243 17320 15255 17323
rect 15286 17320 15292 17332
rect 15243 17292 15292 17320
rect 15243 17289 15255 17292
rect 15197 17283 15255 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17681 17323 17739 17329
rect 17681 17320 17693 17323
rect 17644 17292 17693 17320
rect 17644 17280 17650 17292
rect 17681 17289 17693 17292
rect 17727 17289 17739 17323
rect 20254 17320 20260 17332
rect 17681 17283 17739 17289
rect 17788 17292 20260 17320
rect 13357 17255 13415 17261
rect 11256 17224 12112 17252
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 9048 17184 9076 17224
rect 7745 17147 7803 17153
rect 7852 17156 9076 17184
rect 2774 17076 2780 17128
rect 2832 17076 2838 17128
rect 5258 17116 5264 17128
rect 4908 17088 5264 17116
rect 4908 17057 4936 17088
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 5902 17076 5908 17128
rect 5960 17076 5966 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 7055 17088 7389 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7377 17085 7389 17088
rect 7423 17116 7435 17119
rect 7852 17116 7880 17156
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 9272 17156 9812 17184
rect 9272 17144 9278 17156
rect 7423 17088 7880 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 4893 17051 4951 17057
rect 4893 17017 4905 17051
rect 4939 17017 4951 17051
rect 6840 17048 6868 17079
rect 9306 17076 9312 17128
rect 9364 17076 9370 17128
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17116 9551 17119
rect 9582 17116 9588 17128
rect 9539 17088 9588 17116
rect 9539 17085 9551 17088
rect 9493 17079 9551 17085
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17085 9735 17119
rect 9784 17116 9812 17156
rect 10502 17144 10508 17196
rect 10560 17193 10566 17196
rect 10560 17187 10588 17193
rect 10576 17153 10588 17187
rect 10560 17147 10588 17153
rect 10560 17144 10566 17147
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 10413 17119 10471 17125
rect 10413 17116 10425 17119
rect 9784 17088 10425 17116
rect 9677 17079 9735 17085
rect 10413 17085 10425 17088
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 4893 17011 4951 17017
rect 5276 17020 6868 17048
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 5276 16980 5304 17020
rect 4580 16952 5304 16980
rect 4580 16940 4586 16952
rect 5350 16940 5356 16992
rect 5408 16940 5414 16992
rect 5902 16940 5908 16992
rect 5960 16980 5966 16992
rect 6822 16980 6828 16992
rect 5960 16952 6828 16980
rect 5960 16940 5966 16952
rect 6822 16940 6828 16952
rect 6880 16980 6886 16992
rect 9324 16980 9352 17076
rect 6880 16952 9352 16980
rect 9692 16980 9720 17079
rect 10686 17076 10692 17128
rect 10744 17076 10750 17128
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 11790 17116 11796 17128
rect 10928 17088 11796 17116
rect 10928 17076 10934 17088
rect 11790 17076 11796 17088
rect 11848 17116 11854 17128
rect 12084 17125 12112 17224
rect 13357 17221 13369 17255
rect 13403 17221 13415 17255
rect 13906 17252 13912 17264
rect 13357 17215 13415 17221
rect 13832 17224 13912 17252
rect 13372 17184 13400 17215
rect 13722 17184 13728 17196
rect 13372 17156 13728 17184
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 13832 17193 13860 17224
rect 13906 17212 13912 17224
rect 13964 17212 13970 17264
rect 15930 17212 15936 17264
rect 15988 17252 15994 17264
rect 16390 17252 16396 17264
rect 15988 17224 16396 17252
rect 15988 17212 15994 17224
rect 16390 17212 16396 17224
rect 16448 17252 16454 17264
rect 17788 17252 17816 17292
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 22186 17320 22192 17332
rect 21284 17292 22192 17320
rect 16448 17224 17816 17252
rect 18049 17255 18107 17261
rect 16448 17212 16454 17224
rect 18049 17221 18061 17255
rect 18095 17252 18107 17255
rect 18095 17224 19380 17252
rect 18095 17221 18107 17224
rect 18049 17215 18107 17221
rect 19352 17196 19380 17224
rect 19518 17212 19524 17264
rect 19576 17212 19582 17264
rect 21284 17261 21312 17292
rect 21269 17255 21327 17261
rect 21269 17252 21281 17255
rect 19628 17224 21281 17252
rect 13817 17187 13875 17193
rect 13817 17153 13829 17187
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 14884 17156 15117 17184
rect 14884 17144 14890 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17184 18199 17187
rect 19153 17187 19211 17193
rect 19153 17184 19165 17187
rect 18187 17156 19165 17184
rect 18187 17153 18199 17156
rect 18141 17147 18199 17153
rect 19153 17153 19165 17156
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 19334 17144 19340 17196
rect 19392 17144 19398 17196
rect 19628 17193 19656 17224
rect 21269 17221 21281 17224
rect 21315 17221 21327 17255
rect 21269 17215 21327 17221
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19880 17187 19938 17193
rect 19880 17153 19892 17187
rect 19926 17184 19938 17187
rect 21450 17184 21456 17196
rect 19926 17156 21456 17184
rect 19926 17153 19938 17156
rect 19880 17147 19938 17153
rect 21450 17144 21456 17156
rect 21508 17144 21514 17196
rect 22112 17184 22140 17292
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 23569 17323 23627 17329
rect 23569 17289 23581 17323
rect 23615 17320 23627 17323
rect 23842 17320 23848 17332
rect 23615 17292 23848 17320
rect 23615 17289 23627 17292
rect 23569 17283 23627 17289
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 24121 17323 24179 17329
rect 24121 17289 24133 17323
rect 24167 17320 24179 17323
rect 24486 17320 24492 17332
rect 24167 17292 24492 17320
rect 24167 17289 24179 17292
rect 24121 17283 24179 17289
rect 24486 17280 24492 17292
rect 24544 17280 24550 17332
rect 24762 17280 24768 17332
rect 24820 17320 24826 17332
rect 25869 17323 25927 17329
rect 25869 17320 25881 17323
rect 24820 17292 25881 17320
rect 24820 17280 24826 17292
rect 25869 17289 25881 17292
rect 25915 17320 25927 17323
rect 25915 17292 26004 17320
rect 25915 17289 25927 17292
rect 25869 17283 25927 17289
rect 24026 17212 24032 17264
rect 24084 17212 24090 17264
rect 25314 17252 25320 17264
rect 24504 17224 25320 17252
rect 22189 17187 22247 17193
rect 22189 17184 22201 17187
rect 22112 17156 22201 17184
rect 22189 17153 22201 17156
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22456 17187 22514 17193
rect 22456 17153 22468 17187
rect 22502 17184 22514 17187
rect 23750 17184 23756 17196
rect 22502 17156 23756 17184
rect 22502 17153 22514 17156
rect 22456 17147 22514 17153
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24394 17184 24400 17196
rect 23992 17156 24400 17184
rect 23992 17144 23998 17156
rect 24394 17144 24400 17156
rect 24452 17184 24458 17196
rect 24504 17193 24532 17224
rect 25314 17212 25320 17224
rect 25372 17252 25378 17264
rect 25372 17224 25912 17252
rect 25372 17212 25378 17224
rect 24489 17187 24547 17193
rect 24489 17184 24501 17187
rect 24452 17156 24501 17184
rect 24452 17144 24458 17156
rect 24489 17153 24501 17156
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 24756 17187 24814 17193
rect 24756 17153 24768 17187
rect 24802 17184 24814 17187
rect 25590 17184 25596 17196
rect 24802 17156 25596 17184
rect 24802 17153 24814 17156
rect 24756 17147 24814 17153
rect 25590 17144 25596 17156
rect 25648 17144 25654 17196
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11848 17088 11989 17116
rect 11848 17076 11854 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 12069 17119 12127 17125
rect 12069 17085 12081 17119
rect 12115 17085 12127 17119
rect 12069 17079 12127 17085
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 9824 17020 10149 17048
rect 9824 17008 9830 17020
rect 10137 17017 10149 17020
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 11422 16980 11428 16992
rect 9692 16952 11428 16980
rect 6880 16940 6886 16952
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 12084 16980 12112 17079
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12768 17088 12909 17116
rect 12768 17076 12774 17088
rect 12897 17085 12909 17088
rect 12943 17116 12955 17119
rect 13354 17116 13360 17128
rect 12943 17088 13360 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 13354 17076 13360 17088
rect 13412 17116 13418 17128
rect 13633 17119 13691 17125
rect 13633 17116 13645 17119
rect 13412 17088 13645 17116
rect 13412 17076 13418 17088
rect 13633 17085 13645 17088
rect 13679 17116 13691 17119
rect 13679 17088 14412 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 13998 17048 14004 17060
rect 12728 17020 14004 17048
rect 12158 16980 12164 16992
rect 12084 16952 12164 16980
rect 12158 16940 12164 16952
rect 12216 16980 12222 16992
rect 12728 16980 12756 17020
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 14384 17048 14412 17088
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 15381 17119 15439 17125
rect 15381 17116 15393 17119
rect 14792 17088 15393 17116
rect 14792 17076 14798 17088
rect 15381 17085 15393 17088
rect 15427 17116 15439 17119
rect 16209 17119 16267 17125
rect 16209 17116 16221 17119
rect 15427 17088 16221 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 16209 17085 16221 17088
rect 16255 17085 16267 17119
rect 16209 17079 16267 17085
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17116 17647 17119
rect 18233 17119 18291 17125
rect 18233 17116 18245 17119
rect 17635 17088 18245 17116
rect 17635 17085 17647 17088
rect 17589 17079 17647 17085
rect 18233 17085 18245 17088
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 17604 17048 17632 17079
rect 18598 17076 18604 17128
rect 18656 17076 18662 17128
rect 24302 17076 24308 17128
rect 24360 17076 24366 17128
rect 25884 17116 25912 17224
rect 25976 17193 26004 17292
rect 28626 17280 28632 17332
rect 28684 17320 28690 17332
rect 29181 17323 29239 17329
rect 29181 17320 29193 17323
rect 28684 17292 29193 17320
rect 28684 17280 28690 17292
rect 29181 17289 29193 17292
rect 29227 17289 29239 17323
rect 29181 17283 29239 17289
rect 29362 17280 29368 17332
rect 29420 17280 29426 17332
rect 31846 17320 31852 17332
rect 31726 17292 31852 17320
rect 28068 17255 28126 17261
rect 28068 17221 28080 17255
rect 28114 17252 28126 17255
rect 29380 17252 29408 17280
rect 28114 17224 29408 17252
rect 28114 17221 28126 17224
rect 28068 17215 28126 17221
rect 25961 17187 26019 17193
rect 25961 17153 25973 17187
rect 26007 17153 26019 17187
rect 29733 17187 29791 17193
rect 29733 17184 29745 17187
rect 25961 17147 26019 17153
rect 29564 17156 29745 17184
rect 26234 17116 26240 17128
rect 25884 17088 26240 17116
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 27801 17119 27859 17125
rect 27801 17085 27813 17119
rect 27847 17085 27859 17119
rect 27801 17079 27859 17085
rect 14384 17020 17632 17048
rect 12216 16952 12756 16980
rect 12216 16940 12222 16952
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 14366 16980 14372 16992
rect 13872 16952 14372 16980
rect 13872 16940 13878 16952
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 20993 16983 21051 16989
rect 20993 16980 21005 16983
rect 19852 16952 21005 16980
rect 19852 16940 19858 16952
rect 20993 16949 21005 16952
rect 21039 16949 21051 16983
rect 20993 16943 21051 16949
rect 23658 16940 23664 16992
rect 23716 16940 23722 16992
rect 26602 16940 26608 16992
rect 26660 16940 26666 16992
rect 27249 16983 27307 16989
rect 27249 16949 27261 16983
rect 27295 16980 27307 16983
rect 27338 16980 27344 16992
rect 27295 16952 27344 16980
rect 27295 16949 27307 16952
rect 27249 16943 27307 16949
rect 27338 16940 27344 16952
rect 27396 16980 27402 16992
rect 27816 16980 27844 17079
rect 29564 16992 29592 17156
rect 29733 17153 29745 17156
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 31481 17187 31539 17193
rect 31481 17153 31493 17187
rect 31527 17184 31539 17187
rect 31726 17184 31754 17292
rect 31846 17280 31852 17292
rect 31904 17280 31910 17332
rect 33134 17280 33140 17332
rect 33192 17280 33198 17332
rect 33781 17323 33839 17329
rect 33781 17289 33793 17323
rect 33827 17320 33839 17323
rect 33962 17320 33968 17332
rect 33827 17292 33968 17320
rect 33827 17289 33839 17292
rect 33781 17283 33839 17289
rect 33962 17280 33968 17292
rect 34020 17280 34026 17332
rect 34241 17323 34299 17329
rect 34241 17289 34253 17323
rect 34287 17320 34299 17323
rect 35342 17320 35348 17332
rect 34287 17292 35348 17320
rect 34287 17289 34299 17292
rect 34241 17283 34299 17289
rect 35342 17280 35348 17292
rect 35400 17280 35406 17332
rect 40034 17280 40040 17332
rect 40092 17280 40098 17332
rect 40678 17280 40684 17332
rect 40736 17280 40742 17332
rect 40770 17280 40776 17332
rect 40828 17320 40834 17332
rect 41233 17323 41291 17329
rect 41233 17320 41245 17323
rect 40828 17292 41245 17320
rect 40828 17280 40834 17292
rect 41233 17289 41245 17292
rect 41279 17289 41291 17323
rect 41233 17283 41291 17289
rect 41506 17280 41512 17332
rect 41564 17280 41570 17332
rect 44910 17320 44916 17332
rect 42720 17292 44916 17320
rect 32392 17255 32450 17261
rect 32392 17221 32404 17255
rect 32438 17252 32450 17255
rect 33152 17252 33180 17280
rect 32438 17224 33180 17252
rect 32438 17221 32450 17224
rect 32392 17215 32450 17221
rect 35250 17212 35256 17264
rect 35308 17252 35314 17264
rect 37553 17255 37611 17261
rect 37553 17252 37565 17255
rect 35308 17224 37565 17252
rect 35308 17212 35314 17224
rect 37553 17221 37565 17224
rect 37599 17252 37611 17255
rect 37599 17224 38056 17252
rect 37599 17221 37611 17224
rect 37553 17215 37611 17221
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 31527 17156 32137 17184
rect 31527 17153 31539 17156
rect 31481 17147 31539 17153
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32766 17144 32772 17196
rect 32824 17184 32830 17196
rect 34149 17187 34207 17193
rect 34149 17184 34161 17187
rect 32824 17156 34161 17184
rect 32824 17144 32830 17156
rect 34149 17153 34161 17156
rect 34195 17184 34207 17187
rect 35161 17187 35219 17193
rect 34195 17156 34928 17184
rect 34195 17153 34207 17156
rect 34149 17147 34207 17153
rect 34900 17128 34928 17156
rect 35161 17153 35173 17187
rect 35207 17184 35219 17187
rect 36265 17187 36323 17193
rect 36265 17184 36277 17187
rect 35207 17156 36277 17184
rect 35207 17153 35219 17156
rect 35161 17147 35219 17153
rect 36265 17153 36277 17156
rect 36311 17153 36323 17187
rect 36265 17147 36323 17153
rect 33318 17076 33324 17128
rect 33376 17116 33382 17128
rect 34333 17119 34391 17125
rect 34333 17116 34345 17119
rect 33376 17088 34345 17116
rect 33376 17076 33382 17088
rect 34333 17085 34345 17088
rect 34379 17085 34391 17119
rect 34333 17079 34391 17085
rect 34882 17076 34888 17128
rect 34940 17116 34946 17128
rect 35253 17119 35311 17125
rect 35253 17116 35265 17119
rect 34940 17088 35265 17116
rect 34940 17076 34946 17088
rect 35253 17085 35265 17088
rect 35299 17085 35311 17119
rect 35253 17079 35311 17085
rect 35434 17076 35440 17128
rect 35492 17076 35498 17128
rect 35618 17076 35624 17128
rect 35676 17076 35682 17128
rect 36357 17119 36415 17125
rect 36357 17085 36369 17119
rect 36403 17085 36415 17119
rect 36357 17079 36415 17085
rect 37921 17119 37979 17125
rect 37921 17085 37933 17119
rect 37967 17085 37979 17119
rect 38028 17116 38056 17224
rect 38102 17144 38108 17196
rect 38160 17144 38166 17196
rect 39853 17187 39911 17193
rect 39853 17153 39865 17187
rect 39899 17184 39911 17187
rect 40052 17184 40080 17280
rect 40120 17255 40178 17261
rect 40120 17221 40132 17255
rect 40166 17252 40178 17255
rect 40696 17252 40724 17280
rect 42720 17264 42748 17292
rect 44910 17280 44916 17292
rect 44968 17280 44974 17332
rect 47394 17280 47400 17332
rect 47452 17280 47458 17332
rect 47486 17280 47492 17332
rect 47544 17320 47550 17332
rect 47581 17323 47639 17329
rect 47581 17320 47593 17323
rect 47544 17292 47593 17320
rect 47544 17280 47550 17292
rect 47581 17289 47593 17292
rect 47627 17289 47639 17323
rect 47581 17283 47639 17289
rect 47949 17323 48007 17329
rect 47949 17289 47961 17323
rect 47995 17320 48007 17323
rect 48222 17320 48228 17332
rect 47995 17292 48228 17320
rect 47995 17289 48007 17292
rect 47949 17283 48007 17289
rect 48222 17280 48228 17292
rect 48280 17280 48286 17332
rect 49329 17323 49387 17329
rect 49329 17320 49341 17323
rect 48700 17292 49341 17320
rect 40166 17224 40724 17252
rect 40166 17221 40178 17224
rect 40120 17215 40178 17221
rect 42702 17212 42708 17264
rect 42760 17212 42766 17264
rect 48314 17252 48320 17264
rect 46032 17224 48320 17252
rect 46032 17193 46060 17224
rect 48314 17212 48320 17224
rect 48372 17212 48378 17264
rect 39899 17156 40080 17184
rect 41877 17187 41935 17193
rect 39899 17153 39911 17156
rect 39853 17147 39911 17153
rect 41877 17153 41889 17187
rect 41923 17184 41935 17187
rect 43073 17187 43131 17193
rect 43073 17184 43085 17187
rect 41923 17156 43085 17184
rect 41923 17153 41935 17156
rect 41877 17147 41935 17153
rect 43073 17153 43085 17156
rect 43119 17153 43131 17187
rect 43073 17147 43131 17153
rect 43800 17187 43858 17193
rect 43800 17153 43812 17187
rect 43846 17184 43858 17187
rect 45649 17187 45707 17193
rect 45649 17184 45661 17187
rect 43846 17156 45661 17184
rect 43846 17153 43858 17156
rect 43800 17147 43858 17153
rect 45649 17153 45661 17156
rect 45695 17153 45707 17187
rect 45649 17147 45707 17153
rect 46017 17187 46075 17193
rect 46017 17153 46029 17187
rect 46063 17153 46075 17187
rect 46017 17147 46075 17153
rect 46284 17187 46342 17193
rect 46284 17153 46296 17187
rect 46330 17184 46342 17187
rect 47118 17184 47124 17196
rect 46330 17156 47124 17184
rect 46330 17153 46342 17156
rect 46284 17147 46342 17153
rect 47118 17144 47124 17156
rect 47176 17144 47182 17196
rect 47302 17144 47308 17196
rect 47360 17184 47366 17196
rect 48041 17187 48099 17193
rect 48041 17184 48053 17187
rect 47360 17156 48053 17184
rect 47360 17144 47366 17156
rect 48041 17153 48053 17156
rect 48087 17184 48099 17187
rect 48700 17184 48728 17292
rect 49329 17289 49341 17292
rect 49375 17320 49387 17323
rect 49510 17320 49516 17332
rect 49375 17292 49516 17320
rect 49375 17289 49387 17292
rect 49329 17283 49387 17289
rect 49510 17280 49516 17292
rect 49568 17320 49574 17332
rect 49970 17320 49976 17332
rect 49568 17292 49976 17320
rect 49568 17280 49574 17292
rect 49970 17280 49976 17292
rect 50028 17280 50034 17332
rect 52733 17323 52791 17329
rect 52733 17289 52745 17323
rect 52779 17320 52791 17323
rect 52822 17320 52828 17332
rect 52779 17292 52828 17320
rect 52779 17289 52791 17292
rect 52733 17283 52791 17289
rect 52822 17280 52828 17292
rect 52880 17280 52886 17332
rect 53193 17323 53251 17329
rect 53193 17289 53205 17323
rect 53239 17320 53251 17323
rect 53374 17320 53380 17332
rect 53239 17292 53380 17320
rect 53239 17289 53251 17292
rect 53193 17283 53251 17289
rect 53374 17280 53380 17292
rect 53432 17280 53438 17332
rect 55033 17323 55091 17329
rect 55033 17289 55045 17323
rect 55079 17320 55091 17323
rect 55398 17320 55404 17332
rect 55079 17292 55404 17320
rect 55079 17289 55091 17292
rect 55033 17283 55091 17289
rect 55398 17280 55404 17292
rect 55456 17320 55462 17332
rect 56410 17320 56416 17332
rect 55456 17292 56416 17320
rect 55456 17280 55462 17292
rect 56410 17280 56416 17292
rect 56468 17280 56474 17332
rect 56686 17280 56692 17332
rect 56744 17320 56750 17332
rect 56781 17323 56839 17329
rect 56781 17320 56793 17323
rect 56744 17292 56793 17320
rect 56744 17280 56750 17292
rect 56781 17289 56793 17292
rect 56827 17320 56839 17323
rect 58434 17320 58440 17332
rect 56827 17292 58440 17320
rect 56827 17289 56839 17292
rect 56781 17283 56839 17289
rect 58434 17280 58440 17292
rect 58492 17280 58498 17332
rect 52457 17255 52515 17261
rect 52457 17252 52469 17255
rect 48087 17156 48728 17184
rect 49344 17224 52469 17252
rect 48087 17153 48099 17156
rect 48041 17147 48099 17153
rect 38565 17119 38623 17125
rect 38565 17116 38577 17119
rect 38028 17088 38577 17116
rect 37921 17079 37979 17085
rect 38565 17085 38577 17088
rect 38611 17085 38623 17119
rect 38565 17079 38623 17085
rect 34793 17051 34851 17057
rect 34793 17017 34805 17051
rect 34839 17048 34851 17051
rect 36372 17048 36400 17079
rect 34839 17020 36400 17048
rect 34839 17017 34851 17020
rect 34793 17011 34851 17017
rect 28074 16980 28080 16992
rect 27396 16952 28080 16980
rect 27396 16940 27402 16952
rect 28074 16940 28080 16952
rect 28132 16980 28138 16992
rect 28902 16980 28908 16992
rect 28132 16952 28908 16980
rect 28132 16940 28138 16952
rect 28902 16940 28908 16952
rect 28960 16940 28966 16992
rect 29546 16940 29552 16992
rect 29604 16940 29610 16992
rect 33502 16940 33508 16992
rect 33560 16980 33566 16992
rect 34330 16980 34336 16992
rect 33560 16952 34336 16980
rect 33560 16940 33566 16952
rect 34330 16940 34336 16952
rect 34388 16940 34394 16992
rect 35986 16940 35992 16992
rect 36044 16980 36050 16992
rect 37001 16983 37059 16989
rect 37001 16980 37013 16983
rect 36044 16952 37013 16980
rect 36044 16940 36050 16952
rect 37001 16949 37013 16952
rect 37047 16949 37059 16983
rect 37936 16980 37964 17079
rect 38654 17076 38660 17128
rect 38712 17116 38718 17128
rect 39022 17125 39028 17128
rect 38841 17119 38899 17125
rect 38841 17116 38853 17119
rect 38712 17088 38853 17116
rect 38712 17076 38718 17088
rect 38841 17085 38853 17088
rect 38887 17085 38899 17119
rect 38841 17079 38899 17085
rect 38979 17119 39028 17125
rect 38979 17085 38991 17119
rect 39025 17085 39028 17119
rect 38979 17079 39028 17085
rect 39022 17076 39028 17079
rect 39080 17076 39086 17128
rect 39117 17119 39175 17125
rect 39117 17085 39129 17119
rect 39163 17116 39175 17119
rect 39482 17116 39488 17128
rect 39163 17088 39488 17116
rect 39163 17085 39175 17088
rect 39117 17079 39175 17085
rect 39482 17076 39488 17088
rect 39540 17076 39546 17128
rect 41966 17076 41972 17128
rect 42024 17076 42030 17128
rect 42058 17076 42064 17128
rect 42116 17076 42122 17128
rect 42426 17076 42432 17128
rect 42484 17076 42490 17128
rect 43438 17076 43444 17128
rect 43496 17116 43502 17128
rect 43533 17119 43591 17125
rect 43533 17116 43545 17119
rect 43496 17088 43545 17116
rect 43496 17076 43502 17088
rect 43533 17085 43545 17088
rect 43579 17085 43591 17119
rect 43533 17079 43591 17085
rect 45002 17076 45008 17128
rect 45060 17076 45066 17128
rect 48133 17119 48191 17125
rect 48133 17085 48145 17119
rect 48179 17085 48191 17119
rect 48133 17079 48191 17085
rect 38654 16980 38660 16992
rect 37936 16952 38660 16980
rect 37001 16943 37059 16949
rect 38654 16940 38660 16952
rect 38712 16940 38718 16992
rect 39758 16940 39764 16992
rect 39816 16940 39822 16992
rect 41984 16980 42012 17076
rect 42076 17048 42104 17076
rect 48148 17048 48176 17079
rect 49142 17076 49148 17128
rect 49200 17116 49206 17128
rect 49344 17116 49372 17224
rect 52457 17221 52469 17224
rect 52503 17221 52515 17255
rect 52457 17215 52515 17221
rect 49421 17187 49479 17193
rect 49421 17153 49433 17187
rect 49467 17184 49479 17187
rect 51169 17187 51227 17193
rect 51169 17184 51181 17187
rect 49467 17156 51181 17184
rect 49467 17153 49479 17156
rect 49421 17147 49479 17153
rect 51169 17153 51181 17156
rect 51215 17153 51227 17187
rect 51169 17147 51227 17153
rect 49513 17119 49571 17125
rect 49513 17116 49525 17119
rect 49200 17088 49525 17116
rect 49200 17076 49206 17088
rect 49513 17085 49525 17088
rect 49559 17085 49571 17119
rect 49513 17079 49571 17085
rect 49789 17119 49847 17125
rect 49789 17085 49801 17119
rect 49835 17085 49847 17119
rect 49789 17079 49847 17085
rect 48593 17051 48651 17057
rect 48593 17048 48605 17051
rect 42076 17020 43576 17048
rect 42058 16980 42064 16992
rect 41984 16952 42064 16980
rect 42058 16940 42064 16952
rect 42116 16940 42122 16992
rect 43438 16940 43444 16992
rect 43496 16940 43502 16992
rect 43548 16980 43576 17020
rect 48056 17020 48605 17048
rect 48056 16980 48084 17020
rect 48593 17017 48605 17020
rect 48639 17017 48651 17051
rect 48593 17011 48651 17017
rect 48961 17051 49019 17057
rect 48961 17017 48973 17051
rect 49007 17048 49019 17051
rect 49804 17048 49832 17079
rect 50522 17076 50528 17128
rect 50580 17076 50586 17128
rect 52472 17116 52500 17215
rect 53006 17144 53012 17196
rect 53064 17184 53070 17196
rect 53101 17187 53159 17193
rect 53101 17184 53113 17187
rect 53064 17156 53113 17184
rect 53064 17144 53070 17156
rect 53101 17153 53113 17156
rect 53147 17153 53159 17187
rect 53101 17147 53159 17153
rect 53920 17187 53978 17193
rect 53920 17153 53932 17187
rect 53966 17184 53978 17187
rect 55769 17187 55827 17193
rect 55769 17184 55781 17187
rect 53966 17156 55781 17184
rect 53966 17153 53978 17156
rect 53920 17147 53978 17153
rect 55769 17153 55781 17156
rect 55815 17153 55827 17187
rect 55769 17147 55827 17153
rect 56873 17187 56931 17193
rect 56873 17153 56885 17187
rect 56919 17184 56931 17187
rect 58529 17187 58587 17193
rect 58529 17184 58541 17187
rect 56919 17156 58541 17184
rect 56919 17153 56931 17156
rect 56873 17147 56931 17153
rect 58529 17153 58541 17156
rect 58575 17153 58587 17187
rect 58529 17147 58587 17153
rect 53285 17119 53343 17125
rect 53285 17116 53297 17119
rect 52472 17088 53297 17116
rect 53285 17085 53297 17088
rect 53331 17116 53343 17119
rect 53374 17116 53380 17128
rect 53331 17088 53380 17116
rect 53331 17085 53343 17088
rect 53285 17079 53343 17085
rect 53374 17076 53380 17088
rect 53432 17076 53438 17128
rect 53558 17076 53564 17128
rect 53616 17116 53622 17128
rect 53653 17119 53711 17125
rect 53653 17116 53665 17119
rect 53616 17088 53665 17116
rect 53616 17076 53622 17088
rect 53653 17085 53665 17088
rect 53699 17085 53711 17119
rect 53653 17079 53711 17085
rect 49007 17020 49832 17048
rect 49007 17017 49019 17020
rect 48961 17011 49019 17017
rect 43548 16952 48084 16980
rect 48608 16980 48636 17011
rect 49694 16980 49700 16992
rect 48608 16952 49700 16980
rect 49694 16940 49700 16952
rect 49752 16940 49758 16992
rect 50430 16940 50436 16992
rect 50488 16940 50494 16992
rect 53668 16980 53696 17079
rect 55122 17076 55128 17128
rect 55180 17076 55186 17128
rect 56965 17119 57023 17125
rect 56965 17116 56977 17119
rect 56336 17088 56977 17116
rect 56336 16992 56364 17088
rect 56965 17085 56977 17088
rect 57011 17085 57023 17119
rect 56965 17079 57023 17085
rect 57422 17076 57428 17128
rect 57480 17116 57486 17128
rect 57885 17119 57943 17125
rect 57885 17116 57897 17119
rect 57480 17088 57897 17116
rect 57480 17076 57486 17088
rect 57885 17085 57897 17088
rect 57931 17085 57943 17119
rect 57885 17079 57943 17085
rect 53834 16980 53840 16992
rect 53668 16952 53840 16980
rect 53834 16940 53840 16952
rect 53892 16940 53898 16992
rect 56318 16940 56324 16992
rect 56376 16940 56382 16992
rect 56410 16940 56416 16992
rect 56468 16940 56474 16992
rect 57422 16940 57428 16992
rect 57480 16940 57486 16992
rect 1104 16890 58880 16912
rect 1104 16838 8172 16890
rect 8224 16838 8236 16890
rect 8288 16838 8300 16890
rect 8352 16838 8364 16890
rect 8416 16838 8428 16890
rect 8480 16838 22616 16890
rect 22668 16838 22680 16890
rect 22732 16838 22744 16890
rect 22796 16838 22808 16890
rect 22860 16838 22872 16890
rect 22924 16838 37060 16890
rect 37112 16838 37124 16890
rect 37176 16838 37188 16890
rect 37240 16838 37252 16890
rect 37304 16838 37316 16890
rect 37368 16838 51504 16890
rect 51556 16838 51568 16890
rect 51620 16838 51632 16890
rect 51684 16838 51696 16890
rect 51748 16838 51760 16890
rect 51812 16838 58880 16890
rect 1104 16816 58880 16838
rect 2774 16736 2780 16788
rect 2832 16736 2838 16788
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 4522 16776 4528 16788
rect 3384 16748 4528 16776
rect 3384 16736 3390 16748
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 5902 16736 5908 16788
rect 5960 16776 5966 16788
rect 6089 16779 6147 16785
rect 6089 16776 6101 16779
rect 5960 16748 6101 16776
rect 5960 16736 5966 16748
rect 6089 16745 6101 16748
rect 6135 16745 6147 16779
rect 6089 16739 6147 16745
rect 6914 16736 6920 16788
rect 6972 16736 6978 16788
rect 10686 16776 10692 16788
rect 9324 16748 10692 16776
rect 2869 16711 2927 16717
rect 2869 16708 2881 16711
rect 2240 16680 2881 16708
rect 2240 16649 2268 16680
rect 2869 16677 2881 16680
rect 2915 16677 2927 16711
rect 2869 16671 2927 16677
rect 3344 16649 3372 16736
rect 8570 16708 8576 16720
rect 3712 16680 8576 16708
rect 3712 16652 3740 16680
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 8754 16668 8760 16720
rect 8812 16708 8818 16720
rect 9324 16717 9352 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11422 16736 11428 16788
rect 11480 16736 11486 16788
rect 11882 16736 11888 16788
rect 11940 16736 11946 16788
rect 12158 16736 12164 16788
rect 12216 16736 12222 16788
rect 14090 16776 14096 16788
rect 12360 16748 14096 16776
rect 9309 16711 9367 16717
rect 9309 16708 9321 16711
rect 8812 16680 9321 16708
rect 8812 16668 8818 16680
rect 9309 16677 9321 16680
rect 9355 16677 9367 16711
rect 9309 16671 9367 16677
rect 9490 16668 9496 16720
rect 9548 16708 9554 16720
rect 9677 16711 9735 16717
rect 9677 16708 9689 16711
rect 9548 16680 9689 16708
rect 9548 16668 9554 16680
rect 9677 16677 9689 16680
rect 9723 16708 9735 16711
rect 9766 16708 9772 16720
rect 9723 16680 9772 16708
rect 9723 16677 9735 16680
rect 9677 16671 9735 16677
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 2225 16643 2283 16649
rect 2225 16609 2237 16643
rect 2271 16609 2283 16643
rect 2225 16603 2283 16609
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16609 3387 16643
rect 3329 16603 3387 16609
rect 3513 16643 3571 16649
rect 3513 16609 3525 16643
rect 3559 16640 3571 16643
rect 3694 16640 3700 16652
rect 3559 16612 3700 16640
rect 3559 16609 3571 16612
rect 3513 16603 3571 16609
rect 3694 16600 3700 16612
rect 3752 16600 3758 16652
rect 3881 16643 3939 16649
rect 3881 16609 3893 16643
rect 3927 16640 3939 16643
rect 4890 16640 4896 16652
rect 3927 16612 4896 16640
rect 3927 16609 3939 16612
rect 3881 16603 3939 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 5813 16643 5871 16649
rect 5813 16640 5825 16643
rect 5040 16612 5825 16640
rect 5040 16600 5046 16612
rect 5813 16609 5825 16612
rect 5859 16640 5871 16643
rect 5859 16612 6316 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 6288 16572 6316 16612
rect 6362 16600 6368 16652
rect 6420 16600 6426 16652
rect 8478 16640 8484 16652
rect 6472 16612 8484 16640
rect 6472 16572 6500 16612
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 8588 16640 8616 16668
rect 11333 16643 11391 16649
rect 8588 16612 11008 16640
rect 6288 16544 6500 16572
rect 3237 16507 3295 16513
rect 3237 16473 3249 16507
rect 3283 16504 3295 16507
rect 4433 16507 4491 16513
rect 4433 16504 4445 16507
rect 3283 16476 4445 16504
rect 3283 16473 3295 16476
rect 3237 16467 3295 16473
rect 4433 16473 4445 16476
rect 4479 16473 4491 16507
rect 10980 16504 11008 16612
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 11440 16640 11468 16736
rect 11379 16612 11468 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 12360 16581 12388 16748
rect 14090 16736 14096 16748
rect 14148 16776 14154 16788
rect 18325 16779 18383 16785
rect 14148 16748 16988 16776
rect 14148 16736 14154 16748
rect 13725 16711 13783 16717
rect 13725 16677 13737 16711
rect 13771 16708 13783 16711
rect 13906 16708 13912 16720
rect 13771 16680 13912 16708
rect 13771 16677 13783 16680
rect 13725 16671 13783 16677
rect 13906 16668 13912 16680
rect 13964 16708 13970 16720
rect 13964 16680 14872 16708
rect 13964 16668 13970 16680
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 14182 16640 14188 16652
rect 14139 16612 14188 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16609 14335 16643
rect 14277 16603 14335 16609
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12124 16544 12357 16572
rect 12124 16532 12130 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12612 16575 12670 16581
rect 12612 16541 12624 16575
rect 12658 16572 12670 16575
rect 13446 16572 13452 16584
rect 12658 16544 13452 16572
rect 12658 16541 12670 16544
rect 12612 16535 12670 16541
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 10980 16476 14228 16504
rect 4433 16467 4491 16473
rect 14200 16448 14228 16476
rect 14182 16396 14188 16448
rect 14240 16396 14246 16448
rect 14292 16436 14320 16603
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 14737 16643 14795 16649
rect 14737 16640 14749 16643
rect 14424 16612 14749 16640
rect 14424 16600 14430 16612
rect 14737 16609 14749 16612
rect 14783 16609 14795 16643
rect 14844 16640 14872 16680
rect 16390 16668 16396 16720
rect 16448 16708 16454 16720
rect 16448 16680 16620 16708
rect 16448 16668 16454 16680
rect 15013 16643 15071 16649
rect 15013 16640 15025 16643
rect 14844 16612 15025 16640
rect 14737 16603 14795 16609
rect 15013 16609 15025 16612
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 15286 16600 15292 16652
rect 15344 16600 15350 16652
rect 16592 16649 16620 16680
rect 16960 16652 16988 16748
rect 18325 16745 18337 16779
rect 18371 16776 18383 16779
rect 18598 16776 18604 16788
rect 18371 16748 18604 16776
rect 18371 16745 18383 16748
rect 18325 16739 18383 16745
rect 18598 16736 18604 16748
rect 18656 16776 18662 16788
rect 20162 16776 20168 16788
rect 18656 16748 20168 16776
rect 18656 16736 18662 16748
rect 20162 16736 20168 16748
rect 20220 16736 20226 16788
rect 20254 16736 20260 16788
rect 20312 16776 20318 16788
rect 22189 16779 22247 16785
rect 22189 16776 22201 16779
rect 20312 16748 22201 16776
rect 20312 16736 20318 16748
rect 19260 16680 20024 16708
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 15979 16612 16497 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 16942 16600 16948 16652
rect 17000 16600 17006 16652
rect 19260 16649 19288 16680
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16609 19303 16643
rect 19245 16603 19303 16609
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19794 16640 19800 16652
rect 19475 16612 19800 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 19794 16600 19800 16612
rect 19852 16600 19858 16652
rect 19886 16600 19892 16652
rect 19944 16600 19950 16652
rect 19996 16640 20024 16680
rect 20806 16640 20812 16652
rect 19996 16612 20812 16640
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 21085 16643 21143 16649
rect 21085 16609 21097 16643
rect 21131 16640 21143 16643
rect 21637 16643 21695 16649
rect 21637 16640 21649 16643
rect 21131 16612 21649 16640
rect 21131 16609 21143 16612
rect 21085 16603 21143 16609
rect 21637 16609 21649 16612
rect 21683 16609 21695 16643
rect 21637 16603 21695 16609
rect 21821 16643 21879 16649
rect 21821 16609 21833 16643
rect 21867 16640 21879 16643
rect 22066 16640 22094 16748
rect 22189 16745 22201 16748
rect 22235 16776 22247 16779
rect 23290 16776 23296 16788
rect 22235 16748 23296 16776
rect 22235 16745 22247 16748
rect 22189 16739 22247 16745
rect 23290 16736 23296 16748
rect 23348 16736 23354 16788
rect 23658 16736 23664 16788
rect 23716 16736 23722 16788
rect 23750 16736 23756 16788
rect 23808 16736 23814 16788
rect 24121 16779 24179 16785
rect 24121 16745 24133 16779
rect 24167 16776 24179 16779
rect 24394 16776 24400 16788
rect 24167 16748 24400 16776
rect 24167 16745 24179 16748
rect 24121 16739 24179 16745
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 25682 16776 25688 16788
rect 24912 16748 25688 16776
rect 24912 16736 24918 16748
rect 25682 16736 25688 16748
rect 25740 16776 25746 16788
rect 25740 16748 28856 16776
rect 25740 16736 25746 16748
rect 21867 16612 22094 16640
rect 23201 16643 23259 16649
rect 21867 16609 21879 16612
rect 21821 16603 21879 16609
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 23676 16640 23704 16736
rect 24026 16668 24032 16720
rect 24084 16708 24090 16720
rect 26602 16708 26608 16720
rect 24084 16680 25452 16708
rect 24084 16668 24090 16680
rect 23247 16612 23704 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 24854 16600 24860 16652
rect 24912 16600 24918 16652
rect 15102 16532 15108 16584
rect 15160 16581 15166 16584
rect 15160 16575 15188 16581
rect 15176 16541 15188 16575
rect 15160 16535 15188 16541
rect 15160 16532 15166 16535
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16393 16575 16451 16581
rect 16393 16572 16405 16575
rect 16172 16544 16405 16572
rect 16172 16532 16178 16544
rect 16393 16541 16405 16544
rect 16439 16541 16451 16575
rect 16393 16535 16451 16541
rect 17212 16575 17270 16581
rect 17212 16541 17224 16575
rect 17258 16572 17270 16575
rect 18138 16572 18144 16584
rect 17258 16544 18144 16572
rect 17258 16541 17270 16544
rect 17212 16535 17270 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 18564 16544 19196 16572
rect 18564 16532 18570 16544
rect 15194 16436 15200 16448
rect 14292 16408 15200 16436
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 15286 16396 15292 16448
rect 15344 16436 15350 16448
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 15344 16408 16037 16436
rect 15344 16396 15350 16408
rect 16025 16405 16037 16408
rect 16071 16405 16083 16439
rect 16025 16399 16083 16405
rect 19058 16396 19064 16448
rect 19116 16396 19122 16448
rect 19168 16436 19196 16544
rect 20162 16532 20168 16584
rect 20220 16532 20226 16584
rect 20254 16532 20260 16584
rect 20312 16581 20318 16584
rect 20312 16575 20340 16581
rect 20328 16541 20340 16575
rect 20312 16535 20340 16541
rect 20312 16532 20318 16535
rect 20438 16532 20444 16584
rect 20496 16532 20502 16584
rect 25424 16581 25452 16680
rect 25608 16680 26608 16708
rect 25501 16643 25559 16649
rect 25501 16609 25513 16643
rect 25547 16640 25559 16643
rect 25608 16640 25636 16680
rect 26602 16668 26608 16680
rect 26660 16668 26666 16720
rect 28828 16708 28856 16748
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 29365 16779 29423 16785
rect 29365 16776 29377 16779
rect 28960 16748 29377 16776
rect 28960 16736 28966 16748
rect 29365 16745 29377 16748
rect 29411 16776 29423 16779
rect 29825 16779 29883 16785
rect 29825 16776 29837 16779
rect 29411 16748 29837 16776
rect 29411 16745 29423 16748
rect 29365 16739 29423 16745
rect 29825 16745 29837 16748
rect 29871 16776 29883 16779
rect 31662 16776 31668 16788
rect 29871 16748 31668 16776
rect 29871 16745 29883 16748
rect 29825 16739 29883 16745
rect 29086 16708 29092 16720
rect 28828 16680 29092 16708
rect 29086 16668 29092 16680
rect 29144 16668 29150 16720
rect 25547 16612 25636 16640
rect 25547 16609 25559 16612
rect 25501 16603 25559 16609
rect 25682 16600 25688 16652
rect 25740 16600 25746 16652
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 27338 16640 27344 16652
rect 26292 16612 27344 16640
rect 26292 16600 26298 16612
rect 27338 16600 27344 16612
rect 27396 16600 27402 16652
rect 28350 16600 28356 16652
rect 28408 16640 28414 16652
rect 29362 16640 29368 16652
rect 28408 16612 29368 16640
rect 28408 16600 28414 16612
rect 29362 16600 29368 16612
rect 29420 16600 29426 16652
rect 29932 16649 29960 16748
rect 31662 16736 31668 16748
rect 31720 16776 31726 16788
rect 31846 16776 31852 16788
rect 31720 16748 31852 16776
rect 31720 16736 31726 16748
rect 31846 16736 31852 16748
rect 31904 16776 31910 16788
rect 32953 16779 33011 16785
rect 32953 16776 32965 16779
rect 31904 16748 32965 16776
rect 31904 16736 31910 16748
rect 32953 16745 32965 16748
rect 32999 16776 33011 16779
rect 36449 16779 36507 16785
rect 36449 16776 36461 16779
rect 32999 16748 36461 16776
rect 32999 16745 33011 16748
rect 32953 16739 33011 16745
rect 29917 16643 29975 16649
rect 29917 16609 29929 16643
rect 29963 16609 29975 16643
rect 32968 16640 32996 16739
rect 34514 16668 34520 16720
rect 34572 16668 34578 16720
rect 34716 16652 34744 16748
rect 36449 16745 36461 16748
rect 36495 16745 36507 16779
rect 36449 16739 36507 16745
rect 37660 16748 38240 16776
rect 33137 16643 33195 16649
rect 33137 16640 33149 16643
rect 32968 16612 33149 16640
rect 29917 16603 29975 16609
rect 33137 16609 33149 16612
rect 33183 16609 33195 16643
rect 33137 16603 33195 16609
rect 34698 16600 34704 16652
rect 34756 16600 34762 16652
rect 36464 16640 36492 16739
rect 36630 16640 36636 16652
rect 36464 16612 36636 16640
rect 36630 16600 36636 16612
rect 36688 16600 36694 16652
rect 25409 16575 25467 16581
rect 25409 16572 25421 16575
rect 25367 16544 25421 16572
rect 25409 16541 25421 16544
rect 25455 16572 25467 16575
rect 26142 16572 26148 16584
rect 25455 16544 26148 16572
rect 25455 16541 25467 16544
rect 25409 16535 25467 16541
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26697 16575 26755 16581
rect 26697 16541 26709 16575
rect 26743 16572 26755 16575
rect 27608 16575 27666 16581
rect 26743 16544 27568 16572
rect 26743 16541 26755 16544
rect 26697 16535 26755 16541
rect 21082 16464 21088 16516
rect 21140 16504 21146 16516
rect 21545 16507 21603 16513
rect 21545 16504 21557 16507
rect 21140 16476 21557 16504
rect 21140 16464 21146 16476
rect 21545 16473 21557 16476
rect 21591 16473 21603 16507
rect 21545 16467 21603 16473
rect 26237 16507 26295 16513
rect 26237 16473 26249 16507
rect 26283 16504 26295 16507
rect 26970 16504 26976 16516
rect 26283 16476 26976 16504
rect 26283 16473 26295 16476
rect 26237 16467 26295 16473
rect 26970 16464 26976 16476
rect 27028 16464 27034 16516
rect 27540 16504 27568 16544
rect 27608 16541 27620 16575
rect 27654 16572 27666 16575
rect 27890 16572 27896 16584
rect 27654 16544 27896 16572
rect 27654 16541 27666 16544
rect 27608 16535 27666 16541
rect 27890 16532 27896 16544
rect 27948 16532 27954 16584
rect 30184 16575 30242 16581
rect 30184 16541 30196 16575
rect 30230 16572 30242 16575
rect 30466 16572 30472 16584
rect 30230 16544 30472 16572
rect 30230 16541 30242 16544
rect 30184 16535 30242 16541
rect 30466 16532 30472 16544
rect 30524 16532 30530 16584
rect 32122 16532 32128 16584
rect 32180 16532 32186 16584
rect 33404 16575 33462 16581
rect 33404 16541 33416 16575
rect 33450 16572 33462 16575
rect 34606 16572 34612 16584
rect 33450 16544 34612 16572
rect 33450 16541 33462 16544
rect 33404 16535 33462 16541
rect 34606 16532 34612 16544
rect 34664 16532 34670 16584
rect 34968 16575 35026 16581
rect 34968 16541 34980 16575
rect 35014 16572 35026 16575
rect 35986 16572 35992 16584
rect 35014 16544 35992 16572
rect 35014 16541 35026 16544
rect 34968 16535 35026 16541
rect 35986 16532 35992 16544
rect 36044 16532 36050 16584
rect 37660 16572 37688 16748
rect 38013 16711 38071 16717
rect 38013 16677 38025 16711
rect 38059 16677 38071 16711
rect 38013 16671 38071 16677
rect 36096 16544 37688 16572
rect 38028 16572 38056 16671
rect 38212 16652 38240 16748
rect 38930 16736 38936 16788
rect 38988 16736 38994 16788
rect 39853 16779 39911 16785
rect 39853 16745 39865 16779
rect 39899 16776 39911 16779
rect 40126 16776 40132 16788
rect 39899 16748 40132 16776
rect 39899 16745 39911 16748
rect 39853 16739 39911 16745
rect 40126 16736 40132 16748
rect 40184 16736 40190 16788
rect 42153 16779 42211 16785
rect 40236 16748 41828 16776
rect 40236 16708 40264 16748
rect 39592 16680 40264 16708
rect 38194 16600 38200 16652
rect 38252 16640 38258 16652
rect 38657 16643 38715 16649
rect 38657 16640 38669 16643
rect 38252 16612 38669 16640
rect 38252 16600 38258 16612
rect 38657 16609 38669 16612
rect 38703 16609 38715 16643
rect 38657 16603 38715 16609
rect 39482 16600 39488 16652
rect 39540 16640 39546 16652
rect 39592 16649 39620 16680
rect 41800 16652 41828 16748
rect 42153 16745 42165 16779
rect 42199 16776 42211 16779
rect 42426 16776 42432 16788
rect 42199 16748 42432 16776
rect 42199 16745 42211 16748
rect 42153 16739 42211 16745
rect 42426 16736 42432 16748
rect 42484 16776 42490 16788
rect 42484 16748 43484 16776
rect 42484 16736 42490 16748
rect 39577 16643 39635 16649
rect 39577 16640 39589 16643
rect 39540 16612 39589 16640
rect 39540 16600 39546 16612
rect 39577 16609 39589 16612
rect 39623 16609 39635 16643
rect 39577 16603 39635 16609
rect 40034 16600 40040 16652
rect 40092 16600 40098 16652
rect 40402 16600 40408 16652
rect 40460 16600 40466 16652
rect 41782 16600 41788 16652
rect 41840 16600 41846 16652
rect 42702 16600 42708 16652
rect 42760 16600 42766 16652
rect 43254 16600 43260 16652
rect 43312 16640 43318 16652
rect 43349 16643 43407 16649
rect 43349 16640 43361 16643
rect 43312 16612 43361 16640
rect 43312 16600 43318 16612
rect 43349 16609 43361 16612
rect 43395 16609 43407 16643
rect 43456 16640 43484 16748
rect 44082 16736 44088 16788
rect 44140 16776 44146 16788
rect 44545 16779 44603 16785
rect 44140 16748 44312 16776
rect 44140 16736 44146 16748
rect 44284 16708 44312 16748
rect 44545 16745 44557 16779
rect 44591 16776 44603 16779
rect 44634 16776 44640 16788
rect 44591 16748 44640 16776
rect 44591 16745 44603 16748
rect 44545 16739 44603 16745
rect 44634 16736 44640 16748
rect 44692 16736 44698 16788
rect 45002 16736 45008 16788
rect 45060 16736 45066 16788
rect 47486 16776 47492 16788
rect 46032 16748 47492 16776
rect 46032 16717 46060 16748
rect 47486 16736 47492 16748
rect 47544 16736 47550 16788
rect 48130 16736 48136 16788
rect 48188 16776 48194 16788
rect 49789 16779 49847 16785
rect 49789 16776 49801 16779
rect 48188 16748 49801 16776
rect 48188 16736 48194 16748
rect 49789 16745 49801 16748
rect 49835 16776 49847 16779
rect 50522 16776 50528 16788
rect 49835 16748 50528 16776
rect 49835 16745 49847 16748
rect 49789 16739 49847 16745
rect 50522 16736 50528 16748
rect 50580 16736 50586 16788
rect 51902 16776 51908 16788
rect 51736 16748 51908 16776
rect 46017 16711 46075 16717
rect 46017 16708 46029 16711
rect 44284 16680 46029 16708
rect 43742 16643 43800 16649
rect 43742 16640 43754 16643
rect 43456 16612 43754 16640
rect 43349 16603 43407 16609
rect 43742 16609 43754 16612
rect 43788 16609 43800 16643
rect 44284 16640 44312 16680
rect 46017 16677 46029 16680
rect 46063 16677 46075 16711
rect 46017 16671 46075 16677
rect 43742 16603 43800 16609
rect 43916 16612 44312 16640
rect 39022 16572 39028 16584
rect 38028 16544 39028 16572
rect 27540 16476 28764 16504
rect 20254 16436 20260 16448
rect 19168 16408 20260 16436
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 20956 16408 21189 16436
rect 20956 16396 20962 16408
rect 21177 16405 21189 16408
rect 21223 16405 21235 16439
rect 21177 16399 21235 16405
rect 25038 16396 25044 16448
rect 25096 16396 25102 16448
rect 27249 16439 27307 16445
rect 27249 16405 27261 16439
rect 27295 16436 27307 16439
rect 28074 16436 28080 16448
rect 27295 16408 28080 16436
rect 27295 16405 27307 16408
rect 27249 16399 27307 16405
rect 28074 16396 28080 16408
rect 28132 16396 28138 16448
rect 28736 16445 28764 16476
rect 33502 16464 33508 16516
rect 33560 16504 33566 16516
rect 36096 16504 36124 16544
rect 39022 16532 39028 16544
rect 39080 16532 39086 16584
rect 40052 16572 40080 16600
rect 40773 16575 40831 16581
rect 40773 16572 40785 16575
rect 40052 16544 40785 16572
rect 40773 16541 40785 16544
rect 40819 16541 40831 16575
rect 40773 16535 40831 16541
rect 41040 16575 41098 16581
rect 41040 16541 41052 16575
rect 41086 16572 41098 16575
rect 42150 16572 42156 16584
rect 41086 16544 42156 16572
rect 41086 16541 41098 16544
rect 41040 16535 41098 16541
rect 42150 16532 42156 16544
rect 42208 16532 42214 16584
rect 42889 16575 42947 16581
rect 42889 16541 42901 16575
rect 42935 16541 42947 16575
rect 42889 16535 42947 16541
rect 33560 16476 36124 16504
rect 36900 16507 36958 16513
rect 33560 16464 33566 16476
rect 36900 16473 36912 16507
rect 36946 16504 36958 16507
rect 38194 16504 38200 16516
rect 36946 16476 38200 16504
rect 36946 16473 36958 16476
rect 36900 16467 36958 16473
rect 38194 16464 38200 16476
rect 38252 16464 38258 16516
rect 40221 16507 40279 16513
rect 39316 16476 39528 16504
rect 39316 16448 39344 16476
rect 28721 16439 28779 16445
rect 28721 16405 28733 16439
rect 28767 16436 28779 16439
rect 28810 16436 28816 16448
rect 28767 16408 28816 16436
rect 28767 16405 28779 16408
rect 28721 16399 28779 16405
rect 28810 16396 28816 16408
rect 28868 16396 28874 16448
rect 30374 16396 30380 16448
rect 30432 16436 30438 16448
rect 31110 16436 31116 16448
rect 30432 16408 31116 16436
rect 30432 16396 30438 16408
rect 31110 16396 31116 16408
rect 31168 16436 31174 16448
rect 31297 16439 31355 16445
rect 31297 16436 31309 16439
rect 31168 16408 31309 16436
rect 31168 16396 31174 16408
rect 31297 16405 31309 16408
rect 31343 16405 31355 16439
rect 31297 16399 31355 16405
rect 32674 16396 32680 16448
rect 32732 16396 32738 16448
rect 34606 16396 34612 16448
rect 34664 16436 34670 16448
rect 35618 16436 35624 16448
rect 34664 16408 35624 16436
rect 34664 16396 34670 16408
rect 35618 16396 35624 16408
rect 35676 16436 35682 16448
rect 36081 16439 36139 16445
rect 36081 16436 36093 16439
rect 35676 16408 36093 16436
rect 35676 16396 35682 16408
rect 36081 16405 36093 16408
rect 36127 16405 36139 16439
rect 36081 16399 36139 16405
rect 38102 16396 38108 16448
rect 38160 16396 38166 16448
rect 38470 16396 38476 16448
rect 38528 16396 38534 16448
rect 38565 16439 38623 16445
rect 38565 16405 38577 16439
rect 38611 16436 38623 16439
rect 38838 16436 38844 16448
rect 38611 16408 38844 16436
rect 38611 16405 38623 16408
rect 38565 16399 38623 16405
rect 38838 16396 38844 16408
rect 38896 16436 38902 16448
rect 39298 16436 39304 16448
rect 38896 16408 39304 16436
rect 38896 16396 38902 16408
rect 39298 16396 39304 16408
rect 39356 16396 39362 16448
rect 39390 16396 39396 16448
rect 39448 16396 39454 16448
rect 39500 16436 39528 16476
rect 40221 16473 40233 16507
rect 40267 16504 40279 16507
rect 41414 16504 41420 16516
rect 40267 16476 41420 16504
rect 40267 16473 40279 16476
rect 40221 16467 40279 16473
rect 41414 16464 41420 16476
rect 41472 16464 41478 16516
rect 40313 16439 40371 16445
rect 40313 16436 40325 16439
rect 39500 16408 40325 16436
rect 40313 16405 40325 16408
rect 40359 16405 40371 16439
rect 40313 16399 40371 16405
rect 40954 16396 40960 16448
rect 41012 16436 41018 16448
rect 42518 16436 42524 16448
rect 41012 16408 42524 16436
rect 41012 16396 41018 16408
rect 42518 16396 42524 16408
rect 42576 16396 42582 16448
rect 42904 16436 42932 16535
rect 43622 16532 43628 16584
rect 43680 16532 43686 16584
rect 43916 16581 43944 16612
rect 45462 16600 45468 16652
rect 45520 16600 45526 16652
rect 45649 16643 45707 16649
rect 45649 16609 45661 16643
rect 45695 16640 45707 16643
rect 46382 16640 46388 16652
rect 45695 16612 46388 16640
rect 45695 16609 45707 16612
rect 45649 16603 45707 16609
rect 46382 16600 46388 16612
rect 46440 16600 46446 16652
rect 48314 16600 48320 16652
rect 48372 16640 48378 16652
rect 51736 16649 51764 16748
rect 51902 16736 51908 16748
rect 51960 16776 51966 16788
rect 54205 16779 54263 16785
rect 51960 16748 53880 16776
rect 51960 16736 51966 16748
rect 53852 16652 53880 16748
rect 54205 16745 54217 16779
rect 54251 16776 54263 16779
rect 55122 16776 55128 16788
rect 54251 16748 55128 16776
rect 54251 16745 54263 16748
rect 54205 16739 54263 16745
rect 55122 16736 55128 16748
rect 55180 16736 55186 16788
rect 56410 16736 56416 16788
rect 56468 16736 56474 16788
rect 56686 16736 56692 16788
rect 56744 16736 56750 16788
rect 57054 16736 57060 16788
rect 57112 16736 57118 16788
rect 55953 16711 56011 16717
rect 55953 16708 55965 16711
rect 54680 16680 55965 16708
rect 48409 16643 48467 16649
rect 48409 16640 48421 16643
rect 48372 16612 48421 16640
rect 48372 16600 48378 16612
rect 48409 16609 48421 16612
rect 48455 16609 48467 16643
rect 48409 16603 48467 16609
rect 51721 16643 51779 16649
rect 51721 16609 51733 16643
rect 51767 16609 51779 16643
rect 51721 16603 51779 16609
rect 53834 16600 53840 16652
rect 53892 16600 53898 16652
rect 54680 16649 54708 16680
rect 55953 16677 55965 16680
rect 55999 16677 56011 16711
rect 55953 16671 56011 16677
rect 54665 16643 54723 16649
rect 54665 16609 54677 16643
rect 54711 16609 54723 16643
rect 54665 16603 54723 16609
rect 54754 16600 54760 16652
rect 54812 16600 54818 16652
rect 55398 16600 55404 16652
rect 55456 16600 55462 16652
rect 56428 16649 56456 16736
rect 56413 16643 56471 16649
rect 56413 16609 56425 16643
rect 56459 16609 56471 16643
rect 56704 16640 56732 16736
rect 56413 16603 56471 16609
rect 56520 16612 56732 16640
rect 43901 16575 43959 16581
rect 43901 16541 43913 16575
rect 43947 16541 43959 16575
rect 43901 16535 43959 16541
rect 46477 16575 46535 16581
rect 46477 16541 46489 16575
rect 46523 16572 46535 16575
rect 46566 16572 46572 16584
rect 46523 16544 46572 16572
rect 46523 16541 46535 16544
rect 46477 16535 46535 16541
rect 46566 16532 46572 16544
rect 46624 16532 46630 16584
rect 48676 16575 48734 16581
rect 48676 16541 48688 16575
rect 48722 16572 48734 16575
rect 50430 16572 50436 16584
rect 48722 16544 50436 16572
rect 48722 16541 48734 16544
rect 48676 16535 48734 16541
rect 50430 16532 50436 16544
rect 50488 16532 50494 16584
rect 53190 16532 53196 16584
rect 53248 16532 53254 16584
rect 54573 16575 54631 16581
rect 54573 16541 54585 16575
rect 54619 16572 54631 16575
rect 54846 16572 54852 16584
rect 54619 16544 54852 16572
rect 54619 16541 54631 16544
rect 54573 16535 54631 16541
rect 54846 16532 54852 16544
rect 54904 16572 54910 16584
rect 56520 16572 56548 16612
rect 54904 16544 56548 16572
rect 54904 16532 54910 16544
rect 44634 16464 44640 16516
rect 44692 16504 44698 16516
rect 45373 16507 45431 16513
rect 45373 16504 45385 16507
rect 44692 16476 45385 16504
rect 44692 16464 44698 16476
rect 45373 16473 45385 16476
rect 45419 16473 45431 16507
rect 45373 16467 45431 16473
rect 46744 16507 46802 16513
rect 46744 16473 46756 16507
rect 46790 16504 46802 16507
rect 46934 16504 46940 16516
rect 46790 16476 46940 16504
rect 46790 16473 46802 16476
rect 46744 16467 46802 16473
rect 46934 16464 46940 16476
rect 46992 16464 46998 16516
rect 49050 16464 49056 16516
rect 49108 16464 49114 16516
rect 51988 16507 52046 16513
rect 51988 16473 52000 16507
rect 52034 16504 52046 16507
rect 53837 16507 53895 16513
rect 53837 16504 53849 16507
rect 52034 16476 53849 16504
rect 52034 16473 52046 16476
rect 51988 16467 52046 16473
rect 53837 16473 53849 16476
rect 53883 16473 53895 16507
rect 53837 16467 53895 16473
rect 44910 16436 44916 16448
rect 42904 16408 44916 16436
rect 44910 16396 44916 16408
rect 44968 16396 44974 16448
rect 47857 16439 47915 16445
rect 47857 16405 47869 16439
rect 47903 16436 47915 16439
rect 48314 16436 48320 16448
rect 47903 16408 48320 16436
rect 47903 16405 47915 16408
rect 47857 16399 47915 16405
rect 48314 16396 48320 16408
rect 48372 16436 48378 16448
rect 49068 16436 49096 16464
rect 48372 16408 49096 16436
rect 48372 16396 48378 16408
rect 51902 16396 51908 16448
rect 51960 16436 51966 16448
rect 53101 16439 53159 16445
rect 53101 16436 53113 16439
rect 51960 16408 53113 16436
rect 51960 16396 51966 16408
rect 53101 16405 53113 16408
rect 53147 16405 53159 16439
rect 53101 16399 53159 16405
rect 1104 16346 59040 16368
rect 1104 16294 15394 16346
rect 15446 16294 15458 16346
rect 15510 16294 15522 16346
rect 15574 16294 15586 16346
rect 15638 16294 15650 16346
rect 15702 16294 29838 16346
rect 29890 16294 29902 16346
rect 29954 16294 29966 16346
rect 30018 16294 30030 16346
rect 30082 16294 30094 16346
rect 30146 16294 44282 16346
rect 44334 16294 44346 16346
rect 44398 16294 44410 16346
rect 44462 16294 44474 16346
rect 44526 16294 44538 16346
rect 44590 16294 58726 16346
rect 58778 16294 58790 16346
rect 58842 16294 58854 16346
rect 58906 16294 58918 16346
rect 58970 16294 58982 16346
rect 59034 16294 59040 16346
rect 1104 16272 59040 16294
rect 3694 16192 3700 16244
rect 3752 16192 3758 16244
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7984 16204 8217 16232
rect 7984 16192 7990 16204
rect 8205 16201 8217 16204
rect 8251 16232 8263 16235
rect 11606 16232 11612 16244
rect 8251 16204 11612 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13780 16204 14013 16232
rect 13780 16192 13786 16204
rect 14001 16201 14013 16204
rect 14047 16232 14059 16235
rect 14826 16232 14832 16244
rect 14047 16204 14832 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14826 16192 14832 16204
rect 14884 16232 14890 16244
rect 15930 16232 15936 16244
rect 14884 16204 15936 16232
rect 14884 16192 14890 16204
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 18506 16232 18512 16244
rect 18371 16204 18512 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 18785 16235 18843 16241
rect 18785 16201 18797 16235
rect 18831 16232 18843 16235
rect 19058 16232 19064 16244
rect 18831 16204 19064 16232
rect 18831 16201 18843 16204
rect 18785 16195 18843 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 20806 16192 20812 16244
rect 20864 16232 20870 16244
rect 20901 16235 20959 16241
rect 20901 16232 20913 16235
rect 20864 16204 20913 16232
rect 20864 16192 20870 16204
rect 20901 16201 20913 16204
rect 20947 16201 20959 16235
rect 20901 16195 20959 16201
rect 25590 16192 25596 16244
rect 25648 16192 25654 16244
rect 26326 16192 26332 16244
rect 26384 16232 26390 16244
rect 27430 16232 27436 16244
rect 26384 16204 27436 16232
rect 26384 16192 26390 16204
rect 27430 16192 27436 16204
rect 27488 16192 27494 16244
rect 27614 16192 27620 16244
rect 27672 16192 27678 16244
rect 28074 16192 28080 16244
rect 28132 16192 28138 16244
rect 30374 16232 30380 16244
rect 28644 16204 30380 16232
rect 13170 16164 13176 16176
rect 11072 16136 13176 16164
rect 11072 16105 11100 16136
rect 13170 16124 13176 16136
rect 13228 16164 13234 16176
rect 17954 16164 17960 16176
rect 13228 16136 17960 16164
rect 13228 16124 13234 16136
rect 17954 16124 17960 16136
rect 18012 16124 18018 16176
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16164 18935 16167
rect 19334 16164 19340 16176
rect 18923 16136 19340 16164
rect 18923 16133 18935 16136
rect 18877 16127 18935 16133
rect 19334 16124 19340 16136
rect 19392 16164 19398 16176
rect 20254 16164 20260 16176
rect 19392 16136 20260 16164
rect 19392 16124 19398 16136
rect 20254 16124 20260 16136
rect 20312 16124 20318 16176
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 9079 16068 11069 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 11057 16065 11069 16068
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 12336 16099 12394 16105
rect 12336 16065 12348 16099
rect 12382 16096 12394 16099
rect 13630 16096 13636 16108
rect 12382 16068 13636 16096
rect 12382 16065 12394 16068
rect 12336 16059 12394 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16096 13967 16099
rect 15013 16099 15071 16105
rect 15013 16096 15025 16099
rect 13955 16068 15025 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 15013 16065 15025 16068
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 16942 16056 16948 16108
rect 17000 16056 17006 16108
rect 17212 16099 17270 16105
rect 17212 16065 17224 16099
rect 17258 16096 17270 16099
rect 18506 16096 18512 16108
rect 17258 16068 18512 16096
rect 17258 16065 17270 16068
rect 17212 16059 17270 16065
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 19788 16099 19846 16105
rect 19788 16065 19800 16099
rect 19834 16096 19846 16099
rect 21358 16096 21364 16108
rect 19834 16068 21364 16096
rect 19834 16065 19846 16068
rect 19788 16059 19846 16065
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 25038 16056 25044 16108
rect 25096 16056 25102 16108
rect 27982 16056 27988 16108
rect 28040 16096 28046 16108
rect 28350 16096 28356 16108
rect 28040 16068 28356 16096
rect 28040 16056 28046 16068
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28445 16099 28503 16105
rect 28445 16065 28457 16099
rect 28491 16096 28503 16099
rect 28534 16096 28540 16108
rect 28491 16068 28540 16096
rect 28491 16065 28503 16068
rect 28445 16059 28503 16065
rect 28534 16056 28540 16068
rect 28592 16056 28598 16108
rect 28644 16105 28672 16204
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 30745 16235 30803 16241
rect 30745 16201 30757 16235
rect 30791 16232 30803 16235
rect 30926 16232 30932 16244
rect 30791 16204 30932 16232
rect 30791 16201 30803 16204
rect 30745 16195 30803 16201
rect 30926 16192 30932 16204
rect 30984 16192 30990 16244
rect 32122 16192 32128 16244
rect 32180 16232 32186 16244
rect 32217 16235 32275 16241
rect 32217 16232 32229 16235
rect 32180 16204 32229 16232
rect 32180 16192 32186 16204
rect 32217 16201 32229 16204
rect 32263 16201 32275 16235
rect 32217 16195 32275 16201
rect 32677 16235 32735 16241
rect 32677 16201 32689 16235
rect 32723 16232 32735 16235
rect 32766 16232 32772 16244
rect 32723 16204 32772 16232
rect 32723 16201 32735 16204
rect 32677 16195 32735 16201
rect 32766 16192 32772 16204
rect 32824 16192 32830 16244
rect 33318 16192 33324 16244
rect 33376 16192 33382 16244
rect 34514 16232 34520 16244
rect 33428 16204 34520 16232
rect 28629 16099 28687 16105
rect 28629 16065 28641 16099
rect 28675 16065 28687 16099
rect 28629 16059 28687 16065
rect 28810 16056 28816 16108
rect 28868 16056 28874 16108
rect 29638 16056 29644 16108
rect 29696 16056 29702 16108
rect 32585 16099 32643 16105
rect 32585 16065 32597 16099
rect 32631 16096 32643 16099
rect 33134 16096 33140 16108
rect 32631 16068 33140 16096
rect 32631 16065 32643 16068
rect 32585 16059 32643 16065
rect 33134 16056 33140 16068
rect 33192 16056 33198 16108
rect 33428 16105 33456 16204
rect 34514 16192 34520 16204
rect 34572 16192 34578 16244
rect 35713 16235 35771 16241
rect 35713 16201 35725 16235
rect 35759 16232 35771 16235
rect 36538 16232 36544 16244
rect 35759 16204 36544 16232
rect 35759 16201 35771 16204
rect 35713 16195 35771 16201
rect 36538 16192 36544 16204
rect 36596 16192 36602 16244
rect 36630 16192 36636 16244
rect 36688 16232 36694 16244
rect 37001 16235 37059 16241
rect 37001 16232 37013 16235
rect 36688 16204 37013 16232
rect 36688 16192 36694 16204
rect 37001 16201 37013 16204
rect 37047 16201 37059 16235
rect 37001 16195 37059 16201
rect 33413 16099 33471 16105
rect 33413 16065 33425 16099
rect 33459 16065 33471 16099
rect 33413 16059 33471 16065
rect 34330 16056 34336 16108
rect 34388 16056 34394 16108
rect 36722 16096 36728 16108
rect 35176 16068 36728 16096
rect 5442 15988 5448 16040
rect 5500 15988 5506 16040
rect 12066 16028 12072 16040
rect 11440 16000 12072 16028
rect 11440 15904 11468 16000
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 14182 15988 14188 16040
rect 14240 16028 14246 16040
rect 14240 16000 14403 16028
rect 14240 15988 14246 16000
rect 13449 15963 13507 15969
rect 13449 15929 13461 15963
rect 13495 15960 13507 15963
rect 14375 15960 14403 16000
rect 14458 15988 14464 16040
rect 14516 16028 14522 16040
rect 14516 16000 15056 16028
rect 14516 15988 14522 16000
rect 15028 15972 15056 16000
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 19061 16031 19119 16037
rect 19061 15997 19073 16031
rect 19107 16028 19119 16031
rect 19107 16000 19196 16028
rect 19107 15997 19119 16000
rect 19061 15991 19119 15997
rect 13495 15932 14136 15960
rect 14375 15932 14504 15960
rect 13495 15929 13507 15932
rect 13449 15923 13507 15929
rect 5994 15852 6000 15904
rect 6052 15852 6058 15904
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 10321 15895 10379 15901
rect 10321 15892 10333 15895
rect 9640 15864 10333 15892
rect 9640 15852 9646 15864
rect 10321 15861 10333 15864
rect 10367 15892 10379 15895
rect 11054 15892 11060 15904
rect 10367 15864 11060 15892
rect 10367 15861 10379 15864
rect 10321 15855 10379 15861
rect 11054 15852 11060 15864
rect 11112 15892 11118 15904
rect 11422 15892 11428 15904
rect 11112 15864 11428 15892
rect 11112 15852 11118 15864
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 13538 15852 13544 15904
rect 13596 15852 13602 15904
rect 14108 15892 14136 15932
rect 14274 15892 14280 15904
rect 14108 15864 14280 15892
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14476 15892 14504 15932
rect 15010 15920 15016 15972
rect 15068 15920 15074 15972
rect 19168 15960 19196 16000
rect 19518 15988 19524 16040
rect 19576 15988 19582 16040
rect 20806 15988 20812 16040
rect 20864 16028 20870 16040
rect 20993 16031 21051 16037
rect 20993 16028 21005 16031
rect 20864 16000 21005 16028
rect 20864 15988 20870 16000
rect 20993 15997 21005 16000
rect 21039 15997 21051 16031
rect 22462 16028 22468 16040
rect 20993 15991 21051 15997
rect 22066 16000 22468 16028
rect 22066 15960 22094 16000
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 28169 16031 28227 16037
rect 28169 16028 28181 16031
rect 26620 16000 28181 16028
rect 15120 15932 15884 15960
rect 15120 15892 15148 15932
rect 14476 15864 15148 15892
rect 15746 15852 15752 15904
rect 15804 15852 15810 15904
rect 15856 15892 15884 15932
rect 17880 15932 19196 15960
rect 17880 15892 17908 15932
rect 19168 15904 19196 15932
rect 20456 15932 22094 15960
rect 15856 15864 17908 15892
rect 18414 15852 18420 15904
rect 18472 15852 18478 15904
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 20456 15892 20484 15932
rect 26620 15904 26648 16000
rect 28169 15997 28181 16000
rect 28215 15997 28227 16031
rect 28828 16028 28856 16056
rect 29365 16031 29423 16037
rect 29365 16028 29377 16031
rect 28828 16000 29377 16028
rect 28169 15991 28227 15997
rect 29365 15997 29377 16000
rect 29411 15997 29423 16031
rect 29365 15991 29423 15997
rect 29503 16031 29561 16037
rect 29503 15997 29515 16031
rect 29549 16028 29561 16031
rect 30285 16031 30343 16037
rect 29549 16000 30052 16028
rect 29549 15997 29561 16000
rect 29503 15991 29561 15997
rect 26786 15920 26792 15972
rect 26844 15960 26850 15972
rect 28994 15960 29000 15972
rect 26844 15932 29000 15960
rect 26844 15920 26850 15932
rect 28994 15920 29000 15932
rect 29052 15960 29058 15972
rect 29089 15963 29147 15969
rect 29089 15960 29101 15963
rect 29052 15932 29101 15960
rect 29052 15920 29058 15932
rect 29089 15929 29101 15932
rect 29135 15929 29147 15963
rect 29089 15923 29147 15929
rect 19208 15864 20484 15892
rect 19208 15852 19214 15864
rect 21634 15852 21640 15904
rect 21692 15852 21698 15904
rect 23569 15895 23627 15901
rect 23569 15861 23581 15895
rect 23615 15892 23627 15895
rect 24302 15892 24308 15904
rect 23615 15864 24308 15892
rect 23615 15861 23627 15864
rect 23569 15855 23627 15861
rect 24302 15852 24308 15864
rect 24360 15892 24366 15904
rect 26602 15892 26608 15904
rect 24360 15864 26608 15892
rect 24360 15852 24366 15864
rect 26602 15852 26608 15864
rect 26660 15852 26666 15904
rect 28074 15852 28080 15904
rect 28132 15892 28138 15904
rect 30024 15892 30052 16000
rect 30285 15997 30297 16031
rect 30331 16028 30343 16031
rect 30837 16031 30895 16037
rect 30837 16028 30849 16031
rect 30331 16000 30849 16028
rect 30331 15997 30343 16000
rect 30285 15991 30343 15997
rect 30837 15997 30849 16000
rect 30883 15997 30895 16031
rect 30837 15991 30895 15997
rect 30929 16031 30987 16037
rect 30929 15997 30941 16031
rect 30975 15997 30987 16031
rect 30929 15991 30987 15997
rect 32861 16031 32919 16037
rect 32861 15997 32873 16031
rect 32907 16028 32919 16031
rect 33502 16028 33508 16040
rect 32907 16000 33508 16028
rect 32907 15997 32919 16000
rect 32861 15991 32919 15997
rect 30944 15960 30972 15991
rect 33502 15988 33508 16000
rect 33560 15988 33566 16040
rect 33597 16031 33655 16037
rect 33597 15997 33609 16031
rect 33643 15997 33655 16031
rect 33597 15991 33655 15997
rect 30208 15932 30972 15960
rect 30208 15904 30236 15932
rect 28132 15864 30052 15892
rect 28132 15852 28138 15864
rect 30190 15852 30196 15904
rect 30248 15852 30254 15904
rect 30374 15852 30380 15904
rect 30432 15852 30438 15904
rect 33612 15892 33640 15991
rect 34422 15988 34428 16040
rect 34480 16037 34486 16040
rect 34480 16031 34508 16037
rect 34496 15997 34508 16031
rect 34480 15991 34508 15997
rect 34609 16031 34667 16037
rect 34609 15997 34621 16031
rect 34655 16028 34667 16031
rect 34974 16028 34980 16040
rect 34655 16000 34980 16028
rect 34655 15997 34667 16000
rect 34609 15991 34667 15997
rect 34480 15988 34486 15991
rect 34974 15988 34980 16000
rect 35032 16028 35038 16040
rect 35176 16028 35204 16068
rect 36722 16056 36728 16068
rect 36780 16056 36786 16108
rect 37016 16096 37044 16195
rect 38654 16192 38660 16244
rect 38712 16192 38718 16244
rect 39025 16235 39083 16241
rect 39025 16201 39037 16235
rect 39071 16232 39083 16235
rect 39482 16232 39488 16244
rect 39071 16204 39488 16232
rect 39071 16201 39083 16204
rect 39025 16195 39083 16201
rect 39482 16192 39488 16204
rect 39540 16192 39546 16244
rect 39669 16235 39727 16241
rect 39669 16201 39681 16235
rect 39715 16232 39727 16235
rect 39758 16232 39764 16244
rect 39715 16204 39764 16232
rect 39715 16201 39727 16204
rect 39669 16195 39727 16201
rect 39758 16192 39764 16204
rect 39816 16192 39822 16244
rect 40034 16192 40040 16244
rect 40092 16232 40098 16244
rect 40589 16235 40647 16241
rect 40589 16232 40601 16235
rect 40092 16204 40601 16232
rect 40092 16192 40098 16204
rect 40589 16201 40601 16204
rect 40635 16201 40647 16235
rect 40589 16195 40647 16201
rect 42245 16235 42303 16241
rect 42245 16201 42257 16235
rect 42291 16232 42303 16235
rect 42794 16232 42800 16244
rect 42291 16204 42800 16232
rect 42291 16201 42303 16204
rect 42245 16195 42303 16201
rect 42794 16192 42800 16204
rect 42852 16232 42858 16244
rect 43622 16232 43628 16244
rect 42852 16204 43628 16232
rect 42852 16192 42858 16204
rect 43622 16192 43628 16204
rect 43680 16192 43686 16244
rect 43990 16192 43996 16244
rect 44048 16232 44054 16244
rect 44634 16232 44640 16244
rect 44048 16204 44640 16232
rect 44048 16192 44054 16204
rect 44634 16192 44640 16204
rect 44692 16192 44698 16244
rect 44910 16192 44916 16244
rect 44968 16192 44974 16244
rect 45922 16192 45928 16244
rect 45980 16192 45986 16244
rect 47946 16192 47952 16244
rect 48004 16232 48010 16244
rect 48317 16235 48375 16241
rect 48317 16232 48329 16235
rect 48004 16204 48329 16232
rect 48004 16192 48010 16204
rect 48317 16201 48329 16204
rect 48363 16201 48375 16235
rect 48317 16195 48375 16201
rect 51074 16192 51080 16244
rect 51132 16192 51138 16244
rect 51166 16192 51172 16244
rect 51224 16232 51230 16244
rect 51445 16235 51503 16241
rect 51445 16232 51457 16235
rect 51224 16204 51457 16232
rect 51224 16192 51230 16204
rect 51445 16201 51457 16204
rect 51491 16232 51503 16235
rect 52638 16232 52644 16244
rect 51491 16204 52644 16232
rect 51491 16201 51503 16204
rect 51445 16195 51503 16201
rect 52638 16192 52644 16204
rect 52696 16192 52702 16244
rect 52733 16235 52791 16241
rect 52733 16201 52745 16235
rect 52779 16232 52791 16235
rect 53190 16232 53196 16244
rect 52779 16204 53196 16232
rect 52779 16201 52791 16204
rect 52733 16195 52791 16201
rect 53190 16192 53196 16204
rect 53248 16192 53254 16244
rect 54573 16235 54631 16241
rect 54573 16201 54585 16235
rect 54619 16232 54631 16235
rect 54754 16232 54760 16244
rect 54619 16204 54760 16232
rect 54619 16201 54631 16204
rect 54573 16195 54631 16201
rect 54754 16192 54760 16204
rect 54812 16192 54818 16244
rect 37544 16167 37602 16173
rect 37544 16133 37556 16167
rect 37590 16164 37602 16167
rect 38746 16164 38752 16176
rect 37590 16136 38752 16164
rect 37590 16133 37602 16136
rect 37544 16127 37602 16133
rect 38746 16124 38752 16136
rect 38804 16124 38810 16176
rect 39577 16167 39635 16173
rect 39577 16133 39589 16167
rect 39623 16164 39635 16167
rect 40218 16164 40224 16176
rect 39623 16136 40224 16164
rect 39623 16133 39635 16136
rect 39577 16127 39635 16133
rect 40218 16124 40224 16136
rect 40276 16124 40282 16176
rect 40310 16124 40316 16176
rect 40368 16164 40374 16176
rect 56778 16164 56784 16176
rect 40368 16136 56784 16164
rect 40368 16124 40374 16136
rect 56778 16124 56784 16136
rect 56836 16124 56842 16176
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 37016 16068 37289 16096
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37277 16059 37335 16065
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16096 40923 16099
rect 40954 16096 40960 16108
rect 40911 16068 40960 16096
rect 40911 16065 40923 16068
rect 40865 16059 40923 16065
rect 40954 16056 40960 16068
rect 41012 16056 41018 16108
rect 41132 16099 41190 16105
rect 41132 16065 41144 16099
rect 41178 16096 41190 16099
rect 43073 16099 43131 16105
rect 43073 16096 43085 16099
rect 41178 16068 43085 16096
rect 41178 16065 41190 16068
rect 41132 16059 41190 16065
rect 43073 16065 43085 16068
rect 43119 16065 43131 16099
rect 43073 16059 43131 16065
rect 43800 16099 43858 16105
rect 43800 16065 43812 16099
rect 43846 16096 43858 16099
rect 45649 16099 45707 16105
rect 45649 16096 45661 16099
rect 43846 16068 45661 16096
rect 43846 16065 43858 16068
rect 43800 16059 43858 16065
rect 45649 16065 45661 16068
rect 45695 16065 45707 16099
rect 45649 16059 45707 16065
rect 47765 16099 47823 16105
rect 47765 16065 47777 16099
rect 47811 16096 47823 16099
rect 48314 16096 48320 16108
rect 47811 16068 48320 16096
rect 47811 16065 47823 16068
rect 47765 16059 47823 16065
rect 48314 16056 48320 16068
rect 48372 16056 48378 16108
rect 53101 16099 53159 16105
rect 53101 16065 53113 16099
rect 53147 16096 53159 16099
rect 54205 16099 54263 16105
rect 54205 16096 54217 16099
rect 53147 16068 54217 16096
rect 53147 16065 53159 16068
rect 53101 16059 53159 16065
rect 54205 16065 54217 16068
rect 54251 16065 54263 16099
rect 54205 16059 54263 16065
rect 35032 16000 35204 16028
rect 35253 16031 35311 16037
rect 35032 15988 35038 16000
rect 35253 15997 35265 16031
rect 35299 16028 35311 16031
rect 35805 16031 35863 16037
rect 35805 16028 35817 16031
rect 35299 16000 35817 16028
rect 35299 15997 35311 16000
rect 35253 15991 35311 15997
rect 35805 15997 35817 16000
rect 35851 15997 35863 16031
rect 35805 15991 35863 15997
rect 35989 16031 36047 16037
rect 35989 15997 36001 16031
rect 36035 16028 36047 16031
rect 39853 16031 39911 16037
rect 36035 16000 36400 16028
rect 36035 15997 36047 16000
rect 35989 15991 36047 15997
rect 34054 15920 34060 15972
rect 34112 15920 34118 15972
rect 36372 15904 36400 16000
rect 39853 15997 39865 16031
rect 39899 16028 39911 16031
rect 39899 16000 40356 16028
rect 39899 15997 39911 16000
rect 39853 15991 39911 15997
rect 34606 15892 34612 15904
rect 33612 15864 34612 15892
rect 34606 15852 34612 15864
rect 34664 15852 34670 15904
rect 34790 15852 34796 15904
rect 34848 15892 34854 15904
rect 35345 15895 35403 15901
rect 35345 15892 35357 15895
rect 34848 15864 35357 15892
rect 34848 15852 34854 15864
rect 35345 15861 35357 15864
rect 35391 15861 35403 15895
rect 35345 15855 35403 15861
rect 36354 15852 36360 15904
rect 36412 15852 36418 15904
rect 39209 15895 39267 15901
rect 39209 15861 39221 15895
rect 39255 15892 39267 15895
rect 39482 15892 39488 15904
rect 39255 15864 39488 15892
rect 39255 15861 39267 15864
rect 39209 15855 39267 15861
rect 39482 15852 39488 15864
rect 39540 15852 39546 15904
rect 40328 15901 40356 16000
rect 42426 15988 42432 16040
rect 42484 15988 42490 16040
rect 42518 15988 42524 16040
rect 42576 16028 42582 16040
rect 43533 16031 43591 16037
rect 43533 16028 43545 16031
rect 42576 16000 43545 16028
rect 42576 15988 42582 16000
rect 43456 15904 43484 16000
rect 43533 15997 43545 16000
rect 43579 15997 43591 16031
rect 43533 15991 43591 15997
rect 45002 15988 45008 16040
rect 45060 15988 45066 16040
rect 51902 15988 51908 16040
rect 51960 15988 51966 16040
rect 53006 15988 53012 16040
rect 53064 16028 53070 16040
rect 53190 16028 53196 16040
rect 53064 16000 53196 16028
rect 53064 15988 53070 16000
rect 53190 15988 53196 16000
rect 53248 15988 53254 16040
rect 53377 16031 53435 16037
rect 53377 15997 53389 16031
rect 53423 16028 53435 16031
rect 53466 16028 53472 16040
rect 53423 16000 53472 16028
rect 53423 15997 53435 16000
rect 53377 15991 53435 15997
rect 53466 15988 53472 16000
rect 53524 15988 53530 16040
rect 53561 16031 53619 16037
rect 53561 15997 53573 16031
rect 53607 15997 53619 16031
rect 53561 15991 53619 15997
rect 46566 15920 46572 15972
rect 46624 15960 46630 15972
rect 46753 15963 46811 15969
rect 46753 15960 46765 15963
rect 46624 15932 46765 15960
rect 46624 15920 46630 15932
rect 46753 15929 46765 15932
rect 46799 15960 46811 15963
rect 47394 15960 47400 15972
rect 46799 15932 47400 15960
rect 46799 15929 46811 15932
rect 46753 15923 46811 15929
rect 47394 15920 47400 15932
rect 47452 15920 47458 15972
rect 49786 15920 49792 15972
rect 49844 15960 49850 15972
rect 50706 15960 50712 15972
rect 49844 15932 50712 15960
rect 49844 15920 49850 15932
rect 50706 15920 50712 15932
rect 50764 15960 50770 15972
rect 51920 15960 51948 15988
rect 53576 15960 53604 15991
rect 55674 15988 55680 16040
rect 55732 15988 55738 16040
rect 57882 15988 57888 16040
rect 57940 15988 57946 16040
rect 50764 15932 51856 15960
rect 51920 15932 53604 15960
rect 50764 15920 50770 15932
rect 40313 15895 40371 15901
rect 40313 15861 40325 15895
rect 40359 15892 40371 15895
rect 43346 15892 43352 15904
rect 40359 15864 43352 15892
rect 40359 15861 40371 15864
rect 40313 15855 40371 15861
rect 43346 15852 43352 15864
rect 43404 15852 43410 15904
rect 43438 15852 43444 15904
rect 43496 15852 43502 15904
rect 46382 15852 46388 15904
rect 46440 15892 46446 15904
rect 48869 15895 48927 15901
rect 48869 15892 48881 15895
rect 46440 15864 48881 15892
rect 46440 15852 46446 15864
rect 48869 15861 48881 15864
rect 48915 15892 48927 15895
rect 49050 15892 49056 15904
rect 48915 15864 49056 15892
rect 48915 15861 48927 15864
rect 48869 15855 48927 15861
rect 49050 15852 49056 15864
rect 49108 15852 49114 15904
rect 51828 15892 51856 15932
rect 52549 15895 52607 15901
rect 52549 15892 52561 15895
rect 51828 15864 52561 15892
rect 52549 15861 52561 15864
rect 52595 15892 52607 15895
rect 53466 15892 53472 15904
rect 52595 15864 53472 15892
rect 52595 15861 52607 15864
rect 52549 15855 52607 15861
rect 53466 15852 53472 15864
rect 53524 15852 53530 15904
rect 55214 15852 55220 15904
rect 55272 15852 55278 15904
rect 55858 15852 55864 15904
rect 55916 15892 55922 15904
rect 56229 15895 56287 15901
rect 56229 15892 56241 15895
rect 55916 15864 56241 15892
rect 55916 15852 55922 15864
rect 56229 15861 56241 15864
rect 56275 15861 56287 15895
rect 56229 15855 56287 15861
rect 57974 15852 57980 15904
rect 58032 15892 58038 15904
rect 58529 15895 58587 15901
rect 58529 15892 58541 15895
rect 58032 15864 58541 15892
rect 58032 15852 58038 15864
rect 58529 15861 58541 15864
rect 58575 15861 58587 15895
rect 58529 15855 58587 15861
rect 1104 15802 58880 15824
rect 1104 15750 8172 15802
rect 8224 15750 8236 15802
rect 8288 15750 8300 15802
rect 8352 15750 8364 15802
rect 8416 15750 8428 15802
rect 8480 15750 22616 15802
rect 22668 15750 22680 15802
rect 22732 15750 22744 15802
rect 22796 15750 22808 15802
rect 22860 15750 22872 15802
rect 22924 15750 37060 15802
rect 37112 15750 37124 15802
rect 37176 15750 37188 15802
rect 37240 15750 37252 15802
rect 37304 15750 37316 15802
rect 37368 15750 51504 15802
rect 51556 15750 51568 15802
rect 51620 15750 51632 15802
rect 51684 15750 51696 15802
rect 51748 15750 51760 15802
rect 51812 15750 58880 15802
rect 1104 15728 58880 15750
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 5537 15691 5595 15697
rect 5537 15688 5549 15691
rect 5500 15660 5549 15688
rect 5500 15648 5506 15660
rect 5537 15657 5549 15660
rect 5583 15657 5595 15691
rect 5537 15651 5595 15657
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 11149 15691 11207 15697
rect 11149 15688 11161 15691
rect 9732 15660 11161 15688
rect 9732 15648 9738 15660
rect 11149 15657 11161 15660
rect 11195 15657 11207 15691
rect 11149 15651 11207 15657
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 6089 15555 6147 15561
rect 6089 15552 6101 15555
rect 5868 15524 6101 15552
rect 5868 15512 5874 15524
rect 6089 15521 6101 15524
rect 6135 15552 6147 15555
rect 6546 15552 6552 15564
rect 6135 15524 6552 15552
rect 6135 15521 6147 15524
rect 6089 15515 6147 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 7926 15512 7932 15564
rect 7984 15512 7990 15564
rect 9582 15552 9588 15564
rect 8588 15524 9588 15552
rect 8588 15496 8616 15524
rect 9582 15512 9588 15524
rect 9640 15552 9646 15564
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 9640 15524 9781 15552
rect 9640 15512 9646 15524
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 11164 15552 11192 15651
rect 13538 15648 13544 15700
rect 13596 15648 13602 15700
rect 13630 15648 13636 15700
rect 13688 15648 13694 15700
rect 13998 15648 14004 15700
rect 14056 15688 14062 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 14056 15660 14381 15688
rect 14056 15648 14062 15660
rect 14369 15657 14381 15660
rect 14415 15688 14427 15691
rect 14918 15688 14924 15700
rect 14415 15660 14924 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 15746 15648 15752 15700
rect 15804 15648 15810 15700
rect 18414 15648 18420 15700
rect 18472 15648 18478 15700
rect 18506 15648 18512 15700
rect 18564 15648 18570 15700
rect 19518 15648 19524 15700
rect 19576 15648 19582 15700
rect 21358 15648 21364 15700
rect 21416 15648 21422 15700
rect 21634 15648 21640 15700
rect 21692 15648 21698 15700
rect 27430 15648 27436 15700
rect 27488 15688 27494 15700
rect 27488 15660 28028 15688
rect 27488 15648 27494 15660
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 11164 15524 11989 15552
rect 9769 15515 9827 15521
rect 11977 15521 11989 15524
rect 12023 15521 12035 15555
rect 11977 15515 12035 15521
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13556 15552 13584 15648
rect 13127 15524 13584 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 14090 15512 14096 15564
rect 14148 15552 14154 15564
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 14148 15524 14749 15552
rect 14148 15512 14154 15524
rect 14737 15521 14749 15524
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 6454 15444 6460 15496
rect 6512 15444 6518 15496
rect 8018 15444 8024 15496
rect 8076 15484 8082 15496
rect 8113 15487 8171 15493
rect 8113 15484 8125 15487
rect 8076 15456 8125 15484
rect 8076 15444 8082 15456
rect 8113 15453 8125 15456
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 8938 15444 8944 15496
rect 8996 15444 9002 15496
rect 11238 15444 11244 15496
rect 11296 15444 11302 15496
rect 15004 15487 15062 15493
rect 15004 15453 15016 15487
rect 15050 15484 15062 15487
rect 15764 15484 15792 15648
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15552 18015 15555
rect 18432 15552 18460 15648
rect 19889 15623 19947 15629
rect 19889 15589 19901 15623
rect 19935 15620 19947 15623
rect 19935 15592 20760 15620
rect 19935 15589 19947 15592
rect 19889 15583 19947 15589
rect 18003 15524 18460 15552
rect 20533 15555 20591 15561
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 20622 15552 20628 15564
rect 20579 15524 20628 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 20622 15512 20628 15524
rect 20680 15512 20686 15564
rect 20732 15561 20760 15592
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15050 15456 15792 15484
rect 16132 15456 16221 15484
rect 15050 15453 15062 15456
rect 15004 15447 15062 15453
rect 7653 15419 7711 15425
rect 7653 15416 7665 15419
rect 5920 15388 7665 15416
rect 5810 15308 5816 15360
rect 5868 15348 5874 15360
rect 5920 15357 5948 15388
rect 7653 15385 7665 15388
rect 7699 15416 7711 15419
rect 9398 15416 9404 15428
rect 7699 15388 9404 15416
rect 7699 15385 7711 15388
rect 7653 15379 7711 15385
rect 9398 15376 9404 15388
rect 9456 15376 9462 15428
rect 10036 15419 10094 15425
rect 10036 15385 10048 15419
rect 10082 15416 10094 15419
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 10082 15388 11897 15416
rect 10082 15385 10094 15388
rect 10036 15379 10094 15385
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 11885 15379 11943 15385
rect 15194 15376 15200 15428
rect 15252 15376 15258 15428
rect 5905 15351 5963 15357
rect 5905 15348 5917 15351
rect 5868 15320 5917 15348
rect 5868 15308 5874 15320
rect 5905 15317 5917 15320
rect 5951 15317 5963 15351
rect 5905 15311 5963 15317
rect 5997 15351 6055 15357
rect 5997 15317 6009 15351
rect 6043 15348 6055 15351
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6043 15320 7021 15348
rect 6043 15317 6055 15320
rect 5997 15311 6055 15317
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 7282 15308 7288 15360
rect 7340 15308 7346 15360
rect 7745 15351 7803 15357
rect 7745 15317 7757 15351
rect 7791 15348 7803 15351
rect 8757 15351 8815 15357
rect 8757 15348 8769 15351
rect 7791 15320 8769 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 8757 15317 8769 15320
rect 8803 15317 8815 15351
rect 8757 15311 8815 15317
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 12618 15308 12624 15360
rect 12676 15308 12682 15360
rect 15212 15348 15240 15376
rect 16132 15357 16160 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 21652 15484 21680 15648
rect 28000 15620 28028 15660
rect 28074 15648 28080 15700
rect 28132 15648 28138 15700
rect 32674 15648 32680 15700
rect 32732 15648 32738 15700
rect 33134 15648 33140 15700
rect 33192 15688 33198 15700
rect 33597 15691 33655 15697
rect 33597 15688 33609 15691
rect 33192 15660 33609 15688
rect 33192 15648 33198 15660
rect 33597 15657 33609 15660
rect 33643 15657 33655 15691
rect 33597 15651 33655 15657
rect 34422 15648 34428 15700
rect 34480 15648 34486 15700
rect 34698 15648 34704 15700
rect 34756 15688 34762 15700
rect 34885 15691 34943 15697
rect 34885 15688 34897 15691
rect 34756 15660 34897 15688
rect 34756 15648 34762 15660
rect 34885 15657 34897 15660
rect 34931 15657 34943 15691
rect 34885 15651 34943 15657
rect 38102 15648 38108 15700
rect 38160 15648 38166 15700
rect 38194 15648 38200 15700
rect 38252 15648 38258 15700
rect 38470 15648 38476 15700
rect 38528 15688 38534 15700
rect 38933 15691 38991 15697
rect 38933 15688 38945 15691
rect 38528 15660 38945 15688
rect 38528 15648 38534 15660
rect 38933 15657 38945 15660
rect 38979 15657 38991 15691
rect 38933 15651 38991 15657
rect 39022 15648 39028 15700
rect 39080 15648 39086 15700
rect 39390 15648 39396 15700
rect 39448 15688 39454 15700
rect 39669 15691 39727 15697
rect 39669 15688 39681 15691
rect 39448 15660 39681 15688
rect 39448 15648 39454 15660
rect 39669 15657 39681 15660
rect 39715 15657 39727 15691
rect 39669 15651 39727 15657
rect 40310 15648 40316 15700
rect 40368 15648 40374 15700
rect 41414 15648 41420 15700
rect 41472 15648 41478 15700
rect 41509 15691 41567 15697
rect 41509 15657 41521 15691
rect 41555 15688 41567 15691
rect 42426 15688 42432 15700
rect 41555 15660 42432 15688
rect 41555 15657 41567 15660
rect 41509 15651 41567 15657
rect 42426 15648 42432 15660
rect 42484 15648 42490 15700
rect 43901 15691 43959 15697
rect 43901 15657 43913 15691
rect 43947 15688 43959 15691
rect 45002 15688 45008 15700
rect 43947 15660 45008 15688
rect 43947 15657 43959 15660
rect 43901 15651 43959 15657
rect 45002 15648 45008 15660
rect 45060 15648 45066 15700
rect 45922 15648 45928 15700
rect 45980 15688 45986 15700
rect 46293 15691 46351 15697
rect 46293 15688 46305 15691
rect 45980 15660 46305 15688
rect 45980 15648 45986 15660
rect 46293 15657 46305 15660
rect 46339 15657 46351 15691
rect 46293 15651 46351 15657
rect 29638 15620 29644 15632
rect 28000 15592 29644 15620
rect 29638 15580 29644 15592
rect 29696 15580 29702 15632
rect 26234 15512 26240 15564
rect 26292 15552 26298 15564
rect 26694 15552 26700 15564
rect 26292 15524 26700 15552
rect 26292 15512 26298 15524
rect 26694 15512 26700 15524
rect 26752 15512 26758 15564
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28629 15555 28687 15561
rect 28629 15552 28641 15555
rect 28040 15524 28641 15552
rect 28040 15512 28046 15524
rect 28629 15521 28641 15524
rect 28675 15521 28687 15555
rect 28629 15515 28687 15521
rect 28813 15555 28871 15561
rect 28813 15521 28825 15555
rect 28859 15552 28871 15555
rect 29733 15555 29791 15561
rect 29733 15552 29745 15555
rect 28859 15524 29745 15552
rect 28859 15521 28871 15524
rect 28813 15515 28871 15521
rect 29733 15521 29745 15524
rect 29779 15521 29791 15555
rect 29733 15515 29791 15521
rect 30208 15524 31616 15552
rect 20395 15456 21680 15484
rect 22833 15487 22891 15493
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 22833 15453 22845 15487
rect 22879 15484 22891 15487
rect 23198 15484 23204 15496
rect 22879 15456 23204 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 23198 15444 23204 15456
rect 23256 15444 23262 15496
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15484 25559 15487
rect 25682 15484 25688 15496
rect 25547 15456 25688 15484
rect 25547 15453 25559 15456
rect 25501 15447 25559 15453
rect 25682 15444 25688 15456
rect 25740 15444 25746 15496
rect 27246 15444 27252 15496
rect 27304 15484 27310 15496
rect 27304 15456 28396 15484
rect 27304 15444 27310 15456
rect 26964 15419 27022 15425
rect 26964 15385 26976 15419
rect 27010 15416 27022 15419
rect 28258 15416 28264 15428
rect 27010 15388 28264 15416
rect 27010 15385 27022 15388
rect 26964 15379 27022 15385
rect 28258 15376 28264 15388
rect 28316 15376 28322 15428
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15212 15320 16129 15348
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 16117 15311 16175 15317
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 18877 15351 18935 15357
rect 18877 15348 18889 15351
rect 18564 15320 18889 15348
rect 18564 15308 18570 15320
rect 18877 15317 18889 15320
rect 18923 15348 18935 15351
rect 19886 15348 19892 15360
rect 18923 15320 19892 15348
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 23382 15308 23388 15360
rect 23440 15308 23446 15360
rect 26053 15351 26111 15357
rect 26053 15317 26065 15351
rect 26099 15348 26111 15351
rect 26510 15348 26516 15360
rect 26099 15320 26516 15348
rect 26099 15317 26111 15320
rect 26053 15311 26111 15317
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 28166 15308 28172 15360
rect 28224 15308 28230 15360
rect 28368 15348 28396 15456
rect 28442 15444 28448 15496
rect 28500 15484 28506 15496
rect 28828 15484 28856 15515
rect 30208 15496 30236 15524
rect 30190 15484 30196 15496
rect 28500 15456 28856 15484
rect 29104 15456 30196 15484
rect 28500 15444 28506 15456
rect 28537 15419 28595 15425
rect 28537 15385 28549 15419
rect 28583 15416 28595 15419
rect 28994 15416 29000 15428
rect 28583 15388 29000 15416
rect 28583 15385 28595 15388
rect 28537 15379 28595 15385
rect 28994 15376 29000 15388
rect 29052 15376 29058 15428
rect 29104 15348 29132 15456
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 31481 15487 31539 15493
rect 31481 15484 31493 15487
rect 31312 15456 31493 15484
rect 28368 15320 29132 15348
rect 29270 15308 29276 15360
rect 29328 15308 29334 15360
rect 31018 15308 31024 15360
rect 31076 15348 31082 15360
rect 31312 15357 31340 15456
rect 31481 15453 31493 15456
rect 31527 15453 31539 15487
rect 31481 15447 31539 15453
rect 31588 15416 31616 15524
rect 31748 15487 31806 15493
rect 31748 15453 31760 15487
rect 31794 15484 31806 15487
rect 32692 15484 32720 15648
rect 32861 15623 32919 15629
rect 32861 15589 32873 15623
rect 32907 15620 32919 15623
rect 32907 15592 33088 15620
rect 32907 15589 32919 15592
rect 32861 15583 32919 15589
rect 33060 15561 33088 15592
rect 33045 15555 33103 15561
rect 33045 15521 33057 15555
rect 33091 15552 33103 15555
rect 34440 15552 34468 15648
rect 33091 15524 34468 15552
rect 33091 15521 33103 15524
rect 33045 15515 33103 15521
rect 35434 15512 35440 15564
rect 35492 15552 35498 15564
rect 36722 15552 36728 15564
rect 35492 15524 36728 15552
rect 35492 15512 35498 15524
rect 36722 15512 36728 15524
rect 36780 15512 36786 15564
rect 37645 15555 37703 15561
rect 37645 15521 37657 15555
rect 37691 15552 37703 15555
rect 38120 15552 38148 15648
rect 37691 15524 38148 15552
rect 38381 15555 38439 15561
rect 37691 15521 37703 15524
rect 37645 15515 37703 15521
rect 38381 15521 38393 15555
rect 38427 15552 38439 15555
rect 39040 15552 39068 15648
rect 38427 15524 39068 15552
rect 38427 15521 38439 15524
rect 38381 15515 38439 15521
rect 31794 15456 32720 15484
rect 31794 15453 31806 15456
rect 31748 15447 31806 15453
rect 33318 15444 33324 15496
rect 33376 15484 33382 15496
rect 37826 15484 37832 15496
rect 33376 15456 37832 15484
rect 33376 15444 33382 15456
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 38654 15444 38660 15496
rect 38712 15484 38718 15496
rect 39025 15487 39083 15493
rect 39025 15484 39037 15487
rect 38712 15456 39037 15484
rect 38712 15444 38718 15456
rect 39025 15453 39037 15456
rect 39071 15453 39083 15487
rect 39025 15447 39083 15453
rect 40328 15416 40356 15648
rect 41432 15552 41460 15648
rect 46308 15620 46336 15651
rect 47486 15648 47492 15700
rect 47544 15688 47550 15700
rect 47854 15688 47860 15700
rect 47544 15660 47860 15688
rect 47544 15648 47550 15660
rect 47854 15648 47860 15660
rect 47912 15688 47918 15700
rect 48593 15691 48651 15697
rect 48593 15688 48605 15691
rect 47912 15660 48605 15688
rect 47912 15648 47918 15660
rect 48593 15657 48605 15660
rect 48639 15657 48651 15691
rect 48593 15651 48651 15657
rect 47026 15620 47032 15632
rect 46308 15592 47032 15620
rect 47026 15580 47032 15592
rect 47084 15580 47090 15632
rect 48317 15623 48375 15629
rect 48317 15589 48329 15623
rect 48363 15620 48375 15623
rect 48406 15620 48412 15632
rect 48363 15592 48412 15620
rect 48363 15589 48375 15592
rect 48317 15583 48375 15589
rect 48406 15580 48412 15592
rect 48464 15580 48470 15632
rect 48608 15620 48636 15651
rect 49694 15648 49700 15700
rect 49752 15688 49758 15700
rect 50433 15691 50491 15697
rect 50433 15688 50445 15691
rect 49752 15660 50445 15688
rect 49752 15648 49758 15660
rect 50433 15657 50445 15660
rect 50479 15688 50491 15691
rect 53098 15688 53104 15700
rect 50479 15660 51304 15688
rect 50479 15657 50491 15660
rect 50433 15651 50491 15657
rect 51166 15620 51172 15632
rect 48608 15592 51172 15620
rect 51166 15580 51172 15592
rect 51224 15580 51230 15632
rect 42061 15555 42119 15561
rect 42061 15552 42073 15555
rect 41432 15524 42073 15552
rect 42061 15521 42073 15524
rect 42107 15521 42119 15555
rect 42061 15515 42119 15521
rect 42429 15555 42487 15561
rect 42429 15521 42441 15555
rect 42475 15552 42487 15555
rect 42794 15552 42800 15564
rect 42475 15524 42800 15552
rect 42475 15521 42487 15524
rect 42429 15515 42487 15521
rect 42794 15512 42800 15524
rect 42852 15512 42858 15564
rect 43809 15555 43867 15561
rect 43809 15521 43821 15555
rect 43855 15552 43867 15555
rect 44545 15555 44603 15561
rect 44545 15552 44557 15555
rect 43855 15524 44557 15552
rect 43855 15521 43867 15524
rect 43809 15515 43867 15521
rect 44545 15521 44557 15524
rect 44591 15521 44603 15555
rect 44545 15515 44603 15521
rect 41138 15444 41144 15496
rect 41196 15484 41202 15496
rect 43824 15484 43852 15515
rect 41196 15456 43852 15484
rect 44560 15484 44588 15515
rect 44910 15512 44916 15564
rect 44968 15552 44974 15564
rect 45005 15555 45063 15561
rect 45005 15552 45017 15555
rect 44968 15524 45017 15552
rect 44968 15512 44974 15524
rect 45005 15521 45017 15524
rect 45051 15521 45063 15555
rect 45005 15515 45063 15521
rect 49786 15512 49792 15564
rect 49844 15512 49850 15564
rect 49804 15484 49832 15512
rect 44560 15456 49832 15484
rect 41196 15444 41202 15456
rect 50706 15444 50712 15496
rect 50764 15444 50770 15496
rect 51276 15484 51304 15660
rect 51368 15660 53104 15688
rect 51368 15561 51396 15660
rect 53098 15648 53104 15660
rect 53156 15648 53162 15700
rect 56134 15648 56140 15700
rect 56192 15688 56198 15700
rect 56321 15691 56379 15697
rect 56321 15688 56333 15691
rect 56192 15660 56333 15688
rect 56192 15648 56198 15660
rect 56321 15657 56333 15660
rect 56367 15657 56379 15691
rect 56321 15651 56379 15657
rect 51997 15623 52055 15629
rect 51997 15620 52009 15623
rect 51460 15592 52009 15620
rect 51460 15564 51488 15592
rect 51997 15589 52009 15592
rect 52043 15589 52055 15623
rect 51997 15583 52055 15589
rect 55309 15623 55367 15629
rect 55309 15589 55321 15623
rect 55355 15589 55367 15623
rect 55309 15583 55367 15589
rect 51353 15555 51411 15561
rect 51353 15521 51365 15555
rect 51399 15521 51411 15555
rect 51353 15515 51411 15521
rect 51442 15512 51448 15564
rect 51500 15512 51506 15564
rect 51537 15555 51595 15561
rect 51537 15521 51549 15555
rect 51583 15552 51595 15555
rect 51902 15552 51908 15564
rect 51583 15524 51908 15552
rect 51583 15521 51595 15524
rect 51537 15515 51595 15521
rect 51902 15512 51908 15524
rect 51960 15512 51966 15564
rect 52546 15512 52552 15564
rect 52604 15512 52610 15564
rect 53098 15512 53104 15564
rect 53156 15552 53162 15564
rect 53837 15555 53895 15561
rect 53837 15552 53849 15555
rect 53156 15524 53849 15552
rect 53156 15512 53162 15524
rect 53837 15521 53849 15524
rect 53883 15521 53895 15555
rect 53837 15515 53895 15521
rect 54573 15555 54631 15561
rect 54573 15521 54585 15555
rect 54619 15552 54631 15555
rect 55324 15552 55352 15583
rect 54619 15524 55352 15552
rect 55861 15555 55919 15561
rect 54619 15521 54631 15524
rect 54573 15515 54631 15521
rect 55861 15521 55873 15555
rect 55907 15521 55919 15555
rect 55861 15515 55919 15521
rect 51276 15456 51396 15484
rect 31588 15388 40356 15416
rect 31297 15351 31355 15357
rect 31297 15348 31309 15351
rect 31076 15320 31309 15348
rect 31076 15308 31082 15320
rect 31297 15317 31309 15320
rect 31343 15317 31355 15351
rect 31297 15311 31355 15317
rect 33965 15351 34023 15357
rect 33965 15317 33977 15351
rect 34011 15348 34023 15351
rect 34054 15348 34060 15360
rect 34011 15320 34060 15348
rect 34011 15317 34023 15320
rect 33965 15311 34023 15317
rect 34054 15308 34060 15320
rect 34112 15348 34118 15360
rect 35066 15348 35072 15360
rect 34112 15320 35072 15348
rect 34112 15308 34118 15320
rect 35066 15308 35072 15320
rect 35124 15348 35130 15360
rect 35250 15348 35256 15360
rect 35124 15320 35256 15348
rect 35124 15308 35130 15320
rect 35250 15308 35256 15320
rect 35308 15308 35314 15360
rect 35345 15351 35403 15357
rect 35345 15317 35357 15351
rect 35391 15348 35403 15351
rect 36354 15348 36360 15360
rect 35391 15320 36360 15348
rect 35391 15317 35403 15320
rect 35345 15311 35403 15317
rect 36354 15308 36360 15320
rect 36412 15308 36418 15360
rect 40129 15351 40187 15357
rect 40129 15317 40141 15351
rect 40175 15348 40187 15351
rect 40402 15348 40408 15360
rect 40175 15320 40408 15348
rect 40175 15317 40187 15320
rect 40129 15311 40187 15317
rect 40402 15308 40408 15320
rect 40460 15348 40466 15360
rect 41156 15348 41184 15444
rect 51368 15428 51396 15456
rect 52270 15444 52276 15496
rect 52328 15444 52334 15496
rect 52362 15444 52368 15496
rect 52420 15493 52426 15496
rect 52420 15487 52448 15493
rect 52436 15453 52448 15487
rect 52420 15447 52448 15453
rect 52420 15444 52426 15447
rect 53282 15444 53288 15496
rect 53340 15484 53346 15496
rect 53653 15487 53711 15493
rect 53653 15484 53665 15487
rect 53340 15456 53665 15484
rect 53340 15444 53346 15456
rect 53653 15453 53665 15456
rect 53699 15453 53711 15487
rect 53653 15447 53711 15453
rect 55214 15444 55220 15496
rect 55272 15484 55278 15496
rect 55876 15484 55904 15515
rect 56042 15512 56048 15564
rect 56100 15552 56106 15564
rect 56781 15555 56839 15561
rect 56781 15552 56793 15555
rect 56100 15524 56793 15552
rect 56100 15512 56106 15524
rect 56781 15521 56793 15524
rect 56827 15521 56839 15555
rect 56781 15515 56839 15521
rect 55272 15456 55904 15484
rect 55272 15444 55278 15456
rect 41877 15419 41935 15425
rect 41877 15385 41889 15419
rect 41923 15416 41935 15419
rect 42058 15416 42064 15428
rect 41923 15388 42064 15416
rect 41923 15385 41935 15388
rect 41877 15379 41935 15385
rect 42058 15376 42064 15388
rect 42116 15416 42122 15428
rect 44269 15419 44327 15425
rect 42116 15388 44036 15416
rect 42116 15376 42122 15388
rect 44008 15360 44036 15388
rect 44269 15385 44281 15419
rect 44315 15416 44327 15419
rect 45649 15419 45707 15425
rect 45649 15416 45661 15419
rect 44315 15388 45661 15416
rect 44315 15385 44327 15388
rect 44269 15379 44327 15385
rect 45649 15385 45661 15388
rect 45695 15385 45707 15419
rect 45649 15379 45707 15385
rect 51350 15376 51356 15428
rect 51408 15376 51414 15428
rect 53193 15419 53251 15425
rect 53193 15385 53205 15419
rect 53239 15416 53251 15419
rect 53745 15419 53803 15425
rect 53745 15416 53757 15419
rect 53239 15388 53757 15416
rect 53239 15385 53251 15388
rect 53193 15379 53251 15385
rect 53745 15385 53757 15388
rect 53791 15385 53803 15419
rect 53745 15379 53803 15385
rect 57048 15419 57106 15425
rect 57048 15385 57060 15419
rect 57094 15416 57106 15419
rect 58526 15416 58532 15428
rect 57094 15388 58532 15416
rect 57094 15385 57106 15388
rect 57048 15379 57106 15385
rect 58526 15376 58532 15388
rect 58584 15376 58590 15428
rect 40460 15320 41184 15348
rect 41969 15351 42027 15357
rect 40460 15308 40466 15320
rect 41969 15317 41981 15351
rect 42015 15348 42027 15351
rect 42981 15351 43039 15357
rect 42981 15348 42993 15351
rect 42015 15320 42993 15348
rect 42015 15317 42027 15320
rect 41969 15311 42027 15317
rect 42981 15317 42993 15320
rect 43027 15317 43039 15351
rect 42981 15311 43039 15317
rect 43990 15308 43996 15360
rect 44048 15348 44054 15360
rect 44361 15351 44419 15357
rect 44361 15348 44373 15351
rect 44048 15320 44373 15348
rect 44048 15308 44054 15320
rect 44361 15317 44373 15320
rect 44407 15317 44419 15351
rect 44361 15311 44419 15317
rect 47394 15308 47400 15360
rect 47452 15308 47458 15360
rect 51258 15308 51264 15360
rect 51316 15308 51322 15360
rect 52638 15308 52644 15360
rect 52696 15348 52702 15360
rect 53285 15351 53343 15357
rect 53285 15348 53297 15351
rect 52696 15320 53297 15348
rect 52696 15308 52702 15320
rect 53285 15317 53297 15320
rect 53331 15317 53343 15351
rect 53285 15311 53343 15317
rect 54570 15308 54576 15360
rect 54628 15348 54634 15360
rect 55125 15351 55183 15357
rect 55125 15348 55137 15351
rect 54628 15320 55137 15348
rect 54628 15308 54634 15320
rect 55125 15317 55137 15320
rect 55171 15317 55183 15351
rect 55125 15311 55183 15317
rect 55582 15308 55588 15360
rect 55640 15348 55646 15360
rect 55677 15351 55735 15357
rect 55677 15348 55689 15351
rect 55640 15320 55689 15348
rect 55640 15308 55646 15320
rect 55677 15317 55689 15320
rect 55723 15317 55735 15351
rect 55677 15311 55735 15317
rect 55766 15308 55772 15360
rect 55824 15308 55830 15360
rect 57330 15308 57336 15360
rect 57388 15348 57394 15360
rect 57882 15348 57888 15360
rect 57388 15320 57888 15348
rect 57388 15308 57394 15320
rect 57882 15308 57888 15320
rect 57940 15348 57946 15360
rect 58161 15351 58219 15357
rect 58161 15348 58173 15351
rect 57940 15320 58173 15348
rect 57940 15308 57946 15320
rect 58161 15317 58173 15320
rect 58207 15317 58219 15351
rect 58161 15311 58219 15317
rect 1104 15258 59040 15280
rect 1104 15206 15394 15258
rect 15446 15206 15458 15258
rect 15510 15206 15522 15258
rect 15574 15206 15586 15258
rect 15638 15206 15650 15258
rect 15702 15206 29838 15258
rect 29890 15206 29902 15258
rect 29954 15206 29966 15258
rect 30018 15206 30030 15258
rect 30082 15206 30094 15258
rect 30146 15206 44282 15258
rect 44334 15206 44346 15258
rect 44398 15206 44410 15258
rect 44462 15206 44474 15258
rect 44526 15206 44538 15258
rect 44590 15206 58726 15258
rect 58778 15206 58790 15258
rect 58842 15206 58854 15258
rect 58906 15206 58918 15258
rect 58970 15206 58982 15258
rect 59034 15206 59040 15258
rect 1104 15184 59040 15206
rect 5534 15104 5540 15156
rect 5592 15104 5598 15156
rect 6181 15147 6239 15153
rect 6181 15113 6193 15147
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 5552 15076 5580 15104
rect 4816 15048 5580 15076
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 4816 15017 4844 15048
rect 5994 15036 6000 15088
rect 6052 15036 6058 15088
rect 6196 15076 6224 15107
rect 6546 15104 6552 15156
rect 6604 15104 6610 15156
rect 9858 15144 9864 15156
rect 6932 15116 9864 15144
rect 6454 15076 6460 15088
rect 6196 15048 6460 15076
rect 6454 15036 6460 15048
rect 6512 15076 6518 15088
rect 6512 15048 6868 15076
rect 6512 15036 6518 15048
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4764 14980 4813 15008
rect 4764 14968 4770 14980
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 5068 15011 5126 15017
rect 5068 14977 5080 15011
rect 5114 15008 5126 15011
rect 6012 15008 6040 15036
rect 5114 14980 6040 15008
rect 5114 14977 5126 14980
rect 5068 14971 5126 14977
rect 6733 14943 6791 14949
rect 6733 14909 6745 14943
rect 6779 14909 6791 14943
rect 6840 14940 6868 15048
rect 6932 15017 6960 15116
rect 9858 15104 9864 15116
rect 9916 15144 9922 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9916 15116 10057 15144
rect 9916 15104 9922 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 10045 15107 10103 15113
rect 10229 15147 10287 15153
rect 10229 15113 10241 15147
rect 10275 15113 10287 15147
rect 10229 15107 10287 15113
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 12618 15144 12624 15156
rect 10735 15116 12624 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 8932 15079 8990 15085
rect 8932 15045 8944 15079
rect 8978 15076 8990 15079
rect 9582 15076 9588 15088
rect 8978 15048 9588 15076
rect 8978 15045 8990 15048
rect 8932 15039 8990 15045
rect 9582 15036 9588 15048
rect 9640 15036 9646 15088
rect 10244 15076 10272 15107
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12768 15116 13461 15144
rect 12768 15104 12774 15116
rect 13449 15113 13461 15116
rect 13495 15144 13507 15147
rect 14182 15144 14188 15156
rect 13495 15116 14188 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 15102 15104 15108 15156
rect 15160 15104 15166 15156
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 16850 15144 16856 15156
rect 15519 15116 16856 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18690 15144 18696 15156
rect 18371 15116 18696 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 18690 15104 18696 15116
rect 18748 15144 18754 15156
rect 19150 15144 19156 15156
rect 18748 15116 19156 15144
rect 18748 15104 18754 15116
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 20349 15147 20407 15153
rect 20349 15144 20361 15147
rect 19576 15116 20361 15144
rect 19576 15104 19582 15116
rect 20349 15113 20361 15116
rect 20395 15144 20407 15147
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20395 15116 21189 15144
rect 20395 15113 20407 15116
rect 20349 15107 20407 15113
rect 21177 15113 21189 15116
rect 21223 15144 21235 15147
rect 21545 15147 21603 15153
rect 21545 15144 21557 15147
rect 21223 15116 21557 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21545 15113 21557 15116
rect 21591 15113 21603 15147
rect 21545 15107 21603 15113
rect 11238 15076 11244 15088
rect 10244 15048 11244 15076
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 14977 6975 15011
rect 8754 15008 8760 15020
rect 6917 14971 6975 14977
rect 8496 14980 8760 15008
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 6840 14912 7665 14940
rect 6733 14903 6791 14909
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 6748 14804 6776 14903
rect 7742 14900 7748 14952
rect 7800 14949 7806 14952
rect 7800 14943 7828 14949
rect 7816 14909 7828 14943
rect 7800 14903 7828 14909
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8496 14940 8524 14980
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 10870 15008 10876 15020
rect 10643 14980 10876 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 10870 14968 10876 14980
rect 10928 15008 10934 15020
rect 11054 15008 11060 15020
rect 10928 14980 11060 15008
rect 10928 14968 10934 14980
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 15008 15623 15011
rect 21560 15008 21588 15107
rect 26694 15104 26700 15156
rect 26752 15104 26758 15156
rect 28258 15104 28264 15156
rect 28316 15104 28322 15156
rect 28994 15104 29000 15156
rect 29052 15104 29058 15156
rect 33137 15147 33195 15153
rect 33137 15113 33149 15147
rect 33183 15144 33195 15147
rect 33502 15144 33508 15156
rect 33183 15116 33508 15144
rect 33183 15113 33195 15116
rect 33137 15107 33195 15113
rect 33502 15104 33508 15116
rect 33560 15104 33566 15156
rect 39574 15104 39580 15156
rect 39632 15144 39638 15156
rect 40405 15147 40463 15153
rect 40405 15144 40417 15147
rect 39632 15116 40417 15144
rect 39632 15104 39638 15116
rect 40405 15113 40417 15116
rect 40451 15144 40463 15147
rect 41598 15144 41604 15156
rect 40451 15116 41604 15144
rect 40451 15113 40463 15116
rect 40405 15107 40463 15113
rect 41598 15104 41604 15116
rect 41656 15104 41662 15156
rect 42705 15147 42763 15153
rect 42705 15113 42717 15147
rect 42751 15144 42763 15147
rect 43346 15144 43352 15156
rect 42751 15116 43352 15144
rect 42751 15113 42763 15116
rect 42705 15107 42763 15113
rect 22272 15079 22330 15085
rect 22272 15045 22284 15079
rect 22318 15076 22330 15079
rect 23382 15076 23388 15088
rect 22318 15048 23388 15076
rect 22318 15045 22330 15048
rect 22272 15039 22330 15045
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 23658 15036 23664 15088
rect 23716 15076 23722 15088
rect 24213 15079 24271 15085
rect 24213 15076 24225 15079
rect 23716 15048 24225 15076
rect 23716 15036 23722 15048
rect 24213 15045 24225 15048
rect 24259 15045 24271 15079
rect 24213 15039 24271 15045
rect 38194 15036 38200 15088
rect 38252 15076 38258 15088
rect 38378 15076 38384 15088
rect 38252 15048 38384 15076
rect 38252 15036 38258 15048
rect 38378 15036 38384 15048
rect 38436 15076 38442 15088
rect 42720 15076 42748 15107
rect 43346 15104 43352 15116
rect 43404 15144 43410 15156
rect 45094 15144 45100 15156
rect 43404 15116 45100 15144
rect 43404 15104 43410 15116
rect 45094 15104 45100 15116
rect 45152 15104 45158 15156
rect 48961 15147 49019 15153
rect 48961 15144 48973 15147
rect 46492 15116 48973 15144
rect 46492 15088 46520 15116
rect 48961 15113 48973 15116
rect 49007 15113 49019 15147
rect 48961 15107 49019 15113
rect 38436 15048 42748 15076
rect 45465 15079 45523 15085
rect 38436 15036 38442 15048
rect 45465 15045 45477 15079
rect 45511 15076 45523 15079
rect 46290 15076 46296 15088
rect 45511 15048 46296 15076
rect 45511 15045 45523 15048
rect 45465 15039 45523 15045
rect 46290 15036 46296 15048
rect 46348 15036 46354 15088
rect 46474 15036 46480 15088
rect 46532 15036 46538 15088
rect 21726 15008 21732 15020
rect 15611 14980 15976 15008
rect 21560 14980 21732 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 15948 14952 15976 14980
rect 21726 14968 21732 14980
rect 21784 15008 21790 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21784 14980 22017 15008
rect 21784 14968 21790 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 24302 14968 24308 15020
rect 24360 14968 24366 15020
rect 24572 15011 24630 15017
rect 24572 14977 24584 15011
rect 24618 15008 24630 15011
rect 26421 15011 26479 15017
rect 26421 15008 26433 15011
rect 24618 14980 26433 15008
rect 24618 14977 24630 14980
rect 24572 14971 24630 14977
rect 26421 14977 26433 14980
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 27709 15011 27767 15017
rect 27709 14977 27721 15011
rect 27755 15008 27767 15011
rect 28166 15008 28172 15020
rect 27755 14980 28172 15008
rect 27755 14977 27767 14980
rect 27709 14971 27767 14977
rect 28166 14968 28172 14980
rect 28224 14968 28230 15020
rect 45557 15011 45615 15017
rect 45557 14977 45569 15011
rect 45603 15008 45615 15011
rect 47305 15011 47363 15017
rect 47305 15008 47317 15011
rect 45603 14980 47317 15008
rect 45603 14977 45615 14980
rect 45557 14971 45615 14977
rect 47305 14977 47317 14980
rect 47351 14977 47363 15011
rect 47305 14971 47363 14977
rect 47848 15011 47906 15017
rect 47848 14977 47860 15011
rect 47894 15008 47906 15011
rect 47894 14980 48912 15008
rect 47894 14977 47906 14980
rect 47848 14971 47906 14977
rect 7975 14912 8524 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 7800 14900 7806 14903
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8628 14912 8677 14940
rect 8628 14900 8634 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 9950 14900 9956 14952
rect 10008 14940 10014 14952
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10008 14912 10793 14940
rect 10008 14900 10014 14912
rect 10781 14909 10793 14912
rect 10827 14940 10839 14943
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 10827 14912 11253 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 11241 14909 11253 14912
rect 11287 14940 11299 14943
rect 14734 14940 14740 14952
rect 11287 14912 14740 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15657 14903 15715 14909
rect 7377 14875 7435 14881
rect 7377 14841 7389 14875
rect 7423 14872 7435 14875
rect 7466 14872 7472 14884
rect 7423 14844 7472 14872
rect 7423 14841 7435 14844
rect 7377 14835 7435 14841
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 15672 14872 15700 14903
rect 15930 14900 15936 14952
rect 15988 14900 15994 14952
rect 19150 14900 19156 14952
rect 19208 14900 19214 14952
rect 23661 14943 23719 14949
rect 23661 14909 23673 14943
rect 23707 14940 23719 14943
rect 23707 14912 23796 14940
rect 23707 14909 23719 14912
rect 23661 14903 23719 14909
rect 14936 14844 15700 14872
rect 8018 14804 8024 14816
rect 6748 14776 8024 14804
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 9306 14804 9312 14816
rect 8619 14776 9312 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 14936 14813 14964 14844
rect 23768 14816 23796 14912
rect 25866 14900 25872 14952
rect 25924 14900 25930 14952
rect 28074 14900 28080 14952
rect 28132 14940 28138 14952
rect 28353 14943 28411 14949
rect 28353 14940 28365 14943
rect 28132 14912 28365 14940
rect 28132 14900 28138 14912
rect 28353 14909 28365 14912
rect 28399 14909 28411 14943
rect 28353 14903 28411 14909
rect 36538 14900 36544 14952
rect 36596 14900 36602 14952
rect 43533 14943 43591 14949
rect 43533 14940 43545 14943
rect 42076 14912 43545 14940
rect 26786 14872 26792 14884
rect 25240 14844 26792 14872
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 13964 14776 14933 14804
rect 13964 14764 13970 14776
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 14921 14767 14979 14773
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18380 14776 18889 14804
rect 18380 14764 18386 14776
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 18877 14767 18935 14773
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 19705 14807 19763 14813
rect 19705 14804 19717 14807
rect 19024 14776 19717 14804
rect 19024 14764 19030 14776
rect 19705 14773 19717 14776
rect 19751 14773 19763 14807
rect 19705 14767 19763 14773
rect 20073 14807 20131 14813
rect 20073 14773 20085 14807
rect 20119 14804 20131 14807
rect 20622 14804 20628 14816
rect 20119 14776 20628 14804
rect 20119 14773 20131 14776
rect 20073 14767 20131 14773
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 23385 14807 23443 14813
rect 23385 14773 23397 14807
rect 23431 14804 23443 14807
rect 23750 14804 23756 14816
rect 23431 14776 23756 14804
rect 23431 14773 23443 14776
rect 23385 14767 23443 14773
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 25240 14804 25268 14844
rect 26786 14832 26792 14844
rect 26844 14832 26850 14884
rect 40129 14875 40187 14881
rect 40129 14841 40141 14875
rect 40175 14872 40187 14875
rect 41046 14872 41052 14884
rect 40175 14844 41052 14872
rect 40175 14841 40187 14844
rect 40129 14835 40187 14841
rect 41046 14832 41052 14844
rect 41104 14832 41110 14884
rect 42076 14816 42104 14912
rect 43533 14909 43545 14912
rect 43579 14909 43591 14943
rect 45649 14943 45707 14949
rect 45649 14940 45661 14943
rect 43533 14903 43591 14909
rect 44928 14912 45661 14940
rect 44928 14816 44956 14912
rect 45649 14909 45661 14912
rect 45695 14909 45707 14943
rect 45649 14903 45707 14909
rect 45925 14943 45983 14949
rect 45925 14909 45937 14943
rect 45971 14909 45983 14943
rect 45925 14903 45983 14909
rect 46753 14943 46811 14949
rect 46753 14909 46765 14943
rect 46799 14909 46811 14943
rect 46753 14903 46811 14909
rect 45097 14875 45155 14881
rect 45097 14841 45109 14875
rect 45143 14872 45155 14875
rect 45940 14872 45968 14903
rect 45143 14844 45968 14872
rect 45143 14841 45155 14844
rect 45097 14835 45155 14841
rect 46768 14816 46796 14903
rect 47394 14900 47400 14952
rect 47452 14940 47458 14952
rect 47581 14943 47639 14949
rect 47581 14940 47593 14943
rect 47452 14912 47593 14940
rect 47452 14900 47458 14912
rect 47581 14909 47593 14912
rect 47627 14909 47639 14943
rect 47581 14903 47639 14909
rect 48884 14872 48912 14980
rect 48976 14940 49004 15107
rect 50706 15104 50712 15156
rect 50764 15104 50770 15156
rect 52454 15104 52460 15156
rect 52512 15144 52518 15156
rect 53098 15144 53104 15156
rect 52512 15116 53104 15144
rect 52512 15104 52518 15116
rect 53098 15104 53104 15116
rect 53156 15104 53162 15156
rect 53837 15147 53895 15153
rect 53837 15113 53849 15147
rect 53883 15144 53895 15147
rect 55490 15144 55496 15156
rect 53883 15116 55496 15144
rect 53883 15113 53895 15116
rect 53837 15107 53895 15113
rect 55490 15104 55496 15116
rect 55548 15104 55554 15156
rect 57330 15144 57336 15156
rect 55876 15116 57336 15144
rect 51077 15011 51135 15017
rect 51077 14977 51089 15011
rect 51123 15008 51135 15011
rect 52181 15011 52239 15017
rect 52181 15008 52193 15011
rect 51123 14980 52193 15008
rect 51123 14977 51135 14980
rect 51077 14971 51135 14977
rect 52181 14977 52193 14980
rect 52227 14977 52239 15011
rect 52181 14971 52239 14977
rect 52362 14968 52368 15020
rect 52420 14968 52426 15020
rect 54196 15011 54254 15017
rect 54196 14977 54208 15011
rect 54242 15008 54254 15011
rect 55398 15008 55404 15020
rect 54242 14980 55404 15008
rect 54242 14977 54254 14980
rect 54196 14971 54254 14977
rect 55398 14968 55404 14980
rect 55456 14968 55462 15020
rect 55876 15017 55904 15116
rect 57330 15104 57336 15116
rect 57388 15104 57394 15156
rect 58526 15104 58532 15156
rect 58584 15104 58590 15156
rect 55861 15011 55919 15017
rect 55861 14977 55873 15011
rect 55907 14977 55919 15011
rect 55861 14971 55919 14977
rect 56870 14968 56876 15020
rect 56928 14968 56934 15020
rect 49053 14943 49111 14949
rect 49053 14940 49065 14943
rect 48976 14912 49065 14940
rect 49053 14909 49065 14912
rect 49099 14909 49111 14943
rect 49053 14903 49111 14909
rect 49234 14900 49240 14952
rect 49292 14940 49298 14952
rect 49789 14943 49847 14949
rect 49789 14940 49801 14943
rect 49292 14912 49801 14940
rect 49292 14900 49298 14912
rect 49789 14909 49801 14912
rect 49835 14909 49847 14943
rect 49789 14903 49847 14909
rect 51169 14943 51227 14949
rect 51169 14909 51181 14943
rect 51215 14909 51227 14943
rect 51169 14903 51227 14909
rect 50433 14875 50491 14881
rect 50433 14872 50445 14875
rect 48884 14844 50445 14872
rect 50433 14841 50445 14844
rect 50479 14841 50491 14875
rect 51184 14872 51212 14903
rect 51350 14900 51356 14952
rect 51408 14900 51414 14952
rect 51629 14943 51687 14949
rect 51629 14909 51641 14943
rect 51675 14940 51687 14943
rect 51902 14940 51908 14952
rect 51675 14912 51908 14940
rect 51675 14909 51687 14912
rect 51629 14903 51687 14909
rect 51902 14900 51908 14912
rect 51960 14940 51966 14952
rect 52380 14940 52408 14968
rect 51960 14912 52408 14940
rect 51960 14900 51966 14912
rect 53834 14900 53840 14952
rect 53892 14940 53898 14952
rect 53929 14943 53987 14949
rect 53929 14940 53941 14943
rect 53892 14912 53941 14940
rect 53892 14900 53898 14912
rect 53929 14909 53941 14912
rect 53975 14909 53987 14943
rect 53929 14903 53987 14909
rect 55677 14943 55735 14949
rect 55677 14909 55689 14943
rect 55723 14909 55735 14943
rect 55677 14903 55735 14909
rect 55692 14872 55720 14903
rect 55950 14900 55956 14952
rect 56008 14940 56014 14952
rect 56597 14943 56655 14949
rect 56597 14940 56609 14943
rect 56008 14912 56609 14940
rect 56008 14900 56014 14912
rect 56597 14909 56609 14912
rect 56643 14909 56655 14943
rect 56597 14903 56655 14909
rect 56686 14900 56692 14952
rect 56744 14949 56750 14952
rect 56744 14943 56772 14949
rect 56760 14909 56772 14943
rect 56744 14903 56772 14909
rect 56744 14900 56750 14903
rect 57882 14900 57888 14952
rect 57940 14900 57946 14952
rect 56134 14872 56140 14884
rect 51184 14844 52040 14872
rect 55692 14844 56140 14872
rect 50433 14835 50491 14841
rect 52012 14816 52040 14844
rect 56134 14832 56140 14844
rect 56192 14832 56198 14884
rect 56318 14832 56324 14884
rect 56376 14832 56382 14884
rect 24268 14776 25268 14804
rect 24268 14764 24274 14776
rect 25682 14764 25688 14816
rect 25740 14764 25746 14816
rect 26694 14764 26700 14816
rect 26752 14804 26758 14816
rect 27433 14807 27491 14813
rect 27433 14804 27445 14807
rect 26752 14776 27445 14804
rect 26752 14764 26758 14776
rect 27433 14773 27445 14776
rect 27479 14773 27491 14807
rect 27433 14767 27491 14773
rect 33318 14764 33324 14816
rect 33376 14804 33382 14816
rect 33505 14807 33563 14813
rect 33505 14804 33517 14807
rect 33376 14776 33517 14804
rect 33376 14764 33382 14776
rect 33505 14773 33517 14776
rect 33551 14804 33563 14807
rect 34974 14804 34980 14816
rect 33551 14776 34980 14804
rect 33551 14773 33563 14776
rect 33505 14767 33563 14773
rect 34974 14764 34980 14776
rect 35032 14764 35038 14816
rect 36262 14764 36268 14816
rect 36320 14804 36326 14816
rect 37093 14807 37151 14813
rect 37093 14804 37105 14807
rect 36320 14776 37105 14804
rect 36320 14764 36326 14776
rect 37093 14773 37105 14776
rect 37139 14773 37151 14807
rect 37093 14767 37151 14773
rect 37458 14764 37464 14816
rect 37516 14764 37522 14816
rect 38654 14764 38660 14816
rect 38712 14804 38718 14816
rect 39666 14804 39672 14816
rect 38712 14776 39672 14804
rect 38712 14764 38718 14776
rect 39666 14764 39672 14776
rect 39724 14764 39730 14816
rect 42058 14764 42064 14816
rect 42116 14764 42122 14816
rect 44174 14764 44180 14816
rect 44232 14764 44238 14816
rect 44910 14764 44916 14816
rect 44968 14764 44974 14816
rect 46566 14764 46572 14816
rect 46624 14764 46630 14816
rect 46750 14764 46756 14816
rect 46808 14764 46814 14816
rect 49694 14764 49700 14816
rect 49752 14764 49758 14816
rect 51994 14764 52000 14816
rect 52052 14764 52058 14816
rect 55309 14807 55367 14813
rect 55309 14773 55321 14807
rect 55355 14804 55367 14807
rect 55674 14804 55680 14816
rect 55355 14776 55680 14804
rect 55355 14773 55367 14776
rect 55309 14767 55367 14773
rect 55674 14764 55680 14776
rect 55732 14804 55738 14816
rect 56686 14804 56692 14816
rect 55732 14776 56692 14804
rect 55732 14764 55738 14776
rect 56686 14764 56692 14776
rect 56744 14764 56750 14816
rect 57514 14764 57520 14816
rect 57572 14764 57578 14816
rect 1104 14714 58880 14736
rect 1104 14662 8172 14714
rect 8224 14662 8236 14714
rect 8288 14662 8300 14714
rect 8352 14662 8364 14714
rect 8416 14662 8428 14714
rect 8480 14662 22616 14714
rect 22668 14662 22680 14714
rect 22732 14662 22744 14714
rect 22796 14662 22808 14714
rect 22860 14662 22872 14714
rect 22924 14662 37060 14714
rect 37112 14662 37124 14714
rect 37176 14662 37188 14714
rect 37240 14662 37252 14714
rect 37304 14662 37316 14714
rect 37368 14662 51504 14714
rect 51556 14662 51568 14714
rect 51620 14662 51632 14714
rect 51684 14662 51696 14714
rect 51748 14662 51760 14714
rect 51812 14662 58880 14714
rect 1104 14640 58880 14662
rect 4706 14600 4712 14612
rect 2746 14572 4712 14600
rect 2746 14464 2774 14572
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 6454 14600 6460 14612
rect 6135 14572 6460 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 6454 14560 6460 14572
rect 6512 14600 6518 14612
rect 7742 14600 7748 14612
rect 6512 14572 7748 14600
rect 6512 14560 6518 14572
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 8076 14572 8125 14600
rect 8076 14560 8082 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8938 14560 8944 14612
rect 8996 14560 9002 14612
rect 11146 14600 11152 14612
rect 9508 14572 11152 14600
rect 4724 14473 4752 14560
rect 1964 14436 2774 14464
rect 4709 14467 4767 14473
rect 1964 14408 1992 14436
rect 4709 14433 4721 14467
rect 4755 14433 4767 14467
rect 4709 14427 4767 14433
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 2222 14356 2228 14408
rect 2280 14356 2286 14408
rect 4724 14396 4752 14427
rect 9398 14424 9404 14476
rect 9456 14424 9462 14476
rect 9508 14473 9536 14572
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 19208 14572 19257 14600
rect 19208 14560 19214 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 19245 14563 19303 14569
rect 21652 14572 22692 14600
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 9858 14424 9864 14476
rect 9916 14424 9922 14476
rect 18322 14424 18328 14476
rect 18380 14464 18386 14476
rect 19426 14464 19432 14476
rect 18380 14436 19432 14464
rect 18380 14424 18386 14436
rect 19426 14424 19432 14436
rect 19484 14464 19490 14476
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 19484 14436 19809 14464
rect 19484 14424 19490 14436
rect 19797 14433 19809 14436
rect 19843 14464 19855 14467
rect 21652 14464 21680 14572
rect 22664 14532 22692 14572
rect 23198 14560 23204 14612
rect 23256 14560 23262 14612
rect 23676 14572 25544 14600
rect 23676 14532 23704 14572
rect 22664 14504 23704 14532
rect 25516 14532 25544 14572
rect 25866 14560 25872 14612
rect 25924 14600 25930 14612
rect 26053 14603 26111 14609
rect 26053 14600 26065 14603
rect 25924 14572 26065 14600
rect 25924 14560 25930 14572
rect 26053 14569 26065 14572
rect 26099 14569 26111 14603
rect 26053 14563 26111 14569
rect 29270 14560 29276 14612
rect 29328 14600 29334 14612
rect 31018 14600 31024 14612
rect 29328 14572 31024 14600
rect 29328 14560 29334 14572
rect 31018 14560 31024 14572
rect 31076 14600 31082 14612
rect 31662 14600 31668 14612
rect 31076 14572 31668 14600
rect 31076 14560 31082 14572
rect 31662 14560 31668 14572
rect 31720 14600 31726 14612
rect 32401 14603 32459 14609
rect 32401 14600 32413 14603
rect 31720 14572 32413 14600
rect 31720 14560 31726 14572
rect 32401 14569 32413 14572
rect 32447 14569 32459 14603
rect 32401 14563 32459 14569
rect 34054 14560 34060 14612
rect 34112 14560 34118 14612
rect 41690 14560 41696 14612
rect 41748 14560 41754 14612
rect 44174 14560 44180 14612
rect 44232 14560 44238 14612
rect 46566 14600 46572 14612
rect 46032 14572 46572 14600
rect 26418 14532 26424 14544
rect 25516 14504 26424 14532
rect 26418 14492 26424 14504
rect 26476 14532 26482 14544
rect 26476 14504 26648 14532
rect 26476 14492 26482 14504
rect 19843 14436 21680 14464
rect 19843 14433 19855 14436
rect 19797 14427 19855 14433
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 21784 14436 21864 14464
rect 21784 14424 21790 14436
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 4724 14368 6745 14396
rect 6733 14365 6745 14368
rect 6779 14396 6791 14399
rect 8570 14396 8576 14408
rect 6779 14368 8576 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 12618 14396 12624 14408
rect 12391 14368 12624 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 17589 14399 17647 14405
rect 17589 14365 17601 14399
rect 17635 14396 17647 14399
rect 18046 14396 18052 14408
rect 17635 14368 18052 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18230 14356 18236 14408
rect 18288 14356 18294 14408
rect 19978 14356 19984 14408
rect 20036 14396 20042 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 20036 14368 20085 14396
rect 20036 14356 20042 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 21836 14396 21864 14436
rect 22738 14424 22744 14476
rect 22796 14464 22802 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 22796 14436 23765 14464
rect 22796 14424 22802 14436
rect 23753 14433 23765 14436
rect 23799 14464 23811 14467
rect 23799 14436 24716 14464
rect 23799 14433 23811 14436
rect 23753 14427 23811 14433
rect 24688 14408 24716 14436
rect 26510 14424 26516 14476
rect 26568 14424 26574 14476
rect 26620 14473 26648 14504
rect 31846 14492 31852 14544
rect 31904 14532 31910 14544
rect 34072 14532 34100 14560
rect 39853 14535 39911 14541
rect 39853 14532 39865 14535
rect 31904 14504 34100 14532
rect 39132 14504 39865 14532
rect 31904 14492 31910 14504
rect 26605 14467 26663 14473
rect 26605 14433 26617 14467
rect 26651 14433 26663 14467
rect 26605 14427 26663 14433
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 35618 14464 35624 14476
rect 34848 14436 35624 14464
rect 34848 14424 34854 14436
rect 35618 14424 35624 14436
rect 35676 14424 35682 14476
rect 39132 14473 39160 14504
rect 39853 14501 39865 14504
rect 39899 14501 39911 14535
rect 41708 14532 41736 14560
rect 42705 14535 42763 14541
rect 41708 14504 42472 14532
rect 39853 14495 39911 14501
rect 39117 14467 39175 14473
rect 39117 14433 39129 14467
rect 39163 14433 39175 14467
rect 39117 14427 39175 14433
rect 39666 14424 39672 14476
rect 39724 14464 39730 14476
rect 42444 14473 42472 14504
rect 42705 14501 42717 14535
rect 42751 14532 42763 14535
rect 42751 14504 43576 14532
rect 42751 14501 42763 14504
rect 42705 14495 42763 14501
rect 40405 14467 40463 14473
rect 40405 14464 40417 14467
rect 39724 14436 40417 14464
rect 39724 14424 39730 14436
rect 40405 14433 40417 14436
rect 40451 14433 40463 14467
rect 42429 14467 42487 14473
rect 40405 14427 40463 14433
rect 40512 14436 42288 14464
rect 24486 14396 24492 14408
rect 21836 14368 24492 14396
rect 24486 14356 24492 14368
rect 24544 14396 24550 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24544 14368 24593 14396
rect 24544 14356 24550 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24670 14356 24676 14408
rect 24728 14356 24734 14408
rect 25682 14396 25688 14408
rect 24780 14368 25688 14396
rect 4976 14331 5034 14337
rect 4976 14297 4988 14331
rect 5022 14328 5034 14331
rect 5902 14328 5908 14340
rect 5022 14300 5908 14328
rect 5022 14297 5034 14300
rect 4976 14291 5034 14297
rect 5902 14288 5908 14300
rect 5960 14288 5966 14340
rect 7000 14331 7058 14337
rect 7000 14297 7012 14331
rect 7046 14328 7058 14331
rect 7834 14328 7840 14340
rect 7046 14300 7840 14328
rect 7046 14297 7058 14300
rect 7000 14291 7058 14297
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 9309 14331 9367 14337
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 10413 14331 10471 14337
rect 10413 14328 10425 14331
rect 9355 14300 10425 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 10413 14297 10425 14300
rect 10459 14297 10471 14331
rect 10413 14291 10471 14297
rect 21996 14331 22054 14337
rect 21996 14297 22008 14331
rect 22042 14328 22054 14331
rect 22370 14328 22376 14340
rect 22042 14300 22376 14328
rect 22042 14297 22054 14300
rect 21996 14291 22054 14297
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 23569 14331 23627 14337
rect 23569 14328 23581 14331
rect 23032 14300 23581 14328
rect 23032 14272 23060 14300
rect 23569 14297 23581 14300
rect 23615 14297 23627 14331
rect 23569 14291 23627 14297
rect 23658 14288 23664 14340
rect 23716 14288 23722 14340
rect 23842 14288 23848 14340
rect 23900 14328 23906 14340
rect 24780 14328 24808 14368
rect 25682 14356 25688 14368
rect 25740 14356 25746 14408
rect 26881 14399 26939 14405
rect 26881 14396 26893 14399
rect 25976 14368 26893 14396
rect 23900 14300 24808 14328
rect 24848 14331 24906 14337
rect 23900 14288 23906 14300
rect 24848 14297 24860 14331
rect 24894 14328 24906 14331
rect 25774 14328 25780 14340
rect 24894 14300 25780 14328
rect 24894 14297 24906 14300
rect 24848 14291 24906 14297
rect 25774 14288 25780 14300
rect 25832 14288 25838 14340
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 6178 14220 6184 14272
rect 6236 14260 6242 14272
rect 6641 14263 6699 14269
rect 6641 14260 6653 14263
rect 6236 14232 6653 14260
rect 6236 14220 6242 14232
rect 6641 14229 6653 14232
rect 6687 14260 6699 14263
rect 7466 14260 7472 14272
rect 6687 14232 7472 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 9122 14260 9128 14272
rect 8812 14232 9128 14260
rect 8812 14220 8818 14232
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 12894 14220 12900 14272
rect 12952 14220 12958 14272
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 16540 14232 17325 14260
rect 16540 14220 16546 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 17313 14223 17371 14229
rect 18138 14220 18144 14272
rect 18196 14220 18202 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 18877 14263 18935 14269
rect 18877 14260 18889 14263
rect 18472 14232 18889 14260
rect 18472 14220 18478 14232
rect 18877 14229 18889 14232
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 19610 14220 19616 14272
rect 19668 14220 19674 14272
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 19751 14232 20729 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 21450 14220 21456 14272
rect 21508 14220 21514 14272
rect 23014 14220 23020 14272
rect 23072 14220 23078 14272
rect 23106 14220 23112 14272
rect 23164 14220 23170 14272
rect 23474 14220 23480 14272
rect 23532 14260 23538 14272
rect 25976 14269 26004 14368
rect 26881 14365 26893 14368
rect 26927 14365 26939 14399
rect 26881 14359 26939 14365
rect 28074 14356 28080 14408
rect 28132 14356 28138 14408
rect 28810 14356 28816 14408
rect 28868 14356 28874 14408
rect 29730 14356 29736 14408
rect 29788 14396 29794 14408
rect 29917 14399 29975 14405
rect 29917 14396 29929 14399
rect 29788 14368 29929 14396
rect 29788 14356 29794 14368
rect 29917 14365 29929 14368
rect 29963 14365 29975 14399
rect 29917 14359 29975 14365
rect 35250 14356 35256 14408
rect 35308 14396 35314 14408
rect 35897 14399 35955 14405
rect 35897 14396 35909 14399
rect 35308 14368 35909 14396
rect 35308 14356 35314 14368
rect 35897 14365 35909 14368
rect 35943 14365 35955 14399
rect 35897 14359 35955 14365
rect 36630 14356 36636 14408
rect 36688 14396 36694 14408
rect 37369 14399 37427 14405
rect 37369 14396 37381 14399
rect 36688 14368 37381 14396
rect 36688 14356 36694 14368
rect 37369 14365 37381 14368
rect 37415 14365 37427 14399
rect 40512 14396 40540 14436
rect 37369 14359 37427 14365
rect 40144 14368 40540 14396
rect 36164 14331 36222 14337
rect 36164 14297 36176 14331
rect 36210 14328 36222 14331
rect 38102 14328 38108 14340
rect 36210 14300 38108 14328
rect 36210 14297 36222 14300
rect 36164 14291 36222 14297
rect 38102 14288 38108 14300
rect 38160 14288 38166 14340
rect 40144 14272 40172 14368
rect 40678 14356 40684 14408
rect 40736 14356 40742 14408
rect 42260 14405 42288 14436
rect 42429 14433 42441 14467
rect 42475 14433 42487 14467
rect 42429 14427 42487 14433
rect 43346 14424 43352 14476
rect 43404 14424 43410 14476
rect 43548 14473 43576 14504
rect 43533 14467 43591 14473
rect 43533 14433 43545 14467
rect 43579 14433 43591 14467
rect 43533 14427 43591 14433
rect 42245 14399 42303 14405
rect 42245 14365 42257 14399
rect 42291 14365 42303 14399
rect 42245 14359 42303 14365
rect 43073 14399 43131 14405
rect 43073 14365 43085 14399
rect 43119 14396 43131 14399
rect 44192 14396 44220 14560
rect 45005 14399 45063 14405
rect 45005 14396 45017 14399
rect 43119 14368 44220 14396
rect 44744 14368 45017 14396
rect 43119 14365 43131 14368
rect 43073 14359 43131 14365
rect 40221 14331 40279 14337
rect 40221 14297 40233 14331
rect 40267 14328 40279 14331
rect 41325 14331 41383 14337
rect 41325 14328 41337 14331
rect 40267 14300 41337 14328
rect 40267 14297 40279 14300
rect 40221 14291 40279 14297
rect 41325 14297 41337 14300
rect 41371 14297 41383 14331
rect 42058 14328 42064 14340
rect 41325 14291 41383 14297
rect 41708 14300 42064 14328
rect 25961 14263 26019 14269
rect 25961 14260 25973 14263
rect 23532 14232 25973 14260
rect 23532 14220 23538 14232
rect 25961 14229 25973 14232
rect 26007 14229 26019 14263
rect 25961 14223 26019 14229
rect 26142 14220 26148 14272
rect 26200 14260 26206 14272
rect 26421 14263 26479 14269
rect 26421 14260 26433 14263
rect 26200 14232 26433 14260
rect 26200 14220 26206 14232
rect 26421 14229 26433 14232
rect 26467 14229 26479 14263
rect 26421 14223 26479 14229
rect 27522 14220 27528 14272
rect 27580 14220 27586 14272
rect 28626 14220 28632 14272
rect 28684 14220 28690 14272
rect 28994 14220 29000 14272
rect 29052 14260 29058 14272
rect 29365 14263 29423 14269
rect 29365 14260 29377 14263
rect 29052 14232 29377 14260
rect 29052 14220 29058 14232
rect 29365 14229 29377 14232
rect 29411 14229 29423 14263
rect 29365 14223 29423 14229
rect 30558 14220 30564 14272
rect 30616 14220 30622 14272
rect 30650 14220 30656 14272
rect 30708 14260 30714 14272
rect 31386 14260 31392 14272
rect 30708 14232 31392 14260
rect 30708 14220 30714 14232
rect 31386 14220 31392 14232
rect 31444 14220 31450 14272
rect 35342 14220 35348 14272
rect 35400 14220 35406 14272
rect 37277 14263 37335 14269
rect 37277 14229 37289 14263
rect 37323 14260 37335 14263
rect 37550 14260 37556 14272
rect 37323 14232 37556 14260
rect 37323 14229 37335 14232
rect 37277 14223 37335 14229
rect 37550 14220 37556 14232
rect 37608 14220 37614 14272
rect 38010 14220 38016 14272
rect 38068 14220 38074 14272
rect 39666 14220 39672 14272
rect 39724 14220 39730 14272
rect 40126 14220 40132 14272
rect 40184 14260 40190 14272
rect 40313 14263 40371 14269
rect 40313 14260 40325 14263
rect 40184 14232 40325 14260
rect 40184 14220 40190 14232
rect 40313 14229 40325 14232
rect 40359 14229 40371 14263
rect 40313 14223 40371 14229
rect 40586 14220 40592 14272
rect 40644 14260 40650 14272
rect 41708 14260 41736 14300
rect 42058 14288 42064 14300
rect 42116 14288 42122 14340
rect 42260 14328 42288 14359
rect 43165 14331 43223 14337
rect 43165 14328 43177 14331
rect 42260 14300 43177 14328
rect 43165 14297 43177 14300
rect 43211 14297 43223 14331
rect 43165 14291 43223 14297
rect 44744 14272 44772 14368
rect 45005 14365 45017 14368
rect 45051 14365 45063 14399
rect 45005 14359 45063 14365
rect 45272 14399 45330 14405
rect 45272 14365 45284 14399
rect 45318 14396 45330 14399
rect 46032 14396 46060 14572
rect 46566 14560 46572 14572
rect 46624 14560 46630 14612
rect 49234 14560 49240 14612
rect 49292 14560 49298 14612
rect 49694 14560 49700 14612
rect 49752 14560 49758 14612
rect 51537 14603 51595 14609
rect 51537 14569 51549 14603
rect 51583 14600 51595 14603
rect 51902 14600 51908 14612
rect 51583 14572 51908 14600
rect 51583 14569 51595 14572
rect 51537 14563 51595 14569
rect 51902 14560 51908 14572
rect 51960 14560 51966 14612
rect 54478 14600 54484 14612
rect 52288 14572 54484 14600
rect 46385 14535 46443 14541
rect 46385 14501 46397 14535
rect 46431 14532 46443 14535
rect 46750 14532 46756 14544
rect 46431 14504 46756 14532
rect 46431 14501 46443 14504
rect 46385 14495 46443 14501
rect 46750 14492 46756 14504
rect 46808 14532 46814 14544
rect 46808 14504 47256 14532
rect 46808 14492 46814 14504
rect 47026 14424 47032 14476
rect 47084 14464 47090 14476
rect 47121 14467 47179 14473
rect 47121 14464 47133 14467
rect 47084 14436 47133 14464
rect 47084 14424 47090 14436
rect 47121 14433 47133 14436
rect 47167 14433 47179 14467
rect 47228 14464 47256 14504
rect 47397 14467 47455 14473
rect 47397 14464 47409 14467
rect 47228 14436 47409 14464
rect 47121 14427 47179 14433
rect 47397 14433 47409 14436
rect 47443 14433 47455 14467
rect 47397 14427 47455 14433
rect 47673 14467 47731 14473
rect 47673 14433 47685 14467
rect 47719 14464 47731 14467
rect 47854 14464 47860 14476
rect 47719 14436 47860 14464
rect 47719 14433 47731 14436
rect 47673 14427 47731 14433
rect 47854 14424 47860 14436
rect 47912 14424 47918 14476
rect 48406 14424 48412 14476
rect 48464 14464 48470 14476
rect 49712 14473 49740 14560
rect 48961 14467 49019 14473
rect 48961 14464 48973 14467
rect 48464 14436 48973 14464
rect 48464 14424 48470 14436
rect 48961 14433 48973 14436
rect 49007 14433 49019 14467
rect 48961 14427 49019 14433
rect 49697 14467 49755 14473
rect 49697 14433 49709 14467
rect 49743 14433 49755 14467
rect 49697 14427 49755 14433
rect 49789 14467 49847 14473
rect 49789 14433 49801 14467
rect 49835 14433 49847 14467
rect 49789 14427 49847 14433
rect 45318 14368 46060 14396
rect 45318 14365 45330 14368
rect 45272 14359 45330 14365
rect 46474 14356 46480 14408
rect 46532 14356 46538 14408
rect 46661 14399 46719 14405
rect 46661 14365 46673 14399
rect 46707 14365 46719 14399
rect 46661 14359 46719 14365
rect 40644 14232 41736 14260
rect 40644 14220 40650 14232
rect 41782 14220 41788 14272
rect 41840 14260 41846 14272
rect 41877 14263 41935 14269
rect 41877 14260 41889 14263
rect 41840 14232 41889 14260
rect 41840 14220 41846 14232
rect 41877 14229 41889 14232
rect 41923 14229 41935 14263
rect 41877 14223 41935 14229
rect 42337 14263 42395 14269
rect 42337 14229 42349 14263
rect 42383 14260 42395 14263
rect 43070 14260 43076 14272
rect 42383 14232 43076 14260
rect 42383 14229 42395 14232
rect 42337 14223 42395 14229
rect 43070 14220 43076 14232
rect 43128 14220 43134 14272
rect 44174 14220 44180 14272
rect 44232 14220 44238 14272
rect 44726 14220 44732 14272
rect 44784 14220 44790 14272
rect 46676 14260 46704 14359
rect 47486 14356 47492 14408
rect 47544 14405 47550 14408
rect 47544 14399 47572 14405
rect 47560 14365 47572 14399
rect 47544 14359 47572 14365
rect 47544 14356 47550 14359
rect 49142 14356 49148 14408
rect 49200 14396 49206 14408
rect 49804 14396 49832 14427
rect 51350 14424 51356 14476
rect 51408 14464 51414 14476
rect 52086 14464 52092 14476
rect 51408 14436 52092 14464
rect 51408 14424 51414 14436
rect 52086 14424 52092 14436
rect 52144 14424 52150 14476
rect 52178 14424 52184 14476
rect 52236 14464 52242 14476
rect 52288 14473 52316 14572
rect 54478 14560 54484 14572
rect 54536 14560 54542 14612
rect 55125 14603 55183 14609
rect 55125 14569 55137 14603
rect 55171 14600 55183 14603
rect 55950 14600 55956 14612
rect 55171 14572 55956 14600
rect 55171 14569 55183 14572
rect 55125 14563 55183 14569
rect 55950 14560 55956 14572
rect 56008 14560 56014 14612
rect 56134 14560 56140 14612
rect 56192 14600 56198 14612
rect 57517 14603 57575 14609
rect 57517 14600 57529 14603
rect 56192 14572 57529 14600
rect 56192 14560 56198 14572
rect 57517 14569 57529 14572
rect 57563 14569 57575 14603
rect 57517 14563 57575 14569
rect 57609 14603 57667 14609
rect 57609 14569 57621 14603
rect 57655 14600 57667 14603
rect 57882 14600 57888 14612
rect 57655 14572 57888 14600
rect 57655 14569 57667 14572
rect 57609 14563 57667 14569
rect 57532 14532 57560 14563
rect 57882 14560 57888 14572
rect 57940 14560 57946 14612
rect 57698 14532 57704 14544
rect 54772 14504 55904 14532
rect 57532 14504 57704 14532
rect 54772 14476 54800 14504
rect 52273 14467 52331 14473
rect 52273 14464 52285 14467
rect 52236 14436 52285 14464
rect 52236 14424 52242 14436
rect 52273 14433 52285 14436
rect 52319 14433 52331 14467
rect 53745 14467 53803 14473
rect 53745 14464 53757 14467
rect 52273 14427 52331 14433
rect 52380 14436 53757 14464
rect 49200 14368 49832 14396
rect 50157 14399 50215 14405
rect 49200 14356 49206 14368
rect 50157 14365 50169 14399
rect 50203 14396 50215 14399
rect 50246 14396 50252 14408
rect 50203 14368 50252 14396
rect 50203 14365 50215 14368
rect 50157 14359 50215 14365
rect 50246 14356 50252 14368
rect 50304 14396 50310 14408
rect 52380 14396 52408 14436
rect 53745 14433 53757 14436
rect 53791 14433 53803 14467
rect 53745 14427 53803 14433
rect 50304 14368 52408 14396
rect 52457 14399 52515 14405
rect 50304 14356 50310 14368
rect 52457 14365 52469 14399
rect 52503 14365 52515 14399
rect 53760 14396 53788 14427
rect 54754 14424 54760 14476
rect 54812 14424 54818 14476
rect 55582 14424 55588 14476
rect 55640 14464 55646 14476
rect 55876 14473 55904 14504
rect 57698 14492 57704 14504
rect 57756 14492 57762 14544
rect 55769 14467 55827 14473
rect 55769 14464 55781 14467
rect 55640 14436 55781 14464
rect 55640 14424 55646 14436
rect 55769 14433 55781 14436
rect 55815 14433 55827 14467
rect 55769 14427 55827 14433
rect 55861 14467 55919 14473
rect 55861 14433 55873 14467
rect 55907 14433 55919 14467
rect 55861 14427 55919 14433
rect 57330 14424 57336 14476
rect 57388 14464 57394 14476
rect 58161 14467 58219 14473
rect 58161 14464 58173 14467
rect 57388 14436 58173 14464
rect 57388 14424 57394 14436
rect 58161 14433 58173 14436
rect 58207 14433 58219 14467
rect 58161 14427 58219 14433
rect 53834 14396 53840 14408
rect 53760 14368 53840 14396
rect 52457 14359 52515 14365
rect 50424 14331 50482 14337
rect 50424 14297 50436 14331
rect 50470 14328 50482 14331
rect 51258 14328 51264 14340
rect 50470 14300 51264 14328
rect 50470 14297 50482 14300
rect 50424 14291 50482 14297
rect 51258 14288 51264 14300
rect 51316 14288 51322 14340
rect 51718 14288 51724 14340
rect 51776 14328 51782 14340
rect 52270 14328 52276 14340
rect 51776 14300 52276 14328
rect 51776 14288 51782 14300
rect 52270 14288 52276 14300
rect 52328 14328 52334 14340
rect 52472 14328 52500 14359
rect 53834 14356 53840 14368
rect 53892 14396 53898 14408
rect 56137 14399 56195 14405
rect 56137 14396 56149 14399
rect 53892 14368 56149 14396
rect 53892 14356 53898 14368
rect 56137 14365 56149 14368
rect 56183 14365 56195 14399
rect 56137 14359 56195 14365
rect 57974 14356 57980 14408
rect 58032 14356 58038 14408
rect 52328 14300 52500 14328
rect 54012 14331 54070 14337
rect 52328 14288 52334 14300
rect 54012 14297 54024 14331
rect 54058 14328 54070 14331
rect 54570 14328 54576 14340
rect 54058 14300 54576 14328
rect 54058 14297 54070 14300
rect 54012 14291 54070 14297
rect 54570 14288 54576 14300
rect 54628 14288 54634 14340
rect 55677 14331 55735 14337
rect 55677 14297 55689 14331
rect 55723 14328 55735 14331
rect 55858 14328 55864 14340
rect 55723 14300 55864 14328
rect 55723 14297 55735 14300
rect 55677 14291 55735 14297
rect 55858 14288 55864 14300
rect 55916 14288 55922 14340
rect 56404 14331 56462 14337
rect 56404 14297 56416 14331
rect 56450 14328 56462 14331
rect 57146 14328 57152 14340
rect 56450 14300 57152 14328
rect 56450 14297 56462 14300
rect 56404 14291 56462 14297
rect 57146 14288 57152 14300
rect 57204 14288 57210 14340
rect 48222 14260 48228 14272
rect 46676 14232 48228 14260
rect 48222 14220 48228 14232
rect 48280 14220 48286 14272
rect 48314 14220 48320 14272
rect 48372 14220 48378 14272
rect 48406 14220 48412 14272
rect 48464 14220 48470 14272
rect 48774 14220 48780 14272
rect 48832 14220 48838 14272
rect 48869 14263 48927 14269
rect 48869 14229 48881 14263
rect 48915 14260 48927 14263
rect 48958 14260 48964 14272
rect 48915 14232 48964 14260
rect 48915 14229 48927 14232
rect 48869 14223 48927 14229
rect 48958 14220 48964 14232
rect 49016 14260 49022 14272
rect 49605 14263 49663 14269
rect 49605 14260 49617 14263
rect 49016 14232 49617 14260
rect 49016 14220 49022 14232
rect 49605 14229 49617 14232
rect 49651 14229 49663 14263
rect 49605 14223 49663 14229
rect 51626 14220 51632 14272
rect 51684 14220 51690 14272
rect 51994 14220 52000 14272
rect 52052 14220 52058 14272
rect 52089 14263 52147 14269
rect 52089 14229 52101 14263
rect 52135 14260 52147 14263
rect 53101 14263 53159 14269
rect 53101 14260 53113 14263
rect 52135 14232 53113 14260
rect 52135 14229 52147 14232
rect 52089 14223 52147 14229
rect 53101 14229 53113 14232
rect 53147 14229 53159 14263
rect 53101 14223 53159 14229
rect 55306 14220 55312 14272
rect 55364 14220 55370 14272
rect 56870 14220 56876 14272
rect 56928 14260 56934 14272
rect 58069 14263 58127 14269
rect 58069 14260 58081 14263
rect 56928 14232 58081 14260
rect 56928 14220 56934 14232
rect 58069 14229 58081 14232
rect 58115 14229 58127 14263
rect 58069 14223 58127 14229
rect 1104 14170 59040 14192
rect 1104 14118 15394 14170
rect 15446 14118 15458 14170
rect 15510 14118 15522 14170
rect 15574 14118 15586 14170
rect 15638 14118 15650 14170
rect 15702 14118 29838 14170
rect 29890 14118 29902 14170
rect 29954 14118 29966 14170
rect 30018 14118 30030 14170
rect 30082 14118 30094 14170
rect 30146 14118 44282 14170
rect 44334 14118 44346 14170
rect 44398 14118 44410 14170
rect 44462 14118 44474 14170
rect 44526 14118 44538 14170
rect 44590 14118 58726 14170
rect 58778 14118 58790 14170
rect 58842 14118 58854 14170
rect 58906 14118 58918 14170
rect 58970 14118 58982 14170
rect 59034 14118 59040 14170
rect 1104 14096 59040 14118
rect 2866 14056 2872 14068
rect 2746 14028 2872 14056
rect 2124 13991 2182 13997
rect 2124 13957 2136 13991
rect 2170 13988 2182 13991
rect 2746 13988 2774 14028
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 2170 13960 2774 13988
rect 2170 13957 2182 13960
rect 2124 13951 2182 13957
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 1946 13920 1952 13932
rect 1903 13892 1952 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 3252 13920 3280 14019
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5868 14028 5917 14056
rect 5868 14016 5874 14028
rect 5905 14025 5917 14028
rect 5951 14025 5963 14059
rect 5905 14019 5963 14025
rect 7834 14016 7840 14068
rect 7892 14016 7898 14068
rect 10229 14059 10287 14065
rect 10229 14025 10241 14059
rect 10275 14056 10287 14059
rect 11146 14056 11152 14068
rect 10275 14028 11152 14056
rect 10275 14025 10287 14028
rect 10229 14019 10287 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12894 14056 12900 14068
rect 12406 14028 12900 14056
rect 11784 13991 11842 13997
rect 11784 13957 11796 13991
rect 11830 13988 11842 13991
rect 12406 13988 12434 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 14553 14059 14611 14065
rect 14553 14025 14565 14059
rect 14599 14056 14611 14059
rect 14918 14056 14924 14068
rect 14599 14028 14924 14056
rect 14599 14025 14611 14028
rect 14553 14019 14611 14025
rect 11830 13960 12434 13988
rect 14108 13988 14136 14019
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18230 14056 18236 14068
rect 18095 14028 18236 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18230 14016 18236 14028
rect 18288 14056 18294 14068
rect 18288 14028 18828 14056
rect 18288 14016 18294 14028
rect 14108 13960 15148 13988
rect 11830 13957 11842 13960
rect 11784 13951 11842 13957
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 3252 13892 3341 13920
rect 3329 13889 3341 13892
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 5859 13892 7021 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 7282 13880 7288 13932
rect 7340 13880 7346 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 8018 13920 8024 13932
rect 7524 13892 8024 13920
rect 7524 13880 7530 13892
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 11422 13880 11428 13932
rect 11480 13920 11486 13932
rect 11480 13892 11560 13920
rect 11480 13880 11486 13892
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 6012 13784 6040 13815
rect 6454 13812 6460 13864
rect 6512 13812 6518 13864
rect 9214 13812 9220 13864
rect 9272 13812 9278 13864
rect 11532 13861 11560 13892
rect 14458 13880 14464 13932
rect 14516 13880 14522 13932
rect 15120 13929 15148 13960
rect 16684 13960 18644 13988
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 11517 13855 11575 13861
rect 11517 13821 11529 13855
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13722 13852 13728 13864
rect 13127 13824 13728 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 6086 13784 6092 13796
rect 6012 13756 6092 13784
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 12897 13787 12955 13793
rect 12897 13753 12909 13787
rect 12943 13784 12955 13787
rect 13096 13784 13124 13815
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14734 13852 14740 13864
rect 14047 13824 14740 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16684 13861 16712 13960
rect 16936 13923 16994 13929
rect 16936 13889 16948 13923
rect 16982 13920 16994 13923
rect 18138 13920 18144 13932
rect 16982 13892 18144 13920
rect 16982 13889 16994 13892
rect 16936 13883 16994 13889
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 18616 13929 18644 13960
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18800 13920 18828 14028
rect 18966 14016 18972 14068
rect 19024 14016 19030 14068
rect 19058 14016 19064 14068
rect 19116 14056 19122 14068
rect 19116 14028 19840 14056
rect 19116 14016 19122 14028
rect 18868 13991 18926 13997
rect 18868 13957 18880 13991
rect 18914 13988 18926 13991
rect 18984 13988 19012 14016
rect 18914 13960 19012 13988
rect 19812 13988 19840 14028
rect 19978 14016 19984 14068
rect 20036 14016 20042 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20806 14056 20812 14068
rect 20119 14028 20812 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 24578 14056 24584 14068
rect 23124 14028 24584 14056
rect 23124 14000 23152 14028
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 24670 14016 24676 14068
rect 24728 14056 24734 14068
rect 25777 14059 25835 14065
rect 24728 14028 25176 14056
rect 24728 14016 24734 14028
rect 22281 13991 22339 13997
rect 22281 13988 22293 13991
rect 19812 13960 22293 13988
rect 18914 13957 18926 13960
rect 18868 13951 18926 13957
rect 22281 13957 22293 13960
rect 22327 13988 22339 13991
rect 22738 13988 22744 14000
rect 22327 13960 22744 13988
rect 22327 13957 22339 13960
rect 22281 13951 22339 13957
rect 22738 13948 22744 13960
rect 22796 13948 22802 14000
rect 23106 13948 23112 14000
rect 23164 13948 23170 14000
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 25148 13988 25176 14028
rect 25777 14025 25789 14059
rect 25823 14056 25835 14059
rect 27522 14056 27528 14068
rect 25823 14028 27528 14056
rect 25823 14025 25835 14028
rect 25777 14019 25835 14025
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 28074 14016 28080 14068
rect 28132 14056 28138 14068
rect 28169 14059 28227 14065
rect 28169 14056 28181 14059
rect 28132 14028 28181 14056
rect 28132 14016 28138 14028
rect 28169 14025 28181 14028
rect 28215 14025 28227 14059
rect 28169 14019 28227 14025
rect 28629 14059 28687 14065
rect 28629 14025 28641 14059
rect 28675 14056 28687 14059
rect 28994 14056 29000 14068
rect 28675 14028 29000 14056
rect 28675 14025 28687 14028
rect 28629 14019 28687 14025
rect 28994 14016 29000 14028
rect 29052 14016 29058 14068
rect 29270 14016 29276 14068
rect 29328 14016 29334 14068
rect 30558 14016 30564 14068
rect 30616 14016 30622 14068
rect 31018 14016 31024 14068
rect 31076 14056 31082 14068
rect 31665 14059 31723 14065
rect 31665 14056 31677 14059
rect 31076 14028 31677 14056
rect 31076 14016 31082 14028
rect 31665 14025 31677 14028
rect 31711 14025 31723 14059
rect 31665 14019 31723 14025
rect 33965 14059 34023 14065
rect 33965 14025 33977 14059
rect 34011 14056 34023 14059
rect 34790 14056 34796 14068
rect 34011 14028 34796 14056
rect 34011 14025 34023 14028
rect 33965 14019 34023 14025
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 34974 14016 34980 14068
rect 35032 14056 35038 14068
rect 36078 14056 36084 14068
rect 35032 14028 36084 14056
rect 35032 14016 35038 14028
rect 36078 14016 36084 14028
rect 36136 14016 36142 14068
rect 36538 14016 36544 14068
rect 36596 14056 36602 14068
rect 37277 14059 37335 14065
rect 37277 14056 37289 14059
rect 36596 14028 37289 14056
rect 36596 14016 36602 14028
rect 37277 14025 37289 14028
rect 37323 14025 37335 14059
rect 37277 14019 37335 14025
rect 37737 14059 37795 14065
rect 37737 14025 37749 14059
rect 37783 14056 37795 14059
rect 38010 14056 38016 14068
rect 37783 14028 38016 14056
rect 37783 14025 37795 14028
rect 37737 14019 37795 14025
rect 38010 14016 38016 14028
rect 38068 14016 38074 14068
rect 39853 14059 39911 14065
rect 39853 14025 39865 14059
rect 39899 14056 39911 14059
rect 42058 14056 42064 14068
rect 39899 14028 40356 14056
rect 39899 14025 39911 14028
rect 39853 14019 39911 14025
rect 23532 13960 23704 13988
rect 25148 13960 27384 13988
rect 23532 13948 23538 13960
rect 20162 13920 20168 13932
rect 18800 13892 20168 13920
rect 18601 13883 18659 13889
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 21545 13923 21603 13929
rect 21545 13920 21557 13923
rect 20487 13892 21557 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 21545 13889 21557 13892
rect 21591 13889 21603 13923
rect 21545 13883 21603 13889
rect 22833 13923 22891 13929
rect 22833 13889 22845 13923
rect 22879 13920 22891 13923
rect 23566 13920 23572 13932
rect 22879 13892 23572 13920
rect 22879 13889 22891 13892
rect 22833 13883 22891 13889
rect 23566 13880 23572 13892
rect 23624 13880 23630 13932
rect 23676 13929 23704 13960
rect 24578 13929 24584 13932
rect 23661 13923 23719 13929
rect 23661 13889 23673 13923
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 24535 13923 24584 13929
rect 24535 13889 24547 13923
rect 24581 13889 24584 13923
rect 24535 13883 24584 13889
rect 24578 13880 24584 13883
rect 24636 13880 24642 13932
rect 26142 13920 26148 13932
rect 25884 13892 26148 13920
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16540 13824 16681 13852
rect 16540 13812 16546 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 18506 13812 18512 13864
rect 18564 13812 18570 13864
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 19668 13824 20545 13852
rect 19668 13812 19674 13824
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 20640 13784 20668 13815
rect 20990 13812 20996 13864
rect 21048 13812 21054 13864
rect 22925 13855 22983 13861
rect 22925 13821 22937 13855
rect 22971 13852 22983 13855
rect 23014 13852 23020 13864
rect 22971 13824 23020 13852
rect 22971 13821 22983 13824
rect 22925 13815 22983 13821
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23523 13824 23704 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 21542 13784 21548 13796
rect 12943 13756 13124 13784
rect 20548 13756 21548 13784
rect 12943 13753 12955 13756
rect 12897 13747 12955 13753
rect 3970 13676 3976 13728
rect 4028 13676 4034 13728
rect 5442 13676 5448 13728
rect 5500 13676 5506 13728
rect 9858 13676 9864 13728
rect 9916 13676 9922 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13136 13688 13645 13716
rect 13136 13676 13142 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13633 13679 13691 13685
rect 15746 13676 15752 13728
rect 15804 13676 15810 13728
rect 18966 13676 18972 13728
rect 19024 13716 19030 13728
rect 20548 13716 20576 13756
rect 21542 13744 21548 13756
rect 21600 13784 21606 13796
rect 23124 13784 23152 13815
rect 23382 13784 23388 13796
rect 21600 13756 23060 13784
rect 23124 13756 23388 13784
rect 21600 13744 21606 13756
rect 19024 13688 20576 13716
rect 19024 13676 19030 13688
rect 22462 13676 22468 13728
rect 22520 13676 22526 13728
rect 23032 13716 23060 13756
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 23676 13784 23704 13824
rect 23750 13812 23756 13864
rect 23808 13852 23814 13864
rect 24397 13855 24455 13861
rect 24397 13852 24409 13855
rect 23808 13824 24409 13852
rect 23808 13812 23814 13824
rect 24397 13821 24409 13824
rect 24443 13821 24455 13855
rect 24397 13815 24455 13821
rect 24670 13812 24676 13864
rect 24728 13812 24734 13864
rect 25222 13812 25228 13864
rect 25280 13852 25286 13864
rect 25884 13861 25912 13892
rect 26142 13880 26148 13892
rect 26200 13880 26206 13932
rect 26418 13880 26424 13932
rect 26476 13880 26482 13932
rect 27356 13929 27384 13960
rect 27341 13923 27399 13929
rect 27341 13889 27353 13923
rect 27387 13920 27399 13923
rect 28537 13923 28595 13929
rect 27387 13892 27568 13920
rect 27387 13889 27399 13892
rect 27341 13883 27399 13889
rect 25869 13855 25927 13861
rect 25869 13852 25881 13855
rect 25280 13824 25881 13852
rect 25280 13812 25286 13824
rect 25869 13821 25881 13824
rect 25915 13821 25927 13855
rect 25869 13815 25927 13821
rect 26053 13855 26111 13861
rect 26053 13821 26065 13855
rect 26099 13821 26111 13855
rect 26053 13815 26111 13821
rect 27433 13855 27491 13861
rect 27433 13821 27445 13855
rect 27479 13821 27491 13855
rect 27540 13852 27568 13892
rect 28537 13889 28549 13923
rect 28583 13920 28595 13923
rect 29178 13920 29184 13932
rect 28583 13892 29184 13920
rect 28583 13889 28595 13892
rect 28537 13883 28595 13889
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 29288 13920 29316 14016
rect 29816 13991 29874 13997
rect 29816 13957 29828 13991
rect 29862 13988 29874 13991
rect 30576 13988 30604 14016
rect 36909 13991 36967 13997
rect 36909 13988 36921 13991
rect 29862 13960 30604 13988
rect 35268 13960 36921 13988
rect 29862 13957 29874 13960
rect 29816 13951 29874 13957
rect 29549 13923 29607 13929
rect 29549 13920 29561 13923
rect 29288 13892 29561 13920
rect 29549 13889 29561 13892
rect 29595 13889 29607 13923
rect 29549 13883 29607 13889
rect 30742 13880 30748 13932
rect 30800 13920 30806 13932
rect 30800 13892 31156 13920
rect 30800 13880 30806 13892
rect 28721 13855 28779 13861
rect 28721 13852 28733 13855
rect 27540 13824 28733 13852
rect 27433 13815 27491 13821
rect 28721 13821 28733 13824
rect 28767 13821 28779 13855
rect 31021 13855 31079 13861
rect 31021 13852 31033 13855
rect 28721 13815 28779 13821
rect 30944 13824 31033 13852
rect 23842 13784 23848 13796
rect 23676 13756 23848 13784
rect 23842 13744 23848 13756
rect 23900 13744 23906 13796
rect 24121 13787 24179 13793
rect 24121 13753 24133 13787
rect 24167 13784 24179 13787
rect 24210 13784 24216 13796
rect 24167 13756 24216 13784
rect 24167 13753 24179 13756
rect 24121 13747 24179 13753
rect 24210 13744 24216 13756
rect 24268 13744 24274 13796
rect 25958 13784 25964 13796
rect 25240 13756 25964 13784
rect 25240 13716 25268 13756
rect 25958 13744 25964 13756
rect 26016 13784 26022 13796
rect 26068 13784 26096 13815
rect 26016 13756 26096 13784
rect 27448 13784 27476 13815
rect 30944 13796 30972 13824
rect 31021 13821 31033 13824
rect 31067 13821 31079 13855
rect 31021 13815 31079 13821
rect 28166 13784 28172 13796
rect 27448 13756 28172 13784
rect 26016 13744 26022 13756
rect 28166 13744 28172 13756
rect 28224 13744 28230 13796
rect 30926 13744 30932 13796
rect 30984 13744 30990 13796
rect 23032 13688 25268 13716
rect 25314 13676 25320 13728
rect 25372 13676 25378 13728
rect 25406 13676 25412 13728
rect 25464 13676 25470 13728
rect 28074 13676 28080 13728
rect 28132 13676 28138 13728
rect 29362 13676 29368 13728
rect 29420 13716 29426 13728
rect 30650 13716 30656 13728
rect 29420 13688 30656 13716
rect 29420 13676 29426 13688
rect 30650 13676 30656 13688
rect 30708 13676 30714 13728
rect 31128 13716 31156 13892
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32585 13923 32643 13929
rect 32585 13920 32597 13923
rect 31720 13892 32597 13920
rect 31720 13880 31726 13892
rect 32585 13889 32597 13892
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 32852 13923 32910 13929
rect 32852 13889 32864 13923
rect 32898 13920 32910 13923
rect 34701 13923 34759 13929
rect 34701 13920 34713 13923
rect 32898 13892 34713 13920
rect 32898 13889 32910 13892
rect 32852 13883 32910 13889
rect 34701 13889 34713 13892
rect 34747 13889 34759 13923
rect 34701 13883 34759 13889
rect 35268 13864 35296 13960
rect 36909 13957 36921 13960
rect 36955 13988 36967 13991
rect 37458 13988 37464 14000
rect 36955 13960 37464 13988
rect 36955 13957 36967 13960
rect 36909 13951 36967 13957
rect 37458 13948 37464 13960
rect 37516 13988 37522 14000
rect 38286 13988 38292 14000
rect 37516 13960 38292 13988
rect 37516 13948 37522 13960
rect 38286 13948 38292 13960
rect 38344 13988 38350 14000
rect 38344 13960 38516 13988
rect 38344 13948 38350 13960
rect 35520 13923 35578 13929
rect 35520 13889 35532 13923
rect 35566 13920 35578 13923
rect 36262 13920 36268 13932
rect 35566 13892 36268 13920
rect 35566 13889 35578 13892
rect 35520 13883 35578 13889
rect 36262 13880 36268 13892
rect 36320 13880 36326 13932
rect 37642 13880 37648 13932
rect 37700 13880 37706 13932
rect 38488 13929 38516 13960
rect 38473 13923 38531 13929
rect 38473 13889 38485 13923
rect 38519 13889 38531 13923
rect 38473 13883 38531 13889
rect 38740 13923 38798 13929
rect 38740 13889 38752 13923
rect 38786 13920 38798 13923
rect 39942 13920 39948 13932
rect 38786 13892 39948 13920
rect 38786 13889 38798 13892
rect 38740 13883 38798 13889
rect 34054 13812 34060 13864
rect 34112 13812 34118 13864
rect 34606 13812 34612 13864
rect 34664 13852 34670 13864
rect 35250 13852 35256 13864
rect 34664 13824 35256 13852
rect 34664 13812 34670 13824
rect 35250 13812 35256 13824
rect 35308 13812 35314 13864
rect 37826 13812 37832 13864
rect 37884 13852 37890 13864
rect 38289 13855 38347 13861
rect 38289 13852 38301 13855
rect 37884 13824 38301 13852
rect 37884 13812 37890 13824
rect 38289 13821 38301 13824
rect 38335 13852 38347 13855
rect 38378 13852 38384 13864
rect 38335 13824 38384 13852
rect 38335 13821 38347 13824
rect 38289 13815 38347 13821
rect 38378 13812 38384 13824
rect 38436 13812 38442 13864
rect 31570 13716 31576 13728
rect 31128 13688 31576 13716
rect 31570 13676 31576 13688
rect 31628 13716 31634 13728
rect 32401 13719 32459 13725
rect 32401 13716 32413 13719
rect 31628 13688 32413 13716
rect 31628 13676 31634 13688
rect 32401 13685 32413 13688
rect 32447 13716 32459 13719
rect 33318 13716 33324 13728
rect 32447 13688 33324 13716
rect 32447 13685 32459 13688
rect 32401 13679 32459 13685
rect 33318 13676 33324 13688
rect 33376 13676 33382 13728
rect 36170 13676 36176 13728
rect 36228 13716 36234 13728
rect 36630 13716 36636 13728
rect 36228 13688 36636 13716
rect 36228 13676 36234 13688
rect 36630 13676 36636 13688
rect 36688 13676 36694 13728
rect 38488 13716 38516 13883
rect 39942 13880 39948 13892
rect 40000 13880 40006 13932
rect 40218 13812 40224 13864
rect 40276 13852 40282 13864
rect 40328 13852 40356 14028
rect 40420 14028 42064 14056
rect 40420 13929 40448 14028
rect 42058 14016 42064 14028
rect 42116 14016 42122 14068
rect 42150 14016 42156 14068
rect 42208 14016 42214 14068
rect 42245 14059 42303 14065
rect 42245 14025 42257 14059
rect 42291 14056 42303 14059
rect 42794 14056 42800 14068
rect 42291 14028 42800 14056
rect 42291 14025 42303 14028
rect 42245 14019 42303 14025
rect 42794 14016 42800 14028
rect 42852 14016 42858 14068
rect 44174 14016 44180 14068
rect 44232 14016 44238 14068
rect 45646 14016 45652 14068
rect 45704 14056 45710 14068
rect 46290 14056 46296 14068
rect 45704 14028 46296 14056
rect 45704 14016 45710 14028
rect 46290 14016 46296 14028
rect 46348 14016 46354 14068
rect 48222 14016 48228 14068
rect 48280 14016 48286 14068
rect 48774 14016 48780 14068
rect 48832 14056 48838 14068
rect 49697 14059 49755 14065
rect 49697 14056 49709 14059
rect 48832 14028 49709 14056
rect 48832 14016 48838 14028
rect 49697 14025 49709 14028
rect 49743 14025 49755 14059
rect 49697 14019 49755 14025
rect 50246 14016 50252 14068
rect 50304 14016 50310 14068
rect 51626 14016 51632 14068
rect 51684 14016 51690 14068
rect 51994 14016 52000 14068
rect 52052 14056 52058 14068
rect 53282 14056 53288 14068
rect 52052 14028 53288 14056
rect 52052 14016 52058 14028
rect 53282 14016 53288 14028
rect 53340 14016 53346 14068
rect 55306 14016 55312 14068
rect 55364 14016 55370 14068
rect 55398 14016 55404 14068
rect 55456 14016 55462 14068
rect 55766 14016 55772 14068
rect 55824 14056 55830 14068
rect 56137 14059 56195 14065
rect 56137 14056 56149 14059
rect 55824 14028 56149 14056
rect 55824 14016 55830 14028
rect 56137 14025 56149 14028
rect 56183 14025 56195 14059
rect 56870 14056 56876 14068
rect 56137 14019 56195 14025
rect 56704 14028 56876 14056
rect 40405 13923 40463 13929
rect 40405 13889 40417 13923
rect 40451 13889 40463 13923
rect 40405 13883 40463 13889
rect 40586 13880 40592 13932
rect 40644 13880 40650 13932
rect 42168 13920 42196 14016
rect 42696 13991 42754 13997
rect 42696 13957 42708 13991
rect 42742 13988 42754 13991
rect 44192 13988 44220 14016
rect 42742 13960 44220 13988
rect 46201 13991 46259 13997
rect 42742 13957 42754 13960
rect 42696 13951 42754 13957
rect 46201 13957 46213 13991
rect 46247 13988 46259 13991
rect 47305 13991 47363 13997
rect 47305 13988 47317 13991
rect 46247 13960 47317 13988
rect 46247 13957 46259 13960
rect 46201 13951 46259 13957
rect 47305 13957 47317 13960
rect 47351 13957 47363 13991
rect 48240 13988 48268 14016
rect 48240 13960 49096 13988
rect 47305 13951 47363 13957
rect 44628 13923 44686 13929
rect 42168 13892 43852 13920
rect 41325 13855 41383 13861
rect 41325 13852 41337 13855
rect 40276 13824 41337 13852
rect 40276 13812 40282 13824
rect 41325 13821 41337 13824
rect 41371 13821 41383 13855
rect 41325 13815 41383 13821
rect 41414 13812 41420 13864
rect 41472 13861 41478 13864
rect 41472 13855 41500 13861
rect 41488 13821 41500 13855
rect 41472 13815 41500 13821
rect 41472 13812 41478 13815
rect 41598 13812 41604 13864
rect 41656 13812 41662 13864
rect 42429 13855 42487 13861
rect 42429 13821 42441 13855
rect 42475 13821 42487 13855
rect 42429 13815 42487 13821
rect 41046 13744 41052 13796
rect 41104 13744 41110 13796
rect 42444 13728 42472 13815
rect 43824 13793 43852 13892
rect 44628 13889 44640 13923
rect 44674 13920 44686 13923
rect 45922 13920 45928 13932
rect 44674 13892 45928 13920
rect 44674 13889 44686 13892
rect 44628 13883 44686 13889
rect 45922 13880 45928 13892
rect 45980 13880 45986 13932
rect 46753 13923 46811 13929
rect 46753 13889 46765 13923
rect 46799 13920 46811 13923
rect 47486 13920 47492 13932
rect 46799 13892 47492 13920
rect 46799 13889 46811 13892
rect 46753 13883 46811 13889
rect 44361 13855 44419 13861
rect 44361 13852 44373 13855
rect 44100 13824 44373 13852
rect 43809 13787 43867 13793
rect 43809 13753 43821 13787
rect 43855 13753 43867 13787
rect 43809 13747 43867 13753
rect 44100 13728 44128 13824
rect 44361 13821 44373 13824
rect 44407 13821 44419 13855
rect 44361 13815 44419 13821
rect 46290 13812 46296 13864
rect 46348 13852 46354 13864
rect 46385 13855 46443 13861
rect 46385 13852 46397 13855
rect 46348 13824 46397 13852
rect 46348 13812 46354 13824
rect 46385 13821 46397 13824
rect 46431 13821 46443 13855
rect 46385 13815 46443 13821
rect 45741 13787 45799 13793
rect 45741 13753 45753 13787
rect 45787 13784 45799 13787
rect 46400 13784 46428 13815
rect 46842 13784 46848 13796
rect 45787 13756 46336 13784
rect 46400 13756 46848 13784
rect 45787 13753 45799 13756
rect 45741 13747 45799 13753
rect 40221 13719 40279 13725
rect 40221 13716 40233 13719
rect 38488 13688 40233 13716
rect 40221 13685 40233 13688
rect 40267 13716 40279 13719
rect 40586 13716 40592 13728
rect 40267 13688 40592 13716
rect 40267 13685 40279 13688
rect 40221 13679 40279 13685
rect 40586 13676 40592 13688
rect 40644 13676 40650 13728
rect 42426 13676 42432 13728
rect 42484 13716 42490 13728
rect 43438 13716 43444 13728
rect 42484 13688 43444 13716
rect 42484 13676 42490 13688
rect 43438 13676 43444 13688
rect 43496 13716 43502 13728
rect 44082 13716 44088 13728
rect 43496 13688 44088 13716
rect 43496 13676 43502 13688
rect 44082 13676 44088 13688
rect 44140 13676 44146 13728
rect 45830 13676 45836 13728
rect 45888 13676 45894 13728
rect 46308 13716 46336 13756
rect 46842 13744 46848 13756
rect 46900 13744 46906 13796
rect 46952 13716 46980 13892
rect 47486 13880 47492 13892
rect 47544 13880 47550 13932
rect 47848 13923 47906 13929
rect 47848 13889 47860 13923
rect 47894 13920 47906 13923
rect 48774 13920 48780 13932
rect 47894 13892 48780 13920
rect 47894 13889 47906 13892
rect 47848 13883 47906 13889
rect 48774 13880 48780 13892
rect 48832 13880 48838 13932
rect 49068 13929 49096 13960
rect 50264 13929 50292 14016
rect 49053 13923 49111 13929
rect 49053 13920 49065 13923
rect 48976 13892 49065 13920
rect 47394 13812 47400 13864
rect 47452 13852 47458 13864
rect 47581 13855 47639 13861
rect 47581 13852 47593 13855
rect 47452 13824 47593 13852
rect 47452 13812 47458 13824
rect 47581 13821 47593 13824
rect 47627 13821 47639 13855
rect 47581 13815 47639 13821
rect 48976 13793 49004 13892
rect 49053 13889 49065 13892
rect 49099 13889 49111 13923
rect 49053 13883 49111 13889
rect 50249 13923 50307 13929
rect 50249 13889 50261 13923
rect 50295 13889 50307 13923
rect 50249 13883 50307 13889
rect 50516 13923 50574 13929
rect 50516 13889 50528 13923
rect 50562 13920 50574 13923
rect 51644 13920 51672 14016
rect 52086 13948 52092 14000
rect 52144 13988 52150 14000
rect 52144 13960 54064 13988
rect 52144 13948 52150 13960
rect 54036 13932 54064 13960
rect 51721 13923 51779 13929
rect 51721 13920 51733 13923
rect 50562 13892 51580 13920
rect 51644 13892 51733 13920
rect 50562 13889 50574 13892
rect 50516 13883 50574 13889
rect 51552 13852 51580 13892
rect 51721 13889 51733 13892
rect 51767 13889 51779 13923
rect 51721 13883 51779 13889
rect 52365 13923 52423 13929
rect 52365 13889 52377 13923
rect 52411 13889 52423 13923
rect 52365 13883 52423 13889
rect 52380 13852 52408 13883
rect 54018 13880 54024 13932
rect 54076 13880 54082 13932
rect 54849 13923 54907 13929
rect 54849 13889 54861 13923
rect 54895 13920 54907 13923
rect 55324 13920 55352 14016
rect 55950 13948 55956 14000
rect 56008 13948 56014 14000
rect 54895 13892 55352 13920
rect 55585 13923 55643 13929
rect 54895 13889 54907 13892
rect 54849 13883 54907 13889
rect 55585 13889 55597 13923
rect 55631 13920 55643 13923
rect 55968 13920 55996 13948
rect 55631 13892 55996 13920
rect 55631 13889 55643 13892
rect 55585 13883 55643 13889
rect 56704 13864 56732 14028
rect 56870 14016 56876 14028
rect 56928 14016 56934 14068
rect 56965 13923 57023 13929
rect 56965 13889 56977 13923
rect 57011 13920 57023 13923
rect 58529 13923 58587 13929
rect 58529 13920 58541 13923
rect 57011 13892 58541 13920
rect 57011 13889 57023 13892
rect 56965 13883 57023 13889
rect 58529 13889 58541 13892
rect 58575 13889 58587 13923
rect 58529 13883 58587 13889
rect 51552 13824 52408 13852
rect 53926 13812 53932 13864
rect 53984 13852 53990 13864
rect 54573 13855 54631 13861
rect 54573 13852 54585 13855
rect 53984 13824 54585 13852
rect 53984 13812 53990 13824
rect 54573 13821 54585 13824
rect 54619 13852 54631 13855
rect 54754 13852 54760 13864
rect 54619 13824 54760 13852
rect 54619 13821 54631 13824
rect 54573 13815 54631 13821
rect 54754 13812 54760 13824
rect 54812 13812 54818 13864
rect 55674 13812 55680 13864
rect 55732 13852 55738 13864
rect 56686 13852 56692 13864
rect 55732 13824 56692 13852
rect 55732 13812 55738 13824
rect 56686 13812 56692 13824
rect 56744 13812 56750 13864
rect 57057 13855 57115 13861
rect 57057 13821 57069 13855
rect 57103 13821 57115 13855
rect 57057 13815 57115 13821
rect 48961 13787 49019 13793
rect 48961 13753 48973 13787
rect 49007 13753 49019 13787
rect 48961 13747 49019 13753
rect 51629 13787 51687 13793
rect 51629 13753 51641 13787
rect 51675 13784 51687 13787
rect 51718 13784 51724 13796
rect 51675 13756 51724 13784
rect 51675 13753 51687 13756
rect 51629 13747 51687 13753
rect 51718 13744 51724 13756
rect 51776 13744 51782 13796
rect 57072 13784 57100 13815
rect 57330 13812 57336 13864
rect 57388 13852 57394 13864
rect 57517 13855 57575 13861
rect 57517 13852 57529 13855
rect 57388 13824 57529 13852
rect 57388 13812 57394 13824
rect 57517 13821 57529 13824
rect 57563 13821 57575 13855
rect 57517 13815 57575 13821
rect 57698 13812 57704 13864
rect 57756 13852 57762 13864
rect 57885 13855 57943 13861
rect 57885 13852 57897 13855
rect 57756 13824 57897 13852
rect 57756 13812 57762 13824
rect 57885 13821 57897 13824
rect 57931 13821 57943 13855
rect 57885 13815 57943 13821
rect 56336 13756 57100 13784
rect 56336 13728 56364 13756
rect 46308 13688 46980 13716
rect 56318 13676 56324 13728
rect 56376 13676 56382 13728
rect 56502 13676 56508 13728
rect 56560 13676 56566 13728
rect 1104 13626 58880 13648
rect 1104 13574 8172 13626
rect 8224 13574 8236 13626
rect 8288 13574 8300 13626
rect 8352 13574 8364 13626
rect 8416 13574 8428 13626
rect 8480 13574 22616 13626
rect 22668 13574 22680 13626
rect 22732 13574 22744 13626
rect 22796 13574 22808 13626
rect 22860 13574 22872 13626
rect 22924 13574 37060 13626
rect 37112 13574 37124 13626
rect 37176 13574 37188 13626
rect 37240 13574 37252 13626
rect 37304 13574 37316 13626
rect 37368 13574 51504 13626
rect 51556 13574 51568 13626
rect 51620 13574 51632 13626
rect 51684 13574 51696 13626
rect 51748 13574 51760 13626
rect 51812 13574 58880 13626
rect 1104 13552 58880 13574
rect 5902 13472 5908 13524
rect 5960 13472 5966 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6144 13484 6285 13512
rect 6144 13472 6150 13484
rect 6273 13481 6285 13484
rect 6319 13512 6331 13515
rect 7466 13512 7472 13524
rect 6319 13484 7472 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 11422 13512 11428 13524
rect 11164 13484 11428 13512
rect 3605 13447 3663 13453
rect 3605 13413 3617 13447
rect 3651 13413 3663 13447
rect 3605 13407 3663 13413
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 2004 13348 2237 13376
rect 2004 13336 2010 13348
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 3620 13376 3648 13407
rect 3789 13379 3847 13385
rect 3789 13376 3801 13379
rect 3620 13348 3801 13376
rect 2225 13339 2283 13345
rect 3789 13345 3801 13348
rect 3835 13345 3847 13379
rect 3789 13339 3847 13345
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 5442 13376 5448 13388
rect 5399 13348 5448 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 11164 13385 11192 13484
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 12618 13472 12624 13524
rect 12676 13472 12682 13524
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13412 13484 13645 13512
rect 13412 13472 13418 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 17957 13515 18015 13521
rect 17957 13481 17969 13515
rect 18003 13512 18015 13515
rect 18046 13512 18052 13524
rect 18003 13484 18052 13512
rect 18003 13481 18015 13484
rect 17957 13475 18015 13481
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 19978 13512 19984 13524
rect 19260 13484 19984 13512
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8628 13348 8953 13376
rect 8628 13336 8634 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 11149 13379 11207 13385
rect 11149 13345 11161 13379
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 13078 13336 13084 13388
rect 13136 13336 13142 13388
rect 13265 13379 13323 13385
rect 13265 13345 13277 13379
rect 13311 13376 13323 13379
rect 13372 13376 13400 13472
rect 13311 13348 13400 13376
rect 13311 13345 13323 13348
rect 13265 13339 13323 13345
rect 14090 13336 14096 13388
rect 14148 13336 14154 13388
rect 18414 13336 18420 13388
rect 18472 13336 18478 13388
rect 18598 13336 18604 13388
rect 18656 13376 18662 13388
rect 19058 13376 19064 13388
rect 18656 13348 19064 13376
rect 18656 13336 18662 13348
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 19150 13336 19156 13388
rect 19208 13336 19214 13388
rect 19260 13385 19288 13484
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 22370 13472 22376 13524
rect 22428 13512 22434 13524
rect 22925 13515 22983 13521
rect 22925 13512 22937 13515
rect 22428 13484 22937 13512
rect 22428 13472 22434 13484
rect 22925 13481 22937 13484
rect 22971 13481 22983 13515
rect 22925 13475 22983 13481
rect 23382 13472 23388 13524
rect 23440 13472 23446 13524
rect 23566 13472 23572 13524
rect 23624 13512 23630 13524
rect 23661 13515 23719 13521
rect 23661 13512 23673 13515
rect 23624 13484 23673 13512
rect 23624 13472 23630 13484
rect 23661 13481 23673 13484
rect 23707 13481 23719 13515
rect 23661 13475 23719 13481
rect 25774 13472 25780 13524
rect 25832 13472 25838 13524
rect 25958 13472 25964 13524
rect 26016 13512 26022 13524
rect 26053 13515 26111 13521
rect 26053 13512 26065 13515
rect 26016 13484 26065 13512
rect 26016 13472 26022 13484
rect 26053 13481 26065 13484
rect 26099 13512 26111 13515
rect 29362 13512 29368 13524
rect 26099 13484 29368 13512
rect 26099 13481 26111 13484
rect 26053 13475 26111 13481
rect 29362 13472 29368 13484
rect 29420 13472 29426 13524
rect 30926 13512 30932 13524
rect 29564 13484 30932 13512
rect 22189 13447 22247 13453
rect 19352 13416 20024 13444
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 2492 13243 2550 13249
rect 2492 13209 2504 13243
rect 2538 13240 2550 13243
rect 3326 13240 3332 13252
rect 2538 13212 3332 13240
rect 2538 13209 2550 13212
rect 2492 13203 2550 13209
rect 3326 13200 3332 13212
rect 3384 13200 3390 13252
rect 9208 13243 9266 13249
rect 9208 13209 9220 13243
rect 9254 13240 9266 13243
rect 9858 13240 9864 13252
rect 9254 13212 9864 13240
rect 9254 13209 9266 13212
rect 9208 13203 9266 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 10428 13240 10456 13271
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 13906 13308 13912 13320
rect 11296 13280 13912 13308
rect 11296 13268 11302 13280
rect 13906 13268 13912 13280
rect 13964 13308 13970 13320
rect 14182 13308 14188 13320
rect 13964 13280 14188 13308
rect 13964 13268 13970 13280
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14360 13311 14418 13317
rect 14360 13277 14372 13311
rect 14406 13308 14418 13311
rect 15746 13308 15752 13320
rect 14406 13280 15752 13308
rect 14406 13277 14418 13280
rect 14360 13271 14418 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16482 13268 16488 13320
rect 16540 13268 16546 13320
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 17828 13280 18337 13308
rect 17828 13268 17834 13280
rect 18325 13277 18337 13280
rect 18371 13308 18383 13311
rect 19168 13308 19196 13336
rect 18371 13280 19196 13308
rect 18371 13277 18383 13280
rect 18325 13271 18383 13277
rect 10336 13212 10456 13240
rect 11416 13243 11474 13249
rect 4062 13132 4068 13184
rect 4120 13172 4126 13184
rect 4433 13175 4491 13181
rect 4433 13172 4445 13175
rect 4120 13144 4445 13172
rect 4120 13132 4126 13144
rect 4433 13141 4445 13144
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 10336 13181 10364 13212
rect 11416 13209 11428 13243
rect 11462 13240 11474 13243
rect 12250 13240 12256 13252
rect 11462 13212 12256 13240
rect 11462 13209 11474 13212
rect 11416 13203 11474 13209
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12989 13243 13047 13249
rect 12989 13240 13001 13243
rect 12406 13212 13001 13240
rect 10321 13175 10379 13181
rect 10321 13172 10333 13175
rect 9640 13144 10333 13172
rect 9640 13132 9646 13144
rect 10321 13141 10333 13144
rect 10367 13141 10379 13175
rect 10321 13135 10379 13141
rect 11054 13132 11060 13184
rect 11112 13132 11118 13184
rect 12158 13132 12164 13184
rect 12216 13172 12222 13184
rect 12406 13172 12434 13212
rect 12989 13209 13001 13212
rect 13035 13240 13047 13243
rect 14458 13240 14464 13252
rect 13035 13212 14464 13240
rect 13035 13209 13047 13212
rect 12989 13203 13047 13209
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 16752 13243 16810 13249
rect 16752 13209 16764 13243
rect 16798 13240 16810 13243
rect 17586 13240 17592 13252
rect 16798 13212 17592 13240
rect 16798 13209 16810 13212
rect 16752 13203 16810 13209
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 19352 13240 19380 13416
rect 19886 13336 19892 13388
rect 19944 13336 19950 13388
rect 19996 13376 20024 13416
rect 22189 13413 22201 13447
rect 22235 13444 22247 13447
rect 23400 13444 23428 13472
rect 22235 13416 23428 13444
rect 22235 13413 22247 13416
rect 22189 13407 22247 13413
rect 20282 13379 20340 13385
rect 20282 13376 20294 13379
rect 19996 13348 20294 13376
rect 20282 13345 20294 13348
rect 20328 13345 20340 13379
rect 20282 13339 20340 13345
rect 20438 13336 20444 13388
rect 20496 13336 20502 13388
rect 22373 13379 22431 13385
rect 22373 13345 22385 13379
rect 22419 13376 22431 13379
rect 22462 13376 22468 13388
rect 22419 13348 22468 13376
rect 22419 13345 22431 13348
rect 22373 13339 22431 13345
rect 22462 13336 22468 13348
rect 22520 13336 22526 13388
rect 23106 13336 23112 13388
rect 23164 13336 23170 13388
rect 25225 13379 25283 13385
rect 25225 13345 25237 13379
rect 25271 13376 25283 13379
rect 25406 13376 25412 13388
rect 25271 13348 25412 13376
rect 25271 13345 25283 13348
rect 25225 13339 25283 13345
rect 25406 13336 25412 13348
rect 25464 13336 25470 13388
rect 29564 13385 29592 13484
rect 30926 13472 30932 13484
rect 30984 13472 30990 13524
rect 37550 13512 37556 13524
rect 34900 13484 37556 13512
rect 31846 13444 31852 13456
rect 31312 13416 31852 13444
rect 29549 13379 29607 13385
rect 29549 13345 29561 13379
rect 29595 13345 29607 13379
rect 29549 13339 29607 13345
rect 30193 13379 30251 13385
rect 30193 13345 30205 13379
rect 30239 13376 30251 13379
rect 31312 13376 31340 13416
rect 31846 13404 31852 13416
rect 31904 13404 31910 13456
rect 30239 13348 31340 13376
rect 30239 13345 30251 13348
rect 30193 13339 30251 13345
rect 31386 13336 31392 13388
rect 31444 13376 31450 13388
rect 34900 13385 34928 13484
rect 37550 13472 37556 13484
rect 37608 13472 37614 13524
rect 38102 13472 38108 13524
rect 38160 13472 38166 13524
rect 39669 13515 39727 13521
rect 39669 13481 39681 13515
rect 39715 13512 39727 13515
rect 40678 13512 40684 13524
rect 39715 13484 40684 13512
rect 39715 13481 39727 13484
rect 39669 13475 39727 13481
rect 40678 13472 40684 13484
rect 40736 13512 40742 13524
rect 41322 13512 41328 13524
rect 40736 13484 41328 13512
rect 40736 13472 40742 13484
rect 41322 13472 41328 13484
rect 41380 13472 41386 13524
rect 42058 13472 42064 13524
rect 42116 13472 42122 13524
rect 45922 13472 45928 13524
rect 45980 13472 45986 13524
rect 46290 13472 46296 13524
rect 46348 13472 46354 13524
rect 48774 13472 48780 13524
rect 48832 13472 48838 13524
rect 49142 13472 49148 13524
rect 49200 13472 49206 13524
rect 51537 13515 51595 13521
rect 51537 13512 51549 13515
rect 51046 13484 51549 13512
rect 36633 13447 36691 13453
rect 36633 13413 36645 13447
rect 36679 13444 36691 13447
rect 47670 13444 47676 13456
rect 36679 13416 37504 13444
rect 36679 13413 36691 13416
rect 36633 13407 36691 13413
rect 32033 13379 32091 13385
rect 32033 13376 32045 13379
rect 31444 13348 32045 13376
rect 31444 13336 31450 13348
rect 32033 13345 32045 13348
rect 32079 13345 32091 13379
rect 32033 13339 32091 13345
rect 34885 13379 34943 13385
rect 34885 13345 34897 13379
rect 34931 13345 34943 13379
rect 34885 13339 34943 13345
rect 35066 13336 35072 13388
rect 35124 13376 35130 13388
rect 35345 13379 35403 13385
rect 35345 13376 35357 13379
rect 35124 13348 35357 13376
rect 35124 13336 35130 13348
rect 35345 13345 35357 13348
rect 35391 13345 35403 13379
rect 35345 13339 35403 13345
rect 35618 13336 35624 13388
rect 35676 13336 35682 13388
rect 35710 13336 35716 13388
rect 35768 13385 35774 13388
rect 35768 13379 35817 13385
rect 35768 13345 35771 13379
rect 35805 13345 35817 13379
rect 35768 13339 35817 13345
rect 35895 13379 35953 13385
rect 35895 13345 35907 13379
rect 35941 13376 35953 13379
rect 36078 13376 36084 13388
rect 35941 13348 36084 13376
rect 35941 13345 35953 13348
rect 35895 13339 35953 13345
rect 35768 13336 35774 13339
rect 36078 13336 36084 13348
rect 36136 13336 36142 13388
rect 36722 13336 36728 13388
rect 36780 13376 36786 13388
rect 37476 13385 37504 13416
rect 47504 13416 47676 13444
rect 37185 13379 37243 13385
rect 37185 13376 37197 13379
rect 36780 13348 37197 13376
rect 36780 13336 36786 13348
rect 37185 13345 37197 13348
rect 37231 13345 37243 13379
rect 37185 13339 37243 13345
rect 37461 13379 37519 13385
rect 37461 13345 37473 13379
rect 37507 13345 37519 13379
rect 37461 13339 37519 13345
rect 37642 13336 37648 13388
rect 37700 13336 37706 13388
rect 38286 13336 38292 13388
rect 38344 13336 38350 13388
rect 40405 13379 40463 13385
rect 40405 13376 40417 13379
rect 39776 13348 40417 13376
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 17880 13212 19380 13240
rect 17880 13184 17908 13212
rect 19444 13184 19472 13271
rect 20162 13268 20168 13320
rect 20220 13268 20226 13320
rect 27433 13311 27491 13317
rect 27433 13308 27445 13311
rect 27264 13280 27445 13308
rect 24118 13240 24124 13252
rect 23952 13212 24124 13240
rect 12216 13144 12434 13172
rect 12216 13132 12222 13144
rect 12526 13132 12532 13184
rect 12584 13132 12590 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 14090 13172 14096 13184
rect 13412 13144 14096 13172
rect 13412 13132 13418 13144
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14332 13144 15485 13172
rect 14332 13132 14338 13144
rect 15473 13141 15485 13144
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 17862 13132 17868 13184
rect 17920 13132 17926 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18966 13172 18972 13184
rect 18104 13144 18972 13172
rect 18104 13132 18110 13144
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 19426 13132 19432 13184
rect 19484 13132 19490 13184
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 20772 13144 21097 13172
rect 20772 13132 20778 13144
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21085 13135 21143 13141
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 23952 13181 23980 13212
rect 24118 13200 24124 13212
rect 24176 13240 24182 13252
rect 24670 13240 24676 13252
rect 24176 13212 24676 13240
rect 24176 13200 24182 13212
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 27264 13184 27292 13280
rect 27433 13277 27445 13280
rect 27479 13277 27491 13311
rect 27433 13271 27491 13277
rect 27700 13311 27758 13317
rect 27700 13277 27712 13311
rect 27746 13308 27758 13311
rect 28626 13308 28632 13320
rect 27746 13280 28632 13308
rect 27746 13277 27758 13280
rect 27700 13271 27758 13277
rect 28626 13268 28632 13280
rect 28684 13268 28690 13320
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13277 29791 13311
rect 29733 13271 29791 13277
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 22244 13144 23949 13172
rect 22244 13132 22250 13144
rect 23937 13141 23949 13144
rect 23983 13141 23995 13175
rect 23937 13135 23995 13141
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24544 13144 24593 13172
rect 24544 13132 24550 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 27246 13132 27252 13184
rect 27304 13132 27310 13184
rect 28810 13132 28816 13184
rect 28868 13132 28874 13184
rect 29748 13172 29776 13271
rect 30466 13268 30472 13320
rect 30524 13268 30530 13320
rect 30558 13268 30564 13320
rect 30616 13317 30622 13320
rect 30616 13311 30644 13317
rect 30632 13277 30644 13311
rect 30616 13271 30644 13277
rect 30616 13268 30622 13271
rect 30742 13268 30748 13320
rect 30800 13268 30806 13320
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 32493 13311 32551 13317
rect 32493 13308 32505 13311
rect 32364 13280 32505 13308
rect 32364 13268 32370 13280
rect 32493 13277 32505 13280
rect 32539 13308 32551 13311
rect 34149 13311 34207 13317
rect 34149 13308 34161 13311
rect 32539 13280 34161 13308
rect 32539 13277 32551 13280
rect 32493 13271 32551 13277
rect 34149 13277 34161 13280
rect 34195 13308 34207 13311
rect 34606 13308 34612 13320
rect 34195 13280 34612 13308
rect 34195 13277 34207 13280
rect 34149 13271 34207 13277
rect 34606 13268 34612 13280
rect 34664 13268 34670 13320
rect 34701 13311 34759 13317
rect 34701 13277 34713 13311
rect 34747 13277 34759 13311
rect 34701 13271 34759 13277
rect 31389 13243 31447 13249
rect 31389 13209 31401 13243
rect 31435 13240 31447 13243
rect 31662 13240 31668 13252
rect 31435 13212 31668 13240
rect 31435 13209 31447 13212
rect 31389 13203 31447 13209
rect 31662 13200 31668 13212
rect 31720 13200 31726 13252
rect 32760 13243 32818 13249
rect 31772 13212 31984 13240
rect 30742 13172 30748 13184
rect 29748 13144 30748 13172
rect 30742 13132 30748 13144
rect 30800 13132 30806 13184
rect 31478 13132 31484 13184
rect 31536 13132 31542 13184
rect 31570 13132 31576 13184
rect 31628 13172 31634 13184
rect 31772 13172 31800 13212
rect 31628 13144 31800 13172
rect 31628 13132 31634 13144
rect 31846 13132 31852 13184
rect 31904 13132 31910 13184
rect 31956 13181 31984 13212
rect 32760 13209 32772 13243
rect 32806 13240 32818 13243
rect 33594 13240 33600 13252
rect 32806 13212 33600 13240
rect 32806 13209 32818 13212
rect 32760 13203 32818 13209
rect 33594 13200 33600 13212
rect 33652 13200 33658 13252
rect 31941 13175 31999 13181
rect 31941 13141 31953 13175
rect 31987 13141 31999 13175
rect 31941 13135 31999 13141
rect 33870 13132 33876 13184
rect 33928 13132 33934 13184
rect 34716 13172 34744 13271
rect 36814 13268 36820 13320
rect 36872 13308 36878 13320
rect 37093 13311 37151 13317
rect 37093 13308 37105 13311
rect 36872 13280 37105 13308
rect 36872 13268 36878 13280
rect 37093 13277 37105 13280
rect 37139 13308 37151 13311
rect 37660 13308 37688 13336
rect 37139 13280 37688 13308
rect 38556 13311 38614 13317
rect 37139 13277 37151 13280
rect 37093 13271 37151 13277
rect 38556 13277 38568 13311
rect 38602 13308 38614 13311
rect 39666 13308 39672 13320
rect 38602 13280 39672 13308
rect 38602 13277 38614 13280
rect 38556 13271 38614 13277
rect 39666 13268 39672 13280
rect 39724 13268 39730 13320
rect 39776 13240 39804 13348
rect 40405 13345 40417 13348
rect 40451 13345 40463 13379
rect 40405 13339 40463 13345
rect 40420 13308 40448 13339
rect 40678 13336 40684 13388
rect 40736 13336 40742 13388
rect 44910 13376 44916 13388
rect 41800 13348 44916 13376
rect 41800 13308 41828 13348
rect 44910 13336 44916 13348
rect 44968 13336 44974 13388
rect 45373 13379 45431 13385
rect 45373 13345 45385 13379
rect 45419 13376 45431 13379
rect 45830 13376 45836 13388
rect 45419 13348 45836 13376
rect 45419 13345 45431 13348
rect 45373 13339 45431 13345
rect 45830 13336 45836 13348
rect 45888 13336 45894 13388
rect 47210 13336 47216 13388
rect 47268 13376 47274 13388
rect 47504 13376 47532 13416
rect 47670 13404 47676 13416
rect 47728 13444 47734 13456
rect 51046 13444 51074 13484
rect 51537 13481 51549 13484
rect 51583 13512 51595 13515
rect 52178 13512 52184 13524
rect 51583 13484 52184 13512
rect 51583 13481 51595 13484
rect 51537 13475 51595 13481
rect 52178 13472 52184 13484
rect 52236 13472 52242 13524
rect 57146 13472 57152 13524
rect 57204 13472 57210 13524
rect 47728 13416 51074 13444
rect 47728 13404 47734 13416
rect 47268 13348 47532 13376
rect 48225 13379 48283 13385
rect 47268 13336 47274 13348
rect 48225 13345 48237 13379
rect 48271 13376 48283 13379
rect 48406 13376 48412 13388
rect 48271 13348 48412 13376
rect 48271 13345 48283 13348
rect 48225 13339 48283 13345
rect 48406 13336 48412 13348
rect 48464 13336 48470 13388
rect 56502 13336 56508 13388
rect 56560 13336 56566 13388
rect 40420 13280 41828 13308
rect 41874 13268 41880 13320
rect 41932 13308 41938 13320
rect 42153 13311 42211 13317
rect 42153 13308 42165 13311
rect 41932 13280 42165 13308
rect 41932 13268 41938 13280
rect 42153 13277 42165 13280
rect 42199 13277 42211 13311
rect 42153 13271 42211 13277
rect 39132 13212 39804 13240
rect 40948 13243 41006 13249
rect 39132 13184 39160 13212
rect 40948 13209 40960 13243
rect 40994 13240 41006 13243
rect 41690 13240 41696 13252
rect 40994 13212 41696 13240
rect 40994 13209 41006 13212
rect 40948 13203 41006 13209
rect 41690 13200 41696 13212
rect 41748 13200 41754 13252
rect 43901 13243 43959 13249
rect 43901 13209 43913 13243
rect 43947 13240 43959 13243
rect 44082 13240 44088 13252
rect 43947 13212 44088 13240
rect 43947 13209 43959 13212
rect 43901 13203 43959 13209
rect 44082 13200 44088 13212
rect 44140 13240 44146 13252
rect 44140 13212 44220 13240
rect 44140 13200 44146 13212
rect 36170 13172 36176 13184
rect 34716 13144 36176 13172
rect 36170 13132 36176 13144
rect 36228 13132 36234 13184
rect 36538 13132 36544 13184
rect 36596 13132 36602 13184
rect 36998 13132 37004 13184
rect 37056 13132 37062 13184
rect 39114 13132 39120 13184
rect 39172 13132 39178 13184
rect 39850 13132 39856 13184
rect 39908 13132 39914 13184
rect 40126 13132 40132 13184
rect 40184 13172 40190 13184
rect 40221 13175 40279 13181
rect 40221 13172 40233 13175
rect 40184 13144 40233 13172
rect 40184 13132 40190 13144
rect 40221 13141 40233 13144
rect 40267 13141 40279 13175
rect 40221 13135 40279 13141
rect 40310 13132 40316 13184
rect 40368 13132 40374 13184
rect 44192 13181 44220 13212
rect 44177 13175 44235 13181
rect 44177 13141 44189 13175
rect 44223 13172 44235 13175
rect 44726 13172 44732 13184
rect 44223 13144 44732 13172
rect 44223 13141 44235 13144
rect 44177 13135 44235 13141
rect 44726 13132 44732 13144
rect 44784 13172 44790 13184
rect 47394 13172 47400 13184
rect 44784 13144 47400 13172
rect 44784 13132 44790 13144
rect 47394 13132 47400 13144
rect 47452 13132 47458 13184
rect 55674 13132 55680 13184
rect 55732 13172 55738 13184
rect 56318 13172 56324 13184
rect 55732 13144 56324 13172
rect 55732 13132 55738 13144
rect 56318 13132 56324 13144
rect 56376 13132 56382 13184
rect 1104 13082 59040 13104
rect 1104 13030 15394 13082
rect 15446 13030 15458 13082
rect 15510 13030 15522 13082
rect 15574 13030 15586 13082
rect 15638 13030 15650 13082
rect 15702 13030 29838 13082
rect 29890 13030 29902 13082
rect 29954 13030 29966 13082
rect 30018 13030 30030 13082
rect 30082 13030 30094 13082
rect 30146 13030 44282 13082
rect 44334 13030 44346 13082
rect 44398 13030 44410 13082
rect 44462 13030 44474 13082
rect 44526 13030 44538 13082
rect 44590 13030 58726 13082
rect 58778 13030 58790 13082
rect 58842 13030 58854 13082
rect 58906 13030 58918 13082
rect 58970 13030 58982 13082
rect 59034 13030 59040 13082
rect 1104 13008 59040 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 2222 12968 2228 12980
rect 2179 12940 2228 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 3326 12928 3332 12980
rect 3384 12928 3390 12980
rect 3970 12968 3976 12980
rect 3528 12940 3976 12968
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 3528 12900 3556 12940
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 8754 12968 8760 12980
rect 6880 12940 8760 12968
rect 6880 12928 6886 12940
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9214 12928 9220 12980
rect 9272 12928 9278 12980
rect 9585 12971 9643 12977
rect 9585 12937 9597 12971
rect 9631 12968 9643 12971
rect 11054 12968 11060 12980
rect 9631 12940 11060 12968
rect 9631 12937 9643 12940
rect 9585 12931 9643 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11238 12928 11244 12980
rect 11296 12928 11302 12980
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 12710 12968 12716 12980
rect 11379 12940 12716 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 2547 12872 3556 12900
rect 3697 12903 3755 12909
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 3697 12869 3709 12903
rect 3743 12900 3755 12903
rect 4062 12900 4068 12912
rect 3743 12872 4068 12900
rect 3743 12869 3755 12872
rect 3697 12863 3755 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 7837 12903 7895 12909
rect 7837 12900 7849 12903
rect 7708 12872 7849 12900
rect 7708 12860 7714 12872
rect 7837 12869 7849 12872
rect 7883 12869 7895 12903
rect 7837 12863 7895 12869
rect 10321 12903 10379 12909
rect 10321 12869 10333 12903
rect 10367 12900 10379 12903
rect 11256 12900 11284 12928
rect 10367 12872 11284 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2332 12628 2360 12795
rect 2608 12696 2636 12795
rect 3050 12792 3056 12844
rect 3108 12832 3114 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3108 12804 3433 12832
rect 3108 12792 3114 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3602 12792 3608 12844
rect 3660 12792 3666 12844
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 2823 12736 4016 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3418 12696 3424 12708
rect 2608 12668 3424 12696
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 3988 12705 4016 12736
rect 7006 12724 7012 12776
rect 7064 12724 7070 12776
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9398 12764 9404 12776
rect 8720 12736 9404 12764
rect 8720 12724 8726 12736
rect 9398 12724 9404 12736
rect 9456 12764 9462 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 9456 12736 9689 12764
rect 9456 12724 9462 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 10336 12764 10364 12863
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 9907 12736 10364 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12665 4031 12699
rect 12084 12696 12112 12795
rect 12158 12724 12164 12776
rect 12216 12724 12222 12776
rect 12268 12773 12296 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 14274 12968 14280 12980
rect 12820 12940 14280 12968
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12820 12773 12848 12940
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 14516 12940 15209 12968
rect 14516 12928 14522 12940
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 15197 12931 15255 12937
rect 17589 12971 17647 12977
rect 17589 12937 17601 12971
rect 17635 12968 17647 12971
rect 17770 12968 17776 12980
rect 17635 12940 17776 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18598 12928 18604 12980
rect 18656 12928 18662 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 20990 12968 20996 12980
rect 19484 12940 20996 12968
rect 19484 12928 19490 12940
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 23293 12971 23351 12977
rect 23293 12937 23305 12971
rect 23339 12968 23351 12971
rect 23934 12968 23940 12980
rect 23339 12940 23940 12968
rect 23339 12937 23351 12940
rect 23293 12931 23351 12937
rect 23934 12928 23940 12940
rect 23992 12968 23998 12980
rect 24210 12968 24216 12980
rect 23992 12940 24216 12968
rect 23992 12928 23998 12940
rect 24210 12928 24216 12940
rect 24268 12928 24274 12980
rect 24765 12971 24823 12977
rect 24765 12937 24777 12971
rect 24811 12968 24823 12971
rect 25314 12968 25320 12980
rect 24811 12940 25320 12968
rect 24811 12937 24823 12940
rect 24765 12931 24823 12937
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 28166 12928 28172 12980
rect 28224 12968 28230 12980
rect 28721 12971 28779 12977
rect 28721 12968 28733 12971
rect 28224 12940 28733 12968
rect 28224 12928 28230 12940
rect 28721 12937 28733 12940
rect 28767 12937 28779 12971
rect 28721 12931 28779 12937
rect 28810 12928 28816 12980
rect 28868 12968 28874 12980
rect 30466 12968 30472 12980
rect 28868 12940 30472 12968
rect 28868 12928 28874 12940
rect 30466 12928 30472 12940
rect 30524 12928 30530 12980
rect 30558 12928 30564 12980
rect 30616 12928 30622 12980
rect 31478 12928 31484 12980
rect 31536 12928 31542 12980
rect 33965 12971 34023 12977
rect 33965 12937 33977 12971
rect 34011 12968 34023 12971
rect 34054 12968 34060 12980
rect 34011 12940 34060 12968
rect 34011 12937 34023 12940
rect 33965 12931 34023 12937
rect 34054 12928 34060 12940
rect 34112 12928 34118 12980
rect 34425 12971 34483 12977
rect 34425 12937 34437 12971
rect 34471 12968 34483 12971
rect 35342 12968 35348 12980
rect 34471 12940 35348 12968
rect 34471 12937 34483 12940
rect 34425 12931 34483 12937
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 36998 12928 37004 12980
rect 37056 12968 37062 12980
rect 37093 12971 37151 12977
rect 37093 12968 37105 12971
rect 37056 12940 37105 12968
rect 37056 12928 37062 12940
rect 37093 12937 37105 12940
rect 37139 12937 37151 12971
rect 39850 12968 39856 12980
rect 37093 12931 37151 12937
rect 39408 12940 39856 12968
rect 17037 12903 17095 12909
rect 17037 12869 17049 12903
rect 17083 12900 17095 12903
rect 18616 12900 18644 12928
rect 17083 12872 18644 12900
rect 19880 12903 19938 12909
rect 17083 12869 17095 12872
rect 17037 12863 17095 12869
rect 19880 12869 19892 12903
rect 19926 12900 19938 12903
rect 21450 12900 21456 12912
rect 19926 12872 21456 12900
rect 19926 12869 19938 12872
rect 19880 12863 19938 12869
rect 21450 12860 21456 12872
rect 21508 12860 21514 12912
rect 23106 12860 23112 12912
rect 23164 12900 23170 12912
rect 23382 12900 23388 12912
rect 23164 12872 23388 12900
rect 23164 12860 23170 12872
rect 23382 12860 23388 12872
rect 23440 12900 23446 12912
rect 26326 12900 26332 12912
rect 23440 12872 26332 12900
rect 23440 12860 23446 12872
rect 26326 12860 26332 12872
rect 26384 12860 26390 12912
rect 27516 12903 27574 12909
rect 27516 12869 27528 12903
rect 27562 12900 27574 12903
rect 28074 12900 28080 12912
rect 27562 12872 28080 12900
rect 27562 12869 27574 12872
rect 27516 12863 27574 12869
rect 28074 12860 28080 12872
rect 28132 12860 28138 12912
rect 12912 12804 13124 12832
rect 12805 12767 12863 12773
rect 12492 12736 12756 12764
rect 12492 12724 12498 12736
rect 12526 12696 12532 12708
rect 12084 12668 12532 12696
rect 3973 12659 4031 12665
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12728 12696 12756 12736
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12912 12696 12940 12804
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 13096 12764 13124 12804
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 13998 12792 14004 12844
rect 14056 12792 14062 12844
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 15151 12804 16221 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 16209 12801 16221 12804
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 17543 12804 18613 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19153 12835 19211 12841
rect 19153 12832 19165 12835
rect 18932 12804 19165 12832
rect 18932 12792 18938 12804
rect 19153 12801 19165 12804
rect 19199 12832 19211 12835
rect 20438 12832 20444 12844
rect 19199 12804 20444 12832
rect 19199 12801 19211 12804
rect 19153 12795 19211 12801
rect 20438 12792 20444 12804
rect 20496 12832 20502 12844
rect 24857 12835 24915 12841
rect 20496 12804 22094 12832
rect 20496 12792 20502 12804
rect 13842 12767 13900 12773
rect 13842 12764 13854 12767
rect 13096 12736 13854 12764
rect 12989 12727 13047 12733
rect 13842 12733 13854 12736
rect 13888 12733 13900 12767
rect 13842 12727 13900 12733
rect 12728 12668 12940 12696
rect 3142 12628 3148 12640
rect 2332 12600 3148 12628
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 7558 12588 7564 12640
rect 7616 12588 7622 12640
rect 8297 12631 8355 12637
rect 8297 12597 8309 12631
rect 8343 12628 8355 12631
rect 8570 12628 8576 12640
rect 8343 12600 8576 12628
rect 8343 12597 8355 12600
rect 8297 12591 8355 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 11698 12588 11704 12640
rect 11756 12588 11762 12640
rect 13004 12628 13032 12727
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14550 12764 14556 12776
rect 14240 12736 14556 12764
rect 14240 12724 14246 12736
rect 14550 12724 14556 12736
rect 14608 12764 14614 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 14608 12736 15301 12764
rect 14608 12724 14614 12736
rect 15289 12733 15301 12736
rect 15335 12733 15347 12767
rect 15289 12727 15347 12733
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 13449 12699 13507 12705
rect 13449 12665 13461 12699
rect 13495 12696 13507 12699
rect 13538 12696 13544 12708
rect 13495 12668 13544 12696
rect 13495 12665 13507 12668
rect 13449 12659 13507 12665
rect 13538 12656 13544 12668
rect 13596 12656 13602 12708
rect 15470 12696 15476 12708
rect 14568 12668 15476 12696
rect 14568 12628 14596 12668
rect 15470 12656 15476 12668
rect 15528 12696 15534 12708
rect 15580 12696 15608 12727
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 17681 12767 17739 12773
rect 17681 12764 17693 12767
rect 17460 12736 17693 12764
rect 17460 12724 17466 12736
rect 17681 12733 17693 12736
rect 17727 12764 17739 12767
rect 17770 12764 17776 12776
rect 17727 12736 17776 12764
rect 17727 12733 17739 12736
rect 17681 12727 17739 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 17957 12767 18015 12773
rect 17957 12764 17969 12767
rect 17920 12736 17969 12764
rect 17920 12724 17926 12736
rect 17957 12733 17969 12736
rect 18003 12733 18015 12767
rect 17957 12727 18015 12733
rect 19521 12767 19579 12773
rect 19521 12733 19533 12767
rect 19567 12764 19579 12767
rect 19610 12764 19616 12776
rect 19567 12736 19616 12764
rect 19567 12733 19579 12736
rect 19521 12727 19579 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 15528 12668 15608 12696
rect 15528 12656 15534 12668
rect 13004 12600 14596 12628
rect 14642 12588 14648 12640
rect 14700 12588 14706 12640
rect 14734 12588 14740 12640
rect 14792 12588 14798 12640
rect 17126 12588 17132 12640
rect 17184 12588 17190 12640
rect 22066 12628 22094 12804
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 25130 12832 25136 12844
rect 24903 12804 25136 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 25130 12792 25136 12804
rect 25188 12792 25194 12844
rect 29086 12792 29092 12844
rect 29144 12792 29150 12844
rect 29178 12792 29184 12844
rect 29236 12832 29242 12844
rect 29236 12804 29500 12832
rect 29236 12792 29242 12804
rect 22370 12724 22376 12776
rect 22428 12724 22434 12776
rect 24949 12767 25007 12773
rect 24949 12764 24961 12767
rect 23768 12736 24961 12764
rect 22186 12628 22192 12640
rect 22066 12600 22192 12628
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22925 12631 22983 12637
rect 22925 12628 22937 12631
rect 22520 12600 22937 12628
rect 22520 12588 22526 12600
rect 22925 12597 22937 12600
rect 22971 12597 22983 12631
rect 22925 12591 22983 12597
rect 23474 12588 23480 12640
rect 23532 12628 23538 12640
rect 23768 12628 23796 12736
rect 24949 12733 24961 12736
rect 24995 12733 25007 12767
rect 24949 12727 25007 12733
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 25096 12736 25329 12764
rect 25096 12724 25102 12736
rect 25317 12733 25329 12736
rect 25363 12733 25375 12767
rect 27246 12764 27252 12776
rect 25317 12727 25375 12733
rect 26712 12736 27252 12764
rect 23842 12656 23848 12708
rect 23900 12696 23906 12708
rect 23900 12668 24440 12696
rect 23900 12656 23906 12668
rect 24412 12637 24440 12668
rect 24213 12631 24271 12637
rect 24213 12628 24225 12631
rect 23532 12600 24225 12628
rect 23532 12588 23538 12600
rect 24213 12597 24225 12600
rect 24259 12597 24271 12631
rect 24213 12591 24271 12597
rect 24397 12631 24455 12637
rect 24397 12597 24409 12631
rect 24443 12597 24455 12631
rect 24397 12591 24455 12597
rect 25498 12588 25504 12640
rect 25556 12628 25562 12640
rect 25961 12631 26019 12637
rect 25961 12628 25973 12631
rect 25556 12600 25973 12628
rect 25556 12588 25562 12600
rect 25961 12597 25973 12600
rect 26007 12597 26019 12631
rect 25961 12591 26019 12597
rect 26510 12588 26516 12640
rect 26568 12628 26574 12640
rect 26712 12637 26740 12736
rect 27246 12724 27252 12736
rect 27304 12724 27310 12776
rect 29270 12724 29276 12776
rect 29328 12724 29334 12776
rect 29472 12764 29500 12804
rect 30190 12792 30196 12844
rect 30248 12792 30254 12844
rect 30282 12764 30288 12776
rect 29472 12736 30288 12764
rect 30282 12724 30288 12736
rect 30340 12724 30346 12776
rect 28629 12699 28687 12705
rect 28629 12665 28641 12699
rect 28675 12696 28687 12699
rect 28810 12696 28816 12708
rect 28675 12668 28816 12696
rect 28675 12665 28687 12668
rect 28629 12659 28687 12665
rect 28810 12656 28816 12668
rect 28868 12696 28874 12708
rect 30576 12696 30604 12928
rect 31496 12832 31524 12928
rect 33597 12903 33655 12909
rect 33597 12869 33609 12903
rect 33643 12900 33655 12903
rect 34330 12900 34336 12912
rect 33643 12872 34336 12900
rect 33643 12869 33655 12872
rect 33597 12863 33655 12869
rect 34330 12860 34336 12872
rect 34388 12860 34394 12912
rect 35066 12860 35072 12912
rect 35124 12860 35130 12912
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31496 12804 32137 12832
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 33505 12835 33563 12841
rect 33505 12801 33517 12835
rect 33551 12832 33563 12835
rect 33962 12832 33968 12844
rect 33551 12804 33968 12832
rect 33551 12801 33563 12804
rect 33505 12795 33563 12801
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 34238 12792 34244 12844
rect 34296 12832 34302 12844
rect 35710 12832 35716 12844
rect 34296 12804 35716 12832
rect 34296 12792 34302 12804
rect 34624 12773 34652 12804
rect 35710 12792 35716 12804
rect 35768 12792 35774 12844
rect 36541 12835 36599 12841
rect 36541 12801 36553 12835
rect 36587 12832 36599 12835
rect 37550 12832 37556 12844
rect 36587 12804 37556 12832
rect 36587 12801 36599 12804
rect 36541 12795 36599 12801
rect 37550 12792 37556 12804
rect 37608 12792 37614 12844
rect 39408 12841 39436 12940
rect 39850 12928 39856 12940
rect 39908 12928 39914 12980
rect 39942 12928 39948 12980
rect 40000 12928 40006 12980
rect 40310 12928 40316 12980
rect 40368 12928 40374 12980
rect 40678 12928 40684 12980
rect 40736 12968 40742 12980
rect 40736 12940 41368 12968
rect 40736 12928 40742 12940
rect 40328 12900 40356 12928
rect 41340 12909 41368 12940
rect 41690 12928 41696 12980
rect 41748 12968 41754 12980
rect 42061 12971 42119 12977
rect 42061 12968 42073 12971
rect 41748 12940 42073 12968
rect 41748 12928 41754 12940
rect 42061 12937 42073 12940
rect 42107 12937 42119 12971
rect 42061 12931 42119 12937
rect 42426 12928 42432 12980
rect 42484 12928 42490 12980
rect 43070 12928 43076 12980
rect 43128 12928 43134 12980
rect 47762 12928 47768 12980
rect 47820 12968 47826 12980
rect 47857 12971 47915 12977
rect 47857 12968 47869 12971
rect 47820 12940 47869 12968
rect 47820 12928 47826 12940
rect 47857 12937 47869 12940
rect 47903 12968 47915 12971
rect 48038 12968 48044 12980
rect 47903 12940 48044 12968
rect 47903 12937 47915 12940
rect 47857 12931 47915 12937
rect 48038 12928 48044 12940
rect 48096 12928 48102 12980
rect 53282 12928 53288 12980
rect 53340 12928 53346 12980
rect 53374 12928 53380 12980
rect 53432 12968 53438 12980
rect 55677 12971 55735 12977
rect 55677 12968 55689 12971
rect 53432 12940 55689 12968
rect 53432 12928 53438 12940
rect 55677 12937 55689 12940
rect 55723 12968 55735 12971
rect 56226 12968 56232 12980
rect 55723 12940 56232 12968
rect 55723 12937 55735 12940
rect 55677 12931 55735 12937
rect 56226 12928 56232 12940
rect 56284 12928 56290 12980
rect 56686 12928 56692 12980
rect 56744 12968 56750 12980
rect 56965 12971 57023 12977
rect 56965 12968 56977 12971
rect 56744 12940 56977 12968
rect 56744 12928 56750 12940
rect 56965 12937 56977 12940
rect 57011 12937 57023 12971
rect 56965 12931 57023 12937
rect 40773 12903 40831 12909
rect 40773 12900 40785 12903
rect 40328 12872 40785 12900
rect 40773 12869 40785 12872
rect 40819 12869 40831 12903
rect 40773 12863 40831 12869
rect 41325 12903 41383 12909
rect 41325 12869 41337 12903
rect 41371 12900 41383 12903
rect 42444 12900 42472 12928
rect 41371 12872 42472 12900
rect 41371 12869 41383 12872
rect 41325 12863 41383 12869
rect 39393 12835 39451 12841
rect 39393 12801 39405 12835
rect 39439 12801 39451 12835
rect 39393 12795 39451 12801
rect 40218 12792 40224 12844
rect 40276 12792 40282 12844
rect 41509 12835 41567 12841
rect 41509 12801 41521 12835
rect 41555 12832 41567 12835
rect 41782 12832 41788 12844
rect 41555 12804 41788 12832
rect 41555 12801 41567 12804
rect 41509 12795 41567 12801
rect 41782 12792 41788 12804
rect 41840 12792 41846 12844
rect 42058 12792 42064 12844
rect 42116 12832 42122 12844
rect 42429 12835 42487 12841
rect 42429 12832 42441 12835
rect 42116 12804 42441 12832
rect 42116 12792 42122 12804
rect 42429 12801 42441 12804
rect 42475 12801 42487 12835
rect 42429 12795 42487 12801
rect 47397 12835 47455 12841
rect 47397 12801 47409 12835
rect 47443 12832 47455 12835
rect 49602 12832 49608 12844
rect 47443 12804 49608 12832
rect 47443 12801 47455 12804
rect 47397 12795 47455 12801
rect 49602 12792 49608 12804
rect 49660 12792 49666 12844
rect 53190 12792 53196 12844
rect 53248 12792 53254 12844
rect 33781 12767 33839 12773
rect 33781 12733 33793 12767
rect 33827 12764 33839 12767
rect 34609 12767 34667 12773
rect 33827 12736 33861 12764
rect 33827 12733 33839 12736
rect 33781 12727 33839 12733
rect 34609 12733 34621 12767
rect 34655 12764 34667 12767
rect 34655 12736 34689 12764
rect 34655 12733 34667 12736
rect 34609 12727 34667 12733
rect 28868 12668 30604 12696
rect 28868 12656 28874 12668
rect 33502 12656 33508 12708
rect 33560 12696 33566 12708
rect 33796 12696 33824 12727
rect 47946 12724 47952 12776
rect 48004 12764 48010 12776
rect 48225 12767 48283 12773
rect 48225 12764 48237 12767
rect 48004 12736 48237 12764
rect 48004 12724 48010 12736
rect 48225 12733 48237 12736
rect 48271 12733 48283 12767
rect 48225 12727 48283 12733
rect 50985 12767 51043 12773
rect 50985 12733 50997 12767
rect 51031 12764 51043 12767
rect 51166 12764 51172 12776
rect 51031 12736 51172 12764
rect 51031 12733 51043 12736
rect 50985 12727 51043 12733
rect 51166 12724 51172 12736
rect 51224 12724 51230 12776
rect 51350 12724 51356 12776
rect 51408 12764 51414 12776
rect 51721 12767 51779 12773
rect 51721 12764 51733 12767
rect 51408 12736 51733 12764
rect 51408 12724 51414 12736
rect 51721 12733 51733 12736
rect 51767 12733 51779 12767
rect 51721 12727 51779 12733
rect 53006 12724 53012 12776
rect 53064 12764 53070 12776
rect 53469 12767 53527 12773
rect 53469 12764 53481 12767
rect 53064 12736 53481 12764
rect 53064 12724 53070 12736
rect 53469 12733 53481 12736
rect 53515 12733 53527 12767
rect 53469 12727 53527 12733
rect 55953 12767 56011 12773
rect 55953 12733 55965 12767
rect 55999 12733 56011 12767
rect 56244 12764 56272 12928
rect 57057 12835 57115 12841
rect 57057 12801 57069 12835
rect 57103 12832 57115 12835
rect 58529 12835 58587 12841
rect 58529 12832 58541 12835
rect 57103 12804 58541 12832
rect 57103 12801 57115 12804
rect 57057 12795 57115 12801
rect 58529 12801 58541 12804
rect 58575 12801 58587 12835
rect 58529 12795 58587 12801
rect 57149 12767 57207 12773
rect 57149 12764 57161 12767
rect 56244 12736 57161 12764
rect 55953 12727 56011 12733
rect 57149 12733 57161 12736
rect 57195 12733 57207 12767
rect 57149 12727 57207 12733
rect 35158 12696 35164 12708
rect 33560 12668 35164 12696
rect 33560 12656 33566 12668
rect 35158 12656 35164 12668
rect 35216 12696 35222 12708
rect 35345 12699 35403 12705
rect 35345 12696 35357 12699
rect 35216 12668 35357 12696
rect 35216 12656 35222 12668
rect 35345 12665 35357 12668
rect 35391 12665 35403 12699
rect 35345 12659 35403 12665
rect 36357 12699 36415 12705
rect 36357 12665 36369 12699
rect 36403 12696 36415 12699
rect 36722 12696 36728 12708
rect 36403 12668 36728 12696
rect 36403 12665 36415 12668
rect 36357 12659 36415 12665
rect 36722 12656 36728 12668
rect 36780 12656 36786 12708
rect 55968 12696 55996 12727
rect 57790 12724 57796 12776
rect 57848 12764 57854 12776
rect 57885 12767 57943 12773
rect 57885 12764 57897 12767
rect 57848 12736 57897 12764
rect 57848 12724 57854 12736
rect 57885 12733 57897 12736
rect 57931 12733 57943 12767
rect 57885 12727 57943 12733
rect 56597 12699 56655 12705
rect 56597 12696 56609 12699
rect 55968 12668 56609 12696
rect 56597 12665 56609 12668
rect 56643 12665 56655 12699
rect 56597 12659 56655 12665
rect 26697 12631 26755 12637
rect 26697 12628 26709 12631
rect 26568 12600 26709 12628
rect 26568 12588 26574 12600
rect 26697 12597 26709 12600
rect 26743 12597 26755 12631
rect 26697 12591 26755 12597
rect 31478 12588 31484 12640
rect 31536 12588 31542 12640
rect 32766 12588 32772 12640
rect 32824 12588 32830 12640
rect 33134 12588 33140 12640
rect 33192 12588 33198 12640
rect 34422 12588 34428 12640
rect 34480 12628 34486 12640
rect 39114 12628 39120 12640
rect 34480 12600 39120 12628
rect 34480 12588 34486 12600
rect 39114 12588 39120 12600
rect 39172 12588 39178 12640
rect 48866 12588 48872 12640
rect 48924 12588 48930 12640
rect 51074 12588 51080 12640
rect 51132 12628 51138 12640
rect 51537 12631 51595 12637
rect 51537 12628 51549 12631
rect 51132 12600 51549 12628
rect 51132 12588 51138 12600
rect 51537 12597 51549 12600
rect 51583 12597 51595 12631
rect 51537 12591 51595 12597
rect 52362 12588 52368 12640
rect 52420 12588 52426 12640
rect 54110 12588 54116 12640
rect 54168 12588 54174 12640
rect 56505 12631 56563 12637
rect 56505 12597 56517 12631
rect 56551 12628 56563 12631
rect 56686 12628 56692 12640
rect 56551 12600 56692 12628
rect 56551 12597 56563 12600
rect 56505 12591 56563 12597
rect 56686 12588 56692 12600
rect 56744 12588 56750 12640
rect 1104 12538 58880 12560
rect 1104 12486 8172 12538
rect 8224 12486 8236 12538
rect 8288 12486 8300 12538
rect 8352 12486 8364 12538
rect 8416 12486 8428 12538
rect 8480 12486 22616 12538
rect 22668 12486 22680 12538
rect 22732 12486 22744 12538
rect 22796 12486 22808 12538
rect 22860 12486 22872 12538
rect 22924 12486 37060 12538
rect 37112 12486 37124 12538
rect 37176 12486 37188 12538
rect 37240 12486 37252 12538
rect 37304 12486 37316 12538
rect 37368 12486 51504 12538
rect 51556 12486 51568 12538
rect 51620 12486 51632 12538
rect 51684 12486 51696 12538
rect 51748 12486 51760 12538
rect 51812 12486 58880 12538
rect 1104 12464 58880 12486
rect 4154 12424 4160 12436
rect 3068 12396 4160 12424
rect 3068 12229 3096 12396
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 7006 12384 7012 12436
rect 7064 12384 7070 12436
rect 12250 12384 12256 12436
rect 12308 12384 12314 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12584 12396 13001 12424
rect 12584 12384 12590 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 12989 12387 13047 12393
rect 14108 12396 15424 12424
rect 6178 12316 6184 12368
rect 6236 12356 6242 12368
rect 6822 12356 6828 12368
rect 6236 12328 6828 12356
rect 6236 12316 6242 12328
rect 6822 12316 6828 12328
rect 6880 12356 6886 12368
rect 9122 12356 9128 12368
rect 6880 12328 9128 12356
rect 6880 12316 6886 12328
rect 9122 12316 9128 12328
rect 9180 12356 9186 12368
rect 9398 12356 9404 12368
rect 9180 12328 9404 12356
rect 9180 12316 9186 12328
rect 9398 12316 9404 12328
rect 9456 12316 9462 12368
rect 14108 12356 14136 12396
rect 12268 12328 14136 12356
rect 15396 12356 15424 12396
rect 15470 12384 15476 12436
rect 15528 12384 15534 12436
rect 17586 12384 17592 12436
rect 17644 12384 17650 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 19794 12424 19800 12436
rect 18564 12396 19800 12424
rect 18564 12384 18570 12396
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 22186 12384 22192 12436
rect 22244 12384 22250 12436
rect 22370 12384 22376 12436
rect 22428 12384 22434 12436
rect 24213 12427 24271 12433
rect 24213 12393 24225 12427
rect 24259 12424 24271 12427
rect 24486 12424 24492 12436
rect 24259 12396 24492 12424
rect 24259 12393 24271 12396
rect 24213 12387 24271 12393
rect 24486 12384 24492 12396
rect 24544 12424 24550 12436
rect 26510 12424 26516 12436
rect 24544 12396 26516 12424
rect 24544 12384 24550 12396
rect 26510 12384 26516 12396
rect 26568 12384 26574 12436
rect 29086 12384 29092 12436
rect 29144 12424 29150 12436
rect 29365 12427 29423 12433
rect 29365 12424 29377 12427
rect 29144 12396 29377 12424
rect 29144 12384 29150 12396
rect 29365 12393 29377 12396
rect 29411 12393 29423 12427
rect 30650 12424 30656 12436
rect 29365 12387 29423 12393
rect 29748 12396 30656 12424
rect 16761 12359 16819 12365
rect 16761 12356 16773 12359
rect 15396 12328 16773 12356
rect 12268 12300 12296 12328
rect 16761 12325 16773 12328
rect 16807 12356 16819 12359
rect 17770 12356 17776 12368
rect 16807 12328 17776 12356
rect 16807 12325 16819 12328
rect 16761 12319 16819 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 24762 12356 24768 12368
rect 22940 12328 24768 12356
rect 7650 12248 7656 12300
rect 7708 12248 7714 12300
rect 7760 12260 8708 12288
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3602 12220 3608 12232
rect 3476 12192 3608 12220
rect 3476 12180 3482 12192
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12220 3847 12223
rect 5534 12220 5540 12232
rect 3835 12192 5540 12220
rect 3835 12189 3847 12192
rect 3789 12183 3847 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12220 7435 12223
rect 7760 12220 7788 12260
rect 8680 12232 8708 12260
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 8812 12260 9505 12288
rect 8812 12248 8818 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 11698 12248 11704 12300
rect 11756 12248 11762 12300
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 12345 12291 12403 12297
rect 12345 12257 12357 12291
rect 12391 12288 12403 12291
rect 12434 12288 12440 12300
rect 12391 12260 12440 12288
rect 12391 12257 12403 12260
rect 12345 12251 12403 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 17037 12291 17095 12297
rect 17037 12257 17049 12291
rect 17083 12288 17095 12291
rect 17126 12288 17132 12300
rect 17083 12260 17132 12288
rect 17083 12257 17095 12260
rect 17037 12251 17095 12257
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 21818 12248 21824 12300
rect 21876 12288 21882 12300
rect 22940 12297 22968 12328
rect 24762 12316 24768 12328
rect 24820 12316 24826 12368
rect 25041 12359 25099 12365
rect 25041 12325 25053 12359
rect 25087 12356 25099 12359
rect 25087 12328 26188 12356
rect 25087 12325 25099 12328
rect 25041 12319 25099 12325
rect 22925 12291 22983 12297
rect 22925 12288 22937 12291
rect 21876 12260 22937 12288
rect 21876 12248 21882 12260
rect 22925 12257 22937 12260
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 25222 12288 25228 12300
rect 23072 12260 25228 12288
rect 23072 12248 23078 12260
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 25498 12248 25504 12300
rect 25556 12248 25562 12300
rect 25590 12248 25596 12300
rect 25648 12248 25654 12300
rect 26160 12297 26188 12328
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 28537 12359 28595 12365
rect 28537 12356 28549 12359
rect 26384 12328 28549 12356
rect 26384 12316 26390 12328
rect 28537 12325 28549 12328
rect 28583 12356 28595 12359
rect 29270 12356 29276 12368
rect 28583 12328 29276 12356
rect 28583 12325 28595 12328
rect 28537 12319 28595 12325
rect 29270 12316 29276 12328
rect 29328 12316 29334 12368
rect 26145 12291 26203 12297
rect 26145 12257 26157 12291
rect 26191 12257 26203 12291
rect 26145 12251 26203 12257
rect 28810 12248 28816 12300
rect 28868 12248 28874 12300
rect 7423 12192 7788 12220
rect 7423 12189 7435 12192
rect 7377 12183 7435 12189
rect 7926 12180 7932 12232
rect 7984 12180 7990 12232
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 16482 12220 16488 12232
rect 14139 12192 16488 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 3234 12112 3240 12164
rect 3292 12112 3298 12164
rect 3329 12155 3387 12161
rect 3329 12121 3341 12155
rect 3375 12152 3387 12155
rect 3878 12152 3884 12164
rect 3375 12124 3884 12152
rect 3375 12121 3387 12124
rect 3329 12115 3387 12121
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4056 12155 4114 12161
rect 4056 12121 4068 12155
rect 4102 12152 4114 12155
rect 4982 12152 4988 12164
rect 4102 12124 4988 12152
rect 4102 12121 4114 12124
rect 4056 12115 4114 12121
rect 4982 12112 4988 12124
rect 5040 12112 5046 12164
rect 6917 12155 6975 12161
rect 6917 12121 6929 12155
rect 6963 12152 6975 12155
rect 8018 12152 8024 12164
rect 6963 12124 8024 12152
rect 6963 12121 6975 12124
rect 6917 12115 6975 12121
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 8386 12112 8392 12164
rect 8444 12152 8450 12164
rect 9582 12152 9588 12164
rect 8444 12124 9588 12152
rect 8444 12112 8450 12124
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 14360 12155 14418 12161
rect 14360 12121 14372 12155
rect 14406 12152 14418 12155
rect 15194 12152 15200 12164
rect 14406 12124 15200 12152
rect 14406 12121 14418 12124
rect 14360 12115 14418 12121
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 15856 12096 15884 12192
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 19889 12223 19947 12229
rect 19889 12220 19901 12223
rect 18012 12192 19901 12220
rect 18012 12180 18018 12192
rect 19889 12189 19901 12192
rect 19935 12220 19947 12223
rect 21082 12220 21088 12232
rect 19935 12192 21088 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12220 22799 12223
rect 23032 12220 23060 12248
rect 22787 12192 23060 12220
rect 22787 12189 22799 12192
rect 22741 12183 22799 12189
rect 23290 12180 23296 12232
rect 23348 12180 23354 12232
rect 29748 12220 29776 12396
rect 30650 12384 30656 12396
rect 30708 12384 30714 12436
rect 30742 12384 30748 12436
rect 30800 12424 30806 12436
rect 31389 12427 31447 12433
rect 31389 12424 31401 12427
rect 30800 12396 31401 12424
rect 30800 12384 30806 12396
rect 31389 12393 31401 12396
rect 31435 12393 31447 12427
rect 31389 12387 31447 12393
rect 31404 12288 31432 12387
rect 31846 12384 31852 12436
rect 31904 12424 31910 12436
rect 32125 12427 32183 12433
rect 32125 12424 32137 12427
rect 31904 12396 32137 12424
rect 31904 12384 31910 12396
rect 32125 12393 32137 12396
rect 32171 12393 32183 12427
rect 32125 12387 32183 12393
rect 33594 12384 33600 12436
rect 33652 12384 33658 12436
rect 33962 12384 33968 12436
rect 34020 12424 34026 12436
rect 34425 12427 34483 12433
rect 34425 12424 34437 12427
rect 34020 12396 34437 12424
rect 34020 12384 34026 12396
rect 34425 12393 34437 12396
rect 34471 12393 34483 12427
rect 34425 12387 34483 12393
rect 40129 12427 40187 12433
rect 40129 12393 40141 12427
rect 40175 12424 40187 12427
rect 40497 12427 40555 12433
rect 40497 12424 40509 12427
rect 40175 12396 40509 12424
rect 40175 12393 40187 12396
rect 40129 12387 40187 12393
rect 40497 12393 40509 12396
rect 40543 12424 40555 12427
rect 40678 12424 40684 12436
rect 40543 12396 40684 12424
rect 40543 12393 40555 12396
rect 40497 12387 40555 12393
rect 40678 12384 40684 12396
rect 40736 12384 40742 12436
rect 47854 12384 47860 12436
rect 47912 12424 47918 12436
rect 49326 12424 49332 12436
rect 47912 12396 49332 12424
rect 47912 12384 47918 12396
rect 49326 12384 49332 12396
rect 49384 12424 49390 12436
rect 49384 12396 51396 12424
rect 49384 12384 49390 12396
rect 32766 12356 32772 12368
rect 31726 12328 32772 12356
rect 31481 12291 31539 12297
rect 31481 12288 31493 12291
rect 31404 12260 31493 12288
rect 31481 12257 31493 12260
rect 31527 12257 31539 12291
rect 31481 12251 31539 12257
rect 23492 12192 29776 12220
rect 30009 12223 30067 12229
rect 16500 12152 16528 12180
rect 23492 12164 23520 12192
rect 30009 12189 30021 12223
rect 30055 12220 30067 12223
rect 31110 12220 31116 12232
rect 30055 12192 31116 12220
rect 30055 12189 30067 12192
rect 30009 12183 30067 12189
rect 31110 12180 31116 12192
rect 31168 12180 31174 12232
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 16500 12124 18061 12152
rect 18049 12121 18061 12124
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 20349 12155 20407 12161
rect 20349 12121 20361 12155
rect 20395 12152 20407 12155
rect 20438 12152 20444 12164
rect 20395 12124 20444 12152
rect 20395 12121 20407 12124
rect 20349 12115 20407 12121
rect 20438 12112 20444 12124
rect 20496 12152 20502 12164
rect 23474 12152 23480 12164
rect 20496 12124 23480 12152
rect 20496 12112 20502 12124
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 24762 12112 24768 12164
rect 24820 12152 24826 12164
rect 26694 12152 26700 12164
rect 24820 12124 26700 12152
rect 24820 12112 24826 12124
rect 26694 12112 26700 12124
rect 26752 12112 26758 12164
rect 30276 12155 30334 12161
rect 30276 12121 30288 12155
rect 30322 12152 30334 12155
rect 31726 12152 31754 12328
rect 32766 12316 32772 12328
rect 32824 12316 32830 12368
rect 34330 12316 34336 12368
rect 34388 12356 34394 12368
rect 36814 12356 36820 12368
rect 34388 12328 36820 12356
rect 34388 12316 34394 12328
rect 36814 12316 36820 12328
rect 36872 12316 36878 12368
rect 41690 12316 41696 12368
rect 41748 12356 41754 12368
rect 42334 12356 42340 12368
rect 41748 12328 42340 12356
rect 41748 12316 41754 12328
rect 42334 12316 42340 12328
rect 42392 12356 42398 12368
rect 47762 12356 47768 12368
rect 42392 12328 42748 12356
rect 42392 12316 42398 12328
rect 33045 12291 33103 12297
rect 33045 12257 33057 12291
rect 33091 12288 33103 12291
rect 33134 12288 33140 12300
rect 33091 12260 33140 12288
rect 33091 12257 33103 12260
rect 33045 12251 33103 12257
rect 33134 12248 33140 12260
rect 33192 12248 33198 12300
rect 33870 12248 33876 12300
rect 33928 12288 33934 12300
rect 35802 12288 35808 12300
rect 33928 12260 35808 12288
rect 33928 12248 33934 12260
rect 35802 12248 35808 12260
rect 35860 12248 35866 12300
rect 41414 12248 41420 12300
rect 41472 12288 41478 12300
rect 42720 12297 42748 12328
rect 42996 12328 47768 12356
rect 42996 12300 43024 12328
rect 47762 12316 47768 12328
rect 47820 12356 47826 12368
rect 48409 12359 48467 12365
rect 47820 12328 48176 12356
rect 47820 12316 47826 12328
rect 42705 12291 42763 12297
rect 41472 12260 42564 12288
rect 41472 12248 41478 12260
rect 34606 12180 34612 12232
rect 34664 12220 34670 12232
rect 34701 12223 34759 12229
rect 34701 12220 34713 12223
rect 34664 12192 34713 12220
rect 34664 12180 34670 12192
rect 34701 12189 34713 12192
rect 34747 12189 34759 12223
rect 34701 12183 34759 12189
rect 35986 12180 35992 12232
rect 36044 12180 36050 12232
rect 36354 12180 36360 12232
rect 36412 12220 36418 12232
rect 37001 12223 37059 12229
rect 37001 12220 37013 12223
rect 36412 12192 37013 12220
rect 36412 12180 36418 12192
rect 37001 12189 37013 12192
rect 37047 12220 37059 12223
rect 37458 12220 37464 12232
rect 37047 12192 37464 12220
rect 37047 12189 37059 12192
rect 37001 12183 37059 12189
rect 37458 12180 37464 12192
rect 37516 12220 37522 12232
rect 42242 12220 42248 12232
rect 37516 12192 42248 12220
rect 37516 12180 37522 12192
rect 42242 12180 42248 12192
rect 42300 12180 42306 12232
rect 42536 12229 42564 12260
rect 42705 12257 42717 12291
rect 42751 12257 42763 12291
rect 42705 12251 42763 12257
rect 42978 12248 42984 12300
rect 43036 12248 43042 12300
rect 45646 12248 45652 12300
rect 45704 12288 45710 12300
rect 48148 12297 48176 12328
rect 48409 12325 48421 12359
rect 48455 12356 48467 12359
rect 51368 12356 51396 12396
rect 51442 12384 51448 12436
rect 51500 12424 51506 12436
rect 51813 12427 51871 12433
rect 51813 12424 51825 12427
rect 51500 12396 51825 12424
rect 51500 12384 51506 12396
rect 51813 12393 51825 12396
rect 51859 12393 51871 12427
rect 51813 12387 51871 12393
rect 52181 12427 52239 12433
rect 52181 12393 52193 12427
rect 52227 12424 52239 12427
rect 52914 12424 52920 12436
rect 52227 12396 52920 12424
rect 52227 12393 52239 12396
rect 52181 12387 52239 12393
rect 52196 12356 52224 12387
rect 52914 12384 52920 12396
rect 52972 12384 52978 12436
rect 53742 12384 53748 12436
rect 53800 12424 53806 12436
rect 57330 12424 57336 12436
rect 53800 12396 57336 12424
rect 53800 12384 53806 12396
rect 57330 12384 57336 12396
rect 57388 12424 57394 12436
rect 57388 12396 57928 12424
rect 57388 12384 57394 12396
rect 57900 12368 57928 12396
rect 58434 12384 58440 12436
rect 58492 12384 58498 12436
rect 53834 12356 53840 12368
rect 48455 12328 49280 12356
rect 51368 12328 52224 12356
rect 53484 12328 53840 12356
rect 48455 12325 48467 12328
rect 48409 12319 48467 12325
rect 49252 12297 49280 12328
rect 48133 12291 48191 12297
rect 45704 12260 47348 12288
rect 45704 12248 45710 12260
rect 42521 12223 42579 12229
rect 42521 12189 42533 12223
rect 42567 12189 42579 12223
rect 42521 12183 42579 12189
rect 45278 12180 45284 12232
rect 45336 12180 45342 12232
rect 46014 12180 46020 12232
rect 46072 12180 46078 12232
rect 46845 12223 46903 12229
rect 46845 12189 46857 12223
rect 46891 12189 46903 12223
rect 46845 12183 46903 12189
rect 45002 12152 45008 12164
rect 30322 12124 31754 12152
rect 39040 12124 45008 12152
rect 30322 12121 30334 12124
rect 30276 12115 30334 12121
rect 39040 12096 39068 12124
rect 45002 12112 45008 12124
rect 45060 12112 45066 12164
rect 46860 12096 46888 12183
rect 47320 12152 47348 12260
rect 48133 12257 48145 12291
rect 48179 12257 48191 12291
rect 48133 12251 48191 12257
rect 49053 12291 49111 12297
rect 49053 12257 49065 12291
rect 49099 12257 49111 12291
rect 49053 12251 49111 12257
rect 49237 12291 49295 12297
rect 49237 12257 49249 12291
rect 49283 12257 49295 12291
rect 49237 12251 49295 12257
rect 47949 12223 48007 12229
rect 47949 12189 47961 12223
rect 47995 12220 48007 12223
rect 48314 12220 48320 12232
rect 47995 12192 48320 12220
rect 47995 12189 48007 12192
rect 47949 12183 48007 12189
rect 48314 12180 48320 12192
rect 48372 12180 48378 12232
rect 48777 12223 48835 12229
rect 48777 12189 48789 12223
rect 48823 12220 48835 12223
rect 48866 12220 48872 12232
rect 48823 12192 48872 12220
rect 48823 12189 48835 12192
rect 48777 12183 48835 12189
rect 48866 12180 48872 12192
rect 48924 12180 48930 12232
rect 49068 12220 49096 12251
rect 49602 12248 49608 12300
rect 49660 12248 49666 12300
rect 49620 12220 49648 12248
rect 50433 12223 50491 12229
rect 50433 12220 50445 12223
rect 49068 12192 49648 12220
rect 50172 12192 50445 12220
rect 48958 12152 48964 12164
rect 47320 12124 48964 12152
rect 3602 12044 3608 12096
rect 3660 12044 3666 12096
rect 5166 12044 5172 12096
rect 5224 12044 5230 12096
rect 7469 12087 7527 12093
rect 7469 12053 7481 12087
rect 7515 12084 7527 12087
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 7515 12056 8493 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 8481 12053 8493 12056
rect 8527 12053 8539 12087
rect 8481 12047 8539 12053
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12084 8999 12087
rect 9214 12084 9220 12096
rect 8987 12056 9220 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 9858 12084 9864 12096
rect 9447 12056 9864 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 13722 12084 13728 12096
rect 13320 12056 13728 12084
rect 13320 12044 13326 12056
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 13909 12087 13967 12093
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 14182 12084 14188 12096
rect 13955 12056 14188 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 15838 12044 15844 12096
rect 15896 12044 15902 12096
rect 21818 12044 21824 12096
rect 21876 12044 21882 12096
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12084 22891 12087
rect 23845 12087 23903 12093
rect 23845 12084 23857 12087
rect 22879 12056 23857 12084
rect 22879 12053 22891 12056
rect 22833 12047 22891 12053
rect 23845 12053 23857 12056
rect 23891 12053 23903 12087
rect 23845 12047 23903 12053
rect 24854 12044 24860 12096
rect 24912 12044 24918 12096
rect 25222 12044 25228 12096
rect 25280 12084 25286 12096
rect 25409 12087 25467 12093
rect 25409 12084 25421 12087
rect 25280 12056 25421 12084
rect 25280 12044 25286 12056
rect 25409 12053 25421 12056
rect 25455 12053 25467 12087
rect 25409 12047 25467 12053
rect 26786 12044 26792 12096
rect 26844 12044 26850 12096
rect 30374 12044 30380 12096
rect 30432 12084 30438 12096
rect 31386 12084 31392 12096
rect 30432 12056 31392 12084
rect 30432 12044 30438 12056
rect 31386 12044 31392 12056
rect 31444 12044 31450 12096
rect 35342 12044 35348 12096
rect 35400 12044 35406 12096
rect 36630 12044 36636 12096
rect 36688 12044 36694 12096
rect 39022 12044 39028 12096
rect 39080 12044 39086 12096
rect 42058 12044 42064 12096
rect 42116 12044 42122 12096
rect 42150 12044 42156 12096
rect 42208 12044 42214 12096
rect 42613 12087 42671 12093
rect 42613 12053 42625 12087
rect 42659 12084 42671 12087
rect 43898 12084 43904 12096
rect 42659 12056 43904 12084
rect 42659 12053 42671 12056
rect 42613 12047 42671 12053
rect 43898 12044 43904 12056
rect 43956 12044 43962 12096
rect 45554 12044 45560 12096
rect 45612 12084 45618 12096
rect 45925 12087 45983 12093
rect 45925 12084 45937 12087
rect 45612 12056 45937 12084
rect 45612 12044 45618 12056
rect 45925 12053 45937 12056
rect 45971 12053 45983 12087
rect 45925 12047 45983 12053
rect 46658 12044 46664 12096
rect 46716 12044 46722 12096
rect 46842 12044 46848 12096
rect 46900 12044 46906 12096
rect 47394 12044 47400 12096
rect 47452 12044 47458 12096
rect 47581 12087 47639 12093
rect 47581 12053 47593 12087
rect 47627 12084 47639 12087
rect 47762 12084 47768 12096
rect 47627 12056 47768 12084
rect 47627 12053 47639 12056
rect 47581 12047 47639 12053
rect 47762 12044 47768 12056
rect 47820 12044 47826 12096
rect 48041 12087 48099 12093
rect 48041 12053 48053 12087
rect 48087 12084 48099 12087
rect 48222 12084 48228 12096
rect 48087 12056 48228 12084
rect 48087 12053 48099 12056
rect 48041 12047 48099 12053
rect 48222 12044 48228 12056
rect 48280 12044 48286 12096
rect 48884 12093 48912 12124
rect 48958 12112 48964 12124
rect 49016 12112 49022 12164
rect 50172 12096 50200 12192
rect 50433 12189 50445 12192
rect 50479 12220 50491 12223
rect 52273 12223 52331 12229
rect 52273 12220 52285 12223
rect 50479 12192 52285 12220
rect 50479 12189 50491 12192
rect 50433 12183 50491 12189
rect 52273 12189 52285 12192
rect 52319 12220 52331 12223
rect 53484 12220 53512 12328
rect 53834 12316 53840 12328
rect 53892 12356 53898 12368
rect 53892 12328 54340 12356
rect 53892 12316 53898 12328
rect 54110 12288 54116 12300
rect 52319 12192 53512 12220
rect 53576 12260 54116 12288
rect 52319 12189 52331 12192
rect 52273 12183 52331 12189
rect 50700 12155 50758 12161
rect 50700 12121 50712 12155
rect 50746 12152 50758 12155
rect 51074 12152 51080 12164
rect 50746 12124 51080 12152
rect 50746 12121 50758 12124
rect 50700 12115 50758 12121
rect 51074 12112 51080 12124
rect 51132 12112 51138 12164
rect 52540 12155 52598 12161
rect 52540 12121 52552 12155
rect 52586 12152 52598 12155
rect 53576 12152 53604 12260
rect 54110 12248 54116 12260
rect 54168 12248 54174 12300
rect 54312 12288 54340 12328
rect 54570 12316 54576 12368
rect 54628 12356 54634 12368
rect 55858 12356 55864 12368
rect 54628 12328 55864 12356
rect 54628 12316 54634 12328
rect 55858 12316 55864 12328
rect 55916 12316 55922 12368
rect 57882 12316 57888 12368
rect 57940 12316 57946 12368
rect 54312 12260 56456 12288
rect 53745 12223 53803 12229
rect 53745 12189 53757 12223
rect 53791 12189 53803 12223
rect 53745 12183 53803 12189
rect 52586 12124 53604 12152
rect 52586 12121 52598 12124
rect 52540 12115 52598 12121
rect 48869 12087 48927 12093
rect 48869 12053 48881 12087
rect 48915 12053 48927 12087
rect 48869 12047 48927 12053
rect 49878 12044 49884 12096
rect 49936 12044 49942 12096
rect 50154 12044 50160 12096
rect 50212 12044 50218 12096
rect 52178 12044 52184 12096
rect 52236 12084 52242 12096
rect 53653 12087 53711 12093
rect 53653 12084 53665 12087
rect 52236 12056 53665 12084
rect 52236 12044 52242 12056
rect 53653 12053 53665 12056
rect 53699 12084 53711 12087
rect 53760 12084 53788 12183
rect 54478 12180 54484 12232
rect 54536 12180 54542 12232
rect 55306 12180 55312 12232
rect 55364 12180 55370 12232
rect 56428 12229 56456 12260
rect 56686 12229 56692 12232
rect 56413 12223 56471 12229
rect 56413 12189 56425 12223
rect 56459 12189 56471 12223
rect 56413 12183 56471 12189
rect 56680 12183 56692 12229
rect 56686 12180 56692 12183
rect 56744 12180 56750 12232
rect 57330 12152 57336 12164
rect 57072 12124 57336 12152
rect 53699 12056 53788 12084
rect 53699 12053 53711 12056
rect 53653 12047 53711 12053
rect 54386 12044 54392 12096
rect 54444 12044 54450 12096
rect 55122 12044 55128 12096
rect 55180 12044 55186 12096
rect 55950 12044 55956 12096
rect 56008 12044 56014 12096
rect 56042 12044 56048 12096
rect 56100 12084 56106 12096
rect 56321 12087 56379 12093
rect 56321 12084 56333 12087
rect 56100 12056 56333 12084
rect 56100 12044 56106 12056
rect 56321 12053 56333 12056
rect 56367 12084 56379 12087
rect 57072 12084 57100 12124
rect 57330 12112 57336 12124
rect 57388 12112 57394 12164
rect 58250 12112 58256 12164
rect 58308 12152 58314 12164
rect 58345 12155 58403 12161
rect 58345 12152 58357 12155
rect 58308 12124 58357 12152
rect 58308 12112 58314 12124
rect 58345 12121 58357 12124
rect 58391 12121 58403 12155
rect 58345 12115 58403 12121
rect 56367 12056 57100 12084
rect 56367 12053 56379 12056
rect 56321 12047 56379 12053
rect 57146 12044 57152 12096
rect 57204 12084 57210 12096
rect 57790 12084 57796 12096
rect 57204 12056 57796 12084
rect 57204 12044 57210 12056
rect 57790 12044 57796 12056
rect 57848 12044 57854 12096
rect 1104 11994 59040 12016
rect 1104 11942 15394 11994
rect 15446 11942 15458 11994
rect 15510 11942 15522 11994
rect 15574 11942 15586 11994
rect 15638 11942 15650 11994
rect 15702 11942 29838 11994
rect 29890 11942 29902 11994
rect 29954 11942 29966 11994
rect 30018 11942 30030 11994
rect 30082 11942 30094 11994
rect 30146 11942 44282 11994
rect 44334 11942 44346 11994
rect 44398 11942 44410 11994
rect 44462 11942 44474 11994
rect 44526 11942 44538 11994
rect 44590 11942 58726 11994
rect 58778 11942 58790 11994
rect 58842 11942 58854 11994
rect 58906 11942 58918 11994
rect 58970 11942 58982 11994
rect 59034 11942 59040 11994
rect 1104 11920 59040 11942
rect 2685 11883 2743 11889
rect 2685 11849 2697 11883
rect 2731 11880 2743 11883
rect 3050 11880 3056 11892
rect 2731 11852 3056 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3510 11880 3516 11892
rect 3467 11852 3516 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 3602 11840 3608 11892
rect 3660 11840 3666 11892
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 3936 11852 4261 11880
rect 3936 11840 3942 11852
rect 4249 11849 4261 11852
rect 4295 11849 4307 11883
rect 4249 11843 4307 11849
rect 4982 11840 4988 11892
rect 5040 11840 5046 11892
rect 5166 11840 5172 11892
rect 5224 11840 5230 11892
rect 5534 11840 5540 11892
rect 5592 11840 5598 11892
rect 6178 11840 6184 11892
rect 6236 11840 6242 11892
rect 8570 11880 8576 11892
rect 6472 11852 8576 11880
rect 2884 11784 3280 11812
rect 2884 11753 2912 11784
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 3050 11704 3056 11756
rect 3108 11704 3114 11756
rect 3252 11753 3280 11784
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11713 3203 11747
rect 3145 11707 3203 11713
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3326 11744 3332 11756
rect 3283 11716 3332 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3160 11676 3188 11707
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3620 11744 3648 11840
rect 4341 11747 4399 11753
rect 4341 11744 4353 11747
rect 3620 11716 4353 11744
rect 3421 11707 3479 11713
rect 4341 11713 4353 11716
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 3436 11676 3464 11707
rect 2884 11648 3464 11676
rect 3697 11679 3755 11685
rect 2884 11552 2912 11648
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 5184 11676 5212 11840
rect 5552 11744 5580 11840
rect 6472 11753 6500 11852
rect 8570 11840 8576 11852
rect 8628 11880 8634 11892
rect 10410 11880 10416 11892
rect 8628 11852 10416 11880
rect 8628 11840 8634 11852
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 12710 11880 12716 11892
rect 12575 11852 12716 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 12710 11840 12716 11852
rect 12768 11880 12774 11892
rect 13538 11880 13544 11892
rect 12768 11852 13544 11880
rect 12768 11840 12774 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 15194 11840 15200 11892
rect 15252 11840 15258 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 17589 11883 17647 11889
rect 17589 11880 17601 11883
rect 16540 11852 17601 11880
rect 16540 11840 16546 11852
rect 17589 11849 17601 11852
rect 17635 11880 17647 11883
rect 19334 11880 19340 11892
rect 17635 11852 19340 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 19334 11840 19340 11852
rect 19392 11880 19398 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 19392 11852 21189 11880
rect 19392 11840 19398 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 23201 11883 23259 11889
rect 23201 11849 23213 11883
rect 23247 11880 23259 11883
rect 23290 11880 23296 11892
rect 23247 11852 23296 11880
rect 23247 11849 23259 11852
rect 23201 11843 23259 11849
rect 6724 11815 6782 11821
rect 6724 11781 6736 11815
rect 6770 11812 6782 11815
rect 7558 11812 7564 11824
rect 6770 11784 7564 11812
rect 6770 11781 6782 11784
rect 6724 11775 6782 11781
rect 7558 11772 7564 11784
rect 7616 11772 7622 11824
rect 9858 11772 9864 11824
rect 9916 11772 9922 11824
rect 12802 11772 12808 11824
rect 12860 11812 12866 11824
rect 15565 11815 15623 11821
rect 15565 11812 15577 11815
rect 12860 11784 15577 11812
rect 12860 11772 12866 11784
rect 15565 11781 15577 11784
rect 15611 11812 15623 11815
rect 16298 11812 16304 11824
rect 15611 11784 16304 11812
rect 15611 11781 15623 11784
rect 15565 11775 15623 11781
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18049 11815 18107 11821
rect 18049 11812 18061 11815
rect 18012 11784 18061 11812
rect 18012 11772 18018 11784
rect 18049 11781 18061 11784
rect 18095 11781 18107 11815
rect 18049 11775 18107 11781
rect 20257 11815 20315 11821
rect 20257 11781 20269 11815
rect 20303 11812 20315 11815
rect 20714 11812 20720 11824
rect 20303 11784 20720 11812
rect 20303 11781 20315 11784
rect 20257 11775 20315 11781
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 5552 11716 6469 11744
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8205 11747 8263 11753
rect 7984 11716 8156 11744
rect 7984 11704 7990 11716
rect 3743 11648 5212 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 4246 11608 4252 11620
rect 3068 11580 4252 11608
rect 3068 11552 3096 11580
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 7837 11611 7895 11617
rect 7837 11577 7849 11611
rect 7883 11608 7895 11611
rect 7944 11608 7972 11704
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11645 8079 11679
rect 8128 11676 8156 11716
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8386 11744 8392 11756
rect 8251 11716 8392 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11744 14703 11747
rect 14734 11744 14740 11756
rect 14691 11716 14740 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 21192 11744 21220 11843
rect 23290 11840 23296 11852
rect 23348 11880 23354 11892
rect 24210 11880 24216 11892
rect 23348 11852 24216 11880
rect 23348 11840 23354 11852
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 24486 11840 24492 11892
rect 24544 11880 24550 11892
rect 25590 11880 25596 11892
rect 24544 11852 25268 11880
rect 24544 11840 24550 11852
rect 22088 11815 22146 11821
rect 22088 11781 22100 11815
rect 22134 11812 22146 11815
rect 22462 11812 22468 11824
rect 22134 11784 22468 11812
rect 22134 11781 22146 11784
rect 22088 11775 22146 11781
rect 22462 11772 22468 11784
rect 22520 11772 22526 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 21634 11744 21640 11756
rect 21192 11716 21640 11744
rect 21634 11704 21640 11716
rect 21692 11744 21698 11756
rect 25240 11753 25268 11852
rect 25332 11852 25596 11880
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21692 11716 21833 11744
rect 21692 11704 21698 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 24489 11747 24547 11753
rect 21821 11707 21879 11713
rect 21928 11716 23428 11744
rect 9122 11685 9128 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 8128 11648 8953 11676
rect 8021 11639 8079 11645
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 9079 11679 9128 11685
rect 9079 11645 9091 11679
rect 9125 11645 9128 11679
rect 9079 11639 9128 11645
rect 7883 11580 7972 11608
rect 7883 11577 7895 11580
rect 7837 11571 7895 11577
rect 2866 11500 2872 11552
rect 2924 11500 2930 11552
rect 3050 11500 3056 11552
rect 3108 11500 3114 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4614 11540 4620 11552
rect 3660 11512 4620 11540
rect 3660 11500 3666 11512
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 8036 11540 8064 11639
rect 9122 11636 9128 11639
rect 9180 11636 9186 11688
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9398 11676 9404 11688
rect 9263 11648 9404 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9398 11636 9404 11648
rect 9456 11676 9462 11688
rect 12434 11676 12440 11688
rect 9456 11648 12440 11676
rect 9456 11636 9462 11648
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 16666 11636 16672 11688
rect 16724 11636 16730 11688
rect 20346 11636 20352 11688
rect 20404 11636 20410 11688
rect 20438 11636 20444 11688
rect 20496 11636 20502 11688
rect 21928 11676 21956 11716
rect 23293 11679 23351 11685
rect 23293 11676 23305 11679
rect 21560 11648 21956 11676
rect 23124 11648 23305 11676
rect 8386 11568 8392 11620
rect 8444 11608 8450 11620
rect 8665 11611 8723 11617
rect 8665 11608 8677 11611
rect 8444 11580 8677 11608
rect 8444 11568 8450 11580
rect 8665 11577 8677 11580
rect 8711 11577 8723 11611
rect 8665 11571 8723 11577
rect 19794 11568 19800 11620
rect 19852 11608 19858 11620
rect 20806 11608 20812 11620
rect 19852 11580 20812 11608
rect 19852 11568 19858 11580
rect 20806 11568 20812 11580
rect 20864 11608 20870 11620
rect 21560 11617 21588 11648
rect 21545 11611 21603 11617
rect 21545 11608 21557 11611
rect 20864 11580 21557 11608
rect 20864 11568 20870 11580
rect 21545 11577 21557 11580
rect 21591 11577 21603 11611
rect 21545 11571 21603 11577
rect 10318 11540 10324 11552
rect 8036 11512 10324 11540
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 17310 11500 17316 11552
rect 17368 11500 17374 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 19576 11512 19901 11540
rect 19576 11500 19582 11512
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 23124 11540 23152 11648
rect 23293 11645 23305 11648
rect 23339 11645 23351 11679
rect 23293 11639 23351 11645
rect 23400 11608 23428 11716
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 25225 11747 25283 11753
rect 25225 11713 25237 11747
rect 25271 11713 25283 11747
rect 25225 11707 25283 11713
rect 23474 11636 23480 11688
rect 23532 11636 23538 11688
rect 24210 11636 24216 11688
rect 24268 11636 24274 11688
rect 24302 11636 24308 11688
rect 24360 11685 24366 11688
rect 24360 11679 24388 11685
rect 24376 11645 24388 11679
rect 24504 11676 24532 11707
rect 24670 11676 24676 11688
rect 24504 11648 24676 11676
rect 24360 11639 24388 11645
rect 24360 11636 24366 11639
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 24854 11636 24860 11688
rect 24912 11676 24918 11688
rect 25332 11676 25360 11852
rect 25590 11840 25596 11852
rect 25648 11840 25654 11892
rect 26786 11840 26792 11892
rect 26844 11840 26850 11892
rect 29730 11840 29736 11892
rect 29788 11880 29794 11892
rect 30009 11883 30067 11889
rect 30009 11880 30021 11883
rect 29788 11852 30021 11880
rect 29788 11840 29794 11852
rect 30009 11849 30021 11852
rect 30055 11849 30067 11883
rect 30009 11843 30067 11849
rect 30374 11840 30380 11892
rect 30432 11840 30438 11892
rect 30469 11883 30527 11889
rect 30469 11849 30481 11883
rect 30515 11880 30527 11883
rect 31018 11880 31024 11892
rect 30515 11852 31024 11880
rect 30515 11849 30527 11852
rect 30469 11843 30527 11849
rect 31018 11840 31024 11852
rect 31076 11840 31082 11892
rect 31110 11840 31116 11892
rect 31168 11880 31174 11892
rect 31481 11883 31539 11889
rect 31481 11880 31493 11883
rect 31168 11852 31493 11880
rect 31168 11840 31174 11852
rect 31481 11849 31493 11852
rect 31527 11880 31539 11883
rect 32306 11880 32312 11892
rect 31527 11852 32312 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 32306 11840 32312 11852
rect 32364 11840 32370 11892
rect 34333 11883 34391 11889
rect 34333 11849 34345 11883
rect 34379 11880 34391 11883
rect 35342 11880 35348 11892
rect 34379 11852 35348 11880
rect 34379 11849 34391 11852
rect 34333 11843 34391 11849
rect 35342 11840 35348 11852
rect 35400 11840 35406 11892
rect 35986 11840 35992 11892
rect 36044 11840 36050 11892
rect 36280 11852 38792 11880
rect 25492 11815 25550 11821
rect 25492 11781 25504 11815
rect 25538 11812 25550 11815
rect 26804 11812 26832 11840
rect 25538 11784 26832 11812
rect 33413 11815 33471 11821
rect 25538 11781 25550 11784
rect 25492 11775 25550 11781
rect 33413 11781 33425 11815
rect 33459 11812 33471 11815
rect 35713 11815 35771 11821
rect 33459 11784 35388 11812
rect 33459 11781 33471 11784
rect 33413 11775 33471 11781
rect 26418 11704 26424 11756
rect 26476 11744 26482 11756
rect 29825 11747 29883 11753
rect 29825 11744 29837 11747
rect 26476 11716 29837 11744
rect 26476 11704 26482 11716
rect 29825 11713 29837 11716
rect 29871 11744 29883 11747
rect 33505 11747 33563 11753
rect 29871 11716 30604 11744
rect 29871 11713 29883 11716
rect 29825 11707 29883 11713
rect 24912 11648 25360 11676
rect 28353 11679 28411 11685
rect 24912 11636 24918 11648
rect 28353 11645 28365 11679
rect 28399 11676 28411 11679
rect 28718 11676 28724 11688
rect 28399 11648 28724 11676
rect 28399 11645 28411 11648
rect 28353 11639 28411 11645
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 30576 11685 30604 11716
rect 33505 11713 33517 11747
rect 33551 11744 33563 11747
rect 34241 11747 34299 11753
rect 34241 11744 34253 11747
rect 33551 11716 34253 11744
rect 33551 11713 33563 11716
rect 33505 11707 33563 11713
rect 34241 11713 34253 11716
rect 34287 11744 34299 11747
rect 34330 11744 34336 11756
rect 34287 11716 34336 11744
rect 34287 11713 34299 11716
rect 34241 11707 34299 11713
rect 34330 11704 34336 11716
rect 34388 11704 34394 11756
rect 35360 11753 35388 11784
rect 35713 11781 35725 11815
rect 35759 11812 35771 11815
rect 36280 11812 36308 11852
rect 38764 11824 38792 11852
rect 42150 11840 42156 11892
rect 42208 11840 42214 11892
rect 42429 11883 42487 11889
rect 42429 11849 42441 11883
rect 42475 11849 42487 11883
rect 42429 11843 42487 11849
rect 36814 11812 36820 11824
rect 35759 11784 36308 11812
rect 36372 11784 36820 11812
rect 35759 11781 35771 11784
rect 35713 11775 35771 11781
rect 36372 11756 36400 11784
rect 36814 11772 36820 11784
rect 36872 11772 36878 11824
rect 38746 11772 38752 11824
rect 38804 11772 38810 11824
rect 39669 11815 39727 11821
rect 39669 11781 39681 11815
rect 39715 11812 39727 11815
rect 40218 11812 40224 11824
rect 39715 11784 40224 11812
rect 39715 11781 39727 11784
rect 39669 11775 39727 11781
rect 40218 11772 40224 11784
rect 40276 11772 40282 11824
rect 35345 11747 35403 11753
rect 35345 11713 35357 11747
rect 35391 11713 35403 11747
rect 35345 11707 35403 11713
rect 36354 11704 36360 11756
rect 36412 11704 36418 11756
rect 36449 11747 36507 11753
rect 36449 11713 36461 11747
rect 36495 11744 36507 11747
rect 37921 11747 37979 11753
rect 37921 11744 37933 11747
rect 36495 11716 37933 11744
rect 36495 11713 36507 11716
rect 36449 11707 36507 11713
rect 37921 11713 37933 11716
rect 37967 11713 37979 11747
rect 37921 11707 37979 11713
rect 39577 11747 39635 11753
rect 39577 11713 39589 11747
rect 39623 11744 39635 11747
rect 40494 11744 40500 11756
rect 39623 11716 40500 11744
rect 39623 11713 39635 11716
rect 39577 11707 39635 11713
rect 40494 11704 40500 11716
rect 40552 11704 40558 11756
rect 42168 11744 42196 11840
rect 42444 11812 42472 11843
rect 42794 11840 42800 11892
rect 42852 11840 42858 11892
rect 43898 11840 43904 11892
rect 43956 11840 43962 11892
rect 45002 11840 45008 11892
rect 45060 11840 45066 11892
rect 45189 11883 45247 11889
rect 45189 11849 45201 11883
rect 45235 11880 45247 11883
rect 45278 11880 45284 11892
rect 45235 11852 45284 11880
rect 45235 11849 45247 11852
rect 45189 11843 45247 11849
rect 45278 11840 45284 11852
rect 45336 11840 45342 11892
rect 45646 11840 45652 11892
rect 45704 11880 45710 11892
rect 46382 11880 46388 11892
rect 45704 11852 46388 11880
rect 45704 11840 45710 11852
rect 46382 11840 46388 11852
rect 46440 11840 46446 11892
rect 47121 11883 47179 11889
rect 47121 11849 47133 11883
rect 47167 11880 47179 11883
rect 47210 11880 47216 11892
rect 47167 11852 47216 11880
rect 47167 11849 47179 11852
rect 47121 11843 47179 11849
rect 47210 11840 47216 11852
rect 47268 11840 47274 11892
rect 47394 11840 47400 11892
rect 47452 11840 47458 11892
rect 49326 11840 49332 11892
rect 49384 11840 49390 11892
rect 49878 11840 49884 11892
rect 49936 11840 49942 11892
rect 50617 11883 50675 11889
rect 50617 11849 50629 11883
rect 50663 11880 50675 11883
rect 50982 11880 50988 11892
rect 50663 11852 50988 11880
rect 50663 11849 50675 11852
rect 50617 11843 50675 11849
rect 43162 11812 43168 11824
rect 42444 11784 43168 11812
rect 43162 11772 43168 11784
rect 43220 11772 43226 11824
rect 43993 11747 44051 11753
rect 43993 11744 44005 11747
rect 42168 11716 44005 11744
rect 43993 11713 44005 11716
rect 44039 11713 44051 11747
rect 45020 11744 45048 11840
rect 45557 11815 45615 11821
rect 45557 11781 45569 11815
rect 45603 11812 45615 11815
rect 47412 11812 47440 11840
rect 45603 11784 47440 11812
rect 47848 11815 47906 11821
rect 45603 11781 45615 11784
rect 45557 11775 45615 11781
rect 47848 11781 47860 11815
rect 47894 11812 47906 11815
rect 49896 11812 49924 11840
rect 47894 11784 49924 11812
rect 47894 11781 47906 11784
rect 47848 11775 47906 11781
rect 46477 11747 46535 11753
rect 45020 11716 45784 11744
rect 43993 11707 44051 11713
rect 30561 11679 30619 11685
rect 30561 11645 30573 11679
rect 30607 11645 30619 11679
rect 30561 11639 30619 11645
rect 32401 11679 32459 11685
rect 32401 11645 32413 11679
rect 32447 11676 32459 11679
rect 33689 11679 33747 11685
rect 32447 11648 33088 11676
rect 32447 11645 32459 11648
rect 32401 11639 32459 11645
rect 23937 11611 23995 11617
rect 23937 11608 23949 11611
rect 23400 11580 23949 11608
rect 23937 11577 23949 11580
rect 23983 11608 23995 11611
rect 24026 11608 24032 11620
rect 23983 11580 24032 11608
rect 23983 11577 23995 11580
rect 23937 11571 23995 11577
rect 24026 11568 24032 11580
rect 24084 11568 24090 11620
rect 33060 11617 33088 11648
rect 33689 11645 33701 11679
rect 33735 11676 33747 11679
rect 34146 11676 34152 11688
rect 33735 11648 34152 11676
rect 33735 11645 33747 11648
rect 33689 11639 33747 11645
rect 34146 11636 34152 11648
rect 34204 11636 34210 11688
rect 34422 11636 34428 11688
rect 34480 11636 34486 11688
rect 34701 11679 34759 11685
rect 34701 11645 34713 11679
rect 34747 11645 34759 11679
rect 34701 11639 34759 11645
rect 36633 11679 36691 11685
rect 36633 11645 36645 11679
rect 36679 11676 36691 11679
rect 36679 11648 36860 11676
rect 36679 11645 36691 11648
rect 36633 11639 36691 11645
rect 26605 11611 26663 11617
rect 26605 11577 26617 11611
rect 26651 11577 26663 11611
rect 26605 11571 26663 11577
rect 33045 11611 33103 11617
rect 33045 11577 33057 11611
rect 33091 11577 33103 11611
rect 34716 11608 34744 11639
rect 35066 11608 35072 11620
rect 33045 11571 33103 11577
rect 33796 11580 35072 11608
rect 25038 11540 25044 11552
rect 23124 11512 25044 11540
rect 19889 11503 19947 11509
rect 25038 11500 25044 11512
rect 25096 11540 25102 11552
rect 26620 11540 26648 11571
rect 33796 11552 33824 11580
rect 35066 11568 35072 11580
rect 35124 11568 35130 11620
rect 36832 11552 36860 11648
rect 36906 11636 36912 11688
rect 36964 11676 36970 11688
rect 37277 11679 37335 11685
rect 37277 11676 37289 11679
rect 36964 11648 37289 11676
rect 36964 11636 36970 11648
rect 37277 11645 37289 11648
rect 37323 11645 37335 11679
rect 37277 11639 37335 11645
rect 38565 11679 38623 11685
rect 38565 11645 38577 11679
rect 38611 11645 38623 11679
rect 38565 11639 38623 11645
rect 38580 11608 38608 11639
rect 39022 11636 39028 11688
rect 39080 11676 39086 11688
rect 39761 11679 39819 11685
rect 39761 11676 39773 11679
rect 39080 11648 39773 11676
rect 39080 11636 39086 11648
rect 39761 11645 39773 11648
rect 39807 11645 39819 11679
rect 39761 11639 39819 11645
rect 40034 11636 40040 11688
rect 40092 11636 40098 11688
rect 40773 11679 40831 11685
rect 40773 11676 40785 11679
rect 40236 11648 40785 11676
rect 39209 11611 39267 11617
rect 39209 11608 39221 11611
rect 38580 11580 39221 11608
rect 39209 11577 39221 11580
rect 39255 11577 39267 11611
rect 39209 11571 39267 11577
rect 25096 11512 26648 11540
rect 25096 11500 25102 11512
rect 28902 11500 28908 11552
rect 28960 11500 28966 11552
rect 29270 11500 29276 11552
rect 29328 11500 29334 11552
rect 32950 11500 32956 11552
rect 33008 11500 33014 11552
rect 33778 11500 33784 11552
rect 33836 11500 33842 11552
rect 33870 11500 33876 11552
rect 33928 11500 33934 11552
rect 34514 11500 34520 11552
rect 34572 11540 34578 11552
rect 35434 11540 35440 11552
rect 34572 11512 35440 11540
rect 34572 11500 34578 11512
rect 35434 11500 35440 11512
rect 35492 11500 35498 11552
rect 36814 11500 36820 11552
rect 36872 11540 36878 11552
rect 36998 11540 37004 11552
rect 36872 11512 37004 11540
rect 36872 11500 36878 11512
rect 36998 11500 37004 11512
rect 37056 11500 37062 11552
rect 39114 11500 39120 11552
rect 39172 11500 39178 11552
rect 39666 11500 39672 11552
rect 39724 11540 39730 11552
rect 40236 11540 40264 11648
rect 40773 11645 40785 11648
rect 40819 11676 40831 11679
rect 40819 11648 41920 11676
rect 40819 11645 40831 11648
rect 40773 11639 40831 11645
rect 40310 11568 40316 11620
rect 40368 11608 40374 11620
rect 41417 11611 41475 11617
rect 41417 11608 41429 11611
rect 40368 11580 41429 11608
rect 40368 11568 40374 11580
rect 41417 11577 41429 11580
rect 41463 11577 41475 11611
rect 41417 11571 41475 11577
rect 41892 11552 41920 11648
rect 42794 11636 42800 11688
rect 42852 11676 42858 11688
rect 42889 11679 42947 11685
rect 42889 11676 42901 11679
rect 42852 11648 42901 11676
rect 42852 11636 42858 11648
rect 42889 11645 42901 11648
rect 42935 11645 42947 11679
rect 42889 11639 42947 11645
rect 42978 11636 42984 11688
rect 43036 11636 43042 11688
rect 43349 11679 43407 11685
rect 43349 11645 43361 11679
rect 43395 11676 43407 11679
rect 43806 11676 43812 11688
rect 43395 11648 43812 11676
rect 43395 11645 43407 11648
rect 43349 11639 43407 11645
rect 43806 11636 43812 11648
rect 43864 11636 43870 11688
rect 45756 11685 45784 11716
rect 46477 11713 46489 11747
rect 46523 11744 46535 11747
rect 47026 11744 47032 11756
rect 46523 11716 47032 11744
rect 46523 11713 46535 11716
rect 46477 11707 46535 11713
rect 47026 11704 47032 11716
rect 47084 11704 47090 11756
rect 47302 11704 47308 11756
rect 47360 11744 47366 11756
rect 50632 11744 50660 11843
rect 50982 11840 50988 11852
rect 51040 11840 51046 11892
rect 51077 11883 51135 11889
rect 51077 11849 51089 11883
rect 51123 11880 51135 11883
rect 51166 11880 51172 11892
rect 51123 11852 51172 11880
rect 51123 11849 51135 11852
rect 51077 11843 51135 11849
rect 51166 11840 51172 11852
rect 51224 11840 51230 11892
rect 51537 11883 51595 11889
rect 51537 11849 51549 11883
rect 51583 11880 51595 11883
rect 52362 11880 52368 11892
rect 51583 11852 52368 11880
rect 51583 11849 51595 11852
rect 51537 11843 51595 11849
rect 52362 11840 52368 11852
rect 52420 11840 52426 11892
rect 52733 11883 52791 11889
rect 52733 11849 52745 11883
rect 52779 11880 52791 11883
rect 53006 11880 53012 11892
rect 52779 11852 53012 11880
rect 52779 11849 52791 11852
rect 52733 11843 52791 11849
rect 53006 11840 53012 11852
rect 53064 11840 53070 11892
rect 53101 11883 53159 11889
rect 53101 11849 53113 11883
rect 53147 11880 53159 11883
rect 54386 11880 54392 11892
rect 53147 11852 54392 11880
rect 53147 11849 53159 11852
rect 53101 11843 53159 11849
rect 54386 11840 54392 11852
rect 54444 11840 54450 11892
rect 55122 11840 55128 11892
rect 55180 11840 55186 11892
rect 55309 11883 55367 11889
rect 55309 11849 55321 11883
rect 55355 11849 55367 11883
rect 57698 11880 57704 11892
rect 55309 11843 55367 11849
rect 55968 11852 57704 11880
rect 54196 11815 54254 11821
rect 51920 11784 54064 11812
rect 47360 11716 50660 11744
rect 47360 11704 47366 11716
rect 51258 11704 51264 11756
rect 51316 11744 51322 11756
rect 51445 11747 51503 11753
rect 51445 11744 51457 11747
rect 51316 11716 51457 11744
rect 51316 11704 51322 11716
rect 51445 11713 51457 11716
rect 51491 11713 51503 11747
rect 51920 11744 51948 11784
rect 53193 11747 53251 11753
rect 53193 11744 53205 11747
rect 51445 11707 51503 11713
rect 51736 11716 51948 11744
rect 52104 11716 53205 11744
rect 45741 11679 45799 11685
rect 45741 11645 45753 11679
rect 45787 11645 45799 11679
rect 45741 11639 45799 11645
rect 46661 11679 46719 11685
rect 46661 11645 46673 11679
rect 46707 11676 46719 11679
rect 47210 11676 47216 11688
rect 46707 11648 47216 11676
rect 46707 11645 46719 11648
rect 46661 11639 46719 11645
rect 47210 11636 47216 11648
rect 47268 11636 47274 11688
rect 47578 11676 47584 11688
rect 47320 11648 47584 11676
rect 47320 11608 47348 11648
rect 47578 11636 47584 11648
rect 47636 11636 47642 11688
rect 51736 11685 51764 11716
rect 52104 11688 52132 11716
rect 53193 11713 53205 11716
rect 53239 11744 53251 11747
rect 53466 11744 53472 11756
rect 53239 11716 53472 11744
rect 53239 11713 53251 11716
rect 53193 11707 53251 11713
rect 53466 11704 53472 11716
rect 53524 11704 53530 11756
rect 53742 11704 53748 11756
rect 53800 11704 53806 11756
rect 53834 11704 53840 11756
rect 53892 11744 53898 11756
rect 53929 11747 53987 11753
rect 53929 11744 53941 11747
rect 53892 11716 53941 11744
rect 53892 11704 53898 11716
rect 53929 11713 53941 11716
rect 53975 11713 53987 11747
rect 54036 11744 54064 11784
rect 54196 11781 54208 11815
rect 54242 11812 54254 11815
rect 55140 11812 55168 11840
rect 54242 11784 55168 11812
rect 54242 11781 54254 11784
rect 54196 11775 54254 11781
rect 55324 11756 55352 11843
rect 54036 11716 54984 11744
rect 53929 11707 53987 11713
rect 51721 11679 51779 11685
rect 51721 11645 51733 11679
rect 51767 11645 51779 11679
rect 51721 11639 51779 11645
rect 51736 11608 51764 11639
rect 51994 11636 52000 11688
rect 52052 11636 52058 11688
rect 52086 11636 52092 11688
rect 52144 11636 52150 11688
rect 53374 11636 53380 11688
rect 53432 11676 53438 11688
rect 53760 11676 53788 11704
rect 53432 11648 53788 11676
rect 53432 11636 53438 11648
rect 54956 11608 54984 11716
rect 55306 11704 55312 11756
rect 55364 11704 55370 11756
rect 55968 11753 55996 11852
rect 57698 11840 57704 11852
rect 57756 11840 57762 11892
rect 55953 11747 56011 11753
rect 55953 11713 55965 11747
rect 55999 11713 56011 11747
rect 55953 11707 56011 11713
rect 56686 11704 56692 11756
rect 56744 11704 56750 11756
rect 56778 11704 56784 11756
rect 56836 11753 56842 11756
rect 56836 11747 56864 11753
rect 56852 11713 56864 11747
rect 56836 11707 56864 11713
rect 56836 11704 56842 11707
rect 55674 11636 55680 11688
rect 55732 11636 55738 11688
rect 55769 11679 55827 11685
rect 55769 11645 55781 11679
rect 55815 11676 55827 11679
rect 56965 11679 57023 11685
rect 55815 11648 56573 11676
rect 55815 11645 55827 11648
rect 55769 11639 55827 11645
rect 55692 11608 55720 11636
rect 42904 11580 47348 11608
rect 51046 11580 51764 11608
rect 52288 11580 52684 11608
rect 54956 11580 55720 11608
rect 42904 11552 42932 11580
rect 39724 11512 40264 11540
rect 39724 11500 39730 11512
rect 40678 11500 40684 11552
rect 40736 11500 40742 11552
rect 41874 11500 41880 11552
rect 41932 11500 41938 11552
rect 42242 11500 42248 11552
rect 42300 11540 42306 11552
rect 42610 11540 42616 11552
rect 42300 11512 42616 11540
rect 42300 11500 42306 11512
rect 42610 11500 42616 11512
rect 42668 11500 42674 11552
rect 42886 11500 42892 11552
rect 42944 11500 42950 11552
rect 43622 11500 43628 11552
rect 43680 11540 43686 11552
rect 44637 11543 44695 11549
rect 44637 11540 44649 11543
rect 43680 11512 44649 11540
rect 43680 11500 43686 11512
rect 44637 11509 44649 11512
rect 44683 11509 44695 11543
rect 44637 11503 44695 11509
rect 46014 11500 46020 11552
rect 46072 11500 46078 11552
rect 46934 11500 46940 11552
rect 46992 11540 46998 11552
rect 47946 11540 47952 11552
rect 46992 11512 47952 11540
rect 46992 11500 46998 11512
rect 47946 11500 47952 11512
rect 48004 11540 48010 11552
rect 48961 11543 49019 11549
rect 48961 11540 48973 11543
rect 48004 11512 48973 11540
rect 48004 11500 48010 11512
rect 48961 11509 48973 11512
rect 49007 11509 49019 11543
rect 48961 11503 49019 11509
rect 49142 11500 49148 11552
rect 49200 11540 49206 11552
rect 49602 11540 49608 11552
rect 49200 11512 49608 11540
rect 49200 11500 49206 11512
rect 49602 11500 49608 11512
rect 49660 11540 49666 11552
rect 50893 11543 50951 11549
rect 50893 11540 50905 11543
rect 49660 11512 50905 11540
rect 49660 11500 49666 11512
rect 50893 11509 50905 11512
rect 50939 11540 50951 11543
rect 51046 11540 51074 11580
rect 52288 11552 52316 11580
rect 50939 11512 51074 11540
rect 50939 11509 50951 11512
rect 50893 11503 50951 11509
rect 51166 11500 51172 11552
rect 51224 11540 51230 11552
rect 52270 11540 52276 11552
rect 51224 11512 52276 11540
rect 51224 11500 51230 11512
rect 52270 11500 52276 11512
rect 52328 11500 52334 11552
rect 52546 11500 52552 11552
rect 52604 11500 52610 11552
rect 52656 11540 52684 11580
rect 56134 11568 56140 11620
rect 56192 11608 56198 11620
rect 56413 11611 56471 11617
rect 56413 11608 56425 11611
rect 56192 11580 56425 11608
rect 56192 11568 56198 11580
rect 56413 11577 56425 11580
rect 56459 11577 56471 11611
rect 56413 11571 56471 11577
rect 55582 11540 55588 11552
rect 52656 11512 55588 11540
rect 55582 11500 55588 11512
rect 55640 11500 55646 11552
rect 56545 11540 56573 11648
rect 56965 11645 56977 11679
rect 57011 11676 57023 11679
rect 57330 11676 57336 11688
rect 57011 11648 57336 11676
rect 57011 11645 57023 11648
rect 56965 11639 57023 11645
rect 57330 11636 57336 11648
rect 57388 11636 57394 11688
rect 57146 11540 57152 11552
rect 56545 11512 57152 11540
rect 57146 11500 57152 11512
rect 57204 11500 57210 11552
rect 57606 11500 57612 11552
rect 57664 11500 57670 11552
rect 1104 11450 58880 11472
rect 1104 11398 8172 11450
rect 8224 11398 8236 11450
rect 8288 11398 8300 11450
rect 8352 11398 8364 11450
rect 8416 11398 8428 11450
rect 8480 11398 22616 11450
rect 22668 11398 22680 11450
rect 22732 11398 22744 11450
rect 22796 11398 22808 11450
rect 22860 11398 22872 11450
rect 22924 11398 37060 11450
rect 37112 11398 37124 11450
rect 37176 11398 37188 11450
rect 37240 11398 37252 11450
rect 37304 11398 37316 11450
rect 37368 11398 51504 11450
rect 51556 11398 51568 11450
rect 51620 11398 51632 11450
rect 51684 11398 51696 11450
rect 51748 11398 51760 11450
rect 51812 11398 58880 11450
rect 1104 11376 58880 11398
rect 2866 11296 2872 11348
rect 2924 11296 2930 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 3234 11336 3240 11348
rect 3099 11308 3240 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3970 11296 3976 11348
rect 4028 11296 4034 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4212 11308 4537 11336
rect 4212 11296 4218 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 4614 11296 4620 11348
rect 4672 11296 4678 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8018 11336 8024 11348
rect 7699 11308 8024 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 8018 11296 8024 11308
rect 8076 11336 8082 11348
rect 9122 11336 9128 11348
rect 8076 11308 9128 11336
rect 8076 11296 8082 11308
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 10318 11296 10324 11348
rect 10376 11296 10382 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 10468 11308 11989 11336
rect 10468 11296 10474 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 17310 11296 17316 11348
rect 17368 11296 17374 11348
rect 19061 11339 19119 11345
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19334 11336 19340 11348
rect 19107 11308 19340 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 21634 11296 21640 11348
rect 21692 11296 21698 11348
rect 23109 11339 23167 11345
rect 23109 11305 23121 11339
rect 23155 11336 23167 11339
rect 23382 11336 23388 11348
rect 23155 11308 23388 11336
rect 23155 11305 23167 11308
rect 23109 11299 23167 11305
rect 23382 11296 23388 11308
rect 23440 11336 23446 11348
rect 24302 11336 24308 11348
rect 23440 11308 24308 11336
rect 23440 11296 23446 11308
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 24412 11308 25789 11336
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 3200 11240 3372 11268
rect 3200 11228 3206 11240
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3237 11203 3295 11209
rect 3237 11200 3249 11203
rect 3108 11172 3249 11200
rect 3108 11160 3114 11172
rect 3237 11169 3249 11172
rect 3283 11169 3295 11203
rect 3344 11200 3372 11240
rect 3510 11228 3516 11280
rect 3568 11268 3574 11280
rect 3568 11240 4568 11268
rect 3568 11228 3574 11240
rect 3602 11200 3608 11212
rect 3344 11172 3608 11200
rect 3237 11163 3295 11169
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 3436 11141 3464 11172
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3936 11172 4077 11200
rect 3936 11160 3942 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4304 11172 4476 11200
rect 4304 11160 4310 11172
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3329 11135 3387 11141
rect 3007 11104 3096 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3068 11008 3096 11104
rect 3329 11101 3341 11135
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 3344 11064 3372 11095
rect 3510 11092 3516 11144
rect 3568 11092 3574 11144
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4448 11141 4476 11172
rect 4540 11141 4568 11240
rect 4632 11200 4660 11296
rect 4801 11203 4859 11209
rect 4801 11200 4813 11203
rect 4632 11172 4813 11200
rect 4801 11169 4813 11172
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 8386 11160 8392 11212
rect 8444 11160 8450 11212
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8628 11172 8953 11200
rect 8628 11160 8634 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 10336 11200 10364 11296
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 10336 11172 10425 11200
rect 8941 11163 8999 11169
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 14921 11203 14979 11209
rect 14921 11200 14933 11203
rect 13872 11172 14933 11200
rect 13872 11160 13878 11172
rect 14921 11169 14933 11172
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11132 6331 11135
rect 6914 11132 6920 11144
rect 6319 11104 6920 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 12250 11132 12256 11144
rect 11471 11104 12256 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 14185 11135 14243 11141
rect 14185 11101 14197 11135
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 6540 11067 6598 11073
rect 3200 11036 4660 11064
rect 3200 11024 3206 11036
rect 3050 10956 3056 11008
rect 3108 10956 3114 11008
rect 4338 10956 4344 11008
rect 4396 10956 4402 11008
rect 4632 11005 4660 11036
rect 6540 11033 6552 11067
rect 6586 11064 6598 11067
rect 7834 11064 7840 11076
rect 6586 11036 7840 11064
rect 6586 11033 6598 11036
rect 6540 11027 6598 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8113 11067 8171 11073
rect 8113 11033 8125 11067
rect 8159 11064 8171 11067
rect 8570 11064 8576 11076
rect 8159 11036 8576 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 9208 11067 9266 11073
rect 9208 11033 9220 11067
rect 9254 11064 9266 11067
rect 10502 11064 10508 11076
rect 9254 11036 10508 11064
rect 9254 11033 9266 11036
rect 9208 11027 9266 11033
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 13262 11064 13268 11076
rect 12492 11036 13268 11064
rect 12492 11024 12498 11036
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 4617 10999 4675 11005
rect 4617 10965 4629 10999
rect 4663 10996 4675 10999
rect 4982 10996 4988 11008
rect 4663 10968 4988 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 7742 10956 7748 11008
rect 7800 10956 7806 11008
rect 8205 10999 8263 11005
rect 8205 10965 8217 10999
rect 8251 10996 8263 10999
rect 8662 10996 8668 11008
rect 8251 10968 8668 10996
rect 8251 10965 8263 10968
rect 8205 10959 8263 10965
rect 8662 10956 8668 10968
rect 8720 10996 8726 11008
rect 9398 10996 9404 11008
rect 8720 10968 9404 10996
rect 8720 10956 8726 10968
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 11054 10956 11060 11008
rect 11112 10956 11118 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 14200 10996 14228 11095
rect 15102 11092 15108 11144
rect 15160 11132 15166 11144
rect 15838 11132 15844 11144
rect 15160 11104 15844 11132
rect 15160 11092 15166 11104
rect 15838 11092 15844 11104
rect 15896 11132 15902 11144
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15896 11104 15945 11132
rect 15896 11092 15902 11104
rect 15933 11101 15945 11104
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16200 11135 16258 11141
rect 16200 11101 16212 11135
rect 16246 11132 16258 11135
rect 17328 11132 17356 11296
rect 19352 11209 19380 11296
rect 20438 11228 20444 11280
rect 20496 11268 20502 11280
rect 20717 11271 20775 11277
rect 20717 11268 20729 11271
rect 20496 11240 20729 11268
rect 20496 11228 20502 11240
rect 20717 11237 20729 11240
rect 20763 11237 20775 11271
rect 20717 11231 20775 11237
rect 19337 11203 19395 11209
rect 19337 11169 19349 11203
rect 19383 11169 19395 11203
rect 21652 11200 21680 11296
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24412 11268 24440 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 25777 11299 25835 11305
rect 23532 11240 24440 11268
rect 23532 11228 23538 11240
rect 21729 11203 21787 11209
rect 21729 11200 21741 11203
rect 21652 11172 21741 11200
rect 19337 11163 19395 11169
rect 21729 11169 21741 11172
rect 21775 11169 21787 11203
rect 21729 11163 21787 11169
rect 16246 11104 17356 11132
rect 17497 11135 17555 11141
rect 16246 11101 16258 11104
rect 16200 11095 16258 11101
rect 17497 11101 17509 11135
rect 17543 11132 17555 11135
rect 18782 11132 18788 11144
rect 17543 11104 18788 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 17512 11064 17540 11095
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 21744 11132 21772 11163
rect 23750 11160 23756 11212
rect 23808 11160 23814 11212
rect 25792 11200 25820 11299
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29730 11336 29736 11348
rect 29052 11308 29736 11336
rect 29052 11296 29058 11308
rect 29730 11296 29736 11308
rect 29788 11296 29794 11348
rect 33778 11296 33784 11348
rect 33836 11296 33842 11348
rect 33870 11296 33876 11348
rect 33928 11296 33934 11348
rect 36262 11336 36268 11348
rect 34900 11308 36268 11336
rect 33888 11209 33916 11296
rect 34900 11209 34928 11308
rect 36262 11296 36268 11308
rect 36320 11296 36326 11348
rect 37458 11296 37464 11348
rect 37516 11336 37522 11348
rect 37516 11308 37688 11336
rect 37516 11296 37522 11308
rect 35066 11228 35072 11280
rect 35124 11268 35130 11280
rect 36633 11271 36691 11277
rect 35124 11240 35480 11268
rect 35124 11228 35130 11240
rect 25869 11203 25927 11209
rect 25869 11200 25881 11203
rect 25792 11172 25881 11200
rect 25869 11169 25881 11172
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 33873 11203 33931 11209
rect 33873 11169 33885 11203
rect 33919 11169 33931 11203
rect 33873 11163 33931 11169
rect 34885 11203 34943 11209
rect 34885 11169 34897 11203
rect 34931 11169 34943 11203
rect 34885 11163 34943 11169
rect 34974 11160 34980 11212
rect 35032 11200 35038 11212
rect 35345 11203 35403 11209
rect 35345 11200 35357 11203
rect 35032 11172 35357 11200
rect 35032 11160 35038 11172
rect 35345 11169 35357 11172
rect 35391 11169 35403 11203
rect 35452 11200 35480 11240
rect 36633 11237 36645 11271
rect 36679 11268 36691 11271
rect 37550 11268 37556 11280
rect 36679 11240 37556 11268
rect 36679 11237 36691 11240
rect 36633 11231 36691 11237
rect 37550 11228 37556 11240
rect 37608 11228 37614 11280
rect 35738 11203 35796 11209
rect 35738 11200 35750 11203
rect 35452 11172 35750 11200
rect 35345 11163 35403 11169
rect 35738 11169 35750 11172
rect 35784 11169 35796 11203
rect 35738 11163 35796 11169
rect 35894 11160 35900 11212
rect 35952 11200 35958 11212
rect 36078 11200 36084 11212
rect 35952 11172 36084 11200
rect 35952 11160 35958 11172
rect 36078 11160 36084 11172
rect 36136 11160 36142 11212
rect 36538 11160 36544 11212
rect 36596 11200 36602 11212
rect 37093 11203 37151 11209
rect 37093 11200 37105 11203
rect 36596 11172 37105 11200
rect 36596 11160 36602 11172
rect 37093 11169 37105 11172
rect 37139 11169 37151 11203
rect 37093 11163 37151 11169
rect 37185 11203 37243 11209
rect 37185 11169 37197 11203
rect 37231 11200 37243 11203
rect 37660 11200 37688 11308
rect 39666 11296 39672 11348
rect 39724 11296 39730 11348
rect 39853 11339 39911 11345
rect 39853 11305 39865 11339
rect 39899 11336 39911 11339
rect 40034 11336 40040 11348
rect 39899 11308 40040 11336
rect 39899 11305 39911 11308
rect 39853 11299 39911 11305
rect 40034 11296 40040 11308
rect 40092 11296 40098 11348
rect 40310 11296 40316 11348
rect 40368 11296 40374 11348
rect 40678 11296 40684 11348
rect 40736 11296 40742 11348
rect 40954 11296 40960 11348
rect 41012 11336 41018 11348
rect 41012 11308 41644 11336
rect 41012 11296 41018 11308
rect 37231 11172 37688 11200
rect 37231 11169 37243 11172
rect 37185 11163 37243 11169
rect 38286 11160 38292 11212
rect 38344 11160 38350 11212
rect 40328 11209 40356 11296
rect 40313 11203 40371 11209
rect 40313 11169 40325 11203
rect 40359 11169 40371 11203
rect 40313 11163 40371 11169
rect 40402 11160 40408 11212
rect 40460 11160 40466 11212
rect 24397 11135 24455 11141
rect 24397 11132 24409 11135
rect 21744 11104 24409 11132
rect 24397 11101 24409 11104
rect 24443 11132 24455 11135
rect 24486 11132 24492 11144
rect 24443 11104 24492 11132
rect 24443 11101 24455 11104
rect 24397 11095 24455 11101
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 25222 11132 25228 11144
rect 24596 11104 25228 11132
rect 17328 11036 17540 11064
rect 19604 11067 19662 11073
rect 14274 10996 14280 11008
rect 12676 10968 14280 10996
rect 12676 10956 12682 10968
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 14826 10956 14832 11008
rect 14884 10956 14890 11008
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 17328 11005 17356 11036
rect 19604 11033 19616 11067
rect 19650 11064 19662 11067
rect 21266 11064 21272 11076
rect 19650 11036 21272 11064
rect 19650 11033 19662 11036
rect 19604 11027 19662 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 21996 11067 22054 11073
rect 21996 11033 22008 11067
rect 22042 11064 22054 11067
rect 23290 11064 23296 11076
rect 22042 11036 23296 11064
rect 22042 11033 22054 11036
rect 21996 11027 22054 11033
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 23661 11067 23719 11073
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 24596 11064 24624 11104
rect 25222 11092 25228 11104
rect 25280 11092 25286 11144
rect 27798 11092 27804 11144
rect 27856 11092 27862 11144
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11132 28595 11135
rect 28626 11132 28632 11144
rect 28583 11104 28632 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 32401 11135 32459 11141
rect 32401 11101 32413 11135
rect 32447 11132 32459 11135
rect 32490 11132 32496 11144
rect 32447 11104 32496 11132
rect 32447 11101 32459 11104
rect 32401 11095 32459 11101
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 32668 11135 32726 11141
rect 32668 11101 32680 11135
rect 32714 11132 32726 11135
rect 32950 11132 32956 11144
rect 32714 11104 32956 11132
rect 32714 11101 32726 11104
rect 32668 11095 32726 11101
rect 32950 11092 32956 11104
rect 33008 11092 33014 11144
rect 34701 11135 34759 11141
rect 34701 11101 34713 11135
rect 34747 11132 34759 11135
rect 35066 11132 35072 11144
rect 34747 11104 35072 11132
rect 34747 11101 34759 11104
rect 34701 11095 34759 11101
rect 35066 11092 35072 11104
rect 35124 11092 35130 11144
rect 35618 11092 35624 11144
rect 35676 11092 35682 11144
rect 37458 11092 37464 11144
rect 37516 11092 37522 11144
rect 38556 11135 38614 11141
rect 38556 11101 38568 11135
rect 38602 11132 38614 11135
rect 40696 11132 40724 11296
rect 41616 11277 41644 11308
rect 41708 11308 42564 11336
rect 41601 11271 41659 11277
rect 40972 11240 41414 11268
rect 40972 11209 41000 11240
rect 40957 11203 41015 11209
rect 40957 11169 40969 11203
rect 41003 11169 41015 11203
rect 41386 11200 41414 11240
rect 41601 11237 41613 11271
rect 41647 11237 41659 11271
rect 41601 11231 41659 11237
rect 41708 11200 41736 11308
rect 42536 11268 42564 11308
rect 42794 11296 42800 11348
rect 42852 11296 42858 11348
rect 43806 11336 43812 11348
rect 42904 11308 43812 11336
rect 42904 11268 42932 11308
rect 43806 11296 43812 11308
rect 43864 11296 43870 11348
rect 47578 11296 47584 11348
rect 47636 11336 47642 11348
rect 50154 11336 50160 11348
rect 47636 11308 50160 11336
rect 47636 11296 47642 11308
rect 50154 11296 50160 11308
rect 50212 11296 50218 11348
rect 52546 11336 52552 11348
rect 51276 11308 52552 11336
rect 42536 11240 42932 11268
rect 44082 11228 44088 11280
rect 44140 11268 44146 11280
rect 44269 11271 44327 11277
rect 44269 11268 44281 11271
rect 44140 11240 44281 11268
rect 44140 11228 44146 11240
rect 44269 11237 44281 11240
rect 44315 11237 44327 11271
rect 44269 11231 44327 11237
rect 46385 11271 46443 11277
rect 46385 11237 46397 11271
rect 46431 11268 46443 11271
rect 46842 11268 46848 11280
rect 46431 11240 46848 11268
rect 46431 11237 46443 11240
rect 46385 11231 46443 11237
rect 46842 11228 46848 11240
rect 46900 11268 46906 11280
rect 46900 11240 47348 11268
rect 46900 11228 46906 11240
rect 40957 11163 41015 11169
rect 41064 11172 41276 11200
rect 41386 11172 41736 11200
rect 38602 11104 40724 11132
rect 38602 11101 38614 11104
rect 38556 11095 38614 11101
rect 23707 11036 24624 11064
rect 24664 11067 24722 11073
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 24664 11033 24676 11067
rect 24710 11064 24722 11067
rect 25682 11064 25688 11076
rect 24710 11036 25688 11064
rect 24710 11033 24722 11036
rect 24664 11027 24722 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 28994 11024 29000 11076
rect 29052 11064 29058 11076
rect 29089 11067 29147 11073
rect 29089 11064 29101 11067
rect 29052 11036 29101 11064
rect 29052 11024 29058 11036
rect 29089 11033 29101 11036
rect 29135 11033 29147 11067
rect 29089 11027 29147 11033
rect 30300 11036 33548 11064
rect 30300 11008 30328 11036
rect 15565 10999 15623 11005
rect 15565 10996 15577 10999
rect 15252 10968 15577 10996
rect 15252 10956 15258 10968
rect 15565 10965 15577 10968
rect 15611 10965 15623 10999
rect 15565 10959 15623 10965
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10965 17371 10999
rect 17313 10959 17371 10965
rect 18046 10956 18052 11008
rect 18104 10956 18110 11008
rect 18414 10956 18420 11008
rect 18472 10956 18478 11008
rect 23198 10956 23204 11008
rect 23256 10956 23262 11008
rect 23566 10956 23572 11008
rect 23624 10956 23630 11008
rect 26510 10956 26516 11008
rect 26568 10956 26574 11008
rect 28350 10956 28356 11008
rect 28408 10956 28414 11008
rect 30193 10999 30251 11005
rect 30193 10965 30205 10999
rect 30239 10996 30251 10999
rect 30282 10996 30288 11008
rect 30239 10968 30288 10996
rect 30239 10965 30251 10968
rect 30193 10959 30251 10965
rect 30282 10956 30288 10968
rect 30340 10956 30346 11008
rect 33520 10996 33548 11036
rect 33594 11024 33600 11076
rect 33652 11064 33658 11076
rect 34517 11067 34575 11073
rect 34517 11064 34529 11067
rect 33652 11036 34529 11064
rect 33652 11024 33658 11036
rect 34517 11033 34529 11036
rect 34563 11033 34575 11067
rect 34517 11027 34575 11033
rect 34606 11024 34612 11076
rect 34664 11024 34670 11076
rect 36541 11067 36599 11073
rect 36541 11033 36553 11067
rect 36587 11064 36599 11067
rect 37001 11067 37059 11073
rect 37001 11064 37013 11067
rect 36587 11036 37013 11064
rect 36587 11033 36599 11036
rect 36541 11027 36599 11033
rect 37001 11033 37013 11036
rect 37047 11033 37059 11067
rect 37001 11027 37059 11033
rect 38028 11036 38608 11064
rect 34422 10996 34428 11008
rect 33520 10968 34428 10996
rect 34422 10956 34428 10968
rect 34480 10956 34486 11008
rect 34624 10996 34652 11024
rect 35618 10996 35624 11008
rect 34624 10968 35624 10996
rect 35618 10956 35624 10968
rect 35676 10956 35682 11008
rect 35710 10956 35716 11008
rect 35768 10996 35774 11008
rect 38028 10996 38056 11036
rect 35768 10968 38056 10996
rect 35768 10956 35774 10968
rect 38102 10956 38108 11008
rect 38160 10956 38166 11008
rect 38580 10996 38608 11036
rect 40218 11024 40224 11076
rect 40276 11064 40282 11076
rect 41064 11064 41092 11172
rect 41141 11135 41199 11141
rect 41141 11101 41153 11135
rect 41187 11101 41199 11135
rect 41248 11132 41276 11172
rect 41874 11160 41880 11212
rect 41932 11160 41938 11212
rect 42886 11160 42892 11212
rect 42944 11160 42950 11212
rect 46569 11203 46627 11209
rect 46569 11169 46581 11203
rect 46615 11200 46627 11203
rect 47118 11200 47124 11212
rect 46615 11172 47124 11200
rect 46615 11169 46627 11172
rect 46569 11163 46627 11169
rect 47118 11160 47124 11172
rect 47176 11160 47182 11212
rect 47210 11160 47216 11212
rect 47268 11160 47274 11212
rect 47320 11200 47348 11240
rect 48222 11228 48228 11280
rect 48280 11268 48286 11280
rect 48409 11271 48467 11277
rect 48409 11268 48421 11271
rect 48280 11240 48421 11268
rect 48280 11228 48286 11240
rect 48409 11237 48421 11240
rect 48455 11237 48467 11271
rect 48409 11231 48467 11237
rect 48501 11271 48559 11277
rect 48501 11237 48513 11271
rect 48547 11268 48559 11271
rect 48547 11240 49372 11268
rect 48547 11237 48559 11240
rect 48501 11231 48559 11237
rect 47606 11203 47664 11209
rect 47606 11200 47618 11203
rect 47320 11172 47618 11200
rect 47606 11169 47618 11172
rect 47652 11169 47664 11203
rect 47606 11163 47664 11169
rect 47765 11203 47823 11209
rect 47765 11169 47777 11203
rect 47811 11200 47823 11203
rect 47946 11200 47952 11212
rect 47811 11172 47952 11200
rect 47811 11169 47823 11172
rect 47765 11163 47823 11169
rect 47946 11160 47952 11172
rect 48004 11160 48010 11212
rect 48958 11200 48964 11212
rect 48792 11172 48964 11200
rect 41322 11132 41328 11144
rect 41248 11104 41328 11132
rect 41141 11095 41199 11101
rect 40276 11036 41092 11064
rect 40276 11024 40282 11036
rect 38838 10996 38844 11008
rect 38580 10968 38844 10996
rect 38838 10956 38844 10968
rect 38896 10996 38902 11008
rect 39850 10996 39856 11008
rect 38896 10968 39856 10996
rect 38896 10956 38902 10968
rect 39850 10956 39856 10968
rect 39908 10996 39914 11008
rect 40402 10996 40408 11008
rect 39908 10968 40408 10996
rect 39908 10956 39914 10968
rect 40402 10956 40408 10968
rect 40460 10956 40466 11008
rect 41156 10996 41184 11095
rect 41322 11092 41328 11104
rect 41380 11092 41386 11144
rect 41966 11092 41972 11144
rect 42024 11141 42030 11144
rect 42024 11135 42052 11141
rect 42040 11101 42052 11135
rect 42024 11095 42052 11101
rect 42024 11092 42030 11095
rect 42150 11092 42156 11144
rect 42208 11092 42214 11144
rect 45005 11135 45063 11141
rect 45005 11132 45017 11135
rect 44744 11104 45017 11132
rect 43156 11067 43214 11073
rect 43156 11033 43168 11067
rect 43202 11064 43214 11067
rect 44174 11064 44180 11076
rect 43202 11036 44180 11064
rect 43202 11033 43214 11036
rect 43156 11027 43214 11033
rect 44174 11024 44180 11036
rect 44232 11024 44238 11076
rect 44744 11008 44772 11104
rect 45005 11101 45017 11104
rect 45051 11101 45063 11135
rect 45005 11095 45063 11101
rect 45272 11135 45330 11141
rect 45272 11101 45284 11135
rect 45318 11132 45330 11135
rect 45554 11132 45560 11144
rect 45318 11104 45560 11132
rect 45318 11101 45330 11104
rect 45272 11095 45330 11101
rect 45554 11092 45560 11104
rect 45612 11092 45618 11144
rect 46753 11135 46811 11141
rect 46753 11101 46765 11135
rect 46799 11132 46811 11135
rect 46934 11132 46940 11144
rect 46799 11104 46940 11132
rect 46799 11101 46811 11104
rect 46753 11095 46811 11101
rect 46934 11092 46940 11104
rect 46992 11092 46998 11144
rect 47486 11092 47492 11144
rect 47544 11092 47550 11144
rect 48792 11064 48820 11172
rect 48958 11160 48964 11172
rect 49016 11160 49022 11212
rect 49050 11160 49056 11212
rect 49108 11160 49114 11212
rect 49344 11209 49372 11240
rect 50172 11209 50200 11296
rect 49329 11203 49387 11209
rect 49329 11169 49341 11203
rect 49375 11169 49387 11203
rect 49329 11163 49387 11169
rect 50157 11203 50215 11209
rect 50157 11169 50169 11203
rect 50203 11169 50215 11203
rect 50157 11163 50215 11169
rect 48866 11092 48872 11144
rect 48924 11132 48930 11144
rect 49973 11135 50031 11141
rect 49973 11132 49985 11135
rect 48924 11104 49985 11132
rect 48924 11092 48930 11104
rect 49973 11101 49985 11104
rect 50019 11101 50031 11135
rect 49973 11095 50031 11101
rect 50424 11135 50482 11141
rect 50424 11101 50436 11135
rect 50470 11132 50482 11135
rect 51276 11132 51304 11308
rect 52546 11296 52552 11308
rect 52604 11296 52610 11348
rect 54389 11339 54447 11345
rect 54389 11305 54401 11339
rect 54435 11336 54447 11339
rect 54478 11336 54484 11348
rect 54435 11308 54484 11336
rect 54435 11305 54447 11308
rect 54389 11299 54447 11305
rect 54478 11296 54484 11308
rect 54536 11296 54542 11348
rect 55950 11336 55956 11348
rect 55232 11308 55956 11336
rect 51537 11271 51595 11277
rect 51537 11237 51549 11271
rect 51583 11268 51595 11271
rect 51583 11240 52408 11268
rect 51583 11237 51595 11240
rect 51537 11231 51595 11237
rect 51350 11160 51356 11212
rect 51408 11200 51414 11212
rect 51629 11203 51687 11209
rect 51629 11200 51641 11203
rect 51408 11172 51641 11200
rect 51408 11160 51414 11172
rect 51629 11169 51641 11172
rect 51675 11169 51687 11203
rect 51629 11163 51687 11169
rect 51813 11203 51871 11209
rect 51813 11169 51825 11203
rect 51859 11200 51871 11203
rect 52178 11200 52184 11212
rect 51859 11172 52184 11200
rect 51859 11169 51871 11172
rect 51813 11163 51871 11169
rect 52178 11160 52184 11172
rect 52236 11160 52242 11212
rect 52270 11160 52276 11212
rect 52328 11160 52334 11212
rect 52380 11200 52408 11240
rect 52546 11200 52552 11212
rect 52380 11172 52552 11200
rect 52546 11160 52552 11172
rect 52604 11160 52610 11212
rect 52822 11160 52828 11212
rect 52880 11160 52886 11212
rect 54941 11203 54999 11209
rect 54941 11200 54953 11203
rect 54220 11172 54953 11200
rect 50470 11104 51304 11132
rect 50470 11101 50482 11104
rect 50424 11095 50482 11101
rect 52638 11092 52644 11144
rect 52696 11141 52702 11144
rect 52696 11135 52724 11141
rect 52712 11101 52724 11135
rect 52696 11095 52724 11101
rect 52696 11092 52702 11095
rect 54018 11092 54024 11144
rect 54076 11132 54082 11144
rect 54220 11141 54248 11172
rect 54941 11169 54953 11172
rect 54987 11169 54999 11203
rect 54941 11163 54999 11169
rect 54205 11135 54263 11141
rect 54205 11132 54217 11135
rect 54076 11104 54217 11132
rect 54076 11092 54082 11104
rect 54205 11101 54217 11104
rect 54251 11101 54263 11135
rect 54205 11095 54263 11101
rect 54757 11135 54815 11141
rect 54757 11101 54769 11135
rect 54803 11132 54815 11135
rect 55232 11132 55260 11308
rect 55950 11296 55956 11308
rect 56008 11296 56014 11348
rect 55309 11271 55367 11277
rect 55309 11237 55321 11271
rect 55355 11268 55367 11271
rect 55355 11240 56180 11268
rect 55355 11237 55367 11240
rect 55309 11231 55367 11237
rect 55490 11160 55496 11212
rect 55548 11160 55554 11212
rect 55858 11160 55864 11212
rect 55916 11160 55922 11212
rect 56152 11209 56180 11240
rect 56870 11228 56876 11280
rect 56928 11228 56934 11280
rect 57256 11240 57468 11268
rect 56137 11203 56195 11209
rect 56137 11169 56149 11203
rect 56183 11169 56195 11203
rect 57256 11200 57284 11240
rect 57440 11209 57468 11240
rect 56137 11163 56195 11169
rect 56244 11172 57284 11200
rect 57425 11203 57483 11209
rect 54803 11104 55260 11132
rect 55508 11132 55536 11160
rect 56244 11132 56272 11172
rect 57425 11169 57437 11203
rect 57471 11200 57483 11203
rect 57885 11203 57943 11209
rect 57885 11200 57897 11203
rect 57471 11172 57897 11200
rect 57471 11169 57483 11172
rect 57425 11163 57483 11169
rect 57885 11169 57897 11172
rect 57931 11169 57943 11203
rect 57885 11163 57943 11169
rect 55508 11104 56272 11132
rect 57241 11135 57299 11141
rect 54803 11101 54815 11104
rect 54757 11095 54815 11101
rect 57241 11101 57253 11135
rect 57287 11132 57299 11135
rect 57514 11132 57520 11144
rect 57287 11104 57520 11132
rect 57287 11101 57299 11104
rect 57241 11095 57299 11101
rect 57514 11092 57520 11104
rect 57572 11092 57578 11144
rect 57606 11092 57612 11144
rect 57664 11092 57670 11144
rect 48961 11067 49019 11073
rect 48792 11036 48912 11064
rect 44082 10996 44088 11008
rect 41156 10968 44088 10996
rect 44082 10956 44088 10968
rect 44140 10956 44146 11008
rect 44726 10956 44732 11008
rect 44784 10956 44790 11008
rect 48884 11005 48912 11036
rect 48961 11033 48973 11067
rect 49007 11064 49019 11067
rect 49694 11064 49700 11076
rect 49007 11036 49700 11064
rect 49007 11033 49019 11036
rect 48961 11027 49019 11033
rect 49694 11024 49700 11036
rect 49752 11024 49758 11076
rect 53469 11067 53527 11073
rect 53469 11033 53481 11067
rect 53515 11064 53527 11067
rect 54662 11064 54668 11076
rect 53515 11036 54668 11064
rect 53515 11033 53527 11036
rect 53469 11027 53527 11033
rect 54662 11024 54668 11036
rect 54720 11024 54726 11076
rect 54849 11067 54907 11073
rect 54849 11033 54861 11067
rect 54895 11064 54907 11067
rect 55677 11067 55735 11073
rect 55677 11064 55689 11067
rect 54895 11036 55689 11064
rect 54895 11033 54907 11036
rect 54849 11027 54907 11033
rect 55677 11033 55689 11036
rect 55723 11064 55735 11067
rect 57333 11067 57391 11073
rect 55723 11036 57008 11064
rect 55723 11033 55735 11036
rect 55677 11027 55735 11033
rect 56980 11008 57008 11036
rect 57333 11033 57345 11067
rect 57379 11064 57391 11067
rect 57624 11064 57652 11092
rect 57379 11036 57652 11064
rect 57379 11033 57391 11036
rect 57333 11027 57391 11033
rect 48869 10999 48927 11005
rect 48869 10965 48881 10999
rect 48915 10965 48927 10999
rect 48869 10959 48927 10965
rect 55766 10956 55772 11008
rect 55824 10956 55830 11008
rect 56778 10956 56784 11008
rect 56836 10956 56842 11008
rect 56962 10956 56968 11008
rect 57020 10956 57026 11008
rect 1104 10906 59040 10928
rect 1104 10854 15394 10906
rect 15446 10854 15458 10906
rect 15510 10854 15522 10906
rect 15574 10854 15586 10906
rect 15638 10854 15650 10906
rect 15702 10854 29838 10906
rect 29890 10854 29902 10906
rect 29954 10854 29966 10906
rect 30018 10854 30030 10906
rect 30082 10854 30094 10906
rect 30146 10854 44282 10906
rect 44334 10854 44346 10906
rect 44398 10854 44410 10906
rect 44462 10854 44474 10906
rect 44526 10854 44538 10906
rect 44590 10854 58726 10906
rect 58778 10854 58790 10906
rect 58842 10854 58854 10906
rect 58906 10854 58918 10906
rect 58970 10854 58982 10906
rect 59034 10854 59040 10906
rect 1104 10832 59040 10854
rect 3142 10752 3148 10804
rect 3200 10752 3206 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3384 10764 3617 10792
rect 3384 10752 3390 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 3605 10755 3663 10761
rect 4522 10752 4528 10804
rect 4580 10752 4586 10804
rect 6822 10752 6828 10804
rect 6880 10792 6886 10804
rect 6917 10795 6975 10801
rect 6917 10792 6929 10795
rect 6880 10764 6929 10792
rect 6880 10752 6886 10764
rect 6917 10761 6929 10764
rect 6963 10792 6975 10795
rect 7190 10792 7196 10804
rect 6963 10764 7196 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 7834 10752 7840 10804
rect 7892 10752 7898 10804
rect 8386 10752 8392 10804
rect 8444 10752 8450 10804
rect 8570 10752 8576 10804
rect 8628 10752 8634 10804
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 11054 10792 11060 10804
rect 9539 10764 11060 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11330 10752 11336 10804
rect 11388 10752 11394 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 11756 10764 11989 10792
rect 11756 10752 11762 10764
rect 11977 10761 11989 10764
rect 12023 10792 12035 10795
rect 12158 10792 12164 10804
rect 12023 10764 12164 10792
rect 12023 10761 12035 10764
rect 11977 10755 12035 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12406 10764 13768 10792
rect 3160 10724 3188 10752
rect 8404 10724 8432 10752
rect 8846 10724 8852 10736
rect 2884 10696 3188 10724
rect 3344 10696 4108 10724
rect 2774 10616 2780 10668
rect 2832 10616 2838 10668
rect 2884 10665 2912 10696
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 3344 10656 3372 10696
rect 3108 10628 3372 10656
rect 3421 10659 3479 10665
rect 3108 10616 3114 10628
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 3602 10656 3608 10668
rect 3467 10628 3608 10656
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 2792 10588 2820 10616
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2792 10560 3157 10588
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10588 3295 10591
rect 3326 10588 3332 10600
rect 3283 10560 3332 10588
rect 3283 10557 3295 10560
rect 3237 10551 3295 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 4080 10464 4108 10696
rect 5184 10696 5856 10724
rect 8404 10696 8852 10724
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10656 4951 10659
rect 4982 10656 4988 10668
rect 4939 10628 4988 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 4448 10520 4476 10619
rect 4724 10588 4752 10619
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5184 10665 5212 10696
rect 5828 10668 5856 10696
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 9950 10724 9956 10736
rect 9600 10696 9956 10724
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5323 10659 5381 10665
rect 5323 10625 5335 10659
rect 5369 10656 5381 10659
rect 5442 10656 5448 10668
rect 5369 10628 5448 10656
rect 5369 10625 5381 10628
rect 5323 10619 5381 10625
rect 5442 10616 5448 10628
rect 5500 10656 5506 10668
rect 5810 10665 5816 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5500 10628 5641 10656
rect 5500 10616 5506 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5783 10659 5816 10665
rect 5783 10625 5795 10659
rect 5868 10656 5874 10668
rect 7285 10659 7343 10665
rect 5868 10628 6592 10656
rect 5783 10619 5816 10625
rect 5810 10616 5816 10619
rect 5868 10616 5874 10628
rect 5997 10591 6055 10597
rect 5997 10588 6009 10591
rect 4724 10560 6009 10588
rect 5997 10557 6009 10560
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 5258 10520 5264 10532
rect 4448 10492 5264 10520
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4801 10455 4859 10461
rect 4801 10452 4813 10455
rect 4120 10424 4813 10452
rect 4120 10412 4126 10424
rect 4801 10421 4813 10424
rect 4847 10421 4859 10455
rect 4801 10415 4859 10421
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 6564 10461 6592 10628
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 7742 10656 7748 10668
rect 7331 10628 7748 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 9398 10616 9404 10668
rect 9456 10616 9462 10668
rect 9600 10597 9628 10696
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 10502 10684 10508 10736
rect 10560 10684 10566 10736
rect 11348 10724 11376 10752
rect 12066 10724 12072 10736
rect 11348 10696 12072 10724
rect 12066 10684 12072 10696
rect 12124 10724 12130 10736
rect 12406 10724 12434 10764
rect 12124 10696 12434 10724
rect 12124 10684 12130 10696
rect 13740 10665 13768 10764
rect 13814 10752 13820 10804
rect 13872 10752 13878 10804
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10792 14243 10795
rect 14826 10792 14832 10804
rect 14231 10764 14832 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15749 10795 15807 10801
rect 15749 10761 15761 10795
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 11931 10628 13001 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 15654 10656 15660 10668
rect 13771 10628 15660 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 12161 10591 12219 10597
rect 10827 10560 11560 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10520 9091 10523
rect 9876 10520 9904 10551
rect 11532 10529 11560 10560
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12207 10560 12296 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12268 10532 12296 10560
rect 12342 10548 12348 10600
rect 12400 10548 12406 10600
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14476 10597 14504 10628
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 13872 10560 14289 10588
rect 13872 10548 13878 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10588 15163 10591
rect 15764 10588 15792 10755
rect 16666 10752 16672 10804
rect 16724 10752 16730 10804
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 18046 10792 18052 10804
rect 17175 10764 18052 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 18046 10752 18052 10764
rect 18104 10752 18110 10804
rect 19705 10795 19763 10801
rect 19705 10761 19717 10795
rect 19751 10792 19763 10795
rect 20346 10792 20352 10804
rect 19751 10764 20352 10792
rect 19751 10761 19763 10764
rect 19705 10755 19763 10761
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 22186 10792 22192 10804
rect 21140 10764 22192 10792
rect 21140 10752 21146 10764
rect 22186 10752 22192 10764
rect 22244 10792 22250 10804
rect 29546 10792 29552 10804
rect 22244 10764 29552 10792
rect 22244 10752 22250 10764
rect 29546 10752 29552 10764
rect 29604 10752 29610 10804
rect 30650 10752 30656 10804
rect 30708 10792 30714 10804
rect 31570 10792 31576 10804
rect 30708 10764 31576 10792
rect 30708 10752 30714 10764
rect 31570 10752 31576 10764
rect 31628 10752 31634 10804
rect 33873 10795 33931 10801
rect 33873 10761 33885 10795
rect 33919 10792 33931 10795
rect 34606 10792 34612 10804
rect 33919 10764 34612 10792
rect 33919 10761 33931 10764
rect 33873 10755 33931 10761
rect 34606 10752 34612 10764
rect 34664 10752 34670 10804
rect 34701 10795 34759 10801
rect 34701 10761 34713 10795
rect 34747 10792 34759 10795
rect 34882 10792 34888 10804
rect 34747 10764 34888 10792
rect 34747 10761 34759 10764
rect 34701 10755 34759 10761
rect 34882 10752 34888 10764
rect 34940 10752 34946 10804
rect 35066 10752 35072 10804
rect 35124 10792 35130 10804
rect 36906 10792 36912 10804
rect 35124 10764 36912 10792
rect 35124 10752 35130 10764
rect 36906 10752 36912 10764
rect 36964 10792 36970 10804
rect 37001 10795 37059 10801
rect 37001 10792 37013 10795
rect 36964 10764 37013 10792
rect 36964 10752 36970 10764
rect 37001 10761 37013 10764
rect 37047 10761 37059 10795
rect 37001 10755 37059 10761
rect 37277 10795 37335 10801
rect 37277 10761 37289 10795
rect 37323 10792 37335 10795
rect 37458 10792 37464 10804
rect 37323 10764 37464 10792
rect 37323 10761 37335 10764
rect 37277 10755 37335 10761
rect 37458 10752 37464 10764
rect 37516 10752 37522 10804
rect 38838 10752 38844 10804
rect 38896 10752 38902 10804
rect 40954 10752 40960 10804
rect 41012 10792 41018 10804
rect 41049 10795 41107 10801
rect 41049 10792 41061 10795
rect 41012 10764 41061 10792
rect 41012 10752 41018 10764
rect 41049 10761 41061 10764
rect 41095 10761 41107 10795
rect 41049 10755 41107 10761
rect 41506 10752 41512 10804
rect 41564 10792 41570 10804
rect 42150 10792 42156 10804
rect 41564 10764 42156 10792
rect 41564 10752 41570 10764
rect 42150 10752 42156 10764
rect 42208 10752 42214 10804
rect 43806 10752 43812 10804
rect 43864 10752 43870 10804
rect 44174 10752 44180 10804
rect 44232 10792 44238 10804
rect 44545 10795 44603 10801
rect 44545 10792 44557 10795
rect 44232 10764 44557 10792
rect 44232 10752 44238 10764
rect 44545 10761 44557 10764
rect 44591 10761 44603 10795
rect 44545 10755 44603 10761
rect 47026 10752 47032 10804
rect 47084 10752 47090 10804
rect 47118 10752 47124 10804
rect 47176 10792 47182 10804
rect 48961 10795 49019 10801
rect 48961 10792 48973 10795
rect 47176 10764 48973 10792
rect 47176 10752 47182 10764
rect 48961 10761 48973 10764
rect 49007 10761 49019 10795
rect 48961 10755 49019 10761
rect 16209 10727 16267 10733
rect 16209 10693 16221 10727
rect 16255 10724 16267 10727
rect 19797 10727 19855 10733
rect 16255 10696 17080 10724
rect 16255 10693 16267 10696
rect 16209 10687 16267 10693
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 16758 10656 16764 10668
rect 16163 10628 16764 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 17052 10665 17080 10696
rect 19797 10693 19809 10727
rect 19843 10724 19855 10727
rect 31478 10724 31484 10736
rect 19843 10696 31484 10724
rect 19843 10693 19855 10696
rect 19797 10687 19855 10693
rect 31478 10684 31484 10696
rect 31536 10724 31542 10736
rect 39025 10727 39083 10733
rect 39025 10724 39037 10727
rect 31536 10696 39037 10724
rect 31536 10684 31542 10696
rect 39025 10693 39037 10696
rect 39071 10693 39083 10727
rect 39025 10687 39083 10693
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17678 10656 17684 10668
rect 17083 10628 17684 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17678 10616 17684 10628
rect 17736 10656 17742 10668
rect 17865 10659 17923 10665
rect 17736 10628 17816 10656
rect 17736 10616 17742 10628
rect 15151 10560 15792 10588
rect 15151 10557 15163 10560
rect 15105 10551 15163 10557
rect 16298 10548 16304 10600
rect 16356 10548 16362 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 16960 10560 17233 10588
rect 9079 10492 9904 10520
rect 11517 10523 11575 10529
rect 9079 10489 9091 10492
rect 9033 10483 9091 10489
rect 11517 10489 11529 10523
rect 11563 10489 11575 10523
rect 11517 10483 11575 10489
rect 12250 10480 12256 10532
rect 12308 10520 12314 10532
rect 13538 10520 13544 10532
rect 12308 10492 13544 10520
rect 12308 10480 12314 10492
rect 13538 10480 13544 10492
rect 13596 10480 13602 10532
rect 16960 10520 16988 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17788 10588 17816 10628
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 18230 10656 18236 10668
rect 17911 10628 18236 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 18782 10616 18788 10668
rect 18840 10616 18846 10668
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10656 22799 10659
rect 23198 10656 23204 10668
rect 22787 10628 23204 10656
rect 22787 10625 22799 10628
rect 22741 10619 22799 10625
rect 23198 10616 23204 10628
rect 23256 10616 23262 10668
rect 23290 10616 23296 10668
rect 23348 10616 23354 10668
rect 23382 10616 23388 10668
rect 23440 10616 23446 10668
rect 23566 10616 23572 10668
rect 23624 10656 23630 10668
rect 24029 10659 24087 10665
rect 24029 10656 24041 10659
rect 23624 10628 24041 10656
rect 23624 10616 23630 10628
rect 24029 10625 24041 10628
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10656 24455 10659
rect 24486 10656 24492 10668
rect 24443 10628 24492 10656
rect 24443 10625 24455 10628
rect 24397 10619 24455 10625
rect 24486 10616 24492 10628
rect 24544 10616 24550 10668
rect 25133 10659 25191 10665
rect 25133 10625 25145 10659
rect 25179 10656 25191 10659
rect 26510 10656 26516 10668
rect 25179 10628 26516 10656
rect 25179 10625 25191 10628
rect 25133 10619 25191 10625
rect 26510 10616 26516 10628
rect 26568 10616 26574 10668
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 27338 10656 27344 10668
rect 27295 10628 27344 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 27338 10616 27344 10628
rect 27396 10616 27402 10668
rect 27516 10659 27574 10665
rect 27516 10625 27528 10659
rect 27562 10656 27574 10659
rect 28350 10656 28356 10668
rect 27562 10628 28356 10656
rect 27562 10625 27574 10628
rect 27516 10619 27574 10625
rect 28350 10616 28356 10628
rect 28408 10616 28414 10668
rect 29086 10616 29092 10668
rect 29144 10616 29150 10668
rect 29181 10659 29239 10665
rect 29181 10625 29193 10659
rect 29227 10656 29239 10659
rect 30193 10659 30251 10665
rect 30193 10656 30205 10659
rect 29227 10628 30205 10656
rect 29227 10625 29239 10628
rect 29181 10619 29239 10625
rect 30193 10625 30205 10628
rect 30239 10625 30251 10659
rect 30193 10619 30251 10625
rect 30282 10616 30288 10668
rect 30340 10616 30346 10668
rect 30834 10616 30840 10668
rect 30892 10656 30898 10668
rect 31021 10659 31079 10665
rect 31021 10656 31033 10659
rect 30892 10628 31033 10656
rect 30892 10616 30898 10628
rect 31021 10625 31033 10628
rect 31067 10625 31079 10659
rect 31021 10619 31079 10625
rect 32760 10659 32818 10665
rect 32760 10625 32772 10659
rect 32806 10656 32818 10659
rect 33594 10656 33600 10668
rect 32806 10628 33600 10656
rect 32806 10625 32818 10628
rect 32760 10619 32818 10625
rect 33594 10616 33600 10628
rect 33652 10616 33658 10668
rect 34609 10659 34667 10665
rect 34609 10625 34621 10659
rect 34655 10656 34667 10659
rect 35250 10656 35256 10668
rect 34655 10628 35256 10656
rect 34655 10625 34667 10628
rect 34609 10619 34667 10625
rect 35250 10616 35256 10628
rect 35308 10616 35314 10668
rect 35888 10659 35946 10665
rect 35888 10625 35900 10659
rect 35934 10656 35946 10659
rect 36630 10656 36636 10668
rect 35934 10628 36636 10656
rect 35934 10625 35946 10628
rect 35888 10619 35946 10625
rect 36630 10616 36636 10628
rect 36688 10616 36694 10668
rect 37642 10616 37648 10668
rect 37700 10616 37706 10668
rect 42429 10659 42487 10665
rect 42429 10625 42441 10659
rect 42475 10656 42487 10659
rect 42518 10656 42524 10668
rect 42475 10628 42524 10656
rect 42475 10625 42487 10628
rect 42429 10619 42487 10625
rect 42518 10616 42524 10628
rect 42576 10616 42582 10668
rect 42696 10659 42754 10665
rect 42696 10625 42708 10659
rect 42742 10656 42754 10659
rect 43622 10656 43628 10668
rect 42742 10628 43628 10656
rect 42742 10625 42754 10628
rect 42696 10619 42754 10625
rect 43622 10616 43628 10628
rect 43680 10616 43686 10668
rect 45088 10659 45146 10665
rect 45088 10625 45100 10659
rect 45134 10656 45146 10659
rect 46658 10656 46664 10668
rect 45134 10628 46664 10656
rect 45134 10625 45146 10628
rect 45088 10619 45146 10625
rect 46658 10616 46664 10628
rect 46716 10616 46722 10668
rect 47848 10659 47906 10665
rect 47848 10625 47860 10659
rect 47894 10656 47906 10659
rect 48866 10656 48872 10668
rect 47894 10628 48872 10656
rect 47894 10625 47906 10628
rect 47848 10619 47906 10625
rect 48866 10616 48872 10628
rect 48924 10616 48930 10668
rect 48976 10656 49004 10755
rect 49694 10752 49700 10804
rect 49752 10752 49758 10804
rect 51258 10752 51264 10804
rect 51316 10752 51322 10804
rect 51721 10795 51779 10801
rect 51721 10761 51733 10795
rect 51767 10792 51779 10795
rect 51994 10792 52000 10804
rect 51767 10764 52000 10792
rect 51767 10761 51779 10764
rect 51721 10755 51779 10761
rect 51994 10752 52000 10764
rect 52052 10752 52058 10804
rect 52270 10752 52276 10804
rect 52328 10792 52334 10804
rect 55214 10792 55220 10804
rect 52328 10764 55220 10792
rect 52328 10752 52334 10764
rect 55214 10752 55220 10764
rect 55272 10752 55278 10804
rect 55677 10795 55735 10801
rect 55677 10761 55689 10795
rect 55723 10792 55735 10795
rect 56686 10792 56692 10804
rect 55723 10764 56692 10792
rect 55723 10761 55735 10764
rect 55677 10755 55735 10761
rect 56686 10752 56692 10764
rect 56744 10752 56750 10804
rect 57698 10752 57704 10804
rect 57756 10752 57762 10804
rect 51276 10724 51304 10752
rect 51350 10724 51356 10736
rect 51276 10696 51356 10724
rect 51350 10684 51356 10696
rect 51408 10724 51414 10736
rect 52086 10724 52092 10736
rect 51408 10696 52092 10724
rect 51408 10684 51414 10696
rect 52086 10684 52092 10696
rect 52144 10684 52150 10736
rect 56778 10724 56784 10736
rect 54312 10696 56364 10724
rect 49053 10659 49111 10665
rect 49053 10656 49065 10659
rect 48976 10628 49065 10656
rect 49053 10625 49065 10628
rect 49099 10625 49111 10659
rect 49053 10619 49111 10625
rect 50516 10659 50574 10665
rect 50516 10625 50528 10659
rect 50562 10656 50574 10659
rect 51258 10656 51264 10668
rect 50562 10628 51264 10656
rect 50562 10625 50574 10628
rect 50516 10619 50574 10625
rect 51258 10616 51264 10628
rect 51316 10616 51322 10668
rect 52181 10659 52239 10665
rect 52181 10625 52193 10659
rect 52227 10656 52239 10659
rect 53377 10659 53435 10665
rect 53377 10656 53389 10659
rect 52227 10628 53389 10656
rect 52227 10625 52239 10628
rect 52181 10619 52239 10625
rect 53377 10625 53389 10628
rect 53423 10625 53435 10659
rect 53377 10619 53435 10625
rect 53834 10616 53840 10668
rect 53892 10656 53898 10668
rect 54312 10665 54340 10696
rect 56336 10665 56364 10696
rect 56428 10696 56784 10724
rect 54297 10659 54355 10665
rect 54297 10656 54309 10659
rect 53892 10628 54309 10656
rect 53892 10616 53898 10628
rect 54297 10625 54309 10628
rect 54343 10625 54355 10659
rect 54297 10619 54355 10625
rect 54564 10659 54622 10665
rect 54564 10625 54576 10659
rect 54610 10656 54622 10659
rect 56321 10659 56379 10665
rect 54610 10628 55720 10656
rect 54610 10625 54622 10628
rect 54564 10619 54622 10625
rect 17954 10588 17960 10600
rect 17788 10560 17960 10588
rect 17221 10551 17279 10557
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18095 10560 18184 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 15028 10492 16988 10520
rect 18156 10520 18184 10560
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 18902 10591 18960 10597
rect 18902 10588 18914 10591
rect 18656 10560 18914 10588
rect 18656 10548 18662 10560
rect 18902 10557 18914 10560
rect 18948 10557 18960 10591
rect 18902 10551 18960 10557
rect 19058 10548 19064 10600
rect 19116 10548 19122 10600
rect 25038 10548 25044 10600
rect 25096 10588 25102 10600
rect 25222 10588 25228 10600
rect 25096 10560 25228 10588
rect 25096 10548 25102 10560
rect 25222 10548 25228 10560
rect 25280 10548 25286 10600
rect 25314 10548 25320 10600
rect 25372 10548 25378 10600
rect 25593 10591 25651 10597
rect 25593 10557 25605 10591
rect 25639 10557 25651 10591
rect 25593 10551 25651 10557
rect 18156 10492 18368 10520
rect 15028 10464 15056 10492
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 5040 10424 5365 10452
rect 5040 10412 5046 10424
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5353 10415 5411 10421
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 8018 10452 8024 10464
rect 6595 10424 8024 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 11330 10412 11336 10464
rect 11388 10412 11394 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14148 10424 14933 10452
rect 14148 10412 14154 10424
rect 14921 10421 14933 10424
rect 14967 10452 14979 10455
rect 15010 10452 15016 10464
rect 14967 10424 15016 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 15657 10455 15715 10461
rect 15657 10421 15669 10455
rect 15703 10452 15715 10455
rect 15838 10452 15844 10464
rect 15703 10424 15844 10452
rect 15703 10421 15715 10424
rect 15657 10415 15715 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 17678 10452 17684 10464
rect 16632 10424 17684 10452
rect 16632 10412 16638 10424
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 18340 10452 18368 10492
rect 18414 10480 18420 10532
rect 18472 10520 18478 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 18472 10492 18521 10520
rect 18472 10480 18478 10492
rect 18509 10489 18521 10492
rect 18555 10489 18567 10523
rect 18509 10483 18567 10489
rect 24765 10523 24823 10529
rect 24765 10489 24777 10523
rect 24811 10520 24823 10523
rect 25608 10520 25636 10551
rect 25682 10548 25688 10600
rect 25740 10588 25746 10600
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 25740 10560 26249 10588
rect 25740 10548 25746 10560
rect 26237 10557 26249 10560
rect 26283 10557 26295 10591
rect 29273 10591 29331 10597
rect 29273 10588 29285 10591
rect 26237 10551 26295 10557
rect 28276 10560 29285 10588
rect 24811 10492 25636 10520
rect 24811 10489 24823 10492
rect 24765 10483 24823 10489
rect 20438 10452 20444 10464
rect 18340 10424 20444 10452
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 26694 10412 26700 10464
rect 26752 10452 26758 10464
rect 26789 10455 26847 10461
rect 26789 10452 26801 10455
rect 26752 10424 26801 10452
rect 26752 10412 26758 10424
rect 26789 10421 26801 10424
rect 26835 10452 26847 10455
rect 28276 10452 28304 10560
rect 29273 10557 29285 10560
rect 29319 10557 29331 10591
rect 29273 10551 29331 10557
rect 29641 10591 29699 10597
rect 29641 10557 29653 10591
rect 29687 10557 29699 10591
rect 29641 10551 29699 10557
rect 28626 10480 28632 10532
rect 28684 10520 28690 10532
rect 29656 10520 29684 10551
rect 29914 10548 29920 10600
rect 29972 10588 29978 10600
rect 30300 10588 30328 10616
rect 29972 10560 30328 10588
rect 32493 10591 32551 10597
rect 29972 10548 29978 10560
rect 32493 10557 32505 10591
rect 32539 10557 32551 10591
rect 35621 10591 35679 10597
rect 35621 10588 35633 10591
rect 32493 10551 32551 10557
rect 35452 10560 35633 10588
rect 30282 10520 30288 10532
rect 28684 10492 29040 10520
rect 29656 10492 30288 10520
rect 28684 10480 28690 10492
rect 26835 10424 28304 10452
rect 26835 10421 26847 10424
rect 26789 10415 26847 10421
rect 28718 10412 28724 10464
rect 28776 10412 28782 10464
rect 29012 10452 29040 10492
rect 30282 10480 30288 10492
rect 30340 10480 30346 10532
rect 32508 10464 32536 10551
rect 35452 10529 35480 10560
rect 35621 10557 35633 10560
rect 35667 10557 35679 10591
rect 35621 10551 35679 10557
rect 37737 10591 37795 10597
rect 37737 10557 37749 10591
rect 37783 10557 37795 10591
rect 37737 10551 37795 10557
rect 37921 10591 37979 10597
rect 37921 10557 37933 10591
rect 37967 10588 37979 10591
rect 37967 10560 38240 10588
rect 37967 10557 37979 10560
rect 37921 10551 37979 10557
rect 35437 10523 35495 10529
rect 35437 10520 35449 10523
rect 33428 10492 35449 10520
rect 30558 10452 30564 10464
rect 29012 10424 30564 10452
rect 30558 10412 30564 10424
rect 30616 10412 30622 10464
rect 32490 10412 32496 10464
rect 32548 10452 32554 10464
rect 33428 10452 33456 10492
rect 34256 10464 34284 10492
rect 35437 10489 35449 10492
rect 35483 10489 35495 10523
rect 35437 10483 35495 10489
rect 32548 10424 33456 10452
rect 32548 10412 32554 10424
rect 34238 10412 34244 10464
rect 34296 10412 34302 10464
rect 34330 10412 34336 10464
rect 34388 10452 34394 10464
rect 35069 10455 35127 10461
rect 35069 10452 35081 10455
rect 34388 10424 35081 10452
rect 34388 10412 34394 10424
rect 35069 10421 35081 10424
rect 35115 10421 35127 10455
rect 35069 10415 35127 10421
rect 36354 10412 36360 10464
rect 36412 10452 36418 10464
rect 37752 10452 37780 10551
rect 38212 10464 38240 10560
rect 43898 10548 43904 10600
rect 43956 10548 43962 10600
rect 44821 10591 44879 10597
rect 44821 10557 44833 10591
rect 44867 10557 44879 10591
rect 46477 10591 46535 10597
rect 46477 10588 46489 10591
rect 44821 10551 44879 10557
rect 46216 10560 46489 10588
rect 42058 10520 42064 10532
rect 40328 10492 42064 10520
rect 40328 10464 40356 10492
rect 42058 10480 42064 10492
rect 42116 10520 42122 10532
rect 42116 10492 42472 10520
rect 42116 10480 42122 10492
rect 36412 10424 37780 10452
rect 36412 10412 36418 10424
rect 38194 10412 38200 10464
rect 38252 10452 38258 10464
rect 38289 10455 38347 10461
rect 38289 10452 38301 10455
rect 38252 10424 38301 10452
rect 38252 10412 38258 10424
rect 38289 10421 38301 10424
rect 38335 10421 38347 10455
rect 38289 10415 38347 10421
rect 40310 10412 40316 10464
rect 40368 10412 40374 10464
rect 42444 10452 42472 10492
rect 42702 10452 42708 10464
rect 42444 10424 42708 10452
rect 42702 10412 42708 10424
rect 42760 10412 42766 10464
rect 44726 10412 44732 10464
rect 44784 10452 44790 10464
rect 44836 10452 44864 10551
rect 46216 10529 46244 10560
rect 46477 10557 46489 10560
rect 46523 10588 46535 10591
rect 47486 10588 47492 10600
rect 46523 10560 47492 10588
rect 46523 10557 46535 10560
rect 46477 10551 46535 10557
rect 47486 10548 47492 10560
rect 47544 10548 47550 10600
rect 47581 10591 47639 10597
rect 47581 10557 47593 10591
rect 47627 10557 47639 10591
rect 47581 10551 47639 10557
rect 50157 10591 50215 10597
rect 50157 10557 50169 10591
rect 50203 10588 50215 10591
rect 50249 10591 50307 10597
rect 50249 10588 50261 10591
rect 50203 10560 50261 10588
rect 50203 10557 50215 10560
rect 50157 10551 50215 10557
rect 50249 10557 50261 10560
rect 50295 10557 50307 10591
rect 50249 10551 50307 10557
rect 46201 10523 46259 10529
rect 46201 10489 46213 10523
rect 46247 10489 46259 10523
rect 46201 10483 46259 10489
rect 47397 10523 47455 10529
rect 47397 10489 47409 10523
rect 47443 10520 47455 10523
rect 47596 10520 47624 10551
rect 47443 10492 47624 10520
rect 47443 10489 47455 10492
rect 47397 10483 47455 10489
rect 47596 10452 47624 10492
rect 50172 10452 50200 10551
rect 52270 10548 52276 10600
rect 52328 10548 52334 10600
rect 52546 10548 52552 10600
rect 52604 10588 52610 10600
rect 52733 10591 52791 10597
rect 52733 10588 52745 10591
rect 52604 10560 52745 10588
rect 52604 10548 52610 10560
rect 52733 10557 52745 10560
rect 52779 10557 52791 10591
rect 55692 10588 55720 10628
rect 56321 10625 56333 10659
rect 56367 10625 56379 10659
rect 56321 10619 56379 10625
rect 56428 10588 56456 10696
rect 56778 10684 56784 10696
rect 56836 10684 56842 10736
rect 56588 10659 56646 10665
rect 56588 10625 56600 10659
rect 56634 10656 56646 10659
rect 58529 10659 58587 10665
rect 58529 10656 58541 10659
rect 56634 10628 58541 10656
rect 56634 10625 56646 10628
rect 56588 10619 56646 10625
rect 58529 10625 58541 10628
rect 58575 10625 58587 10659
rect 58529 10619 58587 10625
rect 55692 10560 56456 10588
rect 52733 10551 52791 10557
rect 57882 10548 57888 10600
rect 57940 10548 57946 10600
rect 51629 10523 51687 10529
rect 51629 10489 51641 10523
rect 51675 10520 51687 10523
rect 52638 10520 52644 10532
rect 51675 10492 52644 10520
rect 51675 10489 51687 10492
rect 51629 10483 51687 10489
rect 52638 10480 52644 10492
rect 52696 10480 52702 10532
rect 44784 10424 50200 10452
rect 44784 10412 44790 10424
rect 55306 10412 55312 10464
rect 55364 10452 55370 10464
rect 55858 10452 55864 10464
rect 55364 10424 55864 10452
rect 55364 10412 55370 10424
rect 55858 10412 55864 10424
rect 55916 10452 55922 10464
rect 55953 10455 56011 10461
rect 55953 10452 55965 10455
rect 55916 10424 55965 10452
rect 55916 10412 55922 10424
rect 55953 10421 55965 10424
rect 55999 10421 56011 10455
rect 55953 10415 56011 10421
rect 1104 10362 58880 10384
rect 1104 10310 8172 10362
rect 8224 10310 8236 10362
rect 8288 10310 8300 10362
rect 8352 10310 8364 10362
rect 8416 10310 8428 10362
rect 8480 10310 22616 10362
rect 22668 10310 22680 10362
rect 22732 10310 22744 10362
rect 22796 10310 22808 10362
rect 22860 10310 22872 10362
rect 22924 10310 37060 10362
rect 37112 10310 37124 10362
rect 37176 10310 37188 10362
rect 37240 10310 37252 10362
rect 37304 10310 37316 10362
rect 37368 10310 51504 10362
rect 51556 10310 51568 10362
rect 51620 10310 51632 10362
rect 51684 10310 51696 10362
rect 51748 10310 51760 10362
rect 51812 10310 58880 10362
rect 1104 10288 58880 10310
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 3418 10248 3424 10260
rect 2823 10220 3424 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4157 10251 4215 10257
rect 4157 10217 4169 10251
rect 4203 10248 4215 10251
rect 4246 10248 4252 10260
rect 4203 10220 4252 10248
rect 4203 10217 4215 10220
rect 4157 10211 4215 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 5810 10248 5816 10260
rect 5767 10220 5816 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10778 10248 10784 10260
rect 10008 10220 10784 10248
rect 10008 10208 10014 10220
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12342 10248 12348 10260
rect 12216 10220 12348 10248
rect 12216 10208 12222 10220
rect 12342 10208 12348 10220
rect 12400 10248 12406 10260
rect 12400 10220 13676 10248
rect 12400 10208 12406 10220
rect 11885 10183 11943 10189
rect 2792 10152 3464 10180
rect 2792 10124 2820 10152
rect 2774 10072 2780 10124
rect 2832 10072 2838 10124
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3326 10112 3332 10124
rect 3007 10084 3332 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3436 10044 3464 10152
rect 11885 10149 11897 10183
rect 11931 10180 11943 10183
rect 12066 10180 12072 10192
rect 11931 10152 12072 10180
rect 11931 10149 11943 10152
rect 11885 10143 11943 10149
rect 12066 10140 12072 10152
rect 12124 10180 12130 10192
rect 12124 10152 12848 10180
rect 12124 10140 12130 10152
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 7484 10084 9597 10112
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3099 10016 3372 10044
rect 3436 10016 3801 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 2823 9948 3096 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3068 9908 3096 9948
rect 3142 9936 3148 9988
rect 3200 9936 3206 9988
rect 3344 9976 3372 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4062 10044 4068 10056
rect 4019 10016 4068 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 3602 9976 3608 9988
rect 3344 9948 3608 9976
rect 3602 9936 3608 9948
rect 3660 9936 3666 9988
rect 3988 9908 4016 10007
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 7282 10044 7288 10056
rect 6595 10016 7288 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7484 10053 7512 10084
rect 9585 10081 9597 10084
rect 9631 10081 9643 10115
rect 9585 10075 9643 10081
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10468 10084 10517 10112
rect 10468 10072 10474 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 12253 10115 12311 10121
rect 10505 10075 10563 10081
rect 11992 10084 12204 10112
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8662 10044 8668 10056
rect 8076 10016 8668 10044
rect 8076 10004 8082 10016
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 8803 10016 9045 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9033 10013 9045 10016
rect 9079 10044 9091 10047
rect 9766 10044 9772 10056
rect 9079 10016 9772 10044
rect 9079 10013 9091 10016
rect 9033 10007 9091 10013
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 6822 9936 6828 9988
rect 6880 9936 6886 9988
rect 10772 9979 10830 9985
rect 10772 9945 10784 9979
rect 10818 9976 10830 9979
rect 11790 9976 11796 9988
rect 10818 9948 11796 9976
rect 10818 9945 10830 9948
rect 10772 9939 10830 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 3068 9880 4016 9908
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10226 9908 10232 9920
rect 9732 9880 10232 9908
rect 9732 9868 9738 9880
rect 10226 9868 10232 9880
rect 10284 9908 10290 9920
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10284 9880 10333 9908
rect 10284 9868 10290 9880
rect 10321 9877 10333 9880
rect 10367 9908 10379 9911
rect 11992 9908 12020 10084
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 12176 10044 12204 10084
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12618 10112 12624 10124
rect 12299 10084 12624 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 12710 10072 12716 10124
rect 12768 10072 12774 10124
rect 12820 10112 12848 10152
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12820 10084 13001 10112
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13127 10115 13185 10121
rect 13127 10081 13139 10115
rect 13173 10112 13185 10115
rect 13648 10112 13676 10220
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 14332 10220 15485 10248
rect 14332 10208 14338 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 17034 10208 17040 10260
rect 17092 10208 17098 10260
rect 17310 10208 17316 10260
rect 17368 10248 17374 10260
rect 18046 10248 18052 10260
rect 17368 10220 18052 10248
rect 17368 10208 17374 10220
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 18506 10248 18512 10260
rect 18288 10220 18512 10248
rect 18288 10208 18294 10220
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 21266 10208 21272 10260
rect 21324 10208 21330 10260
rect 28813 10251 28871 10257
rect 28813 10217 28825 10251
rect 28859 10248 28871 10251
rect 34977 10251 35035 10257
rect 28859 10220 30328 10248
rect 28859 10217 28871 10220
rect 28813 10211 28871 10217
rect 19797 10183 19855 10189
rect 19797 10149 19809 10183
rect 19843 10180 19855 10183
rect 23750 10180 23756 10192
rect 19843 10152 20668 10180
rect 19843 10149 19855 10152
rect 19797 10143 19855 10149
rect 13173 10084 13676 10112
rect 19705 10115 19763 10121
rect 13173 10081 13185 10084
rect 13127 10075 13185 10081
rect 19705 10081 19717 10115
rect 19751 10112 19763 10115
rect 19978 10112 19984 10124
rect 19751 10084 19984 10112
rect 19751 10081 19763 10084
rect 19705 10075 19763 10081
rect 19978 10072 19984 10084
rect 20036 10112 20042 10124
rect 20346 10112 20352 10124
rect 20036 10084 20352 10112
rect 20036 10072 20042 10084
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 20640 10121 20668 10152
rect 20732 10152 23756 10180
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10081 20683 10115
rect 20625 10075 20683 10081
rect 12434 10044 12440 10056
rect 12176 10016 12440 10044
rect 12069 10007 12127 10013
rect 10367 9880 12020 9908
rect 12084 9908 12112 10007
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 14056 10016 14105 10044
rect 14056 10004 14062 10016
rect 14093 10013 14105 10016
rect 14139 10044 14151 10047
rect 15102 10044 15108 10056
rect 14139 10016 15108 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 15102 10004 15108 10016
rect 15160 10044 15166 10056
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 15160 10016 15669 10044
rect 15160 10004 15166 10016
rect 15657 10013 15669 10016
rect 15703 10013 15715 10047
rect 15657 10007 15715 10013
rect 15924 10047 15982 10053
rect 15924 10013 15936 10047
rect 15970 10013 15982 10047
rect 15924 10007 15982 10013
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10044 17187 10047
rect 18785 10047 18843 10053
rect 18785 10044 18797 10047
rect 17175 10016 18797 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 18785 10013 18797 10016
rect 18831 10013 18843 10047
rect 18785 10007 18843 10013
rect 14360 9979 14418 9985
rect 13740 9948 14044 9976
rect 13078 9908 13084 9920
rect 12084 9880 13084 9908
rect 10367 9877 10379 9880
rect 10321 9871 10379 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 13740 9908 13768 9948
rect 13320 9880 13768 9908
rect 13320 9868 13326 9880
rect 13906 9868 13912 9920
rect 13964 9868 13970 9920
rect 14016 9908 14044 9948
rect 14360 9945 14372 9979
rect 14406 9976 14418 9979
rect 15194 9976 15200 9988
rect 14406 9948 15200 9976
rect 14406 9945 14418 9948
rect 14360 9939 14418 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 14826 9908 14832 9920
rect 14016 9880 14832 9908
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15672 9908 15700 10007
rect 15838 9936 15844 9988
rect 15896 9976 15902 9988
rect 15948 9976 15976 10007
rect 15896 9948 15976 9976
rect 15896 9936 15902 9948
rect 17144 9908 17172 10007
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 20732 10044 20760 10152
rect 23750 10140 23756 10152
rect 23808 10140 23814 10192
rect 30006 10140 30012 10192
rect 30064 10180 30070 10192
rect 30193 10183 30251 10189
rect 30193 10180 30205 10183
rect 30064 10152 30205 10180
rect 30064 10140 30070 10152
rect 30193 10149 30205 10152
rect 30239 10149 30251 10183
rect 30193 10143 30251 10149
rect 30300 10124 30328 10220
rect 34977 10217 34989 10251
rect 35023 10248 35035 10251
rect 35894 10248 35900 10260
rect 35023 10220 35900 10248
rect 35023 10217 35035 10220
rect 34977 10211 35035 10217
rect 35894 10208 35900 10220
rect 35952 10208 35958 10260
rect 36262 10208 36268 10260
rect 36320 10248 36326 10260
rect 37277 10251 37335 10257
rect 37277 10248 37289 10251
rect 36320 10220 37289 10248
rect 36320 10208 36326 10220
rect 37277 10217 37289 10220
rect 37323 10217 37335 10251
rect 37277 10211 37335 10217
rect 30282 10072 30288 10124
rect 30340 10112 30346 10124
rect 30469 10115 30527 10121
rect 30469 10112 30481 10115
rect 30340 10084 30481 10112
rect 30340 10072 30346 10084
rect 30469 10081 30481 10084
rect 30515 10081 30527 10115
rect 30469 10075 30527 10081
rect 30558 10072 30564 10124
rect 30616 10121 30622 10124
rect 30616 10115 30644 10121
rect 30632 10081 30644 10115
rect 30616 10075 30644 10081
rect 30616 10072 30622 10075
rect 30742 10072 30748 10124
rect 30800 10112 30806 10124
rect 30800 10084 31524 10112
rect 30800 10072 30806 10084
rect 19024 10016 20760 10044
rect 19024 10004 19030 10016
rect 21542 10004 21548 10056
rect 21600 10004 21606 10056
rect 27433 10047 27491 10053
rect 27433 10044 27445 10047
rect 27356 10016 27445 10044
rect 17396 9979 17454 9985
rect 17396 9945 17408 9979
rect 17442 9976 17454 9979
rect 18230 9976 18236 9988
rect 17442 9948 18236 9976
rect 17442 9945 17454 9948
rect 17396 9939 17454 9945
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 20257 9979 20315 9985
rect 20257 9976 20269 9979
rect 18340 9948 20269 9976
rect 17586 9908 17592 9920
rect 15672 9880 17592 9908
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18340 9908 18368 9948
rect 20257 9945 20269 9948
rect 20303 9945 20315 9979
rect 20257 9939 20315 9945
rect 20346 9936 20352 9988
rect 20404 9976 20410 9988
rect 24581 9979 24639 9985
rect 24581 9976 24593 9979
rect 20404 9948 24593 9976
rect 20404 9936 20410 9948
rect 24581 9945 24593 9948
rect 24627 9976 24639 9979
rect 25314 9976 25320 9988
rect 24627 9948 25320 9976
rect 24627 9945 24639 9948
rect 24581 9939 24639 9945
rect 25314 9936 25320 9948
rect 25372 9976 25378 9988
rect 26418 9976 26424 9988
rect 25372 9948 26424 9976
rect 25372 9936 25378 9948
rect 26418 9936 26424 9948
rect 26476 9936 26482 9988
rect 27356 9920 27384 10016
rect 27433 10013 27445 10016
rect 27479 10013 27491 10047
rect 27433 10007 27491 10013
rect 27700 10047 27758 10053
rect 27700 10013 27712 10047
rect 27746 10044 27758 10047
rect 28902 10044 28908 10056
rect 27746 10016 28908 10044
rect 27746 10013 27758 10016
rect 27700 10007 27758 10013
rect 28902 10004 28908 10016
rect 28960 10004 28966 10056
rect 29546 10004 29552 10056
rect 29604 10004 29610 10056
rect 29730 10004 29736 10056
rect 29788 10004 29794 10056
rect 31496 10044 31524 10084
rect 31570 10072 31576 10124
rect 31628 10112 31634 10124
rect 32033 10115 32091 10121
rect 32033 10112 32045 10115
rect 31628 10084 32045 10112
rect 31628 10072 31634 10084
rect 32033 10081 32045 10084
rect 32079 10081 32091 10115
rect 37292 10112 37320 10211
rect 37642 10208 37648 10260
rect 37700 10248 37706 10260
rect 38013 10251 38071 10257
rect 38013 10248 38025 10251
rect 37700 10220 38025 10248
rect 37700 10208 37706 10220
rect 38013 10217 38025 10220
rect 38059 10217 38071 10251
rect 38013 10211 38071 10217
rect 40494 10208 40500 10260
rect 40552 10208 40558 10260
rect 41049 10251 41107 10257
rect 41049 10217 41061 10251
rect 41095 10248 41107 10251
rect 41138 10248 41144 10260
rect 41095 10220 41144 10248
rect 41095 10217 41107 10220
rect 41049 10211 41107 10217
rect 41138 10208 41144 10220
rect 41196 10248 41202 10260
rect 41782 10248 41788 10260
rect 41196 10220 41788 10248
rect 41196 10208 41202 10220
rect 41782 10208 41788 10220
rect 41840 10248 41846 10260
rect 42245 10251 42303 10257
rect 41840 10220 42196 10248
rect 41840 10208 41846 10220
rect 39669 10183 39727 10189
rect 39669 10149 39681 10183
rect 39715 10180 39727 10183
rect 39715 10152 39988 10180
rect 39715 10149 39727 10152
rect 39669 10143 39727 10149
rect 37369 10115 37427 10121
rect 37369 10112 37381 10115
rect 37292 10084 37381 10112
rect 32033 10075 32091 10081
rect 37369 10081 37381 10084
rect 37415 10081 37427 10115
rect 37369 10075 37427 10081
rect 38286 10072 38292 10124
rect 38344 10072 38350 10124
rect 39960 10121 39988 10152
rect 39945 10115 40003 10121
rect 39945 10081 39957 10115
rect 39991 10112 40003 10115
rect 41966 10112 41972 10124
rect 39991 10084 41972 10112
rect 39991 10081 40003 10084
rect 39945 10075 40003 10081
rect 41966 10072 41972 10084
rect 42024 10072 42030 10124
rect 42168 10121 42196 10220
rect 42245 10217 42257 10251
rect 42291 10248 42303 10251
rect 43898 10248 43904 10260
rect 42291 10220 43904 10248
rect 42291 10217 42303 10220
rect 42245 10211 42303 10217
rect 43898 10208 43904 10220
rect 43956 10208 43962 10260
rect 44085 10251 44143 10257
rect 44085 10217 44097 10251
rect 44131 10248 44143 10251
rect 44726 10248 44732 10260
rect 44131 10220 44732 10248
rect 44131 10217 44143 10220
rect 44085 10211 44143 10217
rect 42518 10140 42524 10192
rect 42576 10180 42582 10192
rect 44100 10180 44128 10211
rect 44726 10208 44732 10220
rect 44784 10208 44790 10260
rect 45830 10208 45836 10260
rect 45888 10248 45894 10260
rect 46477 10251 46535 10257
rect 46477 10248 46489 10251
rect 45888 10220 46489 10248
rect 45888 10208 45894 10220
rect 46477 10217 46489 10220
rect 46523 10248 46535 10251
rect 47210 10248 47216 10260
rect 46523 10220 47216 10248
rect 46523 10217 46535 10220
rect 46477 10211 46535 10217
rect 47210 10208 47216 10220
rect 47268 10208 47274 10260
rect 49510 10208 49516 10260
rect 49568 10208 49574 10260
rect 53926 10248 53932 10260
rect 51552 10220 53932 10248
rect 42576 10152 44128 10180
rect 42576 10140 42582 10152
rect 50890 10140 50896 10192
rect 50948 10180 50954 10192
rect 51552 10180 51580 10220
rect 53926 10208 53932 10220
rect 53984 10208 53990 10260
rect 55766 10208 55772 10260
rect 55824 10248 55830 10260
rect 56413 10251 56471 10257
rect 56413 10248 56425 10251
rect 55824 10220 56425 10248
rect 55824 10208 55830 10220
rect 56413 10217 56425 10220
rect 56459 10217 56471 10251
rect 56413 10211 56471 10217
rect 56873 10251 56931 10257
rect 56873 10217 56885 10251
rect 56919 10248 56931 10251
rect 57882 10248 57888 10260
rect 56919 10220 57888 10248
rect 56919 10217 56931 10220
rect 56873 10211 56931 10217
rect 57882 10208 57888 10220
rect 57940 10208 57946 10260
rect 50948 10152 51580 10180
rect 50948 10140 50954 10152
rect 42153 10115 42211 10121
rect 42153 10081 42165 10115
rect 42199 10112 42211 10115
rect 42797 10115 42855 10121
rect 42797 10112 42809 10115
rect 42199 10084 42809 10112
rect 42199 10081 42211 10084
rect 42153 10075 42211 10081
rect 42797 10081 42809 10084
rect 42843 10081 42855 10115
rect 42797 10075 42855 10081
rect 43165 10115 43223 10121
rect 43165 10081 43177 10115
rect 43211 10112 43223 10115
rect 44082 10112 44088 10124
rect 43211 10084 44088 10112
rect 43211 10081 43223 10084
rect 43165 10075 43223 10081
rect 44082 10072 44088 10084
rect 44140 10072 44146 10124
rect 51350 10072 51356 10124
rect 51408 10112 51414 10124
rect 51552 10121 51580 10152
rect 51445 10115 51503 10121
rect 51445 10112 51457 10115
rect 51408 10084 51457 10112
rect 51408 10072 51414 10084
rect 51445 10081 51457 10084
rect 51491 10081 51503 10115
rect 51445 10075 51503 10081
rect 51537 10115 51595 10121
rect 51537 10081 51549 10115
rect 51583 10081 51595 10115
rect 51537 10075 51595 10081
rect 51905 10115 51963 10121
rect 51905 10081 51917 10115
rect 51951 10112 51963 10115
rect 52638 10112 52644 10124
rect 51951 10084 52644 10112
rect 51951 10081 51963 10084
rect 51905 10075 51963 10081
rect 52638 10072 52644 10084
rect 52696 10072 52702 10124
rect 55861 10115 55919 10121
rect 55861 10081 55873 10115
rect 55907 10112 55919 10115
rect 56686 10112 56692 10124
rect 55907 10084 56692 10112
rect 55907 10081 55919 10084
rect 55861 10075 55919 10081
rect 56686 10072 56692 10084
rect 56744 10072 56750 10124
rect 57425 10115 57483 10121
rect 57425 10112 57437 10115
rect 56888 10084 57437 10112
rect 31754 10044 31760 10056
rect 31496 10016 31760 10044
rect 31754 10004 31760 10016
rect 31812 10004 31818 10056
rect 32674 10004 32680 10056
rect 32732 10004 32738 10056
rect 33413 10047 33471 10053
rect 33413 10013 33425 10047
rect 33459 10044 33471 10047
rect 33502 10044 33508 10056
rect 33459 10016 33508 10044
rect 33459 10013 33471 10016
rect 33413 10007 33471 10013
rect 33502 10004 33508 10016
rect 33560 10004 33566 10056
rect 35897 10047 35955 10053
rect 35897 10044 35909 10047
rect 35544 10016 35909 10044
rect 31389 9979 31447 9985
rect 31389 9945 31401 9979
rect 31435 9976 31447 9979
rect 31941 9979 31999 9985
rect 31941 9976 31953 9979
rect 31435 9948 31953 9976
rect 31435 9945 31447 9948
rect 31389 9939 31447 9945
rect 31941 9945 31953 9948
rect 31987 9945 31999 9979
rect 31941 9939 31999 9945
rect 35544 9920 35572 10016
rect 35897 10013 35909 10016
rect 35943 10013 35955 10047
rect 35897 10007 35955 10013
rect 38102 10004 38108 10056
rect 38160 10004 38166 10056
rect 38556 10047 38614 10053
rect 38556 10013 38568 10047
rect 38602 10044 38614 10047
rect 39114 10044 39120 10056
rect 38602 10016 39120 10044
rect 38602 10013 38614 10016
rect 38556 10007 38614 10013
rect 39114 10004 39120 10016
rect 39172 10004 39178 10056
rect 49421 10047 49479 10053
rect 49421 10013 49433 10047
rect 49467 10044 49479 10047
rect 49467 10016 52684 10044
rect 49467 10013 49479 10016
rect 49421 10007 49479 10013
rect 36164 9979 36222 9985
rect 36164 9945 36176 9979
rect 36210 9976 36222 9979
rect 38120 9976 38148 10004
rect 36210 9948 38148 9976
rect 42613 9979 42671 9985
rect 36210 9945 36222 9948
rect 36164 9939 36222 9945
rect 42613 9945 42625 9979
rect 42659 9976 42671 9979
rect 43717 9979 43775 9985
rect 43717 9976 43729 9979
rect 42659 9948 43729 9976
rect 42659 9945 42671 9948
rect 42613 9939 42671 9945
rect 43717 9945 43729 9948
rect 43763 9945 43775 9979
rect 43717 9939 43775 9945
rect 51353 9979 51411 9985
rect 51353 9945 51365 9979
rect 51399 9976 51411 9979
rect 52457 9979 52515 9985
rect 52457 9976 52469 9979
rect 51399 9948 52469 9976
rect 51399 9945 51411 9948
rect 51353 9939 51411 9945
rect 52457 9945 52469 9948
rect 52503 9945 52515 9979
rect 52457 9939 52515 9945
rect 52656 9920 52684 10016
rect 53558 10004 53564 10056
rect 53616 10044 53622 10056
rect 56888 10044 56916 10084
rect 57425 10081 57437 10084
rect 57471 10081 57483 10115
rect 57425 10075 57483 10081
rect 57698 10072 57704 10124
rect 57756 10072 57762 10124
rect 53616 10016 56916 10044
rect 53616 10004 53622 10016
rect 56888 9920 56916 10016
rect 57241 9979 57299 9985
rect 57241 9945 57253 9979
rect 57287 9976 57299 9979
rect 58345 9979 58403 9985
rect 58345 9976 58357 9979
rect 57287 9948 58357 9976
rect 57287 9945 57299 9948
rect 57241 9939 57299 9945
rect 58345 9945 58357 9948
rect 58391 9945 58403 9979
rect 58345 9939 58403 9945
rect 18104 9880 18368 9908
rect 18104 9868 18110 9880
rect 20162 9868 20168 9920
rect 20220 9868 20226 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22189 9911 22247 9917
rect 22189 9908 22201 9911
rect 22152 9880 22201 9908
rect 22152 9868 22158 9880
rect 22189 9877 22201 9880
rect 22235 9877 22247 9911
rect 22189 9871 22247 9877
rect 23109 9911 23167 9917
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23750 9908 23756 9920
rect 23155 9880 23756 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23750 9868 23756 9880
rect 23808 9908 23814 9920
rect 26326 9908 26332 9920
rect 23808 9880 26332 9908
rect 23808 9868 23814 9880
rect 26326 9868 26332 9880
rect 26384 9868 26390 9920
rect 27338 9868 27344 9920
rect 27396 9868 27402 9920
rect 29270 9868 29276 9920
rect 29328 9908 29334 9920
rect 29365 9911 29423 9917
rect 29365 9908 29377 9911
rect 29328 9880 29377 9908
rect 29328 9868 29334 9880
rect 29365 9877 29377 9880
rect 29411 9908 29423 9911
rect 30282 9908 30288 9920
rect 29411 9880 30288 9908
rect 29411 9877 29423 9880
rect 29365 9871 29423 9877
rect 30282 9868 30288 9880
rect 30340 9868 30346 9920
rect 31018 9868 31024 9920
rect 31076 9908 31082 9920
rect 31481 9911 31539 9917
rect 31481 9908 31493 9911
rect 31076 9880 31493 9908
rect 31076 9868 31082 9880
rect 31481 9877 31493 9880
rect 31527 9877 31539 9911
rect 31481 9871 31539 9877
rect 31662 9868 31668 9920
rect 31720 9908 31726 9920
rect 31849 9911 31907 9917
rect 31849 9908 31861 9911
rect 31720 9880 31861 9908
rect 31720 9868 31726 9880
rect 31849 9877 31861 9880
rect 31895 9877 31907 9911
rect 31849 9871 31907 9877
rect 33226 9868 33232 9920
rect 33284 9868 33290 9920
rect 33962 9868 33968 9920
rect 34020 9868 34026 9920
rect 34425 9911 34483 9917
rect 34425 9877 34437 9911
rect 34471 9908 34483 9911
rect 34974 9908 34980 9920
rect 34471 9880 34980 9908
rect 34471 9877 34483 9880
rect 34425 9871 34483 9877
rect 34974 9868 34980 9880
rect 35032 9868 35038 9920
rect 35526 9868 35532 9920
rect 35584 9868 35590 9920
rect 37458 9868 37464 9920
rect 37516 9908 37522 9920
rect 38194 9908 38200 9920
rect 37516 9880 38200 9908
rect 37516 9868 37522 9880
rect 38194 9868 38200 9880
rect 38252 9868 38258 9920
rect 41506 9868 41512 9920
rect 41564 9908 41570 9920
rect 41874 9908 41880 9920
rect 41564 9880 41880 9908
rect 41564 9868 41570 9880
rect 41874 9868 41880 9880
rect 41932 9908 41938 9920
rect 42705 9911 42763 9917
rect 42705 9908 42717 9911
rect 41932 9880 42717 9908
rect 41932 9868 41938 9880
rect 42705 9877 42717 9880
rect 42751 9877 42763 9911
rect 42705 9871 42763 9877
rect 48409 9911 48467 9917
rect 48409 9877 48421 9911
rect 48455 9908 48467 9911
rect 48866 9908 48872 9920
rect 48455 9880 48872 9908
rect 48455 9877 48467 9880
rect 48409 9871 48467 9877
rect 48866 9868 48872 9880
rect 48924 9908 48930 9920
rect 49050 9908 49056 9920
rect 48924 9880 49056 9908
rect 48924 9868 48930 9880
rect 49050 9868 49056 9880
rect 49108 9868 49114 9920
rect 50890 9868 50896 9920
rect 50948 9868 50954 9920
rect 50982 9868 50988 9920
rect 51040 9868 51046 9920
rect 52638 9868 52644 9920
rect 52696 9868 52702 9920
rect 56781 9911 56839 9917
rect 56781 9877 56793 9911
rect 56827 9908 56839 9911
rect 56870 9908 56876 9920
rect 56827 9880 56876 9908
rect 56827 9877 56839 9880
rect 56781 9871 56839 9877
rect 56870 9868 56876 9880
rect 56928 9868 56934 9920
rect 56962 9868 56968 9920
rect 57020 9908 57026 9920
rect 57333 9911 57391 9917
rect 57333 9908 57345 9911
rect 57020 9880 57345 9908
rect 57020 9868 57026 9880
rect 57333 9877 57345 9880
rect 57379 9908 57391 9911
rect 57698 9908 57704 9920
rect 57379 9880 57704 9908
rect 57379 9877 57391 9880
rect 57333 9871 57391 9877
rect 57698 9868 57704 9880
rect 57756 9868 57762 9920
rect 1104 9818 59040 9840
rect 1104 9766 15394 9818
rect 15446 9766 15458 9818
rect 15510 9766 15522 9818
rect 15574 9766 15586 9818
rect 15638 9766 15650 9818
rect 15702 9766 29838 9818
rect 29890 9766 29902 9818
rect 29954 9766 29966 9818
rect 30018 9766 30030 9818
rect 30082 9766 30094 9818
rect 30146 9766 44282 9818
rect 44334 9766 44346 9818
rect 44398 9766 44410 9818
rect 44462 9766 44474 9818
rect 44526 9766 44538 9818
rect 44590 9766 58726 9818
rect 58778 9766 58790 9818
rect 58842 9766 58854 9818
rect 58906 9766 58918 9818
rect 58970 9766 58982 9818
rect 59034 9766 59040 9818
rect 1104 9744 59040 9766
rect 3142 9664 3148 9716
rect 3200 9664 3206 9716
rect 3326 9664 3332 9716
rect 3384 9664 3390 9716
rect 7653 9707 7711 9713
rect 7653 9673 7665 9707
rect 7699 9704 7711 9707
rect 8018 9704 8024 9716
rect 7699 9676 8024 9704
rect 7699 9673 7711 9676
rect 7653 9667 7711 9673
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10468 9676 12434 9704
rect 10468 9664 10474 9676
rect 3160 9636 3188 9664
rect 6181 9639 6239 9645
rect 6181 9636 6193 9639
rect 3160 9608 6193 9636
rect 6181 9605 6193 9608
rect 6227 9636 6239 9639
rect 6270 9636 6276 9648
rect 6227 9608 6276 9636
rect 6227 9605 6239 9608
rect 6181 9599 6239 9605
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 6380 9608 7788 9636
rect 6380 9580 6408 9608
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3053 9571 3111 9577
rect 3053 9568 3065 9571
rect 2976 9540 3065 9568
rect 2774 9460 2780 9512
rect 2832 9460 2838 9512
rect 2792 9432 2820 9460
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 2792 9404 2881 9432
rect 2869 9401 2881 9404
rect 2915 9401 2927 9435
rect 2869 9395 2927 9401
rect 2976 9376 3004 9540
rect 3053 9537 3065 9540
rect 3099 9537 3111 9571
rect 3053 9531 3111 9537
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 3191 9540 3249 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3237 9537 3249 9540
rect 3283 9568 3295 9571
rect 5905 9571 5963 9577
rect 3283 9540 3648 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3620 9376 3648 9540
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6362 9568 6368 9580
rect 5951 9540 6368 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 6503 9540 6868 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 6472 9500 6500 9531
rect 5859 9472 6500 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 5994 9392 6000 9444
rect 6052 9392 6058 9444
rect 6730 9432 6736 9444
rect 6564 9404 6736 9432
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 3789 9367 3847 9373
rect 3789 9333 3801 9367
rect 3835 9364 3847 9367
rect 4706 9364 4712 9376
rect 3835 9336 4712 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9364 6147 9367
rect 6564 9364 6592 9404
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6135 9336 6592 9364
rect 6840 9364 6868 9540
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7466 9528 7472 9580
rect 7524 9528 7530 9580
rect 7760 9577 7788 9608
rect 9766 9596 9772 9648
rect 9824 9596 9830 9648
rect 10220 9639 10278 9645
rect 10220 9605 10232 9639
rect 10266 9636 10278 9639
rect 11330 9636 11336 9648
rect 10266 9608 11336 9636
rect 10266 9605 10278 9608
rect 10220 9599 10278 9605
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 12406 9636 12434 9676
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13817 9707 13875 9713
rect 13817 9704 13829 9707
rect 13136 9676 13829 9704
rect 13136 9664 13142 9676
rect 13817 9673 13829 9676
rect 13863 9673 13875 9707
rect 13817 9667 13875 9673
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 14277 9707 14335 9713
rect 14277 9704 14289 9707
rect 13964 9676 14289 9704
rect 13964 9664 13970 9676
rect 14277 9673 14289 9676
rect 14323 9673 14335 9707
rect 14277 9667 14335 9673
rect 17586 9664 17592 9716
rect 17644 9704 17650 9716
rect 17681 9707 17739 9713
rect 17681 9704 17693 9707
rect 17644 9676 17693 9704
rect 17644 9664 17650 9676
rect 17681 9673 17693 9676
rect 17727 9673 17739 9707
rect 17681 9667 17739 9673
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20441 9707 20499 9713
rect 20441 9704 20453 9707
rect 20220 9676 20453 9704
rect 20220 9664 20226 9676
rect 20441 9673 20453 9676
rect 20487 9673 20499 9707
rect 20441 9667 20499 9673
rect 28261 9707 28319 9713
rect 28261 9673 28273 9707
rect 28307 9704 28319 9707
rect 29086 9704 29092 9716
rect 28307 9676 29092 9704
rect 28307 9673 28319 9676
rect 28261 9667 28319 9673
rect 29086 9664 29092 9676
rect 29144 9664 29150 9716
rect 29546 9664 29552 9716
rect 29604 9704 29610 9716
rect 30009 9707 30067 9713
rect 30009 9704 30021 9707
rect 29604 9676 30021 9704
rect 29604 9664 29610 9676
rect 30009 9673 30021 9676
rect 30055 9673 30067 9707
rect 30009 9667 30067 9673
rect 30098 9664 30104 9716
rect 30156 9704 30162 9716
rect 31478 9704 31484 9716
rect 30156 9676 31484 9704
rect 30156 9664 30162 9676
rect 31478 9664 31484 9676
rect 31536 9664 31542 9716
rect 32401 9707 32459 9713
rect 32401 9673 32413 9707
rect 32447 9704 32459 9707
rect 32490 9704 32496 9716
rect 32447 9676 32496 9704
rect 32447 9673 32459 9676
rect 32401 9667 32459 9673
rect 32490 9664 32496 9676
rect 32548 9664 32554 9716
rect 32674 9664 32680 9716
rect 32732 9664 32738 9716
rect 33962 9664 33968 9716
rect 34020 9664 34026 9716
rect 40494 9664 40500 9716
rect 40552 9704 40558 9716
rect 40954 9704 40960 9716
rect 40552 9676 40960 9704
rect 40552 9664 40558 9676
rect 40954 9664 40960 9676
rect 41012 9704 41018 9716
rect 41012 9676 44128 9704
rect 41012 9664 41018 9676
rect 13998 9636 14004 9648
rect 12406 9608 14004 9636
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 7745 9531 7803 9537
rect 8128 9540 9965 9568
rect 6914 9460 6920 9512
rect 6972 9460 6978 9512
rect 7208 9500 7236 9528
rect 8018 9500 8024 9512
rect 7208 9472 8024 9500
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8128 9509 8156 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 11885 9574 11943 9577
rect 11808 9571 11943 9574
rect 11808 9568 11897 9571
rect 11756 9546 11897 9568
rect 11756 9540 11836 9546
rect 11756 9528 11762 9540
rect 11885 9537 11897 9546
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12452 9577 12480 9608
rect 13998 9596 14004 9608
rect 14056 9636 14062 9648
rect 14921 9639 14979 9645
rect 14921 9636 14933 9639
rect 14056 9608 14933 9636
rect 14056 9596 14062 9608
rect 14921 9605 14933 9608
rect 14967 9636 14979 9639
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 14967 9608 15945 9636
rect 14967 9605 14979 9608
rect 14921 9599 14979 9605
rect 15933 9605 15945 9608
rect 15979 9605 15991 9639
rect 15933 9599 15991 9605
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 27062 9636 27068 9648
rect 16080 9608 27068 9636
rect 16080 9596 16086 9608
rect 27062 9596 27068 9608
rect 27120 9596 27126 9648
rect 27338 9596 27344 9648
rect 27396 9636 27402 9648
rect 33045 9639 33103 9645
rect 27396 9608 30144 9636
rect 27396 9596 27402 9608
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12704 9571 12762 9577
rect 12704 9537 12716 9571
rect 12750 9568 12762 9571
rect 13722 9568 13728 9580
rect 12750 9540 13728 9568
rect 12750 9537 12762 9540
rect 12704 9531 12762 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14642 9568 14648 9580
rect 14415 9540 14648 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9568 15531 9571
rect 15746 9568 15752 9580
rect 15519 9540 15752 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 16816 9540 17325 9568
rect 16816 9528 16822 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 18104 9540 18153 9568
rect 18104 9528 18110 9540
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18141 9531 18199 9537
rect 18233 9571 18291 9577
rect 18233 9537 18245 9571
rect 18279 9568 18291 9571
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 18279 9540 19257 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20438 9568 20444 9580
rect 19935 9540 20444 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 21266 9568 21272 9580
rect 20772 9540 21272 9568
rect 20772 9528 20778 9540
rect 21266 9528 21272 9540
rect 21324 9568 21330 9580
rect 21324 9540 24900 9568
rect 21324 9528 21330 9540
rect 24872 9512 24900 9540
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 26510 9568 26516 9580
rect 25832 9540 26516 9568
rect 25832 9528 25838 9540
rect 26510 9528 26516 9540
rect 26568 9528 26574 9580
rect 26694 9528 26700 9580
rect 26752 9568 26758 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 26752 9540 27445 9568
rect 26752 9528 26758 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 27617 9571 27675 9577
rect 27617 9537 27629 9571
rect 27663 9568 27675 9571
rect 27706 9568 27712 9580
rect 27663 9540 27712 9568
rect 27663 9537 27675 9540
rect 27617 9531 27675 9537
rect 27706 9528 27712 9540
rect 27764 9528 27770 9580
rect 28644 9577 28672 9608
rect 28169 9571 28227 9577
rect 28169 9537 28181 9571
rect 28215 9568 28227 9571
rect 28629 9571 28687 9577
rect 28215 9540 28580 9568
rect 28215 9537 28227 9540
rect 28169 9531 28227 9537
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9469 8171 9503
rect 8113 9463 8171 9469
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8435 9472 9076 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 6932 9432 6960 9460
rect 8128 9432 8156 9463
rect 6932 9404 8156 9432
rect 7190 9364 7196 9376
rect 6840 9336 7196 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7469 9367 7527 9373
rect 7469 9333 7481 9367
rect 7515 9364 7527 9367
rect 9048 9364 9076 9472
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 11480 9472 12081 9500
rect 11480 9460 11486 9472
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 15657 9503 15715 9509
rect 14608 9472 14688 9500
rect 14608 9460 14614 9472
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 12158 9432 12164 9444
rect 11379 9404 12164 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 14660 9432 14688 9472
rect 15657 9469 15669 9503
rect 15703 9500 15715 9503
rect 15930 9500 15936 9512
rect 15703 9472 15936 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9500 16727 9503
rect 17034 9500 17040 9512
rect 16715 9472 17040 9500
rect 16715 9469 16727 9472
rect 16669 9463 16727 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 17920 9472 18337 9500
rect 17920 9460 17926 9472
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 18506 9460 18512 9512
rect 18564 9500 18570 9512
rect 18601 9503 18659 9509
rect 18601 9500 18613 9503
rect 18564 9472 18613 9500
rect 18564 9460 18570 9472
rect 18601 9469 18613 9472
rect 18647 9469 18659 9503
rect 20530 9500 20536 9512
rect 18601 9463 18659 9469
rect 19306 9472 20536 9500
rect 19306 9432 19334 9472
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 20622 9460 20628 9512
rect 20680 9460 20686 9512
rect 21821 9503 21879 9509
rect 21821 9469 21833 9503
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 14660 9404 19334 9432
rect 20070 9392 20076 9444
rect 20128 9432 20134 9444
rect 21836 9432 21864 9463
rect 24210 9460 24216 9512
rect 24268 9460 24274 9512
rect 24854 9460 24860 9512
rect 24912 9500 24918 9512
rect 25498 9500 25504 9512
rect 24912 9472 25504 9500
rect 24912 9460 24918 9472
rect 25498 9460 25504 9472
rect 25556 9500 25562 9512
rect 26142 9500 26148 9512
rect 25556 9472 26148 9500
rect 25556 9460 25562 9472
rect 26142 9460 26148 9472
rect 26200 9460 26206 9512
rect 26234 9460 26240 9512
rect 26292 9460 26298 9512
rect 26326 9460 26332 9512
rect 26384 9500 26390 9512
rect 27154 9500 27160 9512
rect 26384 9472 27160 9500
rect 26384 9460 26390 9472
rect 27154 9460 27160 9472
rect 27212 9500 27218 9512
rect 28350 9500 28356 9512
rect 27212 9472 28356 9500
rect 27212 9460 27218 9472
rect 28350 9460 28356 9472
rect 28408 9460 28414 9512
rect 20128 9404 21864 9432
rect 20128 9392 20134 9404
rect 23106 9392 23112 9444
rect 23164 9432 23170 9444
rect 28258 9432 28264 9444
rect 23164 9404 28264 9432
rect 23164 9392 23170 9404
rect 28258 9392 28264 9404
rect 28316 9392 28322 9444
rect 7515 9336 9076 9364
rect 7515 9333 7527 9336
rect 7469 9327 7527 9333
rect 11514 9324 11520 9376
rect 11572 9324 11578 9376
rect 13906 9324 13912 9376
rect 13964 9324 13970 9376
rect 17770 9324 17776 9376
rect 17828 9324 17834 9376
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20588 9336 21281 9364
rect 20588 9324 20594 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 21634 9324 21640 9376
rect 21692 9364 21698 9376
rect 22094 9364 22100 9376
rect 21692 9336 22100 9364
rect 21692 9324 21698 9336
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 22462 9324 22468 9376
rect 22520 9324 22526 9376
rect 22833 9367 22891 9373
rect 22833 9333 22845 9367
rect 22879 9364 22891 9367
rect 23382 9364 23388 9376
rect 22879 9336 23388 9364
rect 22879 9333 22891 9336
rect 22833 9327 22891 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 24026 9324 24032 9376
rect 24084 9364 24090 9376
rect 24302 9364 24308 9376
rect 24084 9336 24308 9364
rect 24084 9324 24090 9336
rect 24302 9324 24308 9336
rect 24360 9324 24366 9376
rect 24762 9324 24768 9376
rect 24820 9324 24826 9376
rect 25133 9367 25191 9373
rect 25133 9333 25145 9367
rect 25179 9364 25191 9367
rect 25958 9364 25964 9376
rect 25179 9336 25964 9364
rect 25179 9333 25191 9336
rect 25133 9327 25191 9333
rect 25958 9324 25964 9336
rect 26016 9324 26022 9376
rect 26510 9324 26516 9376
rect 26568 9364 26574 9376
rect 26789 9367 26847 9373
rect 26789 9364 26801 9367
rect 26568 9336 26801 9364
rect 26568 9324 26574 9336
rect 26789 9333 26801 9336
rect 26835 9333 26847 9367
rect 26789 9327 26847 9333
rect 27154 9324 27160 9376
rect 27212 9324 27218 9376
rect 27798 9324 27804 9376
rect 27856 9324 27862 9376
rect 28552 9364 28580 9540
rect 28629 9537 28641 9571
rect 28675 9537 28687 9571
rect 28629 9531 28687 9537
rect 28896 9571 28954 9577
rect 28896 9537 28908 9571
rect 28942 9568 28954 9571
rect 29362 9568 29368 9580
rect 28942 9540 29368 9568
rect 28942 9537 28954 9540
rect 28896 9531 28954 9537
rect 29362 9528 29368 9540
rect 29420 9528 29426 9580
rect 30116 9509 30144 9608
rect 33045 9605 33057 9639
rect 33091 9636 33103 9639
rect 33980 9636 34008 9664
rect 33091 9608 34008 9636
rect 33091 9605 33103 9608
rect 33045 9599 33103 9605
rect 34146 9596 34152 9648
rect 34204 9636 34210 9648
rect 34422 9636 34428 9648
rect 34204 9608 34428 9636
rect 34204 9596 34210 9608
rect 34422 9596 34428 9608
rect 34480 9636 34486 9648
rect 35253 9639 35311 9645
rect 35253 9636 35265 9639
rect 34480 9608 35265 9636
rect 34480 9596 34486 9608
rect 35253 9605 35265 9608
rect 35299 9636 35311 9639
rect 38746 9636 38752 9648
rect 35299 9608 38752 9636
rect 35299 9605 35311 9608
rect 35253 9599 35311 9605
rect 38746 9596 38752 9608
rect 38804 9596 38810 9648
rect 39298 9596 39304 9648
rect 39356 9636 39362 9648
rect 39945 9639 40003 9645
rect 39945 9636 39957 9639
rect 39356 9608 39957 9636
rect 39356 9596 39362 9608
rect 39945 9605 39957 9608
rect 39991 9605 40003 9639
rect 39945 9599 40003 9605
rect 40313 9639 40371 9645
rect 40313 9605 40325 9639
rect 40359 9636 40371 9639
rect 42518 9636 42524 9648
rect 40359 9608 42524 9636
rect 40359 9605 40371 9608
rect 40313 9599 40371 9605
rect 42518 9596 42524 9608
rect 42576 9596 42582 9648
rect 43809 9639 43867 9645
rect 43809 9605 43821 9639
rect 43855 9636 43867 9639
rect 43990 9636 43996 9648
rect 43855 9608 43996 9636
rect 43855 9605 43867 9608
rect 43809 9599 43867 9605
rect 43990 9596 43996 9608
rect 44048 9596 44054 9648
rect 44100 9636 44128 9676
rect 51258 9664 51264 9716
rect 51316 9704 51322 9716
rect 51813 9707 51871 9713
rect 51316 9676 51488 9704
rect 51316 9664 51322 9676
rect 44910 9636 44916 9648
rect 44100 9608 44916 9636
rect 44910 9596 44916 9608
rect 44968 9596 44974 9648
rect 46382 9596 46388 9648
rect 46440 9636 46446 9648
rect 51460 9645 51488 9676
rect 51813 9673 51825 9707
rect 51859 9704 51871 9707
rect 52270 9704 52276 9716
rect 51859 9676 52276 9704
rect 51859 9673 51871 9676
rect 51813 9667 51871 9673
rect 52270 9664 52276 9676
rect 52328 9664 52334 9716
rect 53834 9664 53840 9716
rect 53892 9704 53898 9716
rect 54021 9707 54079 9713
rect 54021 9704 54033 9707
rect 53892 9676 54033 9704
rect 53892 9664 53898 9676
rect 54021 9673 54033 9676
rect 54067 9673 54079 9707
rect 54021 9667 54079 9673
rect 46937 9639 46995 9645
rect 46937 9636 46949 9639
rect 46440 9608 46949 9636
rect 46440 9596 46446 9608
rect 46937 9605 46949 9608
rect 46983 9605 46995 9639
rect 46937 9599 46995 9605
rect 51445 9639 51503 9645
rect 51445 9605 51457 9639
rect 51491 9605 51503 9639
rect 51445 9599 51503 9605
rect 52549 9639 52607 9645
rect 52549 9605 52561 9639
rect 52595 9636 52607 9639
rect 52730 9636 52736 9648
rect 52595 9608 52736 9636
rect 52595 9605 52607 9608
rect 52549 9599 52607 9605
rect 30368 9571 30426 9577
rect 30368 9537 30380 9571
rect 30414 9568 30426 9571
rect 30650 9568 30656 9580
rect 30414 9540 30656 9568
rect 30414 9537 30426 9540
rect 30368 9531 30426 9537
rect 30650 9528 30656 9540
rect 30708 9528 30714 9580
rect 33505 9571 33563 9577
rect 33505 9568 33517 9571
rect 31726 9540 33517 9568
rect 30101 9503 30159 9509
rect 30101 9469 30113 9503
rect 30147 9469 30159 9503
rect 30101 9463 30159 9469
rect 28994 9364 29000 9376
rect 28552 9336 29000 9364
rect 28994 9324 29000 9336
rect 29052 9324 29058 9376
rect 30116 9364 30144 9463
rect 31726 9432 31754 9540
rect 33505 9537 33517 9540
rect 33551 9568 33563 9571
rect 34793 9571 34851 9577
rect 34793 9568 34805 9571
rect 33551 9540 34805 9568
rect 33551 9537 33563 9540
rect 33505 9531 33563 9537
rect 34793 9537 34805 9540
rect 34839 9537 34851 9571
rect 34793 9531 34851 9537
rect 35434 9528 35440 9580
rect 35492 9568 35498 9580
rect 35492 9540 37872 9568
rect 35492 9528 35498 9540
rect 33137 9503 33195 9509
rect 33137 9469 33149 9503
rect 33183 9469 33195 9503
rect 33137 9463 33195 9469
rect 33229 9503 33287 9509
rect 33229 9469 33241 9503
rect 33275 9500 33287 9503
rect 34146 9500 34152 9512
rect 33275 9472 34152 9500
rect 33275 9469 33287 9472
rect 33229 9463 33287 9469
rect 31036 9404 31754 9432
rect 33152 9432 33180 9463
rect 34146 9460 34152 9472
rect 34204 9460 34210 9512
rect 34330 9460 34336 9512
rect 34388 9460 34394 9512
rect 35986 9460 35992 9512
rect 36044 9460 36050 9512
rect 33318 9432 33324 9444
rect 33152 9404 33324 9432
rect 30282 9364 30288 9376
rect 30116 9336 30288 9364
rect 30282 9324 30288 9336
rect 30340 9324 30346 9376
rect 30374 9324 30380 9376
rect 30432 9364 30438 9376
rect 31036 9364 31064 9404
rect 33318 9392 33324 9404
rect 33376 9392 33382 9444
rect 35526 9392 35532 9444
rect 35584 9432 35590 9444
rect 35805 9435 35863 9441
rect 35805 9432 35817 9435
rect 35584 9404 35817 9432
rect 35584 9392 35590 9404
rect 35805 9401 35817 9404
rect 35851 9432 35863 9435
rect 37844 9432 37872 9540
rect 39758 9528 39764 9580
rect 39816 9528 39822 9580
rect 43625 9571 43683 9577
rect 43625 9537 43637 9571
rect 43671 9568 43683 9571
rect 44634 9568 44640 9580
rect 43671 9540 44640 9568
rect 43671 9537 43683 9540
rect 43625 9531 43683 9537
rect 44634 9528 44640 9540
rect 44692 9528 44698 9580
rect 46753 9571 46811 9577
rect 46753 9537 46765 9571
rect 46799 9568 46811 9571
rect 47670 9568 47676 9580
rect 46799 9540 47676 9568
rect 46799 9537 46811 9540
rect 46753 9531 46811 9537
rect 47670 9528 47676 9540
rect 47728 9528 47734 9580
rect 50893 9571 50951 9577
rect 50893 9537 50905 9571
rect 50939 9568 50951 9571
rect 50982 9568 50988 9580
rect 50939 9540 50988 9568
rect 50939 9537 50951 9540
rect 50893 9531 50951 9537
rect 50982 9528 50988 9540
rect 51040 9528 51046 9580
rect 40402 9460 40408 9512
rect 40460 9460 40466 9512
rect 41138 9460 41144 9512
rect 41196 9460 41202 9512
rect 42426 9460 42432 9512
rect 42484 9460 42490 9512
rect 44085 9503 44143 9509
rect 44085 9469 44097 9503
rect 44131 9500 44143 9503
rect 44174 9500 44180 9512
rect 44131 9472 44180 9500
rect 44131 9469 44143 9472
rect 44085 9463 44143 9469
rect 44174 9460 44180 9472
rect 44232 9460 44238 9512
rect 45462 9460 45468 9512
rect 45520 9460 45526 9512
rect 48038 9460 48044 9512
rect 48096 9460 48102 9512
rect 48774 9460 48780 9512
rect 48832 9460 48838 9512
rect 49513 9503 49571 9509
rect 49513 9469 49525 9503
rect 49559 9500 49571 9503
rect 49878 9500 49884 9512
rect 49559 9472 49884 9500
rect 49559 9469 49571 9472
rect 49513 9463 49571 9469
rect 49878 9460 49884 9472
rect 49936 9460 49942 9512
rect 41322 9432 41328 9444
rect 35851 9404 37780 9432
rect 37844 9404 41328 9432
rect 35851 9401 35863 9404
rect 35805 9395 35863 9401
rect 37752 9376 37780 9404
rect 41322 9392 41328 9404
rect 41380 9392 41386 9444
rect 42794 9392 42800 9444
rect 42852 9432 42858 9444
rect 43254 9432 43260 9444
rect 42852 9404 43260 9432
rect 42852 9392 42858 9404
rect 43254 9392 43260 9404
rect 43312 9432 43318 9444
rect 52564 9432 52592 9599
rect 52730 9596 52736 9608
rect 52788 9596 52794 9648
rect 57974 9596 57980 9648
rect 58032 9636 58038 9648
rect 58437 9639 58495 9645
rect 58437 9636 58449 9639
rect 58032 9608 58449 9636
rect 58032 9596 58038 9608
rect 58437 9605 58449 9608
rect 58483 9605 58495 9639
rect 58437 9599 58495 9605
rect 54573 9503 54631 9509
rect 54573 9469 54585 9503
rect 54619 9469 54631 9503
rect 54573 9463 54631 9469
rect 43312 9404 52592 9432
rect 43312 9392 43318 9404
rect 54588 9376 54616 9463
rect 56134 9460 56140 9512
rect 56192 9460 56198 9512
rect 55858 9392 55864 9444
rect 55916 9432 55922 9444
rect 55916 9404 58112 9432
rect 55916 9392 55922 9404
rect 58084 9376 58112 9404
rect 30432 9336 31064 9364
rect 30432 9324 30438 9336
rect 31754 9324 31760 9376
rect 31812 9324 31818 9376
rect 36538 9324 36544 9376
rect 36596 9324 36602 9376
rect 36814 9324 36820 9376
rect 36872 9324 36878 9376
rect 37734 9324 37740 9376
rect 37792 9324 37798 9376
rect 40126 9324 40132 9376
rect 40184 9364 40190 9376
rect 41049 9367 41107 9373
rect 41049 9364 41061 9367
rect 40184 9336 41061 9364
rect 40184 9324 40190 9336
rect 41049 9333 41061 9336
rect 41095 9333 41107 9367
rect 41049 9327 41107 9333
rect 41230 9324 41236 9376
rect 41288 9364 41294 9376
rect 41785 9367 41843 9373
rect 41785 9364 41797 9367
rect 41288 9336 41797 9364
rect 41288 9324 41294 9336
rect 41785 9333 41797 9336
rect 41831 9333 41843 9367
rect 41785 9327 41843 9333
rect 43070 9324 43076 9376
rect 43128 9324 43134 9376
rect 43806 9324 43812 9376
rect 43864 9364 43870 9376
rect 44637 9367 44695 9373
rect 44637 9364 44649 9367
rect 43864 9336 44649 9364
rect 43864 9324 43870 9336
rect 44637 9333 44649 9336
rect 44683 9333 44695 9367
rect 44637 9327 44695 9333
rect 46109 9367 46167 9373
rect 46109 9333 46121 9367
rect 46155 9364 46167 9367
rect 46290 9364 46296 9376
rect 46155 9336 46296 9364
rect 46155 9333 46167 9336
rect 46109 9327 46167 9333
rect 46290 9324 46296 9336
rect 46348 9324 46354 9376
rect 46477 9367 46535 9373
rect 46477 9333 46489 9367
rect 46523 9364 46535 9367
rect 46658 9364 46664 9376
rect 46523 9336 46664 9364
rect 46523 9333 46535 9336
rect 46477 9327 46535 9333
rect 46658 9324 46664 9336
rect 46716 9324 46722 9376
rect 48130 9324 48136 9376
rect 48188 9364 48194 9376
rect 48593 9367 48651 9373
rect 48593 9364 48605 9367
rect 48188 9336 48605 9364
rect 48188 9324 48194 9336
rect 48593 9333 48605 9336
rect 48639 9333 48651 9367
rect 48593 9327 48651 9333
rect 49326 9324 49332 9376
rect 49384 9324 49390 9376
rect 50062 9324 50068 9376
rect 50120 9324 50126 9376
rect 54570 9324 54576 9376
rect 54628 9324 54634 9376
rect 55214 9324 55220 9376
rect 55272 9324 55278 9376
rect 56778 9324 56784 9376
rect 56836 9324 56842 9376
rect 56870 9324 56876 9376
rect 56928 9364 56934 9376
rect 57054 9364 57060 9376
rect 56928 9336 57060 9364
rect 56928 9324 56934 9336
rect 57054 9324 57060 9336
rect 57112 9324 57118 9376
rect 57422 9324 57428 9376
rect 57480 9324 57486 9376
rect 58066 9324 58072 9376
rect 58124 9324 58130 9376
rect 1104 9274 58880 9296
rect 1104 9222 8172 9274
rect 8224 9222 8236 9274
rect 8288 9222 8300 9274
rect 8352 9222 8364 9274
rect 8416 9222 8428 9274
rect 8480 9222 22616 9274
rect 22668 9222 22680 9274
rect 22732 9222 22744 9274
rect 22796 9222 22808 9274
rect 22860 9222 22872 9274
rect 22924 9222 37060 9274
rect 37112 9222 37124 9274
rect 37176 9222 37188 9274
rect 37240 9222 37252 9274
rect 37304 9222 37316 9274
rect 37368 9222 51504 9274
rect 51556 9222 51568 9274
rect 51620 9222 51632 9274
rect 51684 9222 51696 9274
rect 51748 9222 51760 9274
rect 51812 9222 58880 9274
rect 1104 9200 58880 9222
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3510 9160 3516 9172
rect 3007 9132 3516 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3694 9120 3700 9172
rect 3752 9160 3758 9172
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 3752 9132 3893 9160
rect 3752 9120 3758 9132
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 3881 9123 3939 9129
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 6825 9163 6883 9169
rect 6825 9160 6837 9163
rect 6420 9132 6837 9160
rect 6420 9120 6426 9132
rect 6825 9129 6837 9132
rect 6871 9129 6883 9163
rect 7098 9160 7104 9172
rect 6825 9123 6883 9129
rect 6932 9132 7104 9160
rect 3602 9092 3608 9104
rect 2700 9064 3608 9092
rect 2700 9033 2728 9064
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 6932 9092 6960 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 7340 9132 8309 9160
rect 7340 9120 7346 9132
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 9490 9160 9496 9172
rect 8536 9132 9496 9160
rect 8536 9120 8542 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 11146 9160 11152 9172
rect 11072 9132 11152 9160
rect 11072 9101 11100 9132
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11514 9120 11520 9172
rect 11572 9120 11578 9172
rect 11790 9120 11796 9172
rect 11848 9120 11854 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12621 9163 12679 9169
rect 12621 9160 12633 9163
rect 12032 9132 12633 9160
rect 12032 9120 12038 9132
rect 12621 9129 12633 9132
rect 12667 9129 12679 9163
rect 12621 9123 12679 9129
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14737 9163 14795 9169
rect 14737 9160 14749 9163
rect 13780 9132 14749 9160
rect 13780 9120 13786 9132
rect 14737 9129 14749 9132
rect 14783 9129 14795 9163
rect 14737 9123 14795 9129
rect 17770 9120 17776 9172
rect 17828 9120 17834 9172
rect 18230 9120 18236 9172
rect 18288 9120 18294 9172
rect 20073 9163 20131 9169
rect 20073 9129 20085 9163
rect 20119 9160 20131 9163
rect 20254 9160 20260 9172
rect 20119 9132 20260 9160
rect 20119 9129 20131 9132
rect 20073 9123 20131 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20714 9120 20720 9172
rect 20772 9120 20778 9172
rect 23382 9160 23388 9172
rect 20824 9132 23388 9160
rect 6380 9064 6960 9092
rect 11057 9095 11115 9101
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3421 9027 3479 9033
rect 3421 9024 3433 9027
rect 3016 8996 3433 9024
rect 3016 8984 3022 8996
rect 3421 8993 3433 8996
rect 3467 9024 3479 9027
rect 3467 8996 4016 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2976 8956 3004 8984
rect 2639 8928 3004 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 3050 8916 3056 8968
rect 3108 8916 3114 8968
rect 3207 8959 3265 8965
rect 3207 8925 3219 8959
rect 3253 8956 3265 8959
rect 3253 8928 3740 8956
rect 3253 8925 3265 8928
rect 3207 8919 3265 8925
rect 3712 8888 3740 8928
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 3988 8965 4016 8996
rect 5092 8996 5304 9024
rect 5092 8968 5120 8996
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 4706 8956 4712 8968
rect 3973 8919 4031 8925
rect 4080 8928 4712 8956
rect 4080 8888 4108 8928
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5074 8916 5080 8968
rect 5132 8916 5138 8968
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 5276 8956 5304 8996
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6380 9024 6408 9064
rect 11057 9061 11069 9095
rect 11103 9061 11115 9095
rect 11057 9055 11115 9061
rect 5960 8996 6408 9024
rect 5960 8984 5966 8996
rect 6380 8956 6408 8996
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 6788 8996 7052 9024
rect 6788 8984 6794 8996
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 5276 8928 6316 8956
rect 6380 8928 6469 8956
rect 5353 8891 5411 8897
rect 5353 8888 5365 8891
rect 3712 8860 4108 8888
rect 4632 8860 5365 8888
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3878 8820 3884 8832
rect 3200 8792 3884 8820
rect 3200 8780 3206 8792
rect 3878 8780 3884 8792
rect 3936 8820 3942 8832
rect 4632 8820 4660 8860
rect 5353 8857 5365 8860
rect 5399 8857 5411 8891
rect 5353 8851 5411 8857
rect 5445 8891 5503 8897
rect 5445 8857 5457 8891
rect 5491 8888 5503 8891
rect 6086 8888 6092 8900
rect 5491 8860 6092 8888
rect 5491 8857 5503 8860
rect 5445 8851 5503 8857
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 6288 8888 6316 8928
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6656 8888 6684 8919
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7024 8956 7052 8996
rect 9508 8996 10609 9024
rect 9508 8968 9536 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 11241 9027 11299 9033
rect 11241 8993 11253 9027
rect 11287 9024 11299 9027
rect 11532 9024 11560 9120
rect 12989 9095 13047 9101
rect 11624 9064 12434 9092
rect 11624 9036 11652 9064
rect 12406 9036 12434 9064
rect 12989 9061 13001 9095
rect 13035 9092 13047 9095
rect 13035 9064 14136 9092
rect 13035 9061 13047 9064
rect 12989 9055 13047 9061
rect 11287 8996 11560 9024
rect 11287 8993 11299 8996
rect 11241 8987 11299 8993
rect 7173 8959 7231 8965
rect 7173 8956 7185 8959
rect 7024 8928 7185 8956
rect 7173 8925 7185 8928
rect 7219 8925 7231 8959
rect 7173 8919 7231 8925
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9490 8916 9496 8968
rect 9548 8916 9554 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 10134 8956 10140 8968
rect 9815 8928 10140 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10612 8956 10640 8987
rect 11606 8984 11612 9036
rect 11664 8984 11670 9036
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 12342 8984 12348 9036
rect 12400 9024 12434 9036
rect 14108 9033 14136 9064
rect 13541 9027 13599 9033
rect 13541 9024 13553 9027
rect 12400 8996 13553 9024
rect 12400 8984 12406 8996
rect 13541 8993 13553 8996
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 17681 9027 17739 9033
rect 17681 8993 17693 9027
rect 17727 9024 17739 9027
rect 17788 9024 17816 9120
rect 19794 9052 19800 9104
rect 19852 9092 19858 9104
rect 20732 9092 20760 9120
rect 19852 9064 20760 9092
rect 19852 9052 19858 9064
rect 20824 9033 20852 9132
rect 23382 9120 23388 9132
rect 23440 9160 23446 9172
rect 24857 9163 24915 9169
rect 24857 9160 24869 9163
rect 23440 9132 24869 9160
rect 23440 9120 23446 9132
rect 24857 9129 24869 9132
rect 24903 9160 24915 9163
rect 26697 9163 26755 9169
rect 26697 9160 26709 9163
rect 24903 9132 26709 9160
rect 24903 9129 24915 9132
rect 24857 9123 24915 9129
rect 22462 9092 22468 9104
rect 22066 9064 22468 9092
rect 17727 8996 17816 9024
rect 20809 9027 20867 9033
rect 17727 8993 17739 8996
rect 17681 8987 17739 8993
rect 20809 8993 20821 9027
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 11422 8956 11428 8968
rect 10612 8928 11428 8956
rect 11422 8916 11428 8928
rect 11480 8956 11486 8968
rect 14642 8956 14648 8968
rect 11480 8928 14648 8956
rect 11480 8916 11486 8928
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 19702 8956 19708 8968
rect 18555 8928 19708 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 19702 8916 19708 8928
rect 19760 8956 19766 8968
rect 20714 8956 20720 8968
rect 19760 8928 20720 8956
rect 19760 8916 19766 8928
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 21076 8959 21134 8965
rect 21076 8925 21088 8959
rect 21122 8956 21134 8959
rect 22066 8956 22094 9064
rect 22462 9052 22468 9064
rect 22520 9052 22526 9104
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 23293 9095 23351 9101
rect 23293 9092 23305 9095
rect 23164 9064 23305 9092
rect 23164 9052 23170 9064
rect 23293 9061 23305 9064
rect 23339 9061 23351 9095
rect 23293 9055 23351 9061
rect 23308 9024 23336 9055
rect 24762 9052 24768 9104
rect 24820 9052 24826 9104
rect 24029 9027 24087 9033
rect 24029 9024 24041 9027
rect 23308 8996 24041 9024
rect 24029 8993 24041 8996
rect 24075 8993 24087 9027
rect 24029 8987 24087 8993
rect 21122 8928 22094 8956
rect 22373 8959 22431 8965
rect 21122 8925 21134 8928
rect 21076 8919 21134 8925
rect 22373 8925 22385 8959
rect 22419 8925 22431 8959
rect 22373 8919 22431 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24780 8956 24808 9052
rect 24964 9033 24992 9132
rect 26697 9129 26709 9132
rect 26743 9160 26755 9163
rect 27338 9160 27344 9172
rect 26743 9132 27344 9160
rect 26743 9129 26755 9132
rect 26697 9123 26755 9129
rect 27338 9120 27344 9132
rect 27396 9120 27402 9172
rect 29362 9120 29368 9172
rect 29420 9120 29426 9172
rect 39853 9163 39911 9169
rect 39853 9129 39865 9163
rect 39899 9160 39911 9163
rect 40402 9160 40408 9172
rect 39899 9132 40408 9160
rect 39899 9129 39911 9132
rect 39853 9123 39911 9129
rect 40402 9120 40408 9132
rect 40460 9120 40466 9172
rect 41230 9160 41236 9172
rect 40512 9132 41236 9160
rect 26329 9095 26387 9101
rect 26329 9092 26341 9095
rect 26068 9064 26341 9092
rect 24949 9027 25007 9033
rect 24949 8993 24961 9027
rect 24995 8993 25007 9027
rect 24949 8987 25007 8993
rect 23891 8928 24808 8956
rect 25216 8959 25274 8965
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 25216 8925 25228 8959
rect 25262 8956 25274 8959
rect 25774 8956 25780 8968
rect 25262 8928 25780 8956
rect 25262 8925 25274 8928
rect 25216 8919 25274 8925
rect 6288 8860 8064 8888
rect 8036 8832 8064 8860
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 10873 8891 10931 8897
rect 8352 8860 10456 8888
rect 8352 8848 8358 8860
rect 3936 8792 4660 8820
rect 3936 8780 3942 8792
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4764 8792 4813 8820
rect 4764 8780 4770 8792
rect 4801 8789 4813 8792
rect 4847 8820 4859 8823
rect 4982 8820 4988 8832
rect 4847 8792 4988 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 5626 8820 5632 8832
rect 5123 8792 5632 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 7834 8820 7840 8832
rect 6604 8792 7840 8820
rect 6604 8780 6610 8792
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 8665 8823 8723 8829
rect 8665 8820 8677 8823
rect 8628 8792 8677 8820
rect 8628 8780 8634 8792
rect 8665 8789 8677 8792
rect 8711 8789 8723 8823
rect 8665 8783 8723 8789
rect 9582 8780 9588 8832
rect 9640 8780 9646 8832
rect 10318 8780 10324 8832
rect 10376 8780 10382 8832
rect 10428 8820 10456 8860
rect 10873 8857 10885 8891
rect 10919 8888 10931 8891
rect 11054 8888 11060 8900
rect 10919 8860 11060 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 11756 8860 13369 8888
rect 11756 8848 11762 8860
rect 13357 8857 13369 8860
rect 13403 8888 13415 8891
rect 13403 8860 13860 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13832 8832 13860 8860
rect 15838 8848 15844 8900
rect 15896 8888 15902 8900
rect 16209 8891 16267 8897
rect 16209 8888 16221 8891
rect 15896 8860 16221 8888
rect 15896 8848 15902 8860
rect 16209 8857 16221 8860
rect 16255 8888 16267 8891
rect 17310 8888 17316 8900
rect 16255 8860 17316 8888
rect 16255 8857 16267 8860
rect 16209 8851 16267 8857
rect 17310 8848 17316 8860
rect 17368 8848 17374 8900
rect 17880 8860 19196 8888
rect 17880 8832 17908 8860
rect 13262 8820 13268 8832
rect 10428 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 13814 8780 13820 8832
rect 13872 8780 13878 8832
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 17276 8792 17417 8820
rect 17276 8780 17282 8792
rect 17405 8789 17417 8792
rect 17451 8820 17463 8823
rect 17862 8820 17868 8832
rect 17451 8792 17868 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 19058 8780 19064 8832
rect 19116 8780 19122 8832
rect 19168 8820 19196 8860
rect 19610 8848 19616 8900
rect 19668 8888 19674 8900
rect 19981 8891 20039 8897
rect 19981 8888 19993 8891
rect 19668 8860 19993 8888
rect 19668 8848 19674 8860
rect 19981 8857 19993 8860
rect 20027 8857 20039 8891
rect 19981 8851 20039 8857
rect 20622 8848 20628 8900
rect 20680 8888 20686 8900
rect 20680 8860 21036 8888
rect 20680 8848 20686 8860
rect 19794 8820 19800 8832
rect 19168 8792 19800 8820
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 20346 8820 20352 8832
rect 19944 8792 20352 8820
rect 19944 8780 19950 8792
rect 20346 8780 20352 8792
rect 20404 8820 20410 8832
rect 20717 8823 20775 8829
rect 20717 8820 20729 8823
rect 20404 8792 20729 8820
rect 20404 8780 20410 8792
rect 20717 8789 20729 8792
rect 20763 8789 20775 8823
rect 21008 8820 21036 8860
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 22388 8888 22416 8919
rect 25774 8916 25780 8928
rect 25832 8916 25838 8968
rect 21232 8860 22416 8888
rect 21232 8848 21238 8860
rect 22189 8823 22247 8829
rect 22189 8820 22201 8823
rect 21008 8792 22201 8820
rect 20717 8783 20775 8789
rect 22189 8789 22201 8792
rect 22235 8789 22247 8823
rect 22189 8783 22247 8789
rect 23014 8780 23020 8832
rect 23072 8780 23078 8832
rect 23474 8780 23480 8832
rect 23532 8780 23538 8832
rect 23937 8823 23995 8829
rect 23937 8789 23949 8823
rect 23983 8820 23995 8823
rect 24486 8820 24492 8832
rect 23983 8792 24492 8820
rect 23983 8789 23995 8792
rect 23937 8783 23995 8789
rect 24486 8780 24492 8792
rect 24544 8780 24550 8832
rect 24762 8780 24768 8832
rect 24820 8820 24826 8832
rect 26068 8820 26096 9064
rect 26329 9061 26341 9064
rect 26375 9061 26387 9095
rect 26329 9055 26387 9061
rect 26344 9024 26372 9055
rect 28810 9052 28816 9104
rect 28868 9092 28874 9104
rect 29549 9095 29607 9101
rect 29549 9092 29561 9095
rect 28868 9064 29561 9092
rect 28868 9052 28874 9064
rect 29549 9061 29561 9064
rect 29595 9061 29607 9095
rect 40512 9092 40540 9132
rect 41230 9120 41236 9132
rect 41288 9120 41294 9172
rect 41322 9120 41328 9172
rect 41380 9160 41386 9172
rect 47394 9160 47400 9172
rect 41380 9132 47400 9160
rect 41380 9120 41386 9132
rect 47394 9120 47400 9132
rect 47452 9120 47458 9172
rect 48038 9120 48044 9172
rect 48096 9120 48102 9172
rect 49326 9120 49332 9172
rect 49384 9120 49390 9172
rect 56045 9163 56103 9169
rect 56045 9129 56057 9163
rect 56091 9160 56103 9163
rect 56134 9160 56140 9172
rect 56091 9132 56140 9160
rect 56091 9129 56103 9132
rect 56045 9123 56103 9129
rect 56134 9120 56140 9132
rect 56192 9120 56198 9172
rect 56870 9120 56876 9172
rect 56928 9120 56934 9172
rect 29549 9055 29607 9061
rect 40420 9064 40540 9092
rect 26881 9027 26939 9033
rect 26881 9024 26893 9027
rect 26344 8996 26893 9024
rect 26881 8993 26893 8996
rect 26927 8993 26939 9027
rect 30101 9027 30159 9033
rect 30101 9024 30113 9027
rect 26881 8987 26939 8993
rect 28736 8996 30113 9024
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8956 28687 8959
rect 28736 8956 28764 8996
rect 30101 8993 30113 8996
rect 30147 9024 30159 9027
rect 30147 8996 30512 9024
rect 30147 8993 30159 8996
rect 30101 8987 30159 8993
rect 28675 8928 28764 8956
rect 28675 8925 28687 8928
rect 28629 8919 28687 8925
rect 26142 8848 26148 8900
rect 26200 8888 26206 8900
rect 28644 8888 28672 8919
rect 28810 8916 28816 8968
rect 28868 8916 28874 8968
rect 28902 8916 28908 8968
rect 28960 8956 28966 8968
rect 30374 8956 30380 8968
rect 28960 8928 30380 8956
rect 28960 8916 28966 8928
rect 30374 8916 30380 8928
rect 30432 8916 30438 8968
rect 30484 8956 30512 8996
rect 30926 8984 30932 9036
rect 30984 8984 30990 9036
rect 31297 9027 31355 9033
rect 31297 8993 31309 9027
rect 31343 9024 31355 9027
rect 31478 9024 31484 9036
rect 31343 8996 31484 9024
rect 31343 8993 31355 8996
rect 31297 8987 31355 8993
rect 31478 8984 31484 8996
rect 31536 8984 31542 9036
rect 40310 9024 40316 9036
rect 34900 8996 40316 9024
rect 32214 8956 32220 8968
rect 30484 8928 32220 8956
rect 32214 8916 32220 8928
rect 32272 8916 32278 8968
rect 34900 8965 34928 8996
rect 40310 8984 40316 8996
rect 40368 8984 40374 9036
rect 32493 8959 32551 8965
rect 32493 8925 32505 8959
rect 32539 8956 32551 8959
rect 34885 8959 34943 8965
rect 34885 8956 34897 8959
rect 32539 8928 34897 8956
rect 32539 8925 32551 8928
rect 32493 8919 32551 8925
rect 34885 8925 34897 8928
rect 34931 8925 34943 8959
rect 35437 8959 35495 8965
rect 35437 8956 35449 8959
rect 34885 8919 34943 8925
rect 35268 8928 35449 8956
rect 26200 8860 28672 8888
rect 26200 8848 26206 8860
rect 29086 8848 29092 8900
rect 29144 8848 29150 8900
rect 29730 8848 29736 8900
rect 29788 8888 29794 8900
rect 30009 8891 30067 8897
rect 30009 8888 30021 8891
rect 29788 8860 30021 8888
rect 29788 8848 29794 8860
rect 30009 8857 30021 8860
rect 30055 8857 30067 8891
rect 30745 8891 30803 8897
rect 30009 8851 30067 8857
rect 30116 8860 30512 8888
rect 24820 8792 26096 8820
rect 24820 8780 24826 8792
rect 27522 8780 27528 8832
rect 27580 8780 27586 8832
rect 29104 8820 29132 8848
rect 29638 8820 29644 8832
rect 29104 8792 29644 8820
rect 29638 8780 29644 8792
rect 29696 8820 29702 8832
rect 29917 8823 29975 8829
rect 29917 8820 29929 8823
rect 29696 8792 29929 8820
rect 29696 8780 29702 8792
rect 29917 8789 29929 8792
rect 29963 8820 29975 8823
rect 30116 8820 30144 8860
rect 29963 8792 30144 8820
rect 29963 8789 29975 8792
rect 29917 8783 29975 8789
rect 30374 8780 30380 8832
rect 30432 8780 30438 8832
rect 30484 8820 30512 8860
rect 30745 8857 30757 8891
rect 30791 8888 30803 8891
rect 31849 8891 31907 8897
rect 31849 8888 31861 8891
rect 30791 8860 31861 8888
rect 30791 8857 30803 8860
rect 30745 8851 30803 8857
rect 31849 8857 31861 8860
rect 31895 8857 31907 8891
rect 31849 8851 31907 8857
rect 30837 8823 30895 8829
rect 30837 8820 30849 8823
rect 30484 8792 30849 8820
rect 30837 8789 30849 8792
rect 30883 8789 30895 8823
rect 30837 8783 30895 8789
rect 33965 8823 34023 8829
rect 33965 8789 33977 8823
rect 34011 8820 34023 8823
rect 34238 8820 34244 8832
rect 34011 8792 34244 8820
rect 34011 8789 34023 8792
rect 33965 8783 34023 8789
rect 34238 8780 34244 8792
rect 34296 8780 34302 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 35268 8829 35296 8928
rect 35437 8925 35449 8928
rect 35483 8925 35495 8959
rect 35437 8919 35495 8925
rect 36078 8916 36084 8968
rect 36136 8956 36142 8968
rect 36541 8959 36599 8965
rect 36541 8956 36553 8959
rect 36136 8928 36553 8956
rect 36136 8916 36142 8928
rect 36541 8925 36553 8928
rect 36587 8956 36599 8959
rect 36814 8956 36820 8968
rect 36587 8928 36820 8956
rect 36587 8925 36599 8928
rect 36541 8919 36599 8925
rect 36814 8916 36820 8928
rect 36872 8916 36878 8968
rect 37645 8959 37703 8965
rect 37645 8925 37657 8959
rect 37691 8925 37703 8959
rect 37645 8919 37703 8925
rect 36265 8891 36323 8897
rect 36265 8857 36277 8891
rect 36311 8888 36323 8891
rect 36906 8888 36912 8900
rect 36311 8860 36912 8888
rect 36311 8857 36323 8860
rect 36265 8851 36323 8857
rect 36906 8848 36912 8860
rect 36964 8848 36970 8900
rect 37369 8891 37427 8897
rect 37369 8857 37381 8891
rect 37415 8888 37427 8891
rect 37458 8888 37464 8900
rect 37415 8860 37464 8888
rect 37415 8857 37427 8860
rect 37369 8851 37427 8857
rect 37458 8848 37464 8860
rect 37516 8848 37522 8900
rect 35253 8823 35311 8829
rect 35253 8820 35265 8823
rect 34572 8792 35265 8820
rect 34572 8780 34578 8792
rect 35253 8789 35265 8792
rect 35299 8789 35311 8823
rect 35253 8783 35311 8789
rect 36722 8780 36728 8832
rect 36780 8820 36786 8832
rect 37660 8820 37688 8919
rect 38838 8916 38844 8968
rect 38896 8916 38902 8968
rect 40313 8891 40371 8897
rect 40313 8857 40325 8891
rect 40359 8888 40371 8891
rect 40420 8888 40448 9064
rect 40770 9052 40776 9104
rect 40828 9092 40834 9104
rect 41141 9095 41199 9101
rect 40828 9064 41092 9092
rect 40828 9052 40834 9064
rect 40497 9027 40555 9033
rect 40497 8993 40509 9027
rect 40543 9024 40555 9027
rect 41064 9024 41092 9064
rect 41141 9061 41153 9095
rect 41187 9092 41199 9095
rect 41187 9064 42012 9092
rect 41187 9061 41199 9064
rect 41141 9055 41199 9061
rect 41601 9027 41659 9033
rect 41601 9024 41613 9027
rect 40543 8996 41000 9024
rect 41064 8996 41613 9024
rect 40543 8993 40555 8996
rect 40497 8987 40555 8993
rect 40359 8860 40448 8888
rect 40359 8857 40371 8860
rect 40313 8851 40371 8857
rect 40770 8848 40776 8900
rect 40828 8848 40834 8900
rect 36780 8792 37688 8820
rect 36780 8780 36786 8792
rect 38286 8780 38292 8832
rect 38344 8780 38350 8832
rect 38654 8780 38660 8832
rect 38712 8820 38718 8832
rect 39393 8823 39451 8829
rect 39393 8820 39405 8823
rect 38712 8792 39405 8820
rect 38712 8780 38718 8792
rect 39393 8789 39405 8792
rect 39439 8789 39451 8823
rect 39393 8783 39451 8789
rect 40218 8780 40224 8832
rect 40276 8820 40282 8832
rect 40788 8820 40816 8848
rect 40972 8829 41000 8996
rect 41601 8993 41613 8996
rect 41647 8993 41659 9027
rect 41601 8987 41659 8993
rect 41782 8984 41788 9036
rect 41840 8984 41846 9036
rect 41984 9033 42012 9064
rect 43070 9052 43076 9104
rect 43128 9052 43134 9104
rect 43349 9095 43407 9101
rect 43349 9061 43361 9095
rect 43395 9092 43407 9095
rect 46109 9095 46167 9101
rect 43395 9064 44220 9092
rect 43395 9061 43407 9064
rect 43349 9055 43407 9061
rect 41969 9027 42027 9033
rect 41969 8993 41981 9027
rect 42015 8993 42027 9027
rect 41969 8987 42027 8993
rect 41509 8959 41567 8965
rect 41509 8925 41521 8959
rect 41555 8956 41567 8959
rect 43088 8956 43116 9052
rect 43806 8984 43812 9036
rect 43864 8984 43870 9036
rect 44192 9033 44220 9064
rect 46109 9061 46121 9095
rect 46155 9092 46167 9095
rect 49344 9092 49372 9120
rect 57330 9092 57336 9104
rect 46155 9064 46980 9092
rect 46155 9061 46167 9064
rect 46109 9055 46167 9061
rect 43993 9027 44051 9033
rect 43993 8993 44005 9027
rect 44039 8993 44051 9027
rect 43993 8987 44051 8993
rect 44177 9027 44235 9033
rect 44177 8993 44189 9027
rect 44223 8993 44235 9027
rect 44177 8987 44235 8993
rect 44284 8996 45508 9024
rect 41555 8928 43116 8956
rect 43257 8959 43315 8965
rect 41555 8925 41567 8928
rect 41509 8919 41567 8925
rect 43257 8925 43269 8959
rect 43303 8956 43315 8959
rect 43346 8956 43352 8968
rect 43303 8928 43352 8956
rect 43303 8925 43315 8928
rect 43257 8919 43315 8925
rect 43346 8916 43352 8928
rect 43404 8956 43410 8968
rect 44008 8956 44036 8987
rect 44284 8956 44312 8996
rect 43404 8928 44312 8956
rect 43404 8916 43410 8928
rect 44910 8916 44916 8968
rect 44968 8956 44974 8968
rect 45005 8959 45063 8965
rect 45005 8956 45017 8959
rect 44968 8928 45017 8956
rect 44968 8916 44974 8928
rect 45005 8925 45017 8928
rect 45051 8925 45063 8959
rect 45480 8956 45508 8996
rect 45830 8984 45836 9036
rect 45888 8984 45894 9036
rect 46290 8984 46296 9036
rect 46348 9024 46354 9036
rect 46569 9027 46627 9033
rect 46569 9024 46581 9027
rect 46348 8996 46581 9024
rect 46348 8984 46354 8996
rect 46569 8993 46581 8996
rect 46615 8993 46627 9027
rect 46569 8987 46627 8993
rect 46658 8984 46664 9036
rect 46716 8984 46722 9036
rect 46952 9033 46980 9064
rect 48516 9064 49372 9092
rect 54128 9064 57336 9092
rect 48516 9033 48544 9064
rect 46937 9027 46995 9033
rect 46937 8993 46949 9027
rect 46983 8993 46995 9027
rect 46937 8987 46995 8993
rect 48501 9027 48559 9033
rect 48501 8993 48513 9027
rect 48547 8993 48559 9027
rect 48501 8987 48559 8993
rect 48685 9027 48743 9033
rect 48685 8993 48697 9027
rect 48731 9024 48743 9027
rect 52270 9024 52276 9036
rect 48731 8996 52276 9024
rect 48731 8993 48743 8996
rect 48685 8987 48743 8993
rect 45480 8928 47900 8956
rect 45005 8919 45063 8925
rect 43717 8891 43775 8897
rect 43717 8857 43729 8891
rect 43763 8888 43775 8891
rect 44726 8888 44732 8900
rect 43763 8860 44732 8888
rect 43763 8857 43775 8860
rect 43717 8851 43775 8857
rect 44726 8848 44732 8860
rect 44784 8888 44790 8900
rect 44784 8860 45232 8888
rect 44784 8848 44790 8860
rect 40276 8792 40816 8820
rect 40957 8823 41015 8829
rect 40276 8780 40282 8792
rect 40957 8789 40969 8823
rect 41003 8820 41015 8823
rect 42334 8820 42340 8832
rect 41003 8792 42340 8820
rect 41003 8789 41015 8792
rect 40957 8783 41015 8789
rect 42334 8780 42340 8792
rect 42392 8780 42398 8832
rect 42610 8780 42616 8832
rect 42668 8780 42674 8832
rect 43898 8780 43904 8832
rect 43956 8820 43962 8832
rect 44821 8823 44879 8829
rect 44821 8820 44833 8823
rect 43956 8792 44833 8820
rect 43956 8780 43962 8792
rect 44821 8789 44833 8792
rect 44867 8789 44879 8823
rect 45204 8820 45232 8860
rect 46658 8848 46664 8900
rect 46716 8888 46722 8900
rect 47872 8897 47900 8928
rect 47946 8916 47952 8968
rect 48004 8956 48010 8968
rect 48869 8959 48927 8965
rect 48869 8956 48881 8959
rect 48004 8928 48881 8956
rect 48004 8916 48010 8928
rect 48869 8925 48881 8928
rect 48915 8925 48927 8959
rect 48869 8919 48927 8925
rect 47857 8891 47915 8897
rect 46716 8860 47808 8888
rect 46716 8848 46722 8860
rect 46477 8823 46535 8829
rect 46477 8820 46489 8823
rect 45204 8792 46489 8820
rect 44821 8783 44879 8789
rect 46477 8789 46489 8792
rect 46523 8789 46535 8823
rect 46477 8783 46535 8789
rect 46566 8780 46572 8832
rect 46624 8820 46630 8832
rect 47581 8823 47639 8829
rect 47581 8820 47593 8823
rect 46624 8792 47593 8820
rect 46624 8780 46630 8792
rect 47581 8789 47593 8792
rect 47627 8789 47639 8823
rect 47780 8820 47808 8860
rect 47857 8857 47869 8891
rect 47903 8888 47915 8891
rect 48976 8888 49004 8996
rect 52270 8984 52276 8996
rect 52328 8984 52334 9036
rect 53834 8984 53840 9036
rect 53892 8984 53898 9036
rect 50154 8916 50160 8968
rect 50212 8916 50218 8968
rect 52546 8916 52552 8968
rect 52604 8956 52610 8968
rect 52825 8959 52883 8965
rect 52825 8956 52837 8959
rect 52604 8928 52837 8956
rect 52604 8916 52610 8928
rect 52825 8925 52837 8928
rect 52871 8956 52883 8959
rect 53852 8956 53880 8984
rect 52871 8928 53880 8956
rect 52871 8925 52883 8928
rect 52825 8919 52883 8925
rect 47903 8860 49004 8888
rect 53092 8891 53150 8897
rect 47903 8857 47915 8860
rect 47857 8851 47915 8857
rect 53092 8857 53104 8891
rect 53138 8888 53150 8891
rect 54018 8888 54024 8900
rect 53138 8860 54024 8888
rect 53138 8857 53150 8860
rect 53092 8851 53150 8857
rect 54018 8848 54024 8860
rect 54076 8848 54082 8900
rect 54128 8832 54156 9064
rect 57330 9052 57336 9064
rect 57388 9092 57394 9104
rect 57388 9064 57744 9092
rect 57388 9052 57394 9064
rect 54941 9027 54999 9033
rect 54941 8993 54953 9027
rect 54987 9024 54999 9027
rect 55490 9024 55496 9036
rect 54987 8996 55496 9024
rect 54987 8993 54999 8996
rect 54941 8987 54999 8993
rect 55490 8984 55496 8996
rect 55548 8984 55554 9036
rect 55953 9027 56011 9033
rect 55953 8993 55965 9027
rect 55999 9024 56011 9027
rect 56226 9024 56232 9036
rect 55999 8996 56232 9024
rect 55999 8993 56011 8996
rect 55953 8987 56011 8993
rect 56226 8984 56232 8996
rect 56284 9024 56290 9036
rect 56597 9027 56655 9033
rect 56597 9024 56609 9027
rect 56284 8996 56609 9024
rect 56284 8984 56290 8996
rect 56597 8993 56609 8996
rect 56643 8993 56655 9027
rect 56597 8987 56655 8993
rect 57054 8984 57060 9036
rect 57112 9024 57118 9036
rect 57716 9033 57744 9064
rect 57425 9027 57483 9033
rect 57425 9024 57437 9027
rect 57112 8996 57437 9024
rect 57112 8984 57118 8996
rect 57425 8993 57437 8996
rect 57471 8993 57483 9027
rect 57425 8987 57483 8993
rect 57701 9027 57759 9033
rect 57701 8993 57713 9027
rect 57747 8993 57759 9027
rect 57701 8987 57759 8993
rect 54662 8916 54668 8968
rect 54720 8916 54726 8968
rect 57241 8959 57299 8965
rect 57241 8925 57253 8959
rect 57287 8956 57299 8959
rect 57606 8956 57612 8968
rect 57287 8928 57612 8956
rect 57287 8925 57299 8928
rect 57241 8919 57299 8925
rect 57606 8916 57612 8928
rect 57664 8916 57670 8968
rect 54757 8891 54815 8897
rect 54220 8860 54616 8888
rect 48314 8820 48320 8832
rect 47780 8792 48320 8820
rect 47581 8783 47639 8789
rect 48314 8780 48320 8792
rect 48372 8780 48378 8832
rect 48406 8780 48412 8832
rect 48464 8780 48470 8832
rect 48682 8780 48688 8832
rect 48740 8820 48746 8832
rect 49513 8823 49571 8829
rect 49513 8820 49525 8823
rect 48740 8792 49525 8820
rect 48740 8780 48746 8792
rect 49513 8789 49525 8792
rect 49559 8789 49571 8823
rect 49513 8783 49571 8789
rect 50798 8780 50804 8832
rect 50856 8780 50862 8832
rect 54110 8780 54116 8832
rect 54168 8780 54174 8832
rect 54220 8829 54248 8860
rect 54588 8832 54616 8860
rect 54757 8857 54769 8891
rect 54803 8888 54815 8891
rect 55766 8888 55772 8900
rect 54803 8860 55772 8888
rect 54803 8857 54815 8860
rect 54757 8851 54815 8857
rect 55766 8848 55772 8860
rect 55824 8848 55830 8900
rect 56505 8891 56563 8897
rect 56505 8857 56517 8891
rect 56551 8888 56563 8891
rect 58345 8891 58403 8897
rect 58345 8888 58357 8891
rect 56551 8860 58357 8888
rect 56551 8857 56563 8860
rect 56505 8851 56563 8857
rect 58345 8857 58357 8860
rect 58391 8857 58403 8891
rect 58345 8851 58403 8857
rect 54205 8823 54263 8829
rect 54205 8789 54217 8823
rect 54251 8789 54263 8823
rect 54205 8783 54263 8789
rect 54294 8780 54300 8832
rect 54352 8780 54358 8832
rect 54570 8780 54576 8832
rect 54628 8780 54634 8832
rect 55490 8780 55496 8832
rect 55548 8780 55554 8832
rect 55582 8780 55588 8832
rect 55640 8820 55646 8832
rect 56413 8823 56471 8829
rect 56413 8820 56425 8823
rect 55640 8792 56425 8820
rect 55640 8780 55646 8792
rect 56413 8789 56425 8792
rect 56459 8820 56471 8823
rect 57333 8823 57391 8829
rect 57333 8820 57345 8823
rect 56459 8792 57345 8820
rect 56459 8789 56471 8792
rect 56413 8783 56471 8789
rect 57333 8789 57345 8792
rect 57379 8789 57391 8823
rect 57333 8783 57391 8789
rect 1104 8730 59040 8752
rect 1104 8678 15394 8730
rect 15446 8678 15458 8730
rect 15510 8678 15522 8730
rect 15574 8678 15586 8730
rect 15638 8678 15650 8730
rect 15702 8678 29838 8730
rect 29890 8678 29902 8730
rect 29954 8678 29966 8730
rect 30018 8678 30030 8730
rect 30082 8678 30094 8730
rect 30146 8678 44282 8730
rect 44334 8678 44346 8730
rect 44398 8678 44410 8730
rect 44462 8678 44474 8730
rect 44526 8678 44538 8730
rect 44590 8678 58726 8730
rect 58778 8678 58790 8730
rect 58842 8678 58854 8730
rect 58906 8678 58918 8730
rect 58970 8678 58982 8730
rect 59034 8678 59040 8730
rect 1104 8656 59040 8678
rect 2866 8576 2872 8628
rect 2924 8576 2930 8628
rect 3602 8576 3608 8628
rect 3660 8576 3666 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8585 4215 8619
rect 4157 8579 4215 8585
rect 2884 8548 2912 8576
rect 4172 8548 4200 8579
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 4439 8619 4497 8625
rect 4439 8585 4451 8619
rect 4485 8616 4497 8619
rect 5166 8616 5172 8628
rect 4485 8588 5172 8616
rect 4485 8585 4497 8588
rect 4439 8579 4497 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7653 8619 7711 8625
rect 7653 8616 7665 8619
rect 7524 8588 7665 8616
rect 7524 8576 7530 8588
rect 7653 8585 7665 8588
rect 7699 8585 7711 8619
rect 7653 8579 7711 8585
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8573 8619 8631 8625
rect 7892 8588 8524 8616
rect 7892 8576 7898 8588
rect 2884 8520 4200 8548
rect 4356 8548 4384 8576
rect 4356 8520 4660 8548
rect 4632 8489 4660 8520
rect 4706 8508 4712 8560
rect 4764 8508 4770 8560
rect 4909 8551 4967 8557
rect 4909 8548 4921 8551
rect 4816 8520 4921 8548
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 4341 8483 4399 8489
rect 3007 8452 3740 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3712 8421 3740 8452
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 4816 8480 4844 8520
rect 4909 8517 4921 8520
rect 4955 8517 4967 8551
rect 4909 8511 4967 8517
rect 5074 8508 5080 8560
rect 5132 8508 5138 8560
rect 6012 8548 6040 8576
rect 8113 8551 8171 8557
rect 8113 8548 8125 8551
rect 6012 8520 8125 8548
rect 8113 8517 8125 8520
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 8294 8508 8300 8560
rect 8352 8508 8358 8560
rect 8496 8548 8524 8588
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8938 8616 8944 8628
rect 8619 8588 8944 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 10318 8616 10324 8628
rect 9079 8588 10324 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11756 8588 13124 8616
rect 11756 8576 11762 8588
rect 8662 8548 8668 8560
rect 8496 8520 8668 8548
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 11977 8551 12035 8557
rect 8956 8520 11836 8548
rect 4663 8452 4844 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 4062 8412 4068 8424
rect 3743 8384 4068 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 3068 8344 3096 8375
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 3602 8344 3608 8356
rect 3068 8316 3608 8344
rect 3602 8304 3608 8316
rect 3660 8344 3666 8356
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 3660 8316 3985 8344
rect 3660 8304 3666 8316
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 4356 8344 4384 8443
rect 4540 8412 4568 8443
rect 4540 8384 4936 8412
rect 4706 8344 4712 8356
rect 4356 8316 4712 8344
rect 3973 8307 4031 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4908 8288 4936 8384
rect 5092 8353 5120 8508
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 6178 8480 6184 8492
rect 5399 8452 6184 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6270 8440 6276 8492
rect 6328 8440 6334 8492
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 6822 8480 6828 8492
rect 6779 8452 6828 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 6822 8440 6828 8452
rect 6880 8480 6886 8492
rect 7006 8480 7012 8492
rect 6880 8452 7012 8480
rect 6880 8440 6886 8452
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7116 8452 7757 8480
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6052 8384 6224 8412
rect 6052 8372 6058 8384
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8313 5135 8347
rect 5077 8307 5135 8313
rect 4890 8236 4896 8288
rect 4948 8236 4954 8288
rect 6196 8276 6224 8384
rect 6288 8344 6316 8440
rect 6380 8412 6408 8440
rect 7116 8412 7144 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7926 8440 7932 8492
rect 7984 8440 7990 8492
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 6380 8384 7144 8412
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 7248 8384 7297 8412
rect 7248 8372 7254 8384
rect 7285 8381 7297 8384
rect 7331 8412 7343 8415
rect 8312 8412 8340 8508
rect 8570 8440 8576 8492
rect 8628 8440 8634 8492
rect 8956 8489 8984 8520
rect 11808 8492 11836 8520
rect 11977 8517 11989 8551
rect 12023 8548 12035 8551
rect 12986 8548 12992 8560
rect 12023 8520 12992 8548
rect 12023 8517 12035 8520
rect 11977 8511 12035 8517
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 13096 8548 13124 8588
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13504 8588 13553 8616
rect 13504 8576 13510 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 14550 8616 14556 8628
rect 13955 8588 14556 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 13924 8548 13952 8579
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 19702 8576 19708 8628
rect 19760 8576 19766 8628
rect 20070 8576 20076 8628
rect 20128 8576 20134 8628
rect 20530 8576 20536 8628
rect 20588 8576 20594 8628
rect 20901 8619 20959 8625
rect 20901 8585 20913 8619
rect 20947 8616 20959 8619
rect 21174 8616 21180 8628
rect 20947 8588 21180 8616
rect 20947 8585 20959 8588
rect 20901 8579 20959 8585
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21634 8616 21640 8628
rect 21315 8588 21640 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 23290 8616 23296 8628
rect 21744 8588 23296 8616
rect 13096 8520 13952 8548
rect 18233 8551 18291 8557
rect 18233 8517 18245 8551
rect 18279 8548 18291 8551
rect 18570 8551 18628 8557
rect 18570 8548 18582 8551
rect 18279 8520 18582 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18570 8517 18582 8520
rect 18616 8517 18628 8551
rect 21744 8548 21772 8588
rect 23290 8576 23296 8588
rect 23348 8576 23354 8628
rect 23382 8576 23388 8628
rect 23440 8576 23446 8628
rect 25774 8616 25780 8628
rect 24228 8588 25780 8616
rect 23400 8548 23428 8576
rect 24228 8560 24256 8588
rect 25774 8576 25780 8588
rect 25832 8576 25838 8628
rect 26234 8576 26240 8628
rect 26292 8616 26298 8628
rect 26973 8619 27031 8625
rect 26973 8616 26985 8619
rect 26292 8588 26985 8616
rect 26292 8576 26298 8588
rect 26973 8585 26985 8588
rect 27019 8585 27031 8619
rect 26973 8579 27031 8585
rect 27433 8619 27491 8625
rect 27433 8585 27445 8619
rect 27479 8616 27491 8619
rect 27522 8616 27528 8628
rect 27479 8588 27528 8616
rect 27479 8585 27491 8588
rect 27433 8579 27491 8585
rect 27522 8576 27528 8588
rect 27580 8576 27586 8628
rect 29181 8619 29239 8625
rect 29181 8585 29193 8619
rect 29227 8616 29239 8619
rect 29454 8616 29460 8628
rect 29227 8588 29460 8616
rect 29227 8585 29239 8588
rect 29181 8579 29239 8585
rect 29454 8576 29460 8588
rect 29512 8576 29518 8628
rect 29730 8576 29736 8628
rect 29788 8616 29794 8628
rect 30285 8619 30343 8625
rect 30285 8616 30297 8619
rect 29788 8588 30297 8616
rect 29788 8576 29794 8588
rect 30285 8585 30297 8588
rect 30331 8585 30343 8619
rect 30285 8579 30343 8585
rect 30650 8576 30656 8628
rect 30708 8616 30714 8628
rect 31021 8619 31079 8625
rect 31021 8616 31033 8619
rect 30708 8588 31033 8616
rect 30708 8576 30714 8588
rect 31021 8585 31033 8588
rect 31067 8585 31079 8619
rect 31021 8579 31079 8585
rect 34882 8576 34888 8628
rect 34940 8616 34946 8628
rect 36722 8616 36728 8628
rect 34940 8588 36728 8616
rect 34940 8576 34946 8588
rect 36722 8576 36728 8588
rect 36780 8576 36786 8628
rect 39209 8619 39267 8625
rect 39209 8585 39221 8619
rect 39255 8616 39267 8619
rect 40034 8616 40040 8628
rect 39255 8588 40040 8616
rect 39255 8585 39267 8588
rect 39209 8579 39267 8585
rect 40034 8576 40040 8588
rect 40092 8576 40098 8628
rect 40402 8576 40408 8628
rect 40460 8616 40466 8628
rect 40681 8619 40739 8625
rect 40681 8616 40693 8619
rect 40460 8588 40693 8616
rect 40460 8576 40466 8588
rect 40681 8585 40693 8588
rect 40727 8616 40739 8619
rect 41138 8616 41144 8628
rect 40727 8588 41144 8616
rect 40727 8585 40739 8588
rect 40681 8579 40739 8585
rect 41138 8576 41144 8588
rect 41196 8576 41202 8628
rect 42610 8616 42616 8628
rect 41524 8588 42616 8616
rect 18570 8511 18628 8517
rect 18708 8520 21772 8548
rect 21836 8520 23428 8548
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 8941 8443 8999 8449
rect 9048 8452 9413 8480
rect 7331 8384 8340 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 8478 8372 8484 8424
rect 8536 8372 8542 8424
rect 8588 8412 8616 8440
rect 9048 8412 9076 8452
rect 9401 8449 9413 8452
rect 9447 8480 9459 8483
rect 9447 8452 11744 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 8588 8384 9076 8412
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8412 9183 8415
rect 9490 8412 9496 8424
rect 9171 8384 9496 8412
rect 9171 8381 9183 8384
rect 9125 8375 9183 8381
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 6288 8316 7481 8344
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 8496 8344 8524 8372
rect 7469 8307 7527 8313
rect 7576 8316 8524 8344
rect 7576 8276 7604 8316
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9140 8344 9168 8375
rect 9490 8372 9496 8384
rect 9548 8412 9554 8424
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9548 8384 9781 8412
rect 9548 8372 9554 8384
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 11716 8412 11744 8452
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11848 8452 11897 8480
rect 11848 8440 11854 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 18708 8480 18736 8520
rect 21836 8489 21864 8520
rect 20441 8483 20499 8489
rect 20441 8480 20453 8483
rect 11885 8443 11943 8449
rect 11992 8452 18736 8480
rect 19904 8452 20453 8480
rect 11992 8412 12020 8452
rect 19904 8424 19932 8452
rect 20441 8449 20453 8452
rect 20487 8480 20499 8483
rect 21361 8483 21419 8489
rect 21361 8480 21373 8483
rect 20487 8452 21373 8480
rect 20487 8449 20499 8452
rect 20441 8443 20499 8449
rect 21361 8449 21373 8452
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22088 8483 22146 8489
rect 22088 8449 22100 8483
rect 22134 8480 22146 8483
rect 23014 8480 23020 8492
rect 22134 8452 23020 8480
rect 22134 8449 22146 8452
rect 22088 8443 22146 8449
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 23293 8483 23351 8489
rect 23293 8449 23305 8483
rect 23339 8480 23351 8483
rect 23400 8480 23428 8520
rect 24210 8508 24216 8560
rect 24268 8508 24274 8560
rect 24302 8508 24308 8560
rect 24360 8548 24366 8560
rect 24360 8520 24900 8548
rect 24360 8508 24366 8520
rect 23339 8452 23428 8480
rect 23560 8483 23618 8489
rect 23339 8449 23351 8452
rect 23293 8443 23351 8449
rect 23560 8449 23572 8483
rect 23606 8480 23618 8483
rect 24670 8480 24676 8492
rect 23606 8452 24676 8480
rect 23606 8449 23618 8452
rect 23560 8443 23618 8449
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 24762 8440 24768 8492
rect 24820 8440 24826 8492
rect 24872 8480 24900 8520
rect 26602 8508 26608 8560
rect 26660 8548 26666 8560
rect 32392 8551 32450 8557
rect 26660 8520 27568 8548
rect 26660 8508 26666 8520
rect 24872 8452 25176 8480
rect 11716 8384 12020 8412
rect 12161 8415 12219 8421
rect 10781 8375 10839 8381
rect 12161 8381 12173 8415
rect 12207 8412 12219 8415
rect 12989 8415 13047 8421
rect 12207 8384 12388 8412
rect 12207 8381 12219 8384
rect 12161 8375 12219 8381
rect 8720 8316 9168 8344
rect 10796 8344 10824 8375
rect 12360 8356 12388 8384
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13078 8412 13084 8424
rect 13035 8384 13084 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13320 8384 15792 8412
rect 13320 8372 13326 8384
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 10796 8316 11529 8344
rect 8720 8304 8726 8316
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 12400 8316 12817 8344
rect 12400 8304 12406 8316
rect 12805 8313 12817 8316
rect 12851 8344 12863 8347
rect 15764 8344 15792 8384
rect 15838 8372 15844 8424
rect 15896 8372 15902 8424
rect 16758 8372 16764 8424
rect 16816 8372 16822 8424
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8412 17739 8415
rect 17954 8412 17960 8424
rect 17727 8384 17960 8412
rect 17727 8381 17739 8384
rect 17681 8375 17739 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 18322 8372 18328 8424
rect 18380 8372 18386 8424
rect 19794 8372 19800 8424
rect 19852 8372 19858 8424
rect 19886 8372 19892 8424
rect 19944 8372 19950 8424
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8412 20775 8415
rect 21266 8412 21272 8424
rect 20763 8384 21272 8412
rect 20763 8381 20775 8384
rect 20717 8375 20775 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21453 8415 21511 8421
rect 21453 8381 21465 8415
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 15930 8344 15936 8356
rect 12851 8316 13952 8344
rect 15764 8316 15936 8344
rect 12851 8313 12863 8316
rect 12805 8307 12863 8313
rect 6196 8248 7604 8276
rect 11330 8236 11336 8288
rect 11388 8236 11394 8288
rect 13924 8276 13952 8316
rect 15930 8304 15936 8316
rect 15988 8344 15994 8356
rect 16390 8344 16396 8356
rect 15988 8316 16396 8344
rect 15988 8304 15994 8316
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 19812 8344 19840 8372
rect 21468 8344 21496 8375
rect 24946 8372 24952 8424
rect 25004 8372 25010 8424
rect 25148 8356 25176 8452
rect 25774 8440 25780 8492
rect 25832 8489 25838 8492
rect 25832 8483 25860 8489
rect 25848 8449 25860 8483
rect 25832 8443 25860 8449
rect 25832 8440 25838 8443
rect 25958 8440 25964 8492
rect 26016 8440 26022 8492
rect 27341 8483 27399 8489
rect 27341 8449 27353 8483
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 25685 8415 25743 8421
rect 25685 8412 25697 8415
rect 25516 8384 25697 8412
rect 23201 8347 23259 8353
rect 23201 8344 23213 8347
rect 19812 8316 21496 8344
rect 22756 8316 23213 8344
rect 15470 8276 15476 8288
rect 13924 8248 15476 8276
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16485 8279 16543 8285
rect 16485 8276 16497 8279
rect 16080 8248 16497 8276
rect 16080 8236 16086 8248
rect 16485 8245 16497 8248
rect 16531 8245 16543 8279
rect 16485 8239 16543 8245
rect 17402 8236 17408 8288
rect 17460 8236 17466 8288
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 21542 8276 21548 8288
rect 20496 8248 21548 8276
rect 20496 8236 20502 8248
rect 21542 8236 21548 8248
rect 21600 8276 21606 8288
rect 22756 8276 22784 8316
rect 23201 8313 23213 8316
rect 23247 8313 23259 8347
rect 23201 8307 23259 8313
rect 24673 8347 24731 8353
rect 24673 8313 24685 8347
rect 24719 8344 24731 8347
rect 24762 8344 24768 8356
rect 24719 8316 24768 8344
rect 24719 8313 24731 8316
rect 24673 8307 24731 8313
rect 24762 8304 24768 8316
rect 24820 8344 24826 8356
rect 24820 8316 25084 8344
rect 24820 8304 24826 8316
rect 21600 8248 22784 8276
rect 25056 8276 25084 8316
rect 25130 8304 25136 8356
rect 25188 8344 25194 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 25188 8316 25421 8344
rect 25188 8304 25194 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 25409 8307 25467 8313
rect 25516 8276 25544 8384
rect 25685 8381 25697 8384
rect 25731 8381 25743 8415
rect 25685 8375 25743 8381
rect 26326 8372 26332 8424
rect 26384 8412 26390 8424
rect 27356 8412 27384 8443
rect 27540 8424 27568 8520
rect 32392 8517 32404 8551
rect 32438 8548 32450 8551
rect 33226 8548 33232 8560
rect 32438 8520 33232 8548
rect 32438 8517 32450 8520
rect 32392 8511 32450 8517
rect 33226 8508 33232 8520
rect 33284 8508 33290 8560
rect 34238 8508 34244 8560
rect 34296 8548 34302 8560
rect 39390 8548 39396 8560
rect 34296 8520 37596 8548
rect 34296 8508 34302 8520
rect 29086 8440 29092 8492
rect 29144 8440 29150 8492
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 29641 8483 29699 8489
rect 29641 8480 29653 8483
rect 29604 8452 29653 8480
rect 29604 8440 29610 8452
rect 29641 8449 29653 8452
rect 29687 8449 29699 8483
rect 29641 8443 29699 8449
rect 30300 8452 31754 8480
rect 30300 8424 30328 8452
rect 26384 8384 27384 8412
rect 26384 8372 26390 8384
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 27985 8415 28043 8421
rect 27985 8412 27997 8415
rect 27580 8384 27997 8412
rect 27580 8372 27586 8384
rect 27985 8381 27997 8384
rect 28031 8381 28043 8415
rect 27985 8375 28043 8381
rect 30282 8372 30288 8424
rect 30340 8372 30346 8424
rect 30374 8372 30380 8424
rect 30432 8372 30438 8424
rect 31726 8412 31754 8452
rect 33410 8440 33416 8492
rect 33468 8480 33474 8492
rect 35360 8489 35388 8520
rect 33597 8483 33655 8489
rect 33597 8480 33609 8483
rect 33468 8452 33609 8480
rect 33468 8440 33474 8452
rect 33597 8449 33609 8452
rect 33643 8480 33655 8483
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 33643 8452 34897 8480
rect 33643 8449 33655 8452
rect 33597 8443 33655 8449
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34885 8443 34943 8449
rect 35345 8483 35403 8489
rect 35345 8449 35357 8483
rect 35391 8449 35403 8483
rect 35345 8443 35403 8449
rect 35612 8483 35670 8489
rect 35612 8449 35624 8483
rect 35658 8480 35670 8483
rect 36538 8480 36544 8492
rect 35658 8452 36544 8480
rect 35658 8449 35670 8452
rect 35612 8443 35670 8449
rect 32122 8412 32128 8424
rect 31726 8384 32128 8412
rect 32122 8372 32128 8384
rect 32180 8372 32186 8424
rect 34422 8372 34428 8424
rect 34480 8372 34486 8424
rect 26602 8304 26608 8356
rect 26660 8304 26666 8356
rect 35360 8288 35388 8443
rect 36538 8440 36544 8452
rect 36596 8440 36602 8492
rect 37568 8489 37596 8520
rect 37844 8520 39396 8548
rect 37553 8483 37611 8489
rect 37553 8449 37565 8483
rect 37599 8480 37611 8483
rect 37734 8480 37740 8492
rect 37599 8452 37740 8480
rect 37599 8449 37611 8452
rect 37553 8443 37611 8449
rect 37734 8440 37740 8452
rect 37792 8480 37798 8492
rect 37844 8489 37872 8520
rect 37829 8483 37887 8489
rect 37829 8480 37841 8483
rect 37792 8452 37841 8480
rect 37792 8440 37798 8452
rect 37829 8449 37841 8452
rect 37875 8449 37887 8483
rect 37829 8443 37887 8449
rect 38096 8483 38154 8489
rect 38096 8449 38108 8483
rect 38142 8480 38154 8483
rect 38654 8480 38660 8492
rect 38142 8452 38660 8480
rect 38142 8449 38154 8452
rect 38096 8443 38154 8449
rect 38654 8440 38660 8452
rect 38712 8440 38718 8492
rect 39316 8489 39344 8520
rect 39390 8508 39396 8520
rect 39448 8548 39454 8560
rect 41414 8548 41420 8560
rect 39448 8520 41420 8548
rect 39448 8508 39454 8520
rect 39301 8483 39359 8489
rect 39301 8449 39313 8483
rect 39347 8449 39359 8483
rect 39301 8443 39359 8449
rect 39568 8483 39626 8489
rect 39568 8449 39580 8483
rect 39614 8480 39626 8483
rect 40126 8480 40132 8492
rect 39614 8452 40132 8480
rect 39614 8449 39626 8452
rect 39568 8443 39626 8449
rect 40126 8440 40132 8452
rect 40184 8440 40190 8492
rect 40880 8489 40908 8520
rect 41414 8508 41420 8520
rect 41472 8508 41478 8560
rect 40865 8483 40923 8489
rect 40865 8449 40877 8483
rect 40911 8449 40923 8483
rect 40865 8443 40923 8449
rect 41132 8483 41190 8489
rect 41132 8449 41144 8483
rect 41178 8480 41190 8483
rect 41524 8480 41552 8588
rect 42610 8576 42616 8588
rect 42668 8576 42674 8628
rect 43898 8576 43904 8628
rect 43956 8576 43962 8628
rect 44453 8619 44511 8625
rect 44453 8585 44465 8619
rect 44499 8616 44511 8619
rect 44818 8616 44824 8628
rect 44499 8588 44824 8616
rect 44499 8585 44511 8588
rect 44453 8579 44511 8585
rect 42150 8508 42156 8560
rect 42208 8548 42214 8560
rect 42972 8551 43030 8557
rect 42208 8520 42932 8548
rect 42208 8508 42214 8520
rect 41178 8452 41552 8480
rect 41178 8449 41190 8452
rect 41132 8443 41190 8449
rect 42518 8440 42524 8492
rect 42576 8440 42582 8492
rect 42904 8480 42932 8520
rect 42972 8517 42984 8551
rect 43018 8548 43030 8551
rect 43916 8548 43944 8576
rect 43018 8520 43944 8548
rect 43018 8517 43030 8520
rect 42972 8511 43030 8517
rect 44560 8489 44588 8588
rect 44818 8576 44824 8588
rect 44876 8576 44882 8628
rect 46474 8616 46480 8628
rect 45848 8588 46480 8616
rect 45848 8548 45876 8588
rect 46474 8576 46480 8588
rect 46532 8576 46538 8628
rect 46566 8576 46572 8628
rect 46624 8576 46630 8628
rect 47305 8619 47363 8625
rect 47305 8585 47317 8619
rect 47351 8616 47363 8619
rect 47394 8616 47400 8628
rect 47351 8588 47400 8616
rect 47351 8585 47363 8588
rect 47305 8579 47363 8585
rect 46584 8548 46612 8576
rect 44652 8520 45876 8548
rect 45940 8520 46612 8548
rect 44545 8483 44603 8489
rect 42904 8452 44496 8480
rect 42536 8412 42564 8440
rect 42705 8415 42763 8421
rect 42705 8412 42717 8415
rect 42536 8384 42717 8412
rect 42705 8381 42717 8384
rect 42751 8381 42763 8415
rect 44468 8412 44496 8452
rect 44545 8449 44557 8483
rect 44591 8449 44603 8483
rect 44545 8443 44603 8449
rect 44652 8412 44680 8520
rect 44812 8483 44870 8489
rect 44812 8449 44824 8483
rect 44858 8480 44870 8483
rect 45940 8480 45968 8520
rect 44858 8452 45968 8480
rect 46017 8483 46075 8489
rect 44858 8449 44870 8452
rect 44812 8443 44870 8449
rect 46017 8449 46029 8483
rect 46063 8480 46075 8483
rect 47320 8480 47348 8579
rect 47394 8576 47400 8588
rect 47452 8576 47458 8628
rect 47854 8616 47860 8628
rect 47504 8588 47860 8616
rect 46063 8452 47348 8480
rect 46063 8449 46075 8452
rect 46017 8443 46075 8449
rect 44468 8384 44680 8412
rect 46845 8415 46903 8421
rect 42705 8375 42763 8381
rect 46845 8381 46857 8415
rect 46891 8412 46903 8415
rect 47210 8412 47216 8424
rect 46891 8384 47216 8412
rect 46891 8381 46903 8384
rect 46845 8375 46903 8381
rect 47210 8372 47216 8384
rect 47268 8412 47274 8424
rect 47504 8412 47532 8588
rect 47854 8576 47860 8588
rect 47912 8576 47918 8628
rect 48961 8619 49019 8625
rect 48961 8585 48973 8619
rect 49007 8616 49019 8619
rect 49878 8616 49884 8628
rect 49007 8588 49884 8616
rect 49007 8585 49019 8588
rect 48961 8579 49019 8585
rect 49878 8576 49884 8588
rect 49936 8576 49942 8628
rect 50798 8576 50804 8628
rect 50856 8576 50862 8628
rect 52270 8576 52276 8628
rect 52328 8576 52334 8628
rect 53466 8576 53472 8628
rect 53524 8576 53530 8628
rect 53834 8576 53840 8628
rect 53892 8616 53898 8628
rect 53892 8588 55996 8616
rect 53892 8576 53898 8588
rect 49596 8551 49654 8557
rect 47596 8520 49372 8548
rect 47596 8492 47624 8520
rect 47578 8440 47584 8492
rect 47636 8440 47642 8492
rect 47848 8483 47906 8489
rect 47848 8449 47860 8483
rect 47894 8480 47906 8483
rect 48682 8480 48688 8492
rect 47894 8452 48688 8480
rect 47894 8449 47906 8452
rect 47848 8443 47906 8449
rect 48682 8440 48688 8452
rect 48740 8440 48746 8492
rect 49344 8489 49372 8520
rect 49596 8517 49608 8551
rect 49642 8548 49654 8551
rect 50816 8548 50844 8576
rect 49642 8520 50844 8548
rect 52288 8548 52316 8576
rect 54202 8548 54208 8560
rect 52288 8520 54208 8548
rect 49642 8517 49654 8520
rect 49596 8511 49654 8517
rect 54202 8508 54208 8520
rect 54260 8508 54266 8560
rect 55766 8508 55772 8560
rect 55824 8548 55830 8560
rect 55861 8551 55919 8557
rect 55861 8548 55873 8551
rect 55824 8520 55873 8548
rect 55824 8508 55830 8520
rect 55861 8517 55873 8520
rect 55907 8517 55919 8551
rect 55861 8511 55919 8517
rect 55968 8492 55996 8588
rect 56778 8576 56784 8628
rect 56836 8576 56842 8628
rect 56870 8576 56876 8628
rect 56928 8576 56934 8628
rect 57330 8576 57336 8628
rect 57388 8576 57394 8628
rect 57701 8619 57759 8625
rect 57701 8585 57713 8619
rect 57747 8616 57759 8619
rect 58066 8616 58072 8628
rect 57747 8588 58072 8616
rect 57747 8585 57759 8588
rect 57701 8579 57759 8585
rect 58066 8576 58072 8588
rect 58124 8576 58130 8628
rect 56220 8551 56278 8557
rect 56220 8517 56232 8551
rect 56266 8548 56278 8551
rect 56796 8548 56824 8576
rect 56266 8520 56824 8548
rect 56266 8517 56278 8520
rect 56220 8511 56278 8517
rect 49329 8483 49387 8489
rect 49329 8449 49341 8483
rect 49375 8449 49387 8483
rect 49329 8443 49387 8449
rect 49418 8440 49424 8492
rect 49476 8480 49482 8492
rect 51445 8483 51503 8489
rect 51445 8480 51457 8483
rect 49476 8452 51457 8480
rect 49476 8440 49482 8452
rect 51445 8449 51457 8452
rect 51491 8449 51503 8483
rect 51445 8443 51503 8449
rect 53377 8483 53435 8489
rect 53377 8449 53389 8483
rect 53423 8480 53435 8483
rect 54386 8480 54392 8492
rect 53423 8452 54392 8480
rect 53423 8449 53435 8452
rect 53377 8443 53435 8449
rect 54386 8440 54392 8452
rect 54444 8440 54450 8492
rect 55950 8440 55956 8492
rect 56008 8440 56014 8492
rect 56042 8440 56048 8492
rect 56100 8440 56106 8492
rect 56888 8480 56916 8576
rect 57885 8483 57943 8489
rect 57885 8480 57897 8483
rect 56888 8452 57897 8480
rect 57885 8449 57897 8452
rect 57931 8449 57943 8483
rect 57885 8443 57943 8449
rect 50801 8415 50859 8421
rect 50801 8412 50813 8415
rect 47268 8384 47532 8412
rect 47268 8372 47274 8384
rect 42245 8347 42303 8353
rect 42245 8313 42257 8347
rect 42291 8344 42303 8347
rect 42426 8344 42432 8356
rect 42291 8316 42432 8344
rect 42291 8313 42303 8316
rect 42245 8307 42303 8313
rect 25056 8248 25544 8276
rect 21600 8236 21606 8248
rect 33502 8236 33508 8288
rect 33560 8236 33566 8288
rect 35342 8236 35348 8288
rect 35400 8236 35406 8288
rect 36814 8236 36820 8288
rect 36872 8276 36878 8288
rect 37001 8279 37059 8285
rect 37001 8276 37013 8279
rect 36872 8248 37013 8276
rect 36872 8236 36878 8248
rect 37001 8245 37013 8248
rect 37047 8245 37059 8279
rect 37001 8239 37059 8245
rect 40770 8236 40776 8288
rect 40828 8276 40834 8288
rect 42260 8276 42288 8307
rect 42426 8304 42432 8316
rect 42484 8304 42490 8356
rect 44085 8347 44143 8353
rect 44085 8313 44097 8347
rect 44131 8344 44143 8347
rect 44174 8344 44180 8356
rect 44131 8316 44180 8344
rect 44131 8313 44143 8316
rect 44085 8307 44143 8313
rect 44174 8304 44180 8316
rect 44232 8344 44238 8356
rect 44542 8344 44548 8356
rect 44232 8316 44548 8344
rect 44232 8304 44238 8316
rect 44542 8304 44548 8316
rect 44600 8304 44606 8356
rect 45925 8347 45983 8353
rect 45925 8344 45937 8347
rect 45480 8316 45937 8344
rect 45480 8288 45508 8316
rect 45925 8313 45937 8316
rect 45971 8313 45983 8347
rect 45925 8307 45983 8313
rect 40828 8248 42288 8276
rect 40828 8236 40834 8248
rect 45462 8236 45468 8288
rect 45520 8236 45526 8288
rect 47504 8276 47532 8384
rect 50724 8384 50813 8412
rect 50724 8288 50752 8384
rect 50801 8381 50813 8384
rect 50847 8381 50859 8415
rect 50801 8375 50859 8381
rect 51350 8372 51356 8424
rect 51408 8412 51414 8424
rect 51537 8415 51595 8421
rect 51537 8412 51549 8415
rect 51408 8384 51549 8412
rect 51408 8372 51414 8384
rect 51537 8381 51549 8384
rect 51583 8381 51595 8415
rect 53561 8415 53619 8421
rect 53561 8412 53573 8415
rect 51537 8375 51595 8381
rect 52472 8384 53573 8412
rect 50246 8276 50252 8288
rect 47504 8248 50252 8276
rect 50246 8236 50252 8248
rect 50304 8276 50310 8288
rect 50614 8276 50620 8288
rect 50304 8248 50620 8276
rect 50304 8236 50310 8248
rect 50614 8236 50620 8248
rect 50672 8236 50678 8288
rect 50706 8236 50712 8288
rect 50764 8236 50770 8288
rect 52178 8236 52184 8288
rect 52236 8236 52242 8288
rect 52270 8236 52276 8288
rect 52328 8276 52334 8288
rect 52472 8285 52500 8384
rect 53561 8381 53573 8384
rect 53607 8412 53619 8415
rect 53926 8412 53932 8424
rect 53607 8384 53932 8412
rect 53607 8381 53619 8384
rect 53561 8375 53619 8381
rect 53926 8372 53932 8384
rect 53984 8372 53990 8424
rect 54021 8415 54079 8421
rect 54021 8381 54033 8415
rect 54067 8412 54079 8415
rect 54110 8412 54116 8424
rect 54067 8384 54116 8412
rect 54067 8381 54079 8384
rect 54021 8375 54079 8381
rect 54110 8372 54116 8384
rect 54168 8372 54174 8424
rect 54205 8415 54263 8421
rect 54205 8381 54217 8415
rect 54251 8381 54263 8415
rect 54205 8375 54263 8381
rect 54220 8344 54248 8375
rect 54570 8372 54576 8424
rect 54628 8412 54634 8424
rect 54941 8415 54999 8421
rect 54941 8412 54953 8415
rect 54628 8384 54953 8412
rect 54628 8372 54634 8384
rect 54941 8381 54953 8384
rect 54987 8381 54999 8415
rect 54941 8375 54999 8381
rect 55030 8372 55036 8424
rect 55088 8421 55094 8424
rect 55088 8415 55116 8421
rect 55104 8381 55116 8415
rect 55088 8375 55116 8381
rect 55217 8415 55275 8421
rect 55217 8381 55229 8415
rect 55263 8412 55275 8415
rect 55398 8412 55404 8424
rect 55263 8384 55404 8412
rect 55263 8381 55275 8384
rect 55217 8375 55275 8381
rect 55088 8372 55094 8375
rect 55398 8372 55404 8384
rect 55456 8412 55462 8424
rect 56060 8412 56088 8440
rect 55456 8384 56088 8412
rect 55456 8372 55462 8384
rect 54220 8316 54616 8344
rect 52457 8279 52515 8285
rect 52457 8276 52469 8279
rect 52328 8248 52469 8276
rect 52328 8236 52334 8248
rect 52457 8245 52469 8248
rect 52503 8245 52515 8279
rect 52457 8239 52515 8245
rect 53006 8236 53012 8288
rect 53064 8236 53070 8288
rect 54588 8276 54616 8316
rect 54662 8304 54668 8356
rect 54720 8304 54726 8356
rect 57514 8304 57520 8356
rect 57572 8344 57578 8356
rect 58529 8347 58587 8353
rect 58529 8344 58541 8347
rect 57572 8316 58541 8344
rect 57572 8304 57578 8316
rect 58529 8313 58541 8316
rect 58575 8313 58587 8347
rect 58529 8307 58587 8313
rect 56318 8276 56324 8288
rect 54588 8248 56324 8276
rect 56318 8236 56324 8248
rect 56376 8236 56382 8288
rect 1104 8186 58880 8208
rect 1104 8134 8172 8186
rect 8224 8134 8236 8186
rect 8288 8134 8300 8186
rect 8352 8134 8364 8186
rect 8416 8134 8428 8186
rect 8480 8134 22616 8186
rect 22668 8134 22680 8186
rect 22732 8134 22744 8186
rect 22796 8134 22808 8186
rect 22860 8134 22872 8186
rect 22924 8134 37060 8186
rect 37112 8134 37124 8186
rect 37176 8134 37188 8186
rect 37240 8134 37252 8186
rect 37304 8134 37316 8186
rect 37368 8134 51504 8186
rect 51556 8134 51568 8186
rect 51620 8134 51632 8186
rect 51684 8134 51696 8186
rect 51748 8134 51760 8186
rect 51812 8134 58880 8186
rect 1104 8112 58880 8134
rect 3145 8075 3203 8081
rect 3145 8041 3157 8075
rect 3191 8072 3203 8075
rect 3786 8072 3792 8084
rect 3191 8044 3792 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4341 8075 4399 8081
rect 4341 8072 4353 8075
rect 4120 8044 4353 8072
rect 4120 8032 4126 8044
rect 4341 8041 4353 8044
rect 4387 8072 4399 8075
rect 5902 8072 5908 8084
rect 4387 8044 5908 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6144 8044 7297 8072
rect 6144 8032 6150 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7984 8044 8217 8072
rect 7984 8032 7990 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 8662 8032 8668 8084
rect 8720 8032 8726 8084
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 10192 8044 10333 8072
rect 10192 8032 10198 8044
rect 10321 8041 10333 8044
rect 10367 8072 10379 8075
rect 10410 8072 10416 8084
rect 10367 8044 10416 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 12986 8032 12992 8084
rect 13044 8032 13050 8084
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 15528 8044 17632 8072
rect 15528 8032 15534 8044
rect 15565 8007 15623 8013
rect 15565 8004 15577 8007
rect 14936 7976 15577 8004
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 4982 7936 4988 7948
rect 2915 7908 4988 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 2976 7877 3004 7908
rect 4982 7896 4988 7908
rect 5040 7936 5046 7948
rect 14936 7945 14964 7976
rect 15565 7973 15577 7976
rect 15611 7973 15623 8007
rect 15565 7967 15623 7973
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 5040 7908 5580 7936
rect 5040 7896 5046 7908
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 5169 7871 5227 7877
rect 3108 7840 3153 7868
rect 3108 7828 3114 7840
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5184 7732 5212 7831
rect 5552 7800 5580 7908
rect 10980 7908 12357 7936
rect 10980 7880 11008 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7905 14979 7939
rect 14921 7899 14979 7905
rect 16022 7896 16028 7948
rect 16080 7896 16086 7948
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7936 16175 7939
rect 16224 7936 16252 8044
rect 16393 8007 16451 8013
rect 16393 7973 16405 8007
rect 16439 8004 16451 8007
rect 17604 8004 17632 8044
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 18012 8044 18337 8072
rect 18012 8032 18018 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 18325 8035 18383 8041
rect 20714 8032 20720 8084
rect 20772 8032 20778 8084
rect 24210 8032 24216 8084
rect 24268 8032 24274 8084
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 27525 8075 27583 8081
rect 27525 8072 27537 8075
rect 25004 8044 27537 8072
rect 25004 8032 25010 8044
rect 27525 8041 27537 8044
rect 27571 8041 27583 8075
rect 27525 8035 27583 8041
rect 29638 8032 29644 8084
rect 29696 8072 29702 8084
rect 29733 8075 29791 8081
rect 29733 8072 29745 8075
rect 29696 8044 29745 8072
rect 29696 8032 29702 8044
rect 29733 8041 29745 8044
rect 29779 8041 29791 8075
rect 29733 8035 29791 8041
rect 33502 8032 33508 8084
rect 33560 8072 33566 8084
rect 35710 8072 35716 8084
rect 33560 8044 35716 8072
rect 33560 8032 33566 8044
rect 35710 8032 35716 8044
rect 35768 8032 35774 8084
rect 39390 8032 39396 8084
rect 39448 8032 39454 8084
rect 40770 8072 40776 8084
rect 40052 8044 40776 8072
rect 18230 8004 18236 8016
rect 16439 7976 17540 8004
rect 17604 7976 18236 8004
rect 16439 7973 16451 7976
rect 16393 7967 16451 7973
rect 16163 7908 16252 7936
rect 17037 7939 17095 7945
rect 16163 7905 16175 7908
rect 16117 7899 16175 7905
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 17310 7936 17316 7948
rect 17083 7908 17316 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 17512 7945 17540 7976
rect 18230 7964 18236 7976
rect 18288 7964 18294 8016
rect 20732 8004 20760 8032
rect 18800 7976 19334 8004
rect 20732 7976 21036 8004
rect 18800 7945 18828 7976
rect 17497 7939 17555 7945
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 18785 7939 18843 7945
rect 18785 7905 18797 7939
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 18966 7896 18972 7948
rect 19024 7896 19030 7948
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 5905 7871 5963 7877
rect 5684 7840 5856 7868
rect 5684 7828 5690 7840
rect 5718 7800 5724 7812
rect 5552 7772 5724 7800
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 5828 7800 5856 7840
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6914 7868 6920 7880
rect 5951 7840 6920 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6914 7828 6920 7840
rect 6972 7868 6978 7880
rect 7374 7868 7380 7880
rect 6972 7840 7380 7868
rect 6972 7828 6978 7840
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9674 7868 9680 7880
rect 8987 7840 9680 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7868 12127 7871
rect 12250 7868 12256 7880
rect 12115 7840 12256 7868
rect 12115 7837 12127 7840
rect 12069 7831 12127 7837
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 13262 7828 13268 7880
rect 13320 7828 13326 7880
rect 14185 7871 14243 7877
rect 14185 7837 14197 7871
rect 14231 7868 14243 7871
rect 14458 7868 14464 7880
rect 14231 7840 14464 7868
rect 14231 7837 14243 7840
rect 14185 7831 14243 7837
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 16206 7868 16212 7880
rect 14884 7840 16212 7868
rect 14884 7828 14890 7840
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7868 16819 7871
rect 17402 7868 17408 7880
rect 16807 7840 17408 7868
rect 16807 7837 16819 7840
rect 16761 7831 16819 7837
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7868 18751 7871
rect 19058 7868 19064 7880
rect 18739 7840 19064 7868
rect 18739 7837 18751 7840
rect 18693 7831 18751 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19306 7868 19334 7976
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 19978 7936 19984 7948
rect 19935 7908 19984 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20257 7939 20315 7945
rect 20257 7905 20269 7939
rect 20303 7936 20315 7939
rect 20622 7936 20628 7948
rect 20303 7908 20628 7936
rect 20303 7905 20315 7908
rect 20257 7899 20315 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20864 7908 20913 7936
rect 20864 7896 20870 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 21008 7936 21036 7976
rect 24486 7964 24492 8016
rect 24544 8004 24550 8016
rect 24544 7976 26004 8004
rect 24544 7964 24550 7976
rect 21294 7939 21352 7945
rect 21294 7936 21306 7939
rect 21008 7908 21306 7936
rect 20901 7899 20959 7905
rect 21294 7905 21306 7908
rect 21340 7905 21352 7939
rect 21294 7899 21352 7905
rect 24578 7896 24584 7948
rect 24636 7936 24642 7948
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24636 7908 24961 7936
rect 24636 7896 24642 7908
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 25866 7896 25872 7948
rect 25924 7896 25930 7948
rect 25976 7936 26004 7976
rect 33778 7964 33784 8016
rect 33836 8004 33842 8016
rect 33836 7976 35480 8004
rect 33836 7964 33842 7976
rect 25976 7908 26280 7936
rect 26252 7880 26280 7908
rect 34882 7896 34888 7948
rect 34940 7896 34946 7948
rect 34974 7896 34980 7948
rect 35032 7936 35038 7948
rect 35345 7939 35403 7945
rect 35345 7936 35357 7939
rect 35032 7908 35357 7936
rect 35032 7896 35038 7908
rect 35345 7905 35357 7908
rect 35391 7905 35403 7939
rect 35452 7936 35480 7976
rect 35621 7939 35679 7945
rect 35621 7936 35633 7939
rect 35452 7908 35633 7936
rect 35345 7899 35403 7905
rect 35621 7905 35633 7908
rect 35667 7905 35679 7939
rect 35621 7899 35679 7905
rect 35710 7896 35716 7948
rect 35768 7945 35774 7948
rect 35768 7939 35796 7945
rect 35784 7905 35796 7939
rect 35768 7899 35796 7905
rect 35768 7896 35774 7899
rect 35894 7896 35900 7948
rect 35952 7936 35958 7948
rect 36262 7936 36268 7948
rect 35952 7908 36268 7936
rect 35952 7896 35958 7908
rect 36262 7896 36268 7908
rect 36320 7936 36326 7948
rect 36814 7936 36820 7948
rect 36320 7908 36820 7936
rect 36320 7896 36326 7908
rect 36814 7896 36820 7908
rect 36872 7896 36878 7948
rect 36906 7896 36912 7948
rect 36964 7936 36970 7948
rect 37185 7939 37243 7945
rect 37185 7936 37197 7939
rect 36964 7908 37197 7936
rect 36964 7896 36970 7908
rect 37185 7905 37197 7908
rect 37231 7905 37243 7939
rect 37185 7899 37243 7905
rect 37734 7896 37740 7948
rect 37792 7896 37798 7948
rect 40052 7945 40080 8044
rect 40770 8032 40776 8044
rect 40828 8032 40834 8084
rect 40954 8032 40960 8084
rect 41012 8072 41018 8084
rect 42150 8072 42156 8084
rect 41012 8044 42156 8072
rect 41012 8032 41018 8044
rect 42150 8032 42156 8044
rect 42208 8032 42214 8084
rect 43809 8075 43867 8081
rect 43809 8041 43821 8075
rect 43855 8072 43867 8075
rect 44082 8072 44088 8084
rect 43855 8044 44088 8072
rect 43855 8041 43867 8044
rect 43809 8035 43867 8041
rect 44082 8032 44088 8044
rect 44140 8072 44146 8084
rect 44140 8044 45784 8072
rect 44140 8032 44146 8044
rect 40126 7964 40132 8016
rect 40184 8004 40190 8016
rect 45462 8004 45468 8016
rect 40184 7976 40632 8004
rect 40184 7964 40190 7976
rect 40037 7939 40095 7945
rect 40037 7905 40049 7939
rect 40083 7905 40095 7939
rect 40402 7936 40408 7948
rect 40037 7899 40095 7905
rect 40236 7908 40408 7936
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19306 7840 19625 7868
rect 19613 7837 19625 7840
rect 19659 7868 19671 7871
rect 19659 7840 19932 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 19904 7812 19932 7840
rect 20438 7828 20444 7880
rect 20496 7828 20502 7880
rect 21174 7828 21180 7880
rect 21232 7828 21238 7880
rect 21450 7828 21456 7880
rect 21508 7828 21514 7880
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 22922 7868 22928 7880
rect 22879 7840 22928 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 22922 7828 22928 7840
rect 22980 7868 22986 7880
rect 26145 7871 26203 7877
rect 26145 7868 26157 7871
rect 22980 7840 26157 7868
rect 22980 7828 22986 7840
rect 26145 7837 26157 7840
rect 26191 7837 26203 7871
rect 26145 7831 26203 7837
rect 26234 7828 26240 7880
rect 26292 7828 26298 7880
rect 28626 7828 28632 7880
rect 28684 7828 28690 7880
rect 29730 7828 29736 7880
rect 29788 7868 29794 7880
rect 30837 7871 30895 7877
rect 30837 7868 30849 7871
rect 29788 7840 30849 7868
rect 29788 7828 29794 7840
rect 30837 7837 30849 7840
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 31849 7871 31907 7877
rect 31849 7837 31861 7871
rect 31895 7868 31907 7871
rect 32122 7868 32128 7880
rect 31895 7840 32128 7868
rect 31895 7837 31907 7840
rect 31849 7831 31907 7837
rect 32122 7828 32128 7840
rect 32180 7868 32186 7880
rect 32217 7871 32275 7877
rect 32217 7868 32229 7871
rect 32180 7840 32229 7868
rect 32180 7828 32186 7840
rect 32217 7837 32229 7840
rect 32263 7868 32275 7871
rect 32401 7871 32459 7877
rect 32401 7868 32413 7871
rect 32263 7840 32413 7868
rect 32263 7837 32275 7840
rect 32217 7831 32275 7837
rect 32401 7837 32413 7840
rect 32447 7868 32459 7871
rect 33042 7868 33048 7880
rect 32447 7840 33048 7868
rect 32447 7837 32459 7840
rect 32401 7831 32459 7837
rect 33042 7828 33048 7840
rect 33100 7828 33106 7880
rect 33870 7828 33876 7880
rect 33928 7828 33934 7880
rect 34698 7828 34704 7880
rect 34756 7828 34762 7880
rect 39853 7871 39911 7877
rect 39853 7837 39865 7871
rect 39899 7868 39911 7871
rect 40236 7868 40264 7908
rect 40402 7896 40408 7908
rect 40460 7896 40466 7948
rect 40494 7896 40500 7948
rect 40552 7896 40558 7948
rect 40604 7936 40632 7976
rect 44560 7976 44956 8004
rect 40773 7939 40831 7945
rect 40773 7936 40785 7939
rect 40604 7908 40785 7936
rect 40773 7905 40785 7908
rect 40819 7905 40831 7939
rect 40773 7899 40831 7905
rect 41414 7896 41420 7948
rect 41472 7936 41478 7948
rect 44560 7945 44588 7976
rect 44928 7948 44956 7976
rect 45020 7976 45468 8004
rect 42245 7939 42303 7945
rect 42245 7936 42257 7939
rect 41472 7908 42257 7936
rect 41472 7896 41478 7908
rect 42245 7905 42257 7908
rect 42291 7936 42303 7939
rect 42429 7939 42487 7945
rect 42429 7936 42441 7939
rect 42291 7908 42441 7936
rect 42291 7905 42303 7908
rect 42245 7899 42303 7905
rect 42429 7905 42441 7908
rect 42475 7905 42487 7939
rect 42429 7899 42487 7905
rect 44545 7939 44603 7945
rect 44545 7905 44557 7939
rect 44591 7905 44603 7939
rect 44545 7899 44603 7905
rect 44726 7896 44732 7948
rect 44784 7896 44790 7948
rect 44910 7896 44916 7948
rect 44968 7896 44974 7948
rect 45020 7945 45048 7976
rect 45462 7964 45468 7976
rect 45520 7964 45526 8016
rect 45646 7964 45652 8016
rect 45704 7964 45710 8016
rect 45005 7939 45063 7945
rect 45005 7905 45017 7939
rect 45051 7905 45063 7939
rect 45005 7899 45063 7905
rect 45189 7939 45247 7945
rect 45189 7905 45201 7939
rect 45235 7936 45247 7939
rect 45554 7936 45560 7948
rect 45235 7908 45560 7936
rect 45235 7905 45247 7908
rect 45189 7899 45247 7905
rect 45554 7896 45560 7908
rect 45612 7896 45618 7948
rect 45756 7936 45784 8044
rect 47210 8032 47216 8084
rect 47268 8032 47274 8084
rect 48774 8032 48780 8084
rect 48832 8072 48838 8084
rect 48869 8075 48927 8081
rect 48869 8072 48881 8075
rect 48832 8044 48881 8072
rect 48832 8032 48838 8044
rect 48869 8041 48881 8044
rect 48915 8041 48927 8075
rect 48869 8035 48927 8041
rect 49237 8075 49295 8081
rect 49237 8041 49249 8075
rect 49283 8072 49295 8075
rect 50154 8072 50160 8084
rect 49283 8044 50160 8072
rect 49283 8041 49295 8044
rect 49237 8035 49295 8041
rect 50154 8032 50160 8044
rect 50212 8032 50218 8084
rect 51350 8032 51356 8084
rect 51408 8072 51414 8084
rect 51537 8075 51595 8081
rect 51537 8072 51549 8075
rect 51408 8044 51549 8072
rect 51408 8032 51414 8044
rect 51537 8041 51549 8044
rect 51583 8041 51595 8075
rect 51537 8035 51595 8041
rect 53837 8075 53895 8081
rect 53837 8041 53849 8075
rect 53883 8072 53895 8075
rect 54478 8072 54484 8084
rect 53883 8044 54484 8072
rect 53883 8041 53895 8044
rect 53837 8035 53895 8041
rect 54478 8032 54484 8044
rect 54536 8072 54542 8084
rect 55030 8072 55036 8084
rect 54536 8044 55036 8072
rect 54536 8032 54542 8044
rect 55030 8032 55036 8044
rect 55088 8032 55094 8084
rect 55398 8032 55404 8084
rect 55456 8072 55462 8084
rect 55493 8075 55551 8081
rect 55493 8072 55505 8075
rect 55456 8044 55505 8072
rect 55456 8032 55462 8044
rect 55493 8041 55505 8044
rect 55539 8041 55551 8075
rect 55493 8035 55551 8041
rect 55953 8075 56011 8081
rect 55953 8041 55965 8075
rect 55999 8072 56011 8075
rect 56042 8072 56048 8084
rect 55999 8044 56048 8072
rect 55999 8041 56011 8044
rect 55953 8035 56011 8041
rect 56042 8032 56048 8044
rect 56100 8072 56106 8084
rect 56226 8072 56232 8084
rect 56100 8044 56232 8072
rect 56100 8032 56106 8044
rect 56226 8032 56232 8044
rect 56284 8032 56290 8084
rect 56318 8032 56324 8084
rect 56376 8072 56382 8084
rect 56376 8044 57376 8072
rect 56376 8032 56382 8044
rect 46042 7939 46100 7945
rect 46042 7936 46054 7939
rect 45756 7908 46054 7936
rect 46042 7905 46054 7908
rect 46088 7905 46100 7939
rect 46042 7899 46100 7905
rect 46201 7939 46259 7945
rect 46201 7905 46213 7939
rect 46247 7936 46259 7939
rect 46382 7936 46388 7948
rect 46247 7908 46388 7936
rect 46247 7905 46259 7908
rect 46201 7899 46259 7905
rect 46382 7896 46388 7908
rect 46440 7936 46446 7948
rect 47228 7936 47256 8032
rect 49142 7964 49148 8016
rect 49200 8004 49206 8016
rect 49602 8004 49608 8016
rect 49200 7976 49608 8004
rect 49200 7964 49206 7976
rect 49602 7964 49608 7976
rect 49660 8004 49666 8016
rect 55582 8004 55588 8016
rect 49660 7976 49832 8004
rect 49660 7964 49666 7976
rect 46440 7908 47256 7936
rect 46440 7896 46446 7908
rect 49418 7896 49424 7948
rect 49476 7936 49482 7948
rect 49804 7945 49832 7976
rect 54312 7976 55588 8004
rect 49697 7939 49755 7945
rect 49697 7936 49709 7939
rect 49476 7908 49709 7936
rect 49476 7896 49482 7908
rect 49697 7905 49709 7908
rect 49743 7905 49755 7939
rect 49697 7899 49755 7905
rect 49789 7939 49847 7945
rect 49789 7905 49801 7939
rect 49835 7905 49847 7939
rect 49789 7899 49847 7905
rect 39899 7840 40264 7868
rect 39899 7837 39911 7840
rect 39853 7831 39911 7837
rect 40862 7828 40868 7880
rect 40920 7877 40926 7880
rect 40920 7871 40948 7877
rect 40936 7837 40948 7871
rect 40920 7831 40948 7837
rect 40920 7828 40926 7831
rect 41046 7828 41052 7880
rect 41104 7828 41110 7880
rect 44361 7871 44419 7877
rect 44361 7837 44373 7871
rect 44407 7868 44419 7871
rect 44744 7868 44772 7896
rect 44407 7840 44772 7868
rect 44407 7837 44419 7840
rect 44361 7831 44419 7837
rect 45922 7828 45928 7880
rect 45980 7828 45986 7880
rect 47489 7871 47547 7877
rect 47489 7837 47501 7871
rect 47535 7868 47547 7871
rect 47578 7868 47584 7880
rect 47535 7840 47584 7868
rect 47535 7837 47547 7840
rect 47489 7831 47547 7837
rect 47578 7828 47584 7840
rect 47636 7868 47642 7880
rect 50157 7871 50215 7877
rect 50157 7868 50169 7871
rect 47636 7840 50169 7868
rect 47636 7828 47642 7840
rect 50157 7837 50169 7840
rect 50203 7837 50215 7871
rect 50157 7831 50215 7837
rect 50798 7828 50804 7880
rect 50856 7868 50862 7880
rect 51629 7871 51687 7877
rect 51629 7868 51641 7871
rect 50856 7840 51641 7868
rect 50856 7828 50862 7840
rect 51629 7837 51641 7840
rect 51675 7837 51687 7871
rect 51629 7831 51687 7837
rect 52457 7871 52515 7877
rect 52457 7837 52469 7871
rect 52503 7868 52515 7871
rect 52546 7868 52552 7880
rect 52503 7840 52552 7868
rect 52503 7837 52515 7840
rect 52457 7831 52515 7837
rect 52546 7828 52552 7840
rect 52604 7828 52610 7880
rect 53466 7828 53472 7880
rect 53524 7868 53530 7880
rect 54312 7877 54340 7976
rect 55582 7964 55588 7976
rect 55640 7964 55646 8016
rect 57348 8004 57376 8044
rect 57606 8032 57612 8084
rect 57664 8072 57670 8084
rect 58529 8075 58587 8081
rect 58529 8072 58541 8075
rect 57664 8044 58541 8072
rect 57664 8032 57670 8044
rect 58529 8041 58541 8044
rect 58575 8041 58587 8075
rect 58529 8035 58587 8041
rect 57793 8007 57851 8013
rect 57793 8004 57805 8007
rect 57348 7976 57805 8004
rect 57793 7973 57805 7976
rect 57839 7973 57851 8007
rect 57793 7967 57851 7973
rect 54570 7896 54576 7948
rect 54628 7936 54634 7948
rect 55306 7936 55312 7948
rect 54628 7908 55312 7936
rect 54628 7896 54634 7908
rect 55306 7896 55312 7908
rect 55364 7896 55370 7948
rect 55950 7896 55956 7948
rect 56008 7936 56014 7948
rect 56410 7936 56416 7948
rect 56008 7908 56416 7936
rect 56008 7896 56014 7908
rect 56410 7896 56416 7908
rect 56468 7896 56474 7948
rect 57808 7936 57836 7967
rect 57885 7939 57943 7945
rect 57885 7936 57897 7939
rect 57808 7908 57897 7936
rect 57885 7905 57897 7908
rect 57931 7905 57943 7939
rect 57885 7899 57943 7905
rect 54297 7871 54355 7877
rect 54297 7868 54309 7871
rect 53524 7840 54309 7868
rect 53524 7828 53530 7840
rect 54297 7837 54309 7840
rect 54343 7837 54355 7871
rect 54297 7831 54355 7837
rect 54389 7871 54447 7877
rect 54389 7837 54401 7871
rect 54435 7868 54447 7871
rect 55214 7868 55220 7880
rect 54435 7840 55220 7868
rect 54435 7837 54447 7840
rect 54389 7831 54447 7837
rect 55214 7828 55220 7840
rect 55272 7828 55278 7880
rect 56680 7871 56738 7877
rect 56680 7837 56692 7871
rect 56726 7868 56738 7871
rect 57514 7868 57520 7880
rect 56726 7840 57520 7868
rect 56726 7837 56738 7840
rect 56680 7831 56738 7837
rect 57514 7828 57520 7840
rect 57572 7828 57578 7880
rect 6150 7803 6208 7809
rect 6150 7800 6162 7803
rect 5828 7772 6162 7800
rect 6150 7769 6162 7772
rect 6196 7769 6208 7803
rect 6150 7763 6208 7769
rect 9208 7803 9266 7809
rect 9208 7769 9220 7803
rect 9254 7800 9266 7803
rect 9582 7800 9588 7812
rect 9254 7772 9588 7800
rect 9254 7769 9266 7772
rect 9208 7763 9266 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 11514 7800 11520 7812
rect 10704 7772 11520 7800
rect 10704 7744 10732 7772
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 12406 7772 19840 7800
rect 5994 7732 6000 7744
rect 5184 7704 6000 7732
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11238 7732 11244 7744
rect 11195 7704 11244 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 11238 7692 11244 7704
rect 11296 7732 11302 7744
rect 12406 7732 12434 7772
rect 11296 7704 12434 7732
rect 11296 7692 11302 7704
rect 13906 7692 13912 7744
rect 13964 7692 13970 7744
rect 14734 7692 14740 7744
rect 14792 7692 14798 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 15344 7704 15485 7732
rect 15344 7692 15350 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15473 7695 15531 7701
rect 15933 7735 15991 7741
rect 15933 7701 15945 7735
rect 15979 7732 15991 7735
rect 16853 7735 16911 7741
rect 16853 7732 16865 7735
rect 15979 7704 16865 7732
rect 15979 7701 15991 7704
rect 15933 7695 15991 7701
rect 16853 7701 16865 7704
rect 16899 7732 16911 7735
rect 17034 7732 17040 7744
rect 16899 7704 17040 7732
rect 16899 7701 16911 7704
rect 16853 7695 16911 7701
rect 17034 7692 17040 7704
rect 17092 7692 17098 7744
rect 18138 7692 18144 7744
rect 18196 7692 18202 7744
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 19702 7692 19708 7744
rect 19760 7692 19766 7744
rect 19812 7732 19840 7772
rect 19886 7760 19892 7812
rect 19944 7760 19950 7812
rect 23100 7803 23158 7809
rect 21928 7772 23060 7800
rect 21928 7732 21956 7772
rect 19812 7704 21956 7732
rect 22097 7735 22155 7741
rect 22097 7701 22109 7735
rect 22143 7732 22155 7735
rect 22278 7732 22284 7744
rect 22143 7704 22284 7732
rect 22143 7701 22155 7704
rect 22097 7695 22155 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 23032 7732 23060 7772
rect 23100 7769 23112 7803
rect 23146 7800 23158 7803
rect 23934 7800 23940 7812
rect 23146 7772 23940 7800
rect 23146 7769 23158 7772
rect 23100 7763 23158 7769
rect 23934 7760 23940 7772
rect 23992 7760 23998 7812
rect 26412 7803 26470 7809
rect 24044 7772 26372 7800
rect 24044 7732 24072 7772
rect 23032 7704 24072 7732
rect 24394 7692 24400 7744
rect 24452 7692 24458 7744
rect 24486 7692 24492 7744
rect 24544 7732 24550 7744
rect 24765 7735 24823 7741
rect 24765 7732 24777 7735
rect 24544 7704 24777 7732
rect 24544 7692 24550 7704
rect 24765 7701 24777 7704
rect 24811 7701 24823 7735
rect 24765 7695 24823 7701
rect 24854 7692 24860 7744
rect 24912 7692 24918 7744
rect 25317 7735 25375 7741
rect 25317 7701 25329 7735
rect 25363 7732 25375 7735
rect 25590 7732 25596 7744
rect 25363 7704 25596 7732
rect 25363 7701 25375 7704
rect 25317 7695 25375 7701
rect 25590 7692 25596 7704
rect 25648 7692 25654 7744
rect 25682 7692 25688 7744
rect 25740 7692 25746 7744
rect 25777 7735 25835 7741
rect 25777 7701 25789 7735
rect 25823 7732 25835 7735
rect 26234 7732 26240 7744
rect 25823 7704 26240 7732
rect 25823 7701 25835 7704
rect 25777 7695 25835 7701
rect 26234 7692 26240 7704
rect 26292 7692 26298 7744
rect 26344 7732 26372 7772
rect 26412 7769 26424 7803
rect 26458 7800 26470 7803
rect 27614 7800 27620 7812
rect 26458 7772 27620 7800
rect 26458 7769 26470 7772
rect 26412 7763 26470 7769
rect 27614 7760 27620 7772
rect 27672 7760 27678 7812
rect 28994 7760 29000 7812
rect 29052 7800 29058 7812
rect 29641 7803 29699 7809
rect 29641 7800 29653 7803
rect 29052 7772 29653 7800
rect 29052 7760 29058 7772
rect 29641 7769 29653 7772
rect 29687 7769 29699 7803
rect 29641 7763 29699 7769
rect 32668 7803 32726 7809
rect 32668 7769 32680 7803
rect 32714 7800 32726 7803
rect 34517 7803 34575 7809
rect 34517 7800 34529 7803
rect 32714 7772 34529 7800
rect 32714 7769 32726 7772
rect 32668 7763 32726 7769
rect 34517 7769 34529 7772
rect 34563 7769 34575 7803
rect 37001 7803 37059 7809
rect 37001 7800 37013 7803
rect 34517 7763 34575 7769
rect 36464 7772 37013 7800
rect 36464 7744 36492 7772
rect 37001 7769 37013 7772
rect 37047 7769 37059 7803
rect 37001 7763 37059 7769
rect 38004 7803 38062 7809
rect 38004 7769 38016 7803
rect 38050 7800 38062 7803
rect 38930 7800 38936 7812
rect 38050 7772 38936 7800
rect 38050 7769 38062 7772
rect 38004 7763 38062 7769
rect 38930 7760 38936 7772
rect 38988 7760 38994 7812
rect 42696 7803 42754 7809
rect 42696 7769 42708 7803
rect 42742 7800 42754 7803
rect 43990 7800 43996 7812
rect 42742 7772 43996 7800
rect 42742 7769 42754 7772
rect 42696 7763 42754 7769
rect 43990 7760 43996 7772
rect 44048 7760 44054 7812
rect 47756 7803 47814 7809
rect 47756 7769 47768 7803
rect 47802 7800 47814 7803
rect 48130 7800 48136 7812
rect 47802 7772 48136 7800
rect 47802 7769 47814 7772
rect 47756 7763 47814 7769
rect 48130 7760 48136 7772
rect 48188 7760 48194 7812
rect 49050 7760 49056 7812
rect 49108 7800 49114 7812
rect 50424 7803 50482 7809
rect 49108 7772 50108 7800
rect 49108 7760 49114 7772
rect 26878 7732 26884 7744
rect 26344 7704 26884 7732
rect 26878 7692 26884 7704
rect 26936 7692 26942 7744
rect 29178 7692 29184 7744
rect 29236 7692 29242 7744
rect 29362 7692 29368 7744
rect 29420 7732 29426 7744
rect 30193 7735 30251 7741
rect 30193 7732 30205 7735
rect 29420 7704 30205 7732
rect 29420 7692 29426 7704
rect 30193 7701 30205 7704
rect 30239 7732 30251 7735
rect 30926 7732 30932 7744
rect 30239 7704 30932 7732
rect 30239 7701 30251 7704
rect 30193 7695 30251 7701
rect 30926 7692 30932 7704
rect 30984 7692 30990 7744
rect 31294 7692 31300 7744
rect 31352 7732 31358 7744
rect 31481 7735 31539 7741
rect 31481 7732 31493 7735
rect 31352 7704 31493 7732
rect 31352 7692 31358 7704
rect 31481 7701 31493 7704
rect 31527 7701 31539 7735
rect 31481 7695 31539 7701
rect 33318 7692 33324 7744
rect 33376 7732 33382 7744
rect 36446 7732 36452 7744
rect 33376 7704 36452 7732
rect 33376 7692 33382 7704
rect 36446 7692 36452 7704
rect 36504 7692 36510 7744
rect 36538 7692 36544 7744
rect 36596 7692 36602 7744
rect 36630 7692 36636 7744
rect 36688 7692 36694 7744
rect 37090 7692 37096 7744
rect 37148 7692 37154 7744
rect 39114 7692 39120 7744
rect 39172 7732 39178 7744
rect 40862 7732 40868 7744
rect 39172 7704 40868 7732
rect 39172 7692 39178 7704
rect 40862 7692 40868 7704
rect 40920 7692 40926 7744
rect 41690 7692 41696 7744
rect 41748 7692 41754 7744
rect 43898 7692 43904 7744
rect 43956 7692 43962 7744
rect 44174 7692 44180 7744
rect 44232 7732 44238 7744
rect 44269 7735 44327 7741
rect 44269 7732 44281 7735
rect 44232 7704 44281 7732
rect 44232 7692 44238 7704
rect 44269 7701 44281 7704
rect 44315 7701 44327 7735
rect 44269 7695 44327 7701
rect 44542 7692 44548 7744
rect 44600 7732 44606 7744
rect 45922 7732 45928 7744
rect 44600 7704 45928 7732
rect 44600 7692 44606 7704
rect 45922 7692 45928 7704
rect 45980 7692 45986 7744
rect 46842 7692 46848 7744
rect 46900 7692 46906 7744
rect 48406 7692 48412 7744
rect 48464 7732 48470 7744
rect 49605 7735 49663 7741
rect 49605 7732 49617 7735
rect 48464 7704 49617 7732
rect 48464 7692 48470 7704
rect 49605 7701 49617 7704
rect 49651 7732 49663 7735
rect 49970 7732 49976 7744
rect 49651 7704 49976 7732
rect 49651 7701 49663 7704
rect 49605 7695 49663 7701
rect 49970 7692 49976 7704
rect 50028 7692 50034 7744
rect 50080 7732 50108 7772
rect 50424 7769 50436 7803
rect 50470 7800 50482 7803
rect 52273 7803 52331 7809
rect 52273 7800 52285 7803
rect 50470 7772 52285 7800
rect 50470 7769 50482 7772
rect 50424 7763 50482 7769
rect 52273 7769 52285 7772
rect 52319 7769 52331 7803
rect 52273 7763 52331 7769
rect 52724 7803 52782 7809
rect 52724 7769 52736 7803
rect 52770 7800 52782 7803
rect 53558 7800 53564 7812
rect 52770 7772 53564 7800
rect 52770 7769 52782 7772
rect 52724 7763 52782 7769
rect 53558 7760 53564 7772
rect 53616 7760 53622 7812
rect 51350 7732 51356 7744
rect 50080 7704 51356 7732
rect 51350 7692 51356 7704
rect 51408 7692 51414 7744
rect 51442 7692 51448 7744
rect 51500 7732 51506 7744
rect 53374 7732 53380 7744
rect 51500 7704 53380 7732
rect 51500 7692 51506 7704
rect 53374 7692 53380 7704
rect 53432 7692 53438 7744
rect 53926 7692 53932 7744
rect 53984 7692 53990 7744
rect 54662 7692 54668 7744
rect 54720 7732 54726 7744
rect 54938 7732 54944 7744
rect 54720 7704 54944 7732
rect 54720 7692 54726 7704
rect 54938 7692 54944 7704
rect 54996 7692 55002 7744
rect 55582 7692 55588 7744
rect 55640 7732 55646 7744
rect 56229 7735 56287 7741
rect 56229 7732 56241 7735
rect 55640 7704 56241 7732
rect 55640 7692 55646 7704
rect 56229 7701 56241 7704
rect 56275 7701 56287 7735
rect 56229 7695 56287 7701
rect 1104 7642 59040 7664
rect 1104 7590 15394 7642
rect 15446 7590 15458 7642
rect 15510 7590 15522 7642
rect 15574 7590 15586 7642
rect 15638 7590 15650 7642
rect 15702 7590 29838 7642
rect 29890 7590 29902 7642
rect 29954 7590 29966 7642
rect 30018 7590 30030 7642
rect 30082 7590 30094 7642
rect 30146 7590 44282 7642
rect 44334 7590 44346 7642
rect 44398 7590 44410 7642
rect 44462 7590 44474 7642
rect 44526 7590 44538 7642
rect 44590 7590 58726 7642
rect 58778 7590 58790 7642
rect 58842 7590 58854 7642
rect 58906 7590 58918 7642
rect 58970 7590 58982 7642
rect 59034 7590 59040 7642
rect 1104 7568 59040 7590
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 4062 7528 4068 7540
rect 3835 7500 4068 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 5994 7528 6000 7540
rect 5859 7500 6000 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6236 7500 13308 7528
rect 6236 7488 6242 7500
rect 6917 7463 6975 7469
rect 6917 7429 6929 7463
rect 6963 7460 6975 7463
rect 7006 7460 7012 7472
rect 6963 7432 7012 7460
rect 6963 7429 6975 7432
rect 6917 7423 6975 7429
rect 7006 7420 7012 7432
rect 7064 7420 7070 7472
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 7193 7463 7251 7469
rect 7193 7460 7205 7463
rect 7156 7432 7205 7460
rect 7156 7420 7162 7432
rect 7193 7429 7205 7432
rect 7239 7460 7251 7463
rect 8754 7460 8760 7472
rect 7239 7432 8760 7460
rect 7239 7429 7251 7432
rect 7193 7423 7251 7429
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 9968 7432 12434 7460
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 9306 7392 9312 7404
rect 7423 7364 9312 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 2590 7284 2596 7336
rect 2648 7284 2654 7336
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 7834 7324 7840 7336
rect 5776 7296 7840 7324
rect 5776 7284 5782 7296
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 9490 7324 9496 7336
rect 9263 7296 9496 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9968 7333 9996 7432
rect 10220 7395 10278 7401
rect 10220 7361 10232 7395
rect 10266 7392 10278 7395
rect 11330 7392 11336 7404
rect 10266 7364 11336 7392
rect 10266 7361 10278 7364
rect 10220 7355 10278 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 12406 7392 12434 7432
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12406 7364 13093 7392
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13280 7392 13308 7500
rect 13906 7488 13912 7540
rect 13964 7488 13970 7540
rect 14016 7500 18552 7528
rect 13348 7463 13406 7469
rect 13348 7429 13360 7463
rect 13394 7460 13406 7463
rect 13924 7460 13952 7488
rect 13394 7432 13952 7460
rect 13394 7429 13406 7432
rect 13348 7423 13406 7429
rect 14016 7392 14044 7500
rect 14826 7420 14832 7472
rect 14884 7420 14890 7472
rect 18322 7460 18328 7472
rect 15028 7432 18328 7460
rect 13280 7364 14044 7392
rect 13081 7355 13139 7361
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 9674 7256 9680 7268
rect 8680 7228 9680 7256
rect 3234 7148 3240 7200
rect 3292 7148 3298 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 8680 7197 8708 7228
rect 9674 7216 9680 7228
rect 9732 7256 9738 7268
rect 9968 7256 9996 7287
rect 9732 7228 9996 7256
rect 9732 7216 9738 7228
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 7432 7160 8677 7188
rect 7432 7148 7438 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 8665 7151 8723 7157
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10962 7188 10968 7200
rect 10008 7160 10968 7188
rect 10008 7148 10014 7160
rect 10962 7148 10968 7160
rect 11020 7188 11026 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11020 7160 11345 7188
rect 11020 7148 11026 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11532 7188 11560 7352
rect 12158 7284 12164 7336
rect 12216 7284 12222 7336
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15028 7333 15056 7432
rect 15286 7401 15292 7404
rect 15280 7392 15292 7401
rect 15247 7364 15292 7392
rect 15280 7355 15292 7364
rect 15286 7352 15292 7355
rect 15344 7352 15350 7404
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15838 7392 15844 7404
rect 15620 7364 15844 7392
rect 15620 7352 15626 7364
rect 15838 7352 15844 7364
rect 15896 7392 15902 7404
rect 16684 7401 16712 7432
rect 18322 7420 18328 7432
rect 18380 7460 18386 7472
rect 18524 7460 18552 7500
rect 19702 7488 19708 7540
rect 19760 7528 19766 7540
rect 20533 7531 20591 7537
rect 20533 7528 20545 7531
rect 19760 7500 20545 7528
rect 19760 7488 19766 7500
rect 20533 7497 20545 7500
rect 20579 7497 20591 7531
rect 20533 7491 20591 7497
rect 23934 7488 23940 7540
rect 23992 7488 23998 7540
rect 24394 7488 24400 7540
rect 24452 7488 24458 7540
rect 24670 7488 24676 7540
rect 24728 7488 24734 7540
rect 24854 7488 24860 7540
rect 24912 7528 24918 7540
rect 25409 7531 25467 7537
rect 25409 7528 25421 7531
rect 24912 7500 25421 7528
rect 24912 7488 24918 7500
rect 25409 7497 25421 7500
rect 25455 7497 25467 7531
rect 25409 7491 25467 7497
rect 25590 7488 25596 7540
rect 25648 7488 25654 7540
rect 25682 7488 25688 7540
rect 25740 7528 25746 7540
rect 26605 7531 26663 7537
rect 26605 7528 26617 7531
rect 25740 7500 26617 7528
rect 25740 7488 25746 7500
rect 26605 7497 26617 7500
rect 26651 7497 26663 7531
rect 26605 7491 26663 7497
rect 27614 7488 27620 7540
rect 27672 7488 27678 7540
rect 28626 7488 28632 7540
rect 28684 7528 28690 7540
rect 28721 7531 28779 7537
rect 28721 7528 28733 7531
rect 28684 7500 28733 7528
rect 28684 7488 28690 7500
rect 28721 7497 28733 7500
rect 28767 7497 28779 7531
rect 28721 7491 28779 7497
rect 29089 7531 29147 7537
rect 29089 7497 29101 7531
rect 29135 7528 29147 7531
rect 29270 7528 29276 7540
rect 29135 7500 29276 7528
rect 29135 7497 29147 7500
rect 29089 7491 29147 7497
rect 29270 7488 29276 7500
rect 29328 7488 29334 7540
rect 33137 7531 33195 7537
rect 33137 7497 33149 7531
rect 33183 7528 33195 7531
rect 33870 7528 33876 7540
rect 33183 7500 33876 7528
rect 33183 7497 33195 7500
rect 33137 7491 33195 7497
rect 33870 7488 33876 7500
rect 33928 7488 33934 7540
rect 34698 7488 34704 7540
rect 34756 7488 34762 7540
rect 35986 7488 35992 7540
rect 36044 7528 36050 7540
rect 36081 7531 36139 7537
rect 36081 7528 36093 7531
rect 36044 7500 36093 7528
rect 36044 7488 36050 7500
rect 36081 7497 36093 7500
rect 36127 7497 36139 7531
rect 36081 7491 36139 7497
rect 36446 7488 36452 7540
rect 36504 7528 36510 7540
rect 36541 7531 36599 7537
rect 36541 7528 36553 7531
rect 36504 7500 36553 7528
rect 36504 7488 36510 7500
rect 36541 7497 36553 7500
rect 36587 7497 36599 7531
rect 36541 7491 36599 7497
rect 37090 7488 37096 7540
rect 37148 7488 37154 7540
rect 37734 7488 37740 7540
rect 37792 7528 37798 7540
rect 38197 7531 38255 7537
rect 38197 7528 38209 7531
rect 37792 7500 38209 7528
rect 37792 7488 37798 7500
rect 38197 7497 38209 7500
rect 38243 7497 38255 7531
rect 38197 7491 38255 7497
rect 38286 7488 38292 7540
rect 38344 7488 38350 7540
rect 38838 7488 38844 7540
rect 38896 7528 38902 7540
rect 39301 7531 39359 7537
rect 39301 7528 39313 7531
rect 38896 7500 39313 7528
rect 38896 7488 38902 7500
rect 39301 7497 39313 7500
rect 39347 7497 39359 7531
rect 39301 7491 39359 7497
rect 39669 7531 39727 7537
rect 39669 7497 39681 7531
rect 39715 7528 39727 7531
rect 40218 7528 40224 7540
rect 39715 7500 40224 7528
rect 39715 7497 39727 7500
rect 39669 7491 39727 7497
rect 18380 7432 18460 7460
rect 18524 7432 20116 7460
rect 18380 7420 18386 7432
rect 16669 7395 16727 7401
rect 15896 7364 16436 7392
rect 15896 7352 15902 7364
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 14884 7296 15025 7324
rect 14884 7284 14890 7296
rect 15013 7293 15025 7296
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 12308 7228 12817 7256
rect 12308 7216 12314 7228
rect 12805 7225 12817 7228
rect 12851 7225 12863 7259
rect 12805 7219 12863 7225
rect 14458 7216 14464 7268
rect 14516 7256 14522 7268
rect 16408 7265 16436 7364
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16936 7395 16994 7401
rect 16936 7361 16948 7395
rect 16982 7392 16994 7395
rect 18138 7392 18144 7404
rect 16982 7364 18144 7392
rect 16982 7361 16994 7364
rect 16936 7355 16994 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18432 7401 18460 7432
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7361 18475 7395
rect 18417 7355 18475 7361
rect 18684 7395 18742 7401
rect 18684 7361 18696 7395
rect 18730 7392 18742 7395
rect 19426 7392 19432 7404
rect 18730 7364 19432 7392
rect 18730 7361 18742 7364
rect 18684 7355 18742 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7293 19947 7327
rect 20088 7324 20116 7432
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7392 23443 7395
rect 23474 7392 23480 7404
rect 23431 7364 23480 7392
rect 23431 7361 23443 7364
rect 23385 7355 23443 7361
rect 23474 7352 23480 7364
rect 23532 7352 23538 7404
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7392 24179 7395
rect 24412 7392 24440 7488
rect 25222 7460 25228 7472
rect 24872 7432 25228 7460
rect 24167 7364 24440 7392
rect 24167 7361 24179 7364
rect 24121 7355 24179 7361
rect 24762 7352 24768 7404
rect 24820 7352 24826 7404
rect 24872 7324 24900 7432
rect 25222 7420 25228 7432
rect 25280 7420 25286 7472
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 25608 7392 25636 7488
rect 25777 7463 25835 7469
rect 25777 7429 25789 7463
rect 25823 7460 25835 7463
rect 25866 7460 25872 7472
rect 25823 7432 25872 7460
rect 25823 7429 25835 7432
rect 25777 7423 25835 7429
rect 25866 7420 25872 7432
rect 25924 7460 25930 7472
rect 26142 7460 26148 7472
rect 25924 7432 26148 7460
rect 25924 7420 25930 7432
rect 26142 7420 26148 7432
rect 26200 7420 26206 7472
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 34514 7460 34520 7472
rect 26936 7432 34520 7460
rect 26936 7420 26942 7432
rect 34514 7420 34520 7432
rect 34572 7420 34578 7472
rect 34716 7460 34744 7488
rect 37108 7460 37136 7488
rect 37921 7463 37979 7469
rect 37921 7460 37933 7463
rect 34716 7432 36032 7460
rect 37108 7432 37933 7460
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 25608 7364 26985 7392
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 29181 7395 29239 7401
rect 29181 7361 29193 7395
rect 29227 7392 29239 7395
rect 30193 7395 30251 7401
rect 30193 7392 30205 7395
rect 29227 7364 30205 7392
rect 29227 7361 29239 7364
rect 29181 7355 29239 7361
rect 30193 7361 30205 7364
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 30552 7395 30610 7401
rect 30552 7361 30564 7395
rect 30598 7392 30610 7395
rect 33134 7392 33140 7404
rect 30598 7364 33140 7392
rect 30598 7361 30610 7364
rect 30552 7355 30610 7361
rect 33134 7352 33140 7364
rect 33192 7352 33198 7404
rect 33318 7352 33324 7404
rect 33376 7392 33382 7404
rect 33505 7395 33563 7401
rect 33505 7392 33517 7395
rect 33376 7364 33517 7392
rect 33376 7352 33382 7364
rect 33505 7361 33517 7364
rect 33551 7361 33563 7395
rect 34330 7392 34336 7404
rect 33505 7355 33563 7361
rect 33796 7364 34336 7392
rect 20088 7296 24900 7324
rect 24964 7324 24992 7352
rect 25961 7327 26019 7333
rect 25961 7324 25973 7327
rect 24964 7296 25973 7324
rect 19889 7287 19947 7293
rect 25961 7293 25973 7296
rect 26007 7293 26019 7327
rect 25961 7287 26019 7293
rect 29273 7327 29331 7333
rect 29273 7293 29285 7327
rect 29319 7293 29331 7327
rect 29273 7287 29331 7293
rect 16393 7259 16451 7265
rect 14516 7228 14964 7256
rect 14516 7216 14522 7228
rect 14550 7188 14556 7200
rect 11532 7160 14556 7188
rect 11333 7151 11391 7157
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 14936 7188 14964 7228
rect 16393 7225 16405 7259
rect 16439 7225 16451 7259
rect 16393 7219 16451 7225
rect 17678 7216 17684 7268
rect 17736 7256 17742 7268
rect 19797 7259 19855 7265
rect 17736 7228 18184 7256
rect 17736 7216 17742 7228
rect 16022 7188 16028 7200
rect 14936 7160 16028 7188
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 16908 7160 18061 7188
rect 16908 7148 16914 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 18156 7188 18184 7228
rect 19797 7225 19809 7259
rect 19843 7256 19855 7259
rect 19904 7256 19932 7287
rect 21174 7256 21180 7268
rect 19843 7228 21180 7256
rect 19843 7225 19855 7228
rect 19797 7219 19855 7225
rect 21174 7216 21180 7228
rect 21232 7216 21238 7268
rect 28537 7259 28595 7265
rect 28537 7256 28549 7259
rect 24596 7228 28549 7256
rect 24596 7200 24624 7228
rect 28537 7225 28549 7228
rect 28583 7256 28595 7259
rect 29288 7256 29316 7287
rect 29638 7284 29644 7336
rect 29696 7284 29702 7336
rect 30282 7284 30288 7336
rect 30340 7284 30346 7336
rect 32122 7284 32128 7336
rect 32180 7284 32186 7336
rect 33594 7284 33600 7336
rect 33652 7284 33658 7336
rect 33796 7333 33824 7364
rect 34330 7352 34336 7364
rect 34388 7392 34394 7404
rect 34698 7392 34704 7404
rect 34388 7364 34704 7392
rect 34388 7352 34394 7364
rect 34698 7352 34704 7364
rect 34756 7352 34762 7404
rect 34876 7395 34934 7401
rect 34876 7361 34888 7395
rect 34922 7392 34934 7395
rect 35894 7392 35900 7404
rect 34922 7364 35900 7392
rect 34922 7361 34934 7364
rect 34876 7355 34934 7361
rect 35894 7352 35900 7364
rect 35952 7352 35958 7404
rect 33781 7327 33839 7333
rect 33781 7293 33793 7327
rect 33827 7293 33839 7327
rect 33781 7287 33839 7293
rect 34241 7327 34299 7333
rect 34241 7293 34253 7327
rect 34287 7324 34299 7327
rect 34609 7327 34667 7333
rect 34609 7324 34621 7327
rect 34287 7296 34621 7324
rect 34287 7293 34299 7296
rect 34241 7287 34299 7293
rect 34609 7293 34621 7296
rect 34655 7293 34667 7327
rect 34609 7287 34667 7293
rect 28583 7228 29316 7256
rect 28583 7225 28595 7228
rect 28537 7219 28595 7225
rect 33042 7216 33048 7268
rect 33100 7256 33106 7268
rect 34256 7256 34284 7287
rect 33100 7228 34284 7256
rect 33100 7216 33106 7228
rect 34624 7200 34652 7287
rect 36004 7265 36032 7432
rect 37921 7429 37933 7432
rect 37967 7429 37979 7463
rect 37921 7423 37979 7429
rect 36449 7395 36507 7401
rect 36449 7361 36461 7395
rect 36495 7392 36507 7395
rect 38304 7392 38332 7488
rect 38933 7463 38991 7469
rect 38933 7429 38945 7463
rect 38979 7460 38991 7463
rect 39684 7460 39712 7491
rect 40218 7488 40224 7500
rect 40276 7488 40282 7540
rect 41414 7488 41420 7540
rect 41472 7488 41478 7540
rect 42150 7488 42156 7540
rect 42208 7488 42214 7540
rect 43254 7488 43260 7540
rect 43312 7488 43318 7540
rect 43898 7528 43904 7540
rect 43456 7500 43904 7528
rect 38979 7432 39712 7460
rect 38979 7429 38991 7432
rect 38933 7423 38991 7429
rect 40126 7420 40132 7472
rect 40184 7460 40190 7472
rect 41046 7460 41052 7472
rect 40184 7432 41052 7460
rect 40184 7420 40190 7432
rect 41046 7420 41052 7432
rect 41104 7420 41110 7472
rect 36495 7364 38332 7392
rect 36495 7361 36507 7364
rect 36449 7355 36507 7361
rect 38838 7352 38844 7404
rect 38896 7352 38902 7404
rect 43456 7401 43484 7500
rect 43898 7488 43904 7500
rect 43956 7488 43962 7540
rect 43990 7488 43996 7540
rect 44048 7488 44054 7540
rect 44082 7488 44088 7540
rect 44140 7488 44146 7540
rect 44174 7488 44180 7540
rect 44232 7488 44238 7540
rect 44450 7488 44456 7540
rect 44508 7528 44514 7540
rect 44910 7528 44916 7540
rect 44508 7500 44916 7528
rect 44508 7488 44514 7500
rect 44910 7488 44916 7500
rect 44968 7488 44974 7540
rect 45554 7488 45560 7540
rect 45612 7528 45618 7540
rect 46290 7528 46296 7540
rect 45612 7500 46296 7528
rect 45612 7488 45618 7500
rect 46290 7488 46296 7500
rect 46348 7528 46354 7540
rect 46477 7531 46535 7537
rect 46477 7528 46489 7531
rect 46348 7500 46489 7528
rect 46348 7488 46354 7500
rect 46477 7497 46489 7500
rect 46523 7497 46535 7531
rect 46477 7491 46535 7497
rect 47946 7488 47952 7540
rect 48004 7488 48010 7540
rect 48406 7488 48412 7540
rect 48464 7488 48470 7540
rect 50706 7528 50712 7540
rect 48884 7500 50712 7528
rect 44100 7401 44128 7488
rect 44192 7460 44220 7488
rect 44729 7463 44787 7469
rect 44729 7460 44741 7463
rect 44192 7432 44741 7460
rect 44729 7429 44741 7432
rect 44775 7429 44787 7463
rect 44729 7423 44787 7429
rect 45646 7420 45652 7472
rect 45704 7460 45710 7472
rect 47765 7463 47823 7469
rect 47765 7460 47777 7463
rect 45704 7432 47777 7460
rect 45704 7420 45710 7432
rect 47765 7429 47777 7432
rect 47811 7460 47823 7463
rect 47811 7432 48452 7460
rect 47811 7429 47823 7432
rect 47765 7423 47823 7429
rect 39761 7395 39819 7401
rect 39761 7361 39773 7395
rect 39807 7392 39819 7395
rect 40773 7395 40831 7401
rect 40773 7392 40785 7395
rect 39807 7364 40785 7392
rect 39807 7361 39819 7364
rect 39761 7355 39819 7361
rect 40773 7361 40785 7364
rect 40819 7361 40831 7395
rect 40773 7355 40831 7361
rect 43441 7395 43499 7401
rect 43441 7361 43453 7395
rect 43487 7361 43499 7395
rect 43441 7355 43499 7361
rect 44085 7395 44143 7401
rect 44085 7361 44097 7395
rect 44131 7361 44143 7395
rect 44085 7355 44143 7361
rect 45097 7395 45155 7401
rect 45097 7361 45109 7395
rect 45143 7392 45155 7395
rect 45186 7392 45192 7404
rect 45143 7364 45192 7392
rect 45143 7361 45155 7364
rect 45097 7355 45155 7361
rect 45186 7352 45192 7364
rect 45244 7352 45250 7404
rect 45364 7395 45422 7401
rect 45364 7361 45376 7395
rect 45410 7392 45422 7395
rect 47213 7395 47271 7401
rect 47213 7392 47225 7395
rect 45410 7364 47225 7392
rect 45410 7361 45422 7364
rect 45364 7355 45422 7361
rect 47213 7361 47225 7364
rect 47259 7361 47271 7395
rect 47213 7355 47271 7361
rect 48317 7395 48375 7401
rect 48317 7361 48329 7395
rect 48363 7361 48375 7395
rect 48317 7355 48375 7361
rect 36725 7327 36783 7333
rect 36725 7293 36737 7327
rect 36771 7324 36783 7327
rect 37182 7324 37188 7336
rect 36771 7296 37188 7324
rect 36771 7293 36783 7296
rect 36725 7287 36783 7293
rect 37182 7284 37188 7296
rect 37240 7284 37246 7336
rect 37277 7327 37335 7333
rect 37277 7293 37289 7327
rect 37323 7293 37335 7327
rect 37277 7287 37335 7293
rect 35989 7259 36047 7265
rect 35989 7225 36001 7259
rect 36035 7256 36047 7259
rect 37292 7256 37320 7287
rect 39022 7284 39028 7336
rect 39080 7284 39086 7336
rect 39850 7284 39856 7336
rect 39908 7284 39914 7336
rect 40034 7284 40040 7336
rect 40092 7324 40098 7336
rect 40129 7327 40187 7333
rect 40129 7324 40141 7327
rect 40092 7296 40141 7324
rect 40092 7284 40098 7296
rect 40129 7293 40141 7296
rect 40175 7293 40187 7327
rect 40129 7287 40187 7293
rect 46566 7284 46572 7336
rect 46624 7284 46630 7336
rect 36035 7228 37320 7256
rect 38396 7228 40080 7256
rect 36035 7225 36047 7228
rect 35989 7219 36047 7225
rect 20070 7188 20076 7200
rect 18156 7160 20076 7188
rect 18049 7151 18107 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20901 7191 20959 7197
rect 20901 7157 20913 7191
rect 20947 7188 20959 7191
rect 20990 7188 20996 7200
rect 20947 7160 20996 7188
rect 20947 7157 20959 7160
rect 20901 7151 20959 7157
rect 20990 7148 20996 7160
rect 21048 7188 21054 7200
rect 21450 7188 21456 7200
rect 21048 7160 21456 7188
rect 21048 7148 21054 7160
rect 21450 7148 21456 7160
rect 21508 7188 21514 7200
rect 24394 7188 24400 7200
rect 21508 7160 24400 7188
rect 21508 7148 21514 7160
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 24578 7148 24584 7200
rect 24636 7148 24642 7200
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 29546 7188 29552 7200
rect 25280 7160 29552 7188
rect 25280 7148 25286 7160
rect 29546 7148 29552 7160
rect 29604 7148 29610 7200
rect 29730 7148 29736 7200
rect 29788 7188 29794 7200
rect 31665 7191 31723 7197
rect 31665 7188 31677 7191
rect 29788 7160 31677 7188
rect 29788 7148 29794 7160
rect 31665 7157 31677 7160
rect 31711 7157 31723 7191
rect 31665 7151 31723 7157
rect 32766 7148 32772 7200
rect 32824 7148 32830 7200
rect 34606 7148 34612 7200
rect 34664 7188 34670 7200
rect 35342 7188 35348 7200
rect 34664 7160 35348 7188
rect 34664 7148 34670 7160
rect 35342 7148 35348 7160
rect 35400 7148 35406 7200
rect 36722 7148 36728 7200
rect 36780 7188 36786 7200
rect 38396 7188 38424 7228
rect 40052 7200 40080 7228
rect 36780 7160 38424 7188
rect 36780 7148 36786 7160
rect 38470 7148 38476 7200
rect 38528 7148 38534 7200
rect 40034 7148 40040 7200
rect 40092 7148 40098 7200
rect 41877 7191 41935 7197
rect 41877 7157 41889 7191
rect 41923 7188 41935 7191
rect 41966 7188 41972 7200
rect 41923 7160 41972 7188
rect 41923 7157 41935 7160
rect 41877 7151 41935 7157
rect 41966 7148 41972 7160
rect 42024 7188 42030 7200
rect 42426 7188 42432 7200
rect 42024 7160 42432 7188
rect 42024 7148 42030 7160
rect 42426 7148 42432 7160
rect 42484 7148 42490 7200
rect 42610 7148 42616 7200
rect 42668 7148 42674 7200
rect 48332 7188 48360 7355
rect 48424 7256 48452 7432
rect 48774 7352 48780 7404
rect 48832 7352 48838 7404
rect 48884 7401 48912 7500
rect 50706 7488 50712 7500
rect 50764 7488 50770 7540
rect 50798 7488 50804 7540
rect 50856 7488 50862 7540
rect 51169 7531 51227 7537
rect 51169 7497 51181 7531
rect 51215 7528 51227 7531
rect 52178 7528 52184 7540
rect 51215 7500 52184 7528
rect 51215 7497 51227 7500
rect 51169 7491 51227 7497
rect 52178 7488 52184 7500
rect 52236 7488 52242 7540
rect 52730 7488 52736 7540
rect 52788 7528 52794 7540
rect 53466 7528 53472 7540
rect 52788 7500 53472 7528
rect 52788 7488 52794 7500
rect 53466 7488 53472 7500
rect 53524 7488 53530 7540
rect 53558 7488 53564 7540
rect 53616 7488 53622 7540
rect 53926 7488 53932 7540
rect 53984 7488 53990 7540
rect 54018 7488 54024 7540
rect 54076 7528 54082 7540
rect 54297 7531 54355 7537
rect 54297 7528 54309 7531
rect 54076 7500 54309 7528
rect 54076 7488 54082 7500
rect 54297 7497 54309 7500
rect 54343 7497 54355 7531
rect 54297 7491 54355 7497
rect 54386 7488 54392 7540
rect 54444 7528 54450 7540
rect 55033 7531 55091 7537
rect 55033 7528 55045 7531
rect 54444 7500 55045 7528
rect 54444 7488 54450 7500
rect 55033 7497 55045 7500
rect 55079 7497 55091 7531
rect 55033 7491 55091 7497
rect 55306 7488 55312 7540
rect 55364 7488 55370 7540
rect 55398 7488 55404 7540
rect 55456 7528 55462 7540
rect 56045 7531 56103 7537
rect 56045 7528 56057 7531
rect 55456 7500 56057 7528
rect 55456 7488 55462 7500
rect 56045 7497 56057 7500
rect 56091 7528 56103 7531
rect 56226 7528 56232 7540
rect 56091 7500 56232 7528
rect 56091 7497 56103 7500
rect 56045 7491 56103 7497
rect 56226 7488 56232 7500
rect 56284 7488 56290 7540
rect 56870 7488 56876 7540
rect 56928 7528 56934 7540
rect 57422 7528 57428 7540
rect 56928 7500 57428 7528
rect 56928 7488 56934 7500
rect 57422 7488 57428 7500
rect 57480 7488 57486 7540
rect 57698 7488 57704 7540
rect 57756 7528 57762 7540
rect 58437 7531 58495 7537
rect 58437 7528 58449 7531
rect 57756 7500 58449 7528
rect 57756 7488 57762 7500
rect 58437 7497 58449 7500
rect 58483 7497 58495 7531
rect 58437 7491 58495 7497
rect 50614 7420 50620 7472
rect 50672 7460 50678 7472
rect 50672 7432 51488 7460
rect 50672 7420 50678 7432
rect 48869 7395 48927 7401
rect 48869 7361 48881 7395
rect 48915 7361 48927 7395
rect 48869 7355 48927 7361
rect 49050 7352 49056 7404
rect 49108 7352 49114 7404
rect 49878 7352 49884 7404
rect 49936 7401 49942 7404
rect 49936 7395 49964 7401
rect 49952 7361 49964 7395
rect 49936 7355 49964 7361
rect 51261 7395 51319 7401
rect 51261 7361 51273 7395
rect 51307 7361 51319 7395
rect 51261 7355 51319 7361
rect 49936 7352 49942 7355
rect 48498 7284 48504 7336
rect 48556 7284 48562 7336
rect 48792 7324 48820 7352
rect 49789 7327 49847 7333
rect 49789 7324 49801 7327
rect 48792 7296 49801 7324
rect 49789 7293 49801 7296
rect 49835 7293 49847 7327
rect 49789 7287 49847 7293
rect 50065 7327 50123 7333
rect 50065 7293 50077 7327
rect 50111 7324 50123 7327
rect 50246 7324 50252 7336
rect 50111 7296 50252 7324
rect 50111 7293 50123 7296
rect 50065 7287 50123 7293
rect 50246 7284 50252 7296
rect 50304 7284 50310 7336
rect 51276 7324 51304 7355
rect 50448 7296 51304 7324
rect 48590 7256 48596 7268
rect 48424 7228 48596 7256
rect 48590 7216 48596 7228
rect 48648 7256 48654 7268
rect 49510 7256 49516 7268
rect 48648 7228 49516 7256
rect 48648 7216 48654 7228
rect 49510 7216 49516 7228
rect 49568 7216 49574 7268
rect 50062 7188 50068 7200
rect 48332 7160 50068 7188
rect 50062 7148 50068 7160
rect 50120 7148 50126 7200
rect 50154 7148 50160 7200
rect 50212 7188 50218 7200
rect 50448 7188 50476 7296
rect 51350 7284 51356 7336
rect 51408 7284 51414 7336
rect 51460 7324 51488 7432
rect 53006 7352 53012 7404
rect 53064 7352 53070 7404
rect 53745 7395 53803 7401
rect 53745 7361 53757 7395
rect 53791 7392 53803 7395
rect 53944 7392 53972 7488
rect 53791 7364 53972 7392
rect 53791 7361 53803 7364
rect 53745 7355 53803 7361
rect 54478 7352 54484 7404
rect 54536 7352 54542 7404
rect 55416 7324 55444 7488
rect 55490 7420 55496 7472
rect 55548 7460 55554 7472
rect 55769 7463 55827 7469
rect 55769 7460 55781 7463
rect 55548 7432 55781 7460
rect 55548 7420 55554 7432
rect 55769 7429 55781 7432
rect 55815 7460 55827 7463
rect 55858 7460 55864 7472
rect 55815 7432 55864 7460
rect 55815 7429 55827 7432
rect 55769 7423 55827 7429
rect 55858 7420 55864 7432
rect 55916 7420 55922 7472
rect 58342 7352 58348 7404
rect 58400 7352 58406 7404
rect 51460 7296 55444 7324
rect 56686 7284 56692 7336
rect 56744 7324 56750 7336
rect 57057 7327 57115 7333
rect 57057 7324 57069 7327
rect 56744 7296 57069 7324
rect 56744 7284 56750 7296
rect 57057 7293 57069 7296
rect 57103 7293 57115 7327
rect 57057 7287 57115 7293
rect 50212 7160 50476 7188
rect 50212 7148 50218 7160
rect 50706 7148 50712 7200
rect 50764 7148 50770 7200
rect 52178 7148 52184 7200
rect 52236 7188 52242 7200
rect 52549 7191 52607 7197
rect 52549 7188 52561 7191
rect 52236 7160 52561 7188
rect 52236 7148 52242 7160
rect 52549 7157 52561 7160
rect 52595 7188 52607 7191
rect 55490 7188 55496 7200
rect 52595 7160 55496 7188
rect 52595 7157 52607 7160
rect 52549 7151 52607 7157
rect 55490 7148 55496 7160
rect 55548 7148 55554 7200
rect 56505 7191 56563 7197
rect 56505 7157 56517 7191
rect 56551 7188 56563 7191
rect 56778 7188 56784 7200
rect 56551 7160 56784 7188
rect 56551 7157 56563 7160
rect 56505 7151 56563 7157
rect 56778 7148 56784 7160
rect 56836 7188 56842 7200
rect 57054 7188 57060 7200
rect 56836 7160 57060 7188
rect 56836 7148 56842 7160
rect 57054 7148 57060 7160
rect 57112 7148 57118 7200
rect 57698 7148 57704 7200
rect 57756 7148 57762 7200
rect 58066 7148 58072 7200
rect 58124 7148 58130 7200
rect 1104 7098 58880 7120
rect 1104 7046 8172 7098
rect 8224 7046 8236 7098
rect 8288 7046 8300 7098
rect 8352 7046 8364 7098
rect 8416 7046 8428 7098
rect 8480 7046 22616 7098
rect 22668 7046 22680 7098
rect 22732 7046 22744 7098
rect 22796 7046 22808 7098
rect 22860 7046 22872 7098
rect 22924 7046 37060 7098
rect 37112 7046 37124 7098
rect 37176 7046 37188 7098
rect 37240 7046 37252 7098
rect 37304 7046 37316 7098
rect 37368 7046 51504 7098
rect 51556 7046 51568 7098
rect 51620 7046 51632 7098
rect 51684 7046 51696 7098
rect 51748 7046 51760 7098
rect 51812 7046 58880 7098
rect 1104 7024 58880 7046
rect 9490 6944 9496 6996
rect 9548 6984 9554 6996
rect 9548 6956 10272 6984
rect 9548 6944 9554 6956
rect 3513 6919 3571 6925
rect 3513 6885 3525 6919
rect 3559 6885 3571 6919
rect 3513 6879 3571 6885
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 9508 6916 9536 6944
rect 9950 6916 9956 6928
rect 8803 6888 9536 6916
rect 9600 6888 9956 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 3528 6848 3556 6879
rect 3528 6820 3924 6848
rect 1762 6740 1768 6792
rect 1820 6780 1826 6792
rect 3896 6789 3924 6820
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 1820 6752 2145 6780
rect 1820 6740 1826 6752
rect 2133 6749 2145 6752
rect 2179 6780 2191 6783
rect 3881 6783 3939 6789
rect 2179 6752 3740 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2400 6715 2458 6721
rect 2400 6681 2412 6715
rect 2446 6712 2458 6715
rect 3326 6712 3332 6724
rect 2446 6684 3332 6712
rect 2446 6681 2458 6684
rect 2400 6675 2458 6681
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 3712 6712 3740 6752
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 5442 6780 5448 6792
rect 3927 6752 5448 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 9600 6780 9628 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 10134 6808 10140 6860
rect 10192 6808 10198 6860
rect 10244 6848 10272 6956
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 13173 6987 13231 6993
rect 10560 6956 11100 6984
rect 10560 6944 10566 6956
rect 10530 6851 10588 6857
rect 10530 6848 10542 6851
rect 10244 6820 10542 6848
rect 10530 6817 10542 6820
rect 10576 6817 10588 6851
rect 10530 6811 10588 6817
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 11072 6848 11100 6956
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13262 6984 13268 6996
rect 13219 6956 13268 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 14608 6956 16620 6984
rect 14608 6944 14614 6956
rect 14090 6876 14096 6928
rect 14148 6876 14154 6928
rect 15286 6876 15292 6928
rect 15344 6916 15350 6928
rect 16592 6916 16620 6956
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 19484 6956 19901 6984
rect 19484 6944 19490 6956
rect 19889 6953 19901 6956
rect 19935 6953 19947 6987
rect 32033 6987 32091 6993
rect 19889 6947 19947 6953
rect 19996 6956 31754 6984
rect 19996 6916 20024 6956
rect 15344 6888 15700 6916
rect 16592 6888 20024 6916
rect 15344 6876 15350 6888
rect 10735 6820 11100 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13596 6820 13737 6848
rect 13596 6808 13602 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 14642 6808 14648 6860
rect 14700 6808 14706 6860
rect 15013 6851 15071 6857
rect 15013 6817 15025 6851
rect 15059 6848 15071 6851
rect 15562 6848 15568 6860
rect 15059 6820 15568 6848
rect 15059 6817 15071 6820
rect 15013 6811 15071 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 15672 6857 15700 6888
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 22370 6916 22376 6928
rect 20128 6888 22376 6916
rect 20128 6876 20134 6888
rect 22370 6876 22376 6888
rect 22428 6876 22434 6928
rect 30282 6876 30288 6928
rect 30340 6916 30346 6928
rect 31726 6916 31754 6956
rect 32033 6953 32045 6987
rect 32079 6984 32091 6987
rect 32122 6984 32128 6996
rect 32079 6956 32128 6984
rect 32079 6953 32091 6956
rect 32033 6947 32091 6953
rect 32122 6944 32128 6956
rect 32180 6944 32186 6996
rect 33134 6944 33140 6996
rect 33192 6984 33198 6996
rect 33505 6987 33563 6993
rect 33505 6984 33517 6987
rect 33192 6956 33517 6984
rect 33192 6944 33198 6956
rect 33505 6953 33517 6956
rect 33551 6953 33563 6987
rect 33505 6947 33563 6953
rect 33594 6944 33600 6996
rect 33652 6984 33658 6996
rect 34333 6987 34391 6993
rect 34333 6984 34345 6987
rect 33652 6956 34345 6984
rect 33652 6944 33658 6956
rect 34333 6953 34345 6956
rect 34379 6953 34391 6987
rect 34333 6947 34391 6953
rect 34977 6987 35035 6993
rect 34977 6953 34989 6987
rect 35023 6984 35035 6987
rect 35342 6984 35348 6996
rect 35023 6956 35348 6984
rect 35023 6953 35035 6956
rect 34977 6947 35035 6953
rect 35342 6944 35348 6956
rect 35400 6944 35406 6996
rect 35894 6944 35900 6996
rect 35952 6984 35958 6996
rect 36725 6987 36783 6993
rect 36725 6984 36737 6987
rect 35952 6956 36737 6984
rect 35952 6944 35958 6956
rect 36725 6953 36737 6956
rect 36771 6953 36783 6987
rect 36725 6947 36783 6953
rect 37734 6944 37740 6996
rect 37792 6944 37798 6996
rect 38838 6944 38844 6996
rect 38896 6984 38902 6996
rect 39669 6987 39727 6993
rect 39669 6984 39681 6987
rect 38896 6956 39681 6984
rect 38896 6944 38902 6956
rect 39669 6953 39681 6956
rect 39715 6953 39727 6987
rect 39669 6947 39727 6953
rect 40129 6987 40187 6993
rect 40129 6953 40141 6987
rect 40175 6984 40187 6987
rect 40494 6984 40500 6996
rect 40175 6956 40500 6984
rect 40175 6953 40187 6956
rect 40129 6947 40187 6953
rect 40494 6944 40500 6956
rect 40552 6984 40558 6996
rect 40678 6984 40684 6996
rect 40552 6956 40684 6984
rect 40552 6944 40558 6956
rect 40678 6944 40684 6956
rect 40736 6944 40742 6996
rect 40954 6944 40960 6996
rect 41012 6944 41018 6996
rect 44450 6944 44456 6996
rect 44508 6944 44514 6996
rect 45465 6987 45523 6993
rect 45465 6953 45477 6987
rect 45511 6984 45523 6987
rect 46566 6984 46572 6996
rect 45511 6956 46572 6984
rect 45511 6953 45523 6956
rect 45465 6947 45523 6953
rect 46566 6944 46572 6956
rect 46624 6944 46630 6996
rect 48314 6944 48320 6996
rect 48372 6944 48378 6996
rect 48590 6944 48596 6996
rect 48648 6944 48654 6996
rect 49513 6987 49571 6993
rect 49513 6953 49525 6987
rect 49559 6984 49571 6987
rect 49602 6984 49608 6996
rect 49559 6956 49608 6984
rect 49559 6953 49571 6956
rect 49513 6947 49571 6953
rect 49602 6944 49608 6956
rect 49660 6984 49666 6996
rect 50246 6984 50252 6996
rect 49660 6956 50252 6984
rect 49660 6944 49666 6956
rect 50246 6944 50252 6956
rect 50304 6944 50310 6996
rect 50709 6987 50767 6993
rect 50709 6953 50721 6987
rect 50755 6984 50767 6987
rect 51350 6984 51356 6996
rect 50755 6956 51356 6984
rect 50755 6953 50767 6956
rect 50709 6947 50767 6953
rect 36078 6916 36084 6928
rect 30340 6888 30420 6916
rect 31726 6888 36084 6916
rect 30340 6876 30346 6888
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 16022 6808 16028 6860
rect 16080 6857 16086 6860
rect 16080 6851 16108 6857
rect 16096 6817 16108 6851
rect 16080 6811 16108 6817
rect 16080 6808 16086 6811
rect 16206 6808 16212 6860
rect 16264 6808 16270 6860
rect 16850 6808 16856 6860
rect 16908 6808 16914 6860
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 18196 6820 18245 6848
rect 18196 6808 18202 6820
rect 18233 6817 18245 6820
rect 18279 6848 18291 6851
rect 18966 6848 18972 6860
rect 18279 6820 18972 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 19242 6808 19248 6860
rect 19300 6808 19306 6860
rect 19978 6808 19984 6860
rect 20036 6848 20042 6860
rect 21818 6848 21824 6860
rect 20036 6820 21824 6848
rect 20036 6808 20042 6820
rect 21818 6808 21824 6820
rect 21876 6848 21882 6860
rect 23382 6848 23388 6860
rect 21876 6820 23388 6848
rect 21876 6808 21882 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 25038 6808 25044 6860
rect 25096 6808 25102 6860
rect 30392 6848 30420 6888
rect 36078 6876 36084 6888
rect 36136 6876 36142 6928
rect 36906 6876 36912 6928
rect 36964 6916 36970 6928
rect 37093 6919 37151 6925
rect 37093 6916 37105 6919
rect 36964 6888 37105 6916
rect 36964 6876 36970 6888
rect 37093 6885 37105 6888
rect 37139 6916 37151 6919
rect 40972 6916 41000 6944
rect 37139 6888 41000 6916
rect 44468 6916 44496 6944
rect 48332 6916 48360 6944
rect 49053 6919 49111 6925
rect 49053 6916 49065 6919
rect 44468 6888 47072 6916
rect 48332 6888 49065 6916
rect 37139 6885 37151 6888
rect 37093 6879 37151 6885
rect 30561 6851 30619 6857
rect 30561 6848 30573 6851
rect 27540 6820 28120 6848
rect 30392 6820 30573 6848
rect 9539 6752 9628 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 14918 6780 14924 6792
rect 11532 6752 14924 6780
rect 7392 6712 7420 6740
rect 7622 6715 7680 6721
rect 7622 6712 7634 6715
rect 3712 6684 7420 6712
rect 7484 6684 7634 6712
rect 4430 6604 4436 6656
rect 4488 6604 4494 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7484 6644 7512 6684
rect 7622 6681 7634 6684
rect 7668 6681 7680 6715
rect 11532 6712 11560 6752
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 7622 6675 7680 6681
rect 11164 6684 11560 6712
rect 11692 6715 11750 6721
rect 7331 6616 7512 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 11164 6644 11192 6684
rect 11692 6681 11704 6715
rect 11738 6712 11750 6715
rect 13078 6712 13084 6724
rect 11738 6684 13084 6712
rect 11738 6681 11750 6684
rect 11692 6675 11750 6681
rect 13078 6672 13084 6684
rect 13136 6672 13142 6724
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 14734 6712 14740 6724
rect 13587 6684 14740 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 9364 6616 11192 6644
rect 11333 6647 11391 6653
rect 9364 6604 9370 6616
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 11514 6644 11520 6656
rect 11379 6616 11520 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 13633 6647 13691 6653
rect 13633 6613 13645 6647
rect 13679 6644 13691 6647
rect 14458 6644 14464 6656
rect 13679 6616 14464 6644
rect 13679 6613 13691 6616
rect 13633 6607 13691 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 15212 6644 15240 6743
rect 15930 6740 15936 6792
rect 15988 6740 15994 6792
rect 16868 6780 16896 6808
rect 19794 6780 19800 6792
rect 16868 6752 19800 6780
rect 19794 6740 19800 6752
rect 19852 6740 19858 6792
rect 18969 6715 19027 6721
rect 18969 6712 18981 6715
rect 17696 6684 18981 6712
rect 17696 6656 17724 6684
rect 18969 6681 18981 6684
rect 19015 6712 19027 6715
rect 19996 6712 20024 6808
rect 27540 6792 27568 6820
rect 27522 6780 27528 6792
rect 22066 6752 27528 6780
rect 20990 6712 20996 6724
rect 19015 6684 20024 6712
rect 20088 6684 20996 6712
rect 19015 6681 19027 6684
rect 18969 6675 19027 6681
rect 16758 6644 16764 6656
rect 15212 6616 16764 6644
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 17402 6644 17408 6656
rect 16899 6616 17408 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17678 6604 17684 6656
rect 17736 6604 17742 6656
rect 18874 6604 18880 6656
rect 18932 6644 18938 6656
rect 20088 6644 20116 6684
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 18932 6616 20116 6644
rect 18932 6604 18938 6616
rect 20254 6604 20260 6656
rect 20312 6604 20318 6656
rect 20625 6647 20683 6653
rect 20625 6613 20637 6647
rect 20671 6644 20683 6647
rect 21082 6644 21088 6656
rect 20671 6616 21088 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 21082 6604 21088 6616
rect 21140 6644 21146 6656
rect 22066 6644 22094 6752
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 27890 6740 27896 6792
rect 27948 6780 27954 6792
rect 27985 6783 28043 6789
rect 27985 6780 27997 6783
rect 27948 6752 27997 6780
rect 27948 6740 27954 6752
rect 27985 6749 27997 6752
rect 28031 6749 28043 6783
rect 27985 6743 28043 6749
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 26510 6712 26516 6724
rect 24903 6684 26516 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 26510 6672 26516 6684
rect 26568 6672 26574 6724
rect 28092 6712 28120 6820
rect 30561 6817 30573 6820
rect 30607 6817 30619 6851
rect 30561 6811 30619 6817
rect 31846 6808 31852 6860
rect 31904 6848 31910 6860
rect 32585 6851 32643 6857
rect 32585 6848 32597 6851
rect 31904 6820 32597 6848
rect 31904 6808 31910 6820
rect 32585 6817 32597 6820
rect 32631 6817 32643 6851
rect 32585 6811 32643 6817
rect 33778 6808 33784 6860
rect 33836 6808 33842 6860
rect 36173 6851 36231 6857
rect 36173 6817 36185 6851
rect 36219 6848 36231 6851
rect 36630 6848 36636 6860
rect 36219 6820 36636 6848
rect 36219 6817 36231 6820
rect 36173 6811 36231 6817
rect 36630 6808 36636 6820
rect 36688 6808 36694 6860
rect 38381 6851 38439 6857
rect 38381 6817 38393 6851
rect 38427 6848 38439 6851
rect 38470 6848 38476 6860
rect 38427 6820 38476 6848
rect 38427 6817 38439 6820
rect 38381 6811 38439 6817
rect 38470 6808 38476 6820
rect 38528 6808 38534 6860
rect 38930 6808 38936 6860
rect 38988 6808 38994 6860
rect 39114 6808 39120 6860
rect 39172 6808 39178 6860
rect 39850 6808 39856 6860
rect 39908 6848 39914 6860
rect 40405 6851 40463 6857
rect 40405 6848 40417 6851
rect 39908 6820 40417 6848
rect 39908 6808 39914 6820
rect 40405 6817 40417 6820
rect 40451 6848 40463 6851
rect 41506 6848 41512 6860
rect 40451 6820 41512 6848
rect 40451 6817 40463 6820
rect 40405 6811 40463 6817
rect 41506 6808 41512 6820
rect 41564 6808 41570 6860
rect 41874 6808 41880 6860
rect 41932 6808 41938 6860
rect 42245 6851 42303 6857
rect 42245 6817 42257 6851
rect 42291 6848 42303 6851
rect 43346 6848 43352 6860
rect 42291 6820 43352 6848
rect 42291 6817 42303 6820
rect 42245 6811 42303 6817
rect 28252 6783 28310 6789
rect 28252 6749 28264 6783
rect 28298 6780 28310 6783
rect 29178 6780 29184 6792
rect 28298 6752 29184 6780
rect 28298 6749 28310 6752
rect 28252 6743 28310 6749
rect 29178 6740 29184 6752
rect 29236 6740 29242 6792
rect 30650 6780 30656 6792
rect 29288 6752 30656 6780
rect 29288 6712 29316 6752
rect 30650 6740 30656 6752
rect 30708 6740 30714 6792
rect 30828 6783 30886 6789
rect 30828 6749 30840 6783
rect 30874 6780 30886 6783
rect 32766 6780 32772 6792
rect 30874 6752 32772 6780
rect 30874 6749 30886 6752
rect 30828 6743 30886 6749
rect 32766 6740 32772 6752
rect 32824 6740 32830 6792
rect 32858 6740 32864 6792
rect 32916 6740 32922 6792
rect 35989 6783 36047 6789
rect 35989 6749 36001 6783
rect 36035 6780 36047 6783
rect 36354 6780 36360 6792
rect 36035 6752 36360 6780
rect 36035 6749 36047 6752
rect 35989 6743 36047 6749
rect 36354 6740 36360 6752
rect 36412 6740 36418 6792
rect 37458 6740 37464 6792
rect 37516 6740 37522 6792
rect 40494 6780 40500 6792
rect 37568 6752 40500 6780
rect 29638 6712 29644 6724
rect 28092 6684 29316 6712
rect 29380 6684 29644 6712
rect 21140 6616 22094 6644
rect 21140 6604 21146 6616
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 24578 6644 24584 6656
rect 22888 6616 24584 6644
rect 22888 6604 22894 6616
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 27154 6644 27160 6656
rect 25188 6616 27160 6644
rect 25188 6604 25194 6616
rect 27154 6604 27160 6616
rect 27212 6604 27218 6656
rect 29380 6653 29408 6684
rect 29638 6672 29644 6684
rect 29696 6712 29702 6724
rect 32493 6715 32551 6721
rect 32493 6712 32505 6715
rect 29696 6684 30880 6712
rect 29696 6672 29702 6684
rect 30852 6656 30880 6684
rect 31220 6684 32505 6712
rect 31220 6656 31248 6684
rect 32493 6681 32505 6684
rect 32539 6681 32551 6715
rect 32493 6675 32551 6681
rect 35802 6672 35808 6724
rect 35860 6672 35866 6724
rect 29365 6647 29423 6653
rect 29365 6613 29377 6647
rect 29411 6613 29423 6647
rect 29365 6607 29423 6613
rect 30101 6647 30159 6653
rect 30101 6613 30113 6647
rect 30147 6644 30159 6647
rect 30282 6644 30288 6656
rect 30147 6616 30288 6644
rect 30147 6613 30159 6616
rect 30101 6607 30159 6613
rect 30282 6604 30288 6616
rect 30340 6604 30346 6656
rect 30466 6604 30472 6656
rect 30524 6604 30530 6656
rect 30834 6604 30840 6656
rect 30892 6604 30898 6656
rect 31202 6604 31208 6656
rect 31260 6604 31266 6656
rect 31938 6604 31944 6656
rect 31996 6604 32002 6656
rect 32398 6604 32404 6656
rect 32456 6604 32462 6656
rect 34698 6604 34704 6656
rect 34756 6644 34762 6656
rect 35345 6647 35403 6653
rect 35345 6644 35357 6647
rect 34756 6616 35357 6644
rect 34756 6604 34762 6616
rect 35345 6613 35357 6616
rect 35391 6644 35403 6647
rect 37568 6644 37596 6752
rect 40494 6740 40500 6752
rect 40552 6740 40558 6792
rect 41598 6740 41604 6792
rect 41656 6780 41662 6792
rect 42260 6780 42288 6811
rect 43346 6808 43352 6820
rect 43404 6808 43410 6860
rect 44453 6851 44511 6857
rect 44453 6817 44465 6851
rect 44499 6848 44511 6851
rect 44818 6848 44824 6860
rect 44499 6820 44824 6848
rect 44499 6817 44511 6820
rect 44453 6811 44511 6817
rect 44818 6808 44824 6820
rect 44876 6808 44882 6860
rect 46106 6848 46112 6860
rect 44928 6820 46112 6848
rect 41656 6752 42288 6780
rect 41656 6740 41662 6752
rect 42426 6740 42432 6792
rect 42484 6780 42490 6792
rect 44729 6783 44787 6789
rect 44729 6780 44741 6783
rect 42484 6752 44741 6780
rect 42484 6740 42490 6752
rect 44729 6749 44741 6752
rect 44775 6780 44787 6783
rect 44928 6780 44956 6820
rect 46106 6808 46112 6820
rect 46164 6808 46170 6860
rect 46937 6851 46995 6857
rect 46937 6848 46949 6851
rect 46216 6820 46949 6848
rect 44775 6752 44956 6780
rect 45833 6783 45891 6789
rect 44775 6749 44787 6752
rect 44729 6743 44787 6749
rect 45833 6749 45845 6783
rect 45879 6780 45891 6783
rect 46216 6780 46244 6820
rect 46937 6817 46949 6820
rect 46983 6817 46995 6851
rect 47044 6848 47072 6888
rect 49053 6885 49065 6888
rect 49099 6916 49111 6919
rect 49142 6916 49148 6928
rect 49099 6888 49148 6916
rect 49099 6885 49111 6888
rect 49053 6879 49111 6885
rect 49142 6876 49148 6888
rect 49200 6876 49206 6928
rect 49878 6876 49884 6928
rect 49936 6916 49942 6928
rect 50724 6916 50752 6947
rect 51350 6944 51356 6956
rect 51408 6944 51414 6996
rect 51626 6944 51632 6996
rect 51684 6984 51690 6996
rect 53098 6984 53104 6996
rect 51684 6956 53104 6984
rect 51684 6944 51690 6956
rect 53098 6944 53104 6956
rect 53156 6984 53162 6996
rect 54570 6984 54576 6996
rect 53156 6956 54576 6984
rect 53156 6944 53162 6956
rect 54570 6944 54576 6956
rect 54628 6944 54634 6996
rect 54938 6944 54944 6996
rect 54996 6984 55002 6996
rect 55398 6984 55404 6996
rect 54996 6956 55404 6984
rect 54996 6944 55002 6956
rect 55398 6944 55404 6956
rect 55456 6984 55462 6996
rect 55861 6987 55919 6993
rect 55861 6984 55873 6987
rect 55456 6956 55873 6984
rect 55456 6944 55462 6956
rect 55861 6953 55873 6956
rect 55907 6984 55919 6987
rect 56597 6987 56655 6993
rect 56597 6984 56609 6987
rect 55907 6956 56609 6984
rect 55907 6953 55919 6956
rect 55861 6947 55919 6953
rect 56597 6953 56609 6956
rect 56643 6953 56655 6987
rect 56597 6947 56655 6953
rect 49936 6888 50752 6916
rect 49936 6876 49942 6888
rect 50890 6876 50896 6928
rect 50948 6876 50954 6928
rect 52733 6919 52791 6925
rect 52733 6885 52745 6919
rect 52779 6916 52791 6919
rect 52822 6916 52828 6928
rect 52779 6888 52828 6916
rect 52779 6885 52791 6888
rect 52733 6879 52791 6885
rect 52822 6876 52828 6888
rect 52880 6876 52886 6928
rect 56226 6876 56232 6928
rect 56284 6876 56290 6928
rect 47765 6851 47823 6857
rect 47765 6848 47777 6851
rect 47044 6820 47777 6848
rect 46937 6811 46995 6817
rect 47765 6817 47777 6820
rect 47811 6848 47823 6851
rect 48498 6848 48504 6860
rect 47811 6820 48504 6848
rect 47811 6817 47823 6820
rect 47765 6811 47823 6817
rect 48498 6808 48504 6820
rect 48556 6848 48562 6860
rect 50908 6848 50936 6876
rect 51997 6851 52055 6857
rect 51997 6848 52009 6851
rect 48556 6820 52009 6848
rect 48556 6808 48562 6820
rect 51997 6817 52009 6820
rect 52043 6848 52055 6851
rect 53377 6851 53435 6857
rect 53377 6848 53389 6851
rect 52043 6820 53389 6848
rect 52043 6817 52055 6820
rect 51997 6811 52055 6817
rect 53377 6817 53389 6820
rect 53423 6817 53435 6851
rect 53377 6811 53435 6817
rect 54202 6808 54208 6860
rect 54260 6808 54266 6860
rect 54938 6808 54944 6860
rect 54996 6848 55002 6860
rect 54996 6820 56364 6848
rect 54996 6808 55002 6820
rect 45879 6752 46244 6780
rect 45879 6749 45891 6752
rect 45833 6743 45891 6749
rect 46290 6740 46296 6792
rect 46348 6740 46354 6792
rect 52181 6783 52239 6789
rect 52181 6749 52193 6783
rect 52227 6780 52239 6783
rect 52227 6752 52868 6780
rect 52227 6749 52239 6752
rect 52181 6743 52239 6749
rect 38746 6672 38752 6724
rect 38804 6712 38810 6724
rect 39390 6712 39396 6724
rect 38804 6684 39396 6712
rect 38804 6672 38810 6684
rect 39390 6672 39396 6684
rect 39448 6712 39454 6724
rect 40865 6715 40923 6721
rect 40865 6712 40877 6715
rect 39448 6684 40877 6712
rect 39448 6672 39454 6684
rect 40865 6681 40877 6684
rect 40911 6712 40923 6715
rect 41693 6715 41751 6721
rect 40911 6684 41414 6712
rect 40911 6681 40923 6684
rect 40865 6675 40923 6681
rect 35391 6616 37596 6644
rect 35391 6613 35403 6616
rect 35345 6607 35403 6613
rect 38194 6604 38200 6656
rect 38252 6644 38258 6656
rect 39022 6644 39028 6656
rect 38252 6616 39028 6644
rect 38252 6604 38258 6616
rect 39022 6604 39028 6616
rect 39080 6604 39086 6656
rect 40034 6604 40040 6656
rect 40092 6644 40098 6656
rect 41138 6644 41144 6656
rect 40092 6616 41144 6644
rect 40092 6604 40098 6616
rect 41138 6604 41144 6616
rect 41196 6604 41202 6656
rect 41386 6644 41414 6684
rect 41693 6681 41705 6715
rect 41739 6712 41751 6715
rect 42242 6712 42248 6724
rect 41739 6684 42248 6712
rect 41739 6681 41751 6684
rect 41693 6675 41751 6681
rect 42242 6672 42248 6684
rect 42300 6672 42306 6724
rect 42444 6684 42656 6712
rect 42444 6644 42472 6684
rect 41386 6616 42472 6644
rect 42518 6604 42524 6656
rect 42576 6604 42582 6656
rect 42628 6644 42656 6684
rect 42702 6672 42708 6724
rect 42760 6712 42766 6724
rect 42981 6715 43039 6721
rect 42981 6712 42993 6715
rect 42760 6684 42993 6712
rect 42760 6672 42766 6684
rect 42981 6681 42993 6684
rect 43027 6712 43039 6715
rect 43349 6715 43407 6721
rect 43349 6712 43361 6715
rect 43027 6684 43361 6712
rect 43027 6681 43039 6684
rect 42981 6675 43039 6681
rect 43349 6681 43361 6684
rect 43395 6712 43407 6715
rect 45186 6712 45192 6724
rect 43395 6684 45192 6712
rect 43395 6681 43407 6684
rect 43349 6675 43407 6681
rect 45186 6672 45192 6684
rect 45244 6712 45250 6724
rect 45281 6715 45339 6721
rect 45281 6712 45293 6715
rect 45244 6684 45293 6712
rect 45244 6672 45250 6684
rect 45281 6681 45293 6684
rect 45327 6712 45339 6715
rect 45327 6684 46980 6712
rect 45327 6681 45339 6684
rect 45281 6675 45339 6681
rect 46952 6656 46980 6684
rect 43717 6647 43775 6653
rect 43717 6644 43729 6647
rect 42628 6616 43729 6644
rect 43717 6613 43729 6616
rect 43763 6644 43775 6647
rect 44450 6644 44456 6656
rect 43763 6616 44456 6644
rect 43763 6613 43775 6616
rect 43717 6607 43775 6613
rect 44450 6604 44456 6616
rect 44508 6604 44514 6656
rect 44726 6604 44732 6656
rect 44784 6644 44790 6656
rect 45462 6644 45468 6656
rect 44784 6616 45468 6644
rect 44784 6604 44790 6616
rect 45462 6604 45468 6616
rect 45520 6644 45526 6656
rect 45925 6647 45983 6653
rect 45925 6644 45937 6647
rect 45520 6616 45937 6644
rect 45520 6604 45526 6616
rect 45925 6613 45937 6616
rect 45971 6613 45983 6647
rect 45925 6607 45983 6613
rect 46934 6604 46940 6656
rect 46992 6644 46998 6656
rect 47213 6647 47271 6653
rect 47213 6644 47225 6647
rect 46992 6616 47225 6644
rect 46992 6604 46998 6616
rect 47213 6613 47225 6616
rect 47259 6613 47271 6647
rect 47213 6607 47271 6613
rect 48222 6604 48228 6656
rect 48280 6604 48286 6656
rect 52840 6653 52868 6752
rect 53282 6740 53288 6792
rect 53340 6780 53346 6792
rect 54021 6783 54079 6789
rect 54021 6780 54033 6783
rect 53340 6752 54033 6780
rect 53340 6740 53346 6752
rect 54021 6749 54033 6752
rect 54067 6749 54079 6783
rect 54021 6743 54079 6749
rect 54573 6783 54631 6789
rect 54573 6749 54585 6783
rect 54619 6780 54631 6783
rect 56336 6780 56364 6820
rect 56410 6808 56416 6860
rect 56468 6848 56474 6860
rect 56781 6851 56839 6857
rect 56781 6848 56793 6851
rect 56468 6820 56793 6848
rect 56468 6808 56474 6820
rect 56781 6817 56793 6820
rect 56827 6817 56839 6851
rect 56781 6811 56839 6817
rect 56686 6780 56692 6792
rect 54619 6752 55812 6780
rect 56336 6752 56692 6780
rect 54619 6749 54631 6752
rect 54573 6743 54631 6749
rect 53193 6715 53251 6721
rect 53193 6681 53205 6715
rect 53239 6712 53251 6715
rect 55125 6715 55183 6721
rect 55125 6712 55137 6715
rect 53239 6684 55137 6712
rect 53239 6681 53251 6684
rect 53193 6675 53251 6681
rect 55125 6681 55137 6684
rect 55171 6681 55183 6715
rect 55125 6675 55183 6681
rect 55784 6656 55812 6752
rect 56686 6740 56692 6752
rect 56744 6740 56750 6792
rect 57330 6740 57336 6792
rect 57388 6780 57394 6792
rect 58066 6780 58072 6792
rect 57388 6752 58072 6780
rect 57388 6740 57394 6752
rect 58066 6740 58072 6752
rect 58124 6740 58130 6792
rect 58434 6740 58440 6792
rect 58492 6740 58498 6792
rect 52825 6647 52883 6653
rect 52825 6613 52837 6647
rect 52871 6613 52883 6647
rect 52825 6607 52883 6613
rect 53653 6647 53711 6653
rect 53653 6613 53665 6647
rect 53699 6644 53711 6647
rect 53926 6644 53932 6656
rect 53699 6616 53932 6644
rect 53699 6613 53711 6616
rect 53653 6607 53711 6613
rect 53926 6604 53932 6616
rect 53984 6604 53990 6656
rect 54110 6604 54116 6656
rect 54168 6604 54174 6656
rect 54202 6604 54208 6656
rect 54260 6644 54266 6656
rect 55493 6647 55551 6653
rect 55493 6644 55505 6647
rect 54260 6616 55505 6644
rect 54260 6604 54266 6616
rect 55493 6613 55505 6616
rect 55539 6613 55551 6647
rect 55493 6607 55551 6613
rect 55766 6604 55772 6656
rect 55824 6604 55830 6656
rect 56704 6644 56732 6740
rect 57048 6715 57106 6721
rect 57048 6681 57060 6715
rect 57094 6712 57106 6715
rect 58526 6712 58532 6724
rect 57094 6684 58532 6712
rect 57094 6681 57106 6684
rect 57048 6675 57106 6681
rect 58526 6672 58532 6684
rect 58584 6672 58590 6724
rect 58161 6647 58219 6653
rect 58161 6644 58173 6647
rect 56704 6616 58173 6644
rect 58161 6613 58173 6616
rect 58207 6613 58219 6647
rect 58161 6607 58219 6613
rect 58250 6604 58256 6656
rect 58308 6604 58314 6656
rect 1104 6554 59040 6576
rect 1104 6502 15394 6554
rect 15446 6502 15458 6554
rect 15510 6502 15522 6554
rect 15574 6502 15586 6554
rect 15638 6502 15650 6554
rect 15702 6502 29838 6554
rect 29890 6502 29902 6554
rect 29954 6502 29966 6554
rect 30018 6502 30030 6554
rect 30082 6502 30094 6554
rect 30146 6502 44282 6554
rect 44334 6502 44346 6554
rect 44398 6502 44410 6554
rect 44462 6502 44474 6554
rect 44526 6502 44538 6554
rect 44590 6502 58726 6554
rect 58778 6502 58790 6554
rect 58842 6502 58854 6554
rect 58906 6502 58918 6554
rect 58970 6502 58982 6554
rect 59034 6502 59040 6554
rect 1104 6480 59040 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 2590 6440 2596 6452
rect 2271 6412 2596 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 3326 6400 3332 6452
rect 3384 6400 3390 6452
rect 4430 6440 4436 6452
rect 3804 6412 4436 6440
rect 3804 6381 3832 6412
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 6788 6412 7665 6440
rect 6788 6400 6794 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 8021 6443 8079 6449
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 9858 6440 9864 6452
rect 8067 6412 9864 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 11480 6412 13032 6440
rect 11480 6400 11486 6412
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 2240 6344 3801 6372
rect 2240 6313 2268 6344
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3789 6335 3847 6341
rect 5442 6332 5448 6384
rect 5500 6332 5506 6384
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 5822 6375 5880 6381
rect 5822 6372 5834 6375
rect 5684 6344 5834 6372
rect 5684 6332 5690 6344
rect 5822 6341 5834 6344
rect 5868 6341 5880 6375
rect 5822 6335 5880 6341
rect 8754 6332 8760 6384
rect 8812 6332 8818 6384
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 10229 6375 10287 6381
rect 10229 6372 10241 6375
rect 9456 6344 10241 6372
rect 9456 6332 9462 6344
rect 10229 6341 10241 6344
rect 10275 6341 10287 6375
rect 10229 6335 10287 6341
rect 11790 6332 11796 6384
rect 11848 6372 11854 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11848 6344 11989 6372
rect 11848 6332 11854 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 13004 6372 13032 6412
rect 13078 6400 13084 6452
rect 13136 6400 13142 6452
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 15289 6443 15347 6449
rect 15289 6440 15301 6443
rect 14608 6412 15301 6440
rect 14608 6400 14614 6412
rect 15289 6409 15301 6412
rect 15335 6409 15347 6443
rect 15289 6403 15347 6409
rect 15930 6400 15936 6452
rect 15988 6400 15994 6452
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 19245 6443 19303 6449
rect 19245 6440 19257 6443
rect 18104 6412 19257 6440
rect 18104 6400 18110 6412
rect 19245 6409 19257 6412
rect 19291 6409 19303 6443
rect 19245 6403 19303 6409
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 21542 6440 21548 6452
rect 20772 6412 21548 6440
rect 20772 6400 20778 6412
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 22186 6400 22192 6452
rect 22244 6400 22250 6452
rect 24305 6443 24363 6449
rect 24305 6409 24317 6443
rect 24351 6440 24363 6443
rect 24394 6440 24400 6452
rect 24351 6412 24400 6440
rect 24351 6409 24363 6412
rect 24305 6403 24363 6409
rect 24394 6400 24400 6412
rect 24452 6440 24458 6452
rect 25590 6440 25596 6452
rect 24452 6412 25596 6440
rect 24452 6400 24458 6412
rect 25590 6400 25596 6412
rect 25648 6440 25654 6452
rect 25958 6440 25964 6452
rect 25648 6412 25964 6440
rect 25648 6400 25654 6412
rect 25958 6400 25964 6412
rect 26016 6400 26022 6452
rect 26418 6400 26424 6452
rect 26476 6440 26482 6452
rect 29362 6440 29368 6452
rect 26476 6412 29368 6440
rect 26476 6400 26482 6412
rect 29362 6400 29368 6412
rect 29420 6400 29426 6452
rect 29546 6400 29552 6452
rect 29604 6400 29610 6452
rect 30282 6400 30288 6452
rect 30340 6440 30346 6452
rect 31662 6440 31668 6452
rect 30340 6412 31668 6440
rect 30340 6400 30346 6412
rect 31662 6400 31668 6412
rect 31720 6440 31726 6452
rect 33413 6443 33471 6449
rect 33413 6440 33425 6443
rect 31720 6412 33425 6440
rect 31720 6400 31726 6412
rect 33413 6409 33425 6412
rect 33459 6440 33471 6443
rect 34422 6440 34428 6452
rect 33459 6412 34428 6440
rect 33459 6409 33471 6412
rect 33413 6403 33471 6409
rect 34422 6400 34428 6412
rect 34480 6400 34486 6452
rect 37553 6443 37611 6449
rect 37553 6409 37565 6443
rect 37599 6440 37611 6443
rect 37734 6440 37740 6452
rect 37599 6412 37740 6440
rect 37599 6409 37611 6412
rect 37553 6403 37611 6409
rect 37734 6400 37740 6412
rect 37792 6400 37798 6452
rect 39485 6443 39543 6449
rect 39485 6409 39497 6443
rect 39531 6440 39543 6443
rect 39850 6440 39856 6452
rect 39531 6412 39856 6440
rect 39531 6409 39543 6412
rect 39485 6403 39543 6409
rect 14826 6372 14832 6384
rect 13004 6344 14832 6372
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2056 6100 2084 6267
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 3234 6304 3240 6316
rect 2639 6276 3240 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6304 6147 6307
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 6135 6276 7573 6304
rect 6135 6273 6147 6276
rect 6089 6267 6147 6273
rect 7561 6273 7573 6276
rect 7607 6304 7619 6307
rect 8662 6304 8668 6316
rect 7607 6276 8668 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 2685 6239 2743 6245
rect 2685 6236 2697 6239
rect 2608 6208 2697 6236
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6168 2375 6171
rect 2608 6168 2636 6208
rect 2685 6205 2697 6208
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 3620 6168 3648 6267
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8772 6304 8800 6332
rect 9582 6304 9588 6316
rect 8772 6276 9588 6304
rect 9582 6264 9588 6276
rect 9640 6304 9646 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9640 6276 9781 6304
rect 9640 6264 9646 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 7742 6196 7748 6248
rect 7800 6236 7806 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7800 6208 8125 6236
rect 7800 6196 7806 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8251 6208 8861 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 9784 6236 9812 6267
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 13004 6304 13032 6344
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 13173 6307 13231 6313
rect 13173 6304 13185 6307
rect 13004 6276 13185 6304
rect 13173 6273 13185 6276
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 13440 6307 13498 6313
rect 13440 6273 13452 6307
rect 13486 6304 13498 6307
rect 14734 6304 14740 6316
rect 13486 6276 14740 6304
rect 13486 6273 13498 6276
rect 13440 6267 13498 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 10502 6236 10508 6248
rect 9784 6208 10508 6236
rect 8849 6199 8907 6205
rect 2363 6140 2636 6168
rect 2746 6140 3648 6168
rect 2363 6137 2375 6140
rect 2317 6131 2375 6137
rect 2222 6100 2228 6112
rect 2056 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6100 2286 6112
rect 2746 6100 2774 6140
rect 7558 6128 7564 6180
rect 7616 6168 7622 6180
rect 8018 6168 8024 6180
rect 7616 6140 8024 6168
rect 7616 6128 7622 6140
rect 8018 6128 8024 6140
rect 8076 6168 8082 6180
rect 8220 6168 8248 6199
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 12158 6196 12164 6248
rect 12216 6196 12222 6248
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6236 14703 6239
rect 15948 6236 15976 6400
rect 18874 6372 18880 6384
rect 16684 6344 18880 6372
rect 16684 6248 16712 6344
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 22830 6372 22836 6384
rect 19628 6344 22836 6372
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 19153 6307 19211 6313
rect 19153 6304 19165 6307
rect 18564 6276 19165 6304
rect 18564 6264 18570 6276
rect 19153 6273 19165 6276
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 14691 6208 15976 6236
rect 14691 6205 14703 6208
rect 14645 6199 14703 6205
rect 8076 6140 8248 6168
rect 11517 6171 11575 6177
rect 8076 6128 8082 6140
rect 11517 6137 11529 6171
rect 11563 6168 11575 6171
rect 12452 6168 12480 6199
rect 11563 6140 12480 6168
rect 14553 6171 14611 6177
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 14553 6137 14565 6171
rect 14599 6168 14611 6171
rect 14660 6168 14688 6199
rect 16666 6196 16672 6248
rect 16724 6196 16730 6248
rect 19426 6236 19432 6248
rect 17420 6208 19432 6236
rect 17420 6168 17448 6208
rect 19426 6196 19432 6208
rect 19484 6236 19490 6248
rect 19628 6245 19656 6344
rect 22830 6332 22836 6344
rect 22888 6332 22894 6384
rect 32398 6332 32404 6384
rect 32456 6372 32462 6384
rect 32769 6375 32827 6381
rect 32769 6372 32781 6375
rect 32456 6344 32781 6372
rect 32456 6332 32462 6344
rect 32769 6341 32781 6344
rect 32815 6341 32827 6375
rect 32769 6335 32827 6341
rect 33318 6332 33324 6384
rect 33376 6372 33382 6384
rect 34054 6372 34060 6384
rect 33376 6344 34060 6372
rect 33376 6332 33382 6344
rect 34054 6332 34060 6344
rect 34112 6372 34118 6384
rect 34149 6375 34207 6381
rect 34149 6372 34161 6375
rect 34112 6344 34161 6372
rect 34112 6332 34118 6344
rect 34149 6341 34161 6344
rect 34195 6341 34207 6375
rect 34149 6335 34207 6341
rect 35066 6332 35072 6384
rect 35124 6372 35130 6384
rect 35713 6375 35771 6381
rect 35713 6372 35725 6375
rect 35124 6344 35725 6372
rect 35124 6332 35130 6344
rect 35713 6341 35725 6344
rect 35759 6372 35771 6375
rect 39500 6372 39528 6403
rect 39850 6400 39856 6412
rect 39908 6400 39914 6452
rect 40218 6400 40224 6452
rect 40276 6440 40282 6452
rect 40957 6443 41015 6449
rect 40957 6440 40969 6443
rect 40276 6412 40969 6440
rect 40276 6400 40282 6412
rect 40957 6409 40969 6412
rect 41003 6409 41015 6443
rect 40957 6403 41015 6409
rect 41230 6400 41236 6452
rect 41288 6440 41294 6452
rect 41325 6443 41383 6449
rect 41325 6440 41337 6443
rect 41288 6412 41337 6440
rect 41288 6400 41294 6412
rect 41325 6409 41337 6412
rect 41371 6409 41383 6443
rect 41325 6403 41383 6409
rect 41506 6400 41512 6452
rect 41564 6440 41570 6452
rect 42153 6443 42211 6449
rect 41564 6412 41736 6440
rect 41564 6400 41570 6412
rect 35759 6344 39528 6372
rect 35759 6341 35771 6344
rect 35713 6335 35771 6341
rect 40494 6332 40500 6384
rect 40552 6372 40558 6384
rect 41598 6372 41604 6384
rect 40552 6344 41604 6372
rect 40552 6332 40558 6344
rect 41598 6332 41604 6344
rect 41656 6332 41662 6384
rect 20714 6264 20720 6316
rect 20772 6264 20778 6316
rect 23106 6304 23112 6316
rect 22848 6276 23112 6304
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19484 6208 19625 6236
rect 19484 6196 19490 6208
rect 19613 6205 19625 6208
rect 19659 6205 19671 6239
rect 19613 6199 19671 6205
rect 19702 6196 19708 6248
rect 19760 6236 19766 6248
rect 19797 6239 19855 6245
rect 19797 6236 19809 6239
rect 19760 6208 19809 6236
rect 19760 6196 19766 6208
rect 19797 6205 19809 6208
rect 19843 6205 19855 6239
rect 19797 6199 19855 6205
rect 20533 6239 20591 6245
rect 20533 6205 20545 6239
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 14599 6140 14688 6168
rect 15580 6140 17448 6168
rect 14599 6137 14611 6140
rect 14553 6131 14611 6137
rect 2280 6072 2774 6100
rect 2280 6060 2286 6072
rect 3970 6060 3976 6112
rect 4028 6060 4034 6112
rect 5166 6060 5172 6112
rect 5224 6100 5230 6112
rect 5813 6103 5871 6109
rect 5813 6100 5825 6103
rect 5224 6072 5825 6100
rect 5224 6060 5230 6072
rect 5813 6069 5825 6072
rect 5859 6069 5871 6103
rect 5813 6063 5871 6069
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15580 6109 15608 6140
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 20070 6168 20076 6180
rect 17828 6140 20076 6168
rect 17828 6128 17834 6140
rect 20070 6128 20076 6140
rect 20128 6168 20134 6180
rect 20548 6168 20576 6199
rect 22848 6177 22876 6276
rect 23106 6264 23112 6276
rect 23164 6304 23170 6316
rect 24581 6307 24639 6313
rect 24581 6304 24593 6307
rect 23164 6276 24593 6304
rect 23164 6264 23170 6276
rect 24581 6273 24593 6276
rect 24627 6273 24639 6307
rect 24581 6267 24639 6273
rect 27801 6307 27859 6313
rect 27801 6273 27813 6307
rect 27847 6304 27859 6307
rect 27890 6304 27896 6316
rect 27847 6276 27896 6304
rect 27847 6273 27859 6276
rect 27801 6267 27859 6273
rect 27890 6264 27896 6276
rect 27948 6264 27954 6316
rect 28068 6307 28126 6313
rect 28068 6273 28080 6307
rect 28114 6304 28126 6307
rect 28902 6304 28908 6316
rect 28114 6276 28908 6304
rect 28114 6273 28126 6276
rect 28068 6267 28126 6273
rect 28902 6264 28908 6276
rect 28960 6264 28966 6316
rect 29730 6264 29736 6316
rect 29788 6304 29794 6316
rect 29917 6307 29975 6313
rect 29917 6304 29929 6307
rect 29788 6276 29929 6304
rect 29788 6264 29794 6276
rect 29917 6273 29929 6276
rect 29963 6273 29975 6307
rect 29917 6267 29975 6273
rect 30024 6276 30236 6304
rect 24394 6196 24400 6248
rect 24452 6196 24458 6248
rect 25041 6239 25099 6245
rect 25041 6205 25053 6239
rect 25087 6236 25099 6239
rect 25130 6236 25136 6248
rect 25087 6208 25136 6236
rect 25087 6205 25099 6208
rect 25041 6199 25099 6205
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 25409 6239 25467 6245
rect 25409 6205 25421 6239
rect 25455 6205 25467 6239
rect 25409 6199 25467 6205
rect 21177 6171 21235 6177
rect 21177 6168 21189 6171
rect 20128 6140 21189 6168
rect 20128 6128 20134 6140
rect 21177 6137 21189 6140
rect 21223 6137 21235 6171
rect 22833 6171 22891 6177
rect 22833 6168 22845 6171
rect 21177 6131 21235 6137
rect 22296 6140 22845 6168
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 14700 6072 15577 6100
rect 14700 6060 14706 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 16758 6100 16764 6112
rect 15712 6072 16764 6100
rect 15712 6060 15718 6072
rect 16758 6060 16764 6072
rect 16816 6100 16822 6112
rect 16853 6103 16911 6109
rect 16853 6100 16865 6103
rect 16816 6072 16865 6100
rect 16816 6060 16822 6072
rect 16853 6069 16865 6072
rect 16899 6069 16911 6103
rect 16853 6063 16911 6069
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 18509 6103 18567 6109
rect 18509 6100 18521 6103
rect 17000 6072 18521 6100
rect 17000 6060 17006 6072
rect 18509 6069 18521 6072
rect 18555 6100 18567 6103
rect 19334 6100 19340 6112
rect 18555 6072 19340 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20441 6103 20499 6109
rect 20441 6100 20453 6103
rect 19852 6072 20453 6100
rect 19852 6060 19858 6072
rect 20441 6069 20453 6072
rect 20487 6069 20499 6103
rect 20441 6063 20499 6069
rect 20898 6060 20904 6112
rect 20956 6060 20962 6112
rect 21192 6100 21220 6131
rect 22296 6100 22324 6140
rect 22833 6137 22845 6140
rect 22879 6137 22891 6171
rect 24412 6168 24440 6196
rect 25424 6168 25452 6199
rect 24412 6140 25452 6168
rect 29181 6171 29239 6177
rect 22833 6131 22891 6137
rect 29181 6137 29193 6171
rect 29227 6168 29239 6171
rect 29638 6168 29644 6180
rect 29227 6140 29644 6168
rect 29227 6137 29239 6140
rect 29181 6131 29239 6137
rect 29638 6128 29644 6140
rect 29696 6168 29702 6180
rect 30024 6168 30052 6276
rect 30101 6239 30159 6245
rect 30101 6205 30113 6239
rect 30147 6205 30159 6239
rect 30208 6236 30236 6276
rect 30834 6264 30840 6316
rect 30892 6264 30898 6316
rect 33502 6264 33508 6316
rect 33560 6304 33566 6316
rect 33965 6307 34023 6313
rect 33965 6304 33977 6307
rect 33560 6276 33977 6304
rect 33560 6264 33566 6276
rect 33965 6273 33977 6276
rect 34011 6273 34023 6307
rect 33965 6267 34023 6273
rect 34882 6264 34888 6316
rect 34940 6304 34946 6316
rect 36173 6307 36231 6313
rect 36173 6304 36185 6307
rect 34940 6276 36185 6304
rect 34940 6264 34946 6276
rect 36173 6273 36185 6276
rect 36219 6273 36231 6307
rect 40678 6304 40684 6316
rect 36173 6267 36231 6273
rect 37844 6276 40684 6304
rect 30954 6239 31012 6245
rect 30954 6236 30966 6239
rect 30208 6208 30966 6236
rect 30101 6199 30159 6205
rect 30954 6205 30966 6208
rect 31000 6205 31012 6239
rect 30954 6199 31012 6205
rect 31113 6239 31171 6245
rect 31113 6205 31125 6239
rect 31159 6236 31171 6239
rect 31478 6236 31484 6248
rect 31159 6208 31484 6236
rect 31159 6205 31171 6208
rect 31113 6199 31171 6205
rect 29696 6140 30052 6168
rect 29696 6128 29702 6140
rect 21192 6072 22324 6100
rect 22370 6060 22376 6112
rect 22428 6100 22434 6112
rect 22465 6103 22523 6109
rect 22465 6100 22477 6103
rect 22428 6072 22477 6100
rect 22428 6060 22434 6072
rect 22465 6069 22477 6072
rect 22511 6069 22523 6103
rect 22465 6063 22523 6069
rect 23382 6060 23388 6112
rect 23440 6100 23446 6112
rect 24118 6100 24124 6112
rect 23440 6072 24124 6100
rect 23440 6060 23446 6072
rect 24118 6060 24124 6072
rect 24176 6060 24182 6112
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 26053 6103 26111 6109
rect 26053 6100 26065 6103
rect 25096 6072 26065 6100
rect 25096 6060 25102 6072
rect 26053 6069 26065 6072
rect 26099 6069 26111 6103
rect 26053 6063 26111 6069
rect 26142 6060 26148 6112
rect 26200 6100 26206 6112
rect 30006 6100 30012 6112
rect 26200 6072 30012 6100
rect 26200 6060 26206 6072
rect 30006 6060 30012 6072
rect 30064 6060 30070 6112
rect 30116 6100 30144 6199
rect 31478 6196 31484 6208
rect 31536 6196 31542 6248
rect 31938 6236 31944 6248
rect 31588 6208 31944 6236
rect 30558 6128 30564 6180
rect 30616 6128 30622 6180
rect 31588 6100 31616 6208
rect 31938 6196 31944 6208
rect 31996 6236 32002 6248
rect 32125 6239 32183 6245
rect 32125 6236 32137 6239
rect 31996 6208 32137 6236
rect 31996 6196 32002 6208
rect 32125 6205 32137 6208
rect 32171 6205 32183 6239
rect 34974 6236 34980 6248
rect 32125 6199 32183 6205
rect 34440 6208 34980 6236
rect 30116 6072 31616 6100
rect 31754 6060 31760 6112
rect 31812 6060 31818 6112
rect 32950 6060 32956 6112
rect 33008 6100 33014 6112
rect 34440 6109 34468 6208
rect 34974 6196 34980 6208
rect 35032 6236 35038 6248
rect 35618 6236 35624 6248
rect 35032 6208 35624 6236
rect 35032 6196 35038 6208
rect 35618 6196 35624 6208
rect 35676 6236 35682 6248
rect 37844 6245 37872 6276
rect 40678 6264 40684 6276
rect 40736 6264 40742 6316
rect 40865 6307 40923 6313
rect 40865 6273 40877 6307
rect 40911 6304 40923 6307
rect 41506 6304 41512 6316
rect 40911 6276 41512 6304
rect 40911 6273 40923 6276
rect 40865 6267 40923 6273
rect 41506 6264 41512 6276
rect 41564 6264 41570 6316
rect 41708 6304 41736 6412
rect 42153 6409 42165 6443
rect 42199 6440 42211 6443
rect 42702 6440 42708 6452
rect 42199 6412 42708 6440
rect 42199 6409 42211 6412
rect 42153 6403 42211 6409
rect 42702 6400 42708 6412
rect 42760 6440 42766 6452
rect 42981 6443 43039 6449
rect 42981 6440 42993 6443
rect 42760 6412 42993 6440
rect 42760 6400 42766 6412
rect 42981 6409 42993 6412
rect 43027 6440 43039 6443
rect 43349 6443 43407 6449
rect 43349 6440 43361 6443
rect 43027 6412 43361 6440
rect 43027 6409 43039 6412
rect 42981 6403 43039 6409
rect 43349 6409 43361 6412
rect 43395 6409 43407 6443
rect 43349 6403 43407 6409
rect 45462 6400 45468 6452
rect 45520 6440 45526 6452
rect 46017 6443 46075 6449
rect 46017 6440 46029 6443
rect 45520 6412 46029 6440
rect 45520 6400 45526 6412
rect 46017 6409 46029 6412
rect 46063 6409 46075 6443
rect 46017 6403 46075 6409
rect 48590 6400 48596 6452
rect 48648 6440 48654 6452
rect 48869 6443 48927 6449
rect 48869 6440 48881 6443
rect 48648 6412 48881 6440
rect 48648 6400 48654 6412
rect 48869 6409 48881 6412
rect 48915 6440 48927 6443
rect 49142 6440 49148 6452
rect 48915 6412 49148 6440
rect 48915 6409 48927 6412
rect 48869 6403 48927 6409
rect 49142 6400 49148 6412
rect 49200 6440 49206 6452
rect 49237 6443 49295 6449
rect 49237 6440 49249 6443
rect 49200 6412 49249 6440
rect 49200 6400 49206 6412
rect 49237 6409 49249 6412
rect 49283 6409 49295 6443
rect 49237 6403 49295 6409
rect 51169 6443 51227 6449
rect 51169 6409 51181 6443
rect 51215 6440 51227 6443
rect 51537 6443 51595 6449
rect 51537 6440 51549 6443
rect 51215 6412 51549 6440
rect 51215 6409 51227 6412
rect 51169 6403 51227 6409
rect 51537 6409 51549 6412
rect 51583 6440 51595 6443
rect 52178 6440 52184 6452
rect 51583 6412 52184 6440
rect 51583 6409 51595 6412
rect 51537 6403 51595 6409
rect 52178 6400 52184 6412
rect 52236 6400 52242 6452
rect 53742 6400 53748 6452
rect 53800 6440 53806 6452
rect 54481 6443 54539 6449
rect 54481 6440 54493 6443
rect 53800 6412 54493 6440
rect 53800 6400 53806 6412
rect 54481 6409 54493 6412
rect 54527 6440 54539 6443
rect 56870 6440 56876 6452
rect 54527 6412 56876 6440
rect 54527 6409 54539 6412
rect 54481 6403 54539 6409
rect 56870 6400 56876 6412
rect 56928 6400 56934 6452
rect 46106 6332 46112 6384
rect 46164 6372 46170 6384
rect 49878 6372 49884 6384
rect 46164 6344 49884 6372
rect 46164 6332 46170 6344
rect 49878 6332 49884 6344
rect 49936 6332 49942 6384
rect 51626 6332 51632 6384
rect 51684 6332 51690 6384
rect 52822 6332 52828 6384
rect 52880 6372 52886 6384
rect 52978 6375 53036 6381
rect 52978 6372 52990 6375
rect 52880 6344 52990 6372
rect 52880 6332 52886 6344
rect 52978 6341 52990 6344
rect 53024 6341 53036 6375
rect 52978 6335 53036 6341
rect 41708 6276 43760 6304
rect 37829 6239 37887 6245
rect 37829 6236 37841 6239
rect 35676 6208 37841 6236
rect 35676 6196 35682 6208
rect 37829 6205 37841 6208
rect 37875 6205 37887 6239
rect 37829 6199 37887 6205
rect 38562 6196 38568 6248
rect 38620 6196 38626 6248
rect 40126 6196 40132 6248
rect 40184 6236 40190 6248
rect 42613 6239 42671 6245
rect 42613 6236 42625 6239
rect 40184 6208 42625 6236
rect 40184 6196 40190 6208
rect 42613 6205 42625 6208
rect 42659 6205 42671 6239
rect 43732 6236 43760 6276
rect 45554 6264 45560 6316
rect 45612 6304 45618 6316
rect 45925 6307 45983 6313
rect 45925 6304 45937 6307
rect 45612 6276 45937 6304
rect 45612 6264 45618 6276
rect 45925 6273 45937 6276
rect 45971 6273 45983 6307
rect 45925 6267 45983 6273
rect 48222 6264 48228 6316
rect 48280 6304 48286 6316
rect 48280 6276 50016 6304
rect 48280 6264 48286 6276
rect 43898 6236 43904 6248
rect 43732 6208 43904 6236
rect 42613 6199 42671 6205
rect 43898 6196 43904 6208
rect 43956 6236 43962 6248
rect 44177 6239 44235 6245
rect 44177 6236 44189 6239
rect 43956 6208 44189 6236
rect 43956 6196 43962 6208
rect 44177 6205 44189 6208
rect 44223 6205 44235 6239
rect 44177 6199 44235 6205
rect 44910 6196 44916 6248
rect 44968 6196 44974 6248
rect 47118 6196 47124 6248
rect 47176 6196 47182 6248
rect 49602 6196 49608 6248
rect 49660 6196 49666 6248
rect 49988 6236 50016 6276
rect 50062 6264 50068 6316
rect 50120 6304 50126 6316
rect 51644 6304 51672 6332
rect 50120 6276 51672 6304
rect 52365 6307 52423 6313
rect 50120 6264 50126 6276
rect 52365 6273 52377 6307
rect 52411 6304 52423 6307
rect 52411 6276 52500 6304
rect 52411 6273 52423 6276
rect 52365 6267 52423 6273
rect 52089 6239 52147 6245
rect 52089 6236 52101 6239
rect 49988 6208 52101 6236
rect 52089 6205 52101 6208
rect 52135 6236 52147 6239
rect 52270 6236 52276 6248
rect 52135 6208 52276 6236
rect 52135 6205 52147 6208
rect 52089 6199 52147 6205
rect 52270 6196 52276 6208
rect 52328 6196 52334 6248
rect 36541 6171 36599 6177
rect 36541 6168 36553 6171
rect 34716 6140 36553 6168
rect 34716 6112 34744 6140
rect 36541 6137 36553 6140
rect 36587 6137 36599 6171
rect 38194 6168 38200 6180
rect 36541 6131 36599 6137
rect 36648 6140 38200 6168
rect 33045 6103 33103 6109
rect 33045 6100 33057 6103
rect 33008 6072 33057 6100
rect 33008 6060 33014 6072
rect 33045 6069 33057 6072
rect 33091 6100 33103 6103
rect 34425 6103 34483 6109
rect 34425 6100 34437 6103
rect 33091 6072 34437 6100
rect 33091 6069 33103 6072
rect 33045 6063 33103 6069
rect 34425 6069 34437 6072
rect 34471 6069 34483 6103
rect 34425 6063 34483 6069
rect 34698 6060 34704 6112
rect 34756 6060 34762 6112
rect 35158 6060 35164 6112
rect 35216 6100 35222 6112
rect 35526 6100 35532 6112
rect 35216 6072 35532 6100
rect 35216 6060 35222 6072
rect 35526 6060 35532 6072
rect 35584 6100 35590 6112
rect 36648 6100 36676 6140
rect 38194 6128 38200 6140
rect 38252 6128 38258 6180
rect 41230 6168 41236 6180
rect 38396 6140 41236 6168
rect 38396 6112 38424 6140
rect 41230 6128 41236 6140
rect 41288 6168 41294 6180
rect 42334 6168 42340 6180
rect 41288 6140 42340 6168
rect 41288 6128 41294 6140
rect 42334 6128 42340 6140
rect 42392 6168 42398 6180
rect 46845 6171 46903 6177
rect 42392 6140 45692 6168
rect 42392 6128 42398 6140
rect 45664 6112 45692 6140
rect 46845 6137 46857 6171
rect 46891 6168 46903 6171
rect 46934 6168 46940 6180
rect 46891 6140 46940 6168
rect 46891 6137 46903 6140
rect 46845 6131 46903 6137
rect 46934 6128 46940 6140
rect 46992 6168 46998 6180
rect 47857 6171 47915 6177
rect 47857 6168 47869 6171
rect 46992 6140 47869 6168
rect 46992 6128 46998 6140
rect 47857 6137 47869 6140
rect 47903 6168 47915 6171
rect 48225 6171 48283 6177
rect 48225 6168 48237 6171
rect 47903 6140 48237 6168
rect 47903 6137 47915 6140
rect 47857 6131 47915 6137
rect 48225 6137 48237 6140
rect 48271 6168 48283 6171
rect 48593 6171 48651 6177
rect 48593 6168 48605 6171
rect 48271 6140 48605 6168
rect 48271 6137 48283 6140
rect 48225 6131 48283 6137
rect 48593 6137 48605 6140
rect 48639 6168 48651 6171
rect 48639 6140 50568 6168
rect 48639 6137 48651 6140
rect 48593 6131 48651 6137
rect 50540 6112 50568 6140
rect 35584 6072 36676 6100
rect 35584 6060 35590 6072
rect 36722 6060 36728 6112
rect 36780 6100 36786 6112
rect 36909 6103 36967 6109
rect 36909 6100 36921 6103
rect 36780 6072 36921 6100
rect 36780 6060 36786 6072
rect 36909 6069 36921 6072
rect 36955 6069 36967 6103
rect 36909 6063 36967 6069
rect 38378 6060 38384 6112
rect 38436 6060 38442 6112
rect 39114 6060 39120 6112
rect 39172 6060 39178 6112
rect 39853 6103 39911 6109
rect 39853 6069 39865 6103
rect 39899 6100 39911 6103
rect 39942 6100 39948 6112
rect 39899 6072 39948 6100
rect 39899 6069 39911 6072
rect 39853 6063 39911 6069
rect 39942 6060 39948 6072
rect 40000 6060 40006 6112
rect 40221 6103 40279 6109
rect 40221 6069 40233 6103
rect 40267 6100 40279 6103
rect 40589 6103 40647 6109
rect 40589 6100 40601 6103
rect 40267 6072 40601 6100
rect 40267 6069 40279 6072
rect 40221 6063 40279 6069
rect 40589 6069 40601 6072
rect 40635 6100 40647 6103
rect 41322 6100 41328 6112
rect 40635 6072 41328 6100
rect 40635 6069 40647 6072
rect 40589 6063 40647 6069
rect 41322 6060 41328 6072
rect 41380 6100 41386 6112
rect 41693 6103 41751 6109
rect 41693 6100 41705 6103
rect 41380 6072 41705 6100
rect 41380 6060 41386 6072
rect 41693 6069 41705 6072
rect 41739 6100 41751 6103
rect 42610 6100 42616 6112
rect 41739 6072 42616 6100
rect 41739 6069 41751 6072
rect 41693 6063 41751 6069
rect 42610 6060 42616 6072
rect 42668 6100 42674 6112
rect 43717 6103 43775 6109
rect 43717 6100 43729 6103
rect 42668 6072 43729 6100
rect 42668 6060 42674 6072
rect 43717 6069 43729 6072
rect 43763 6100 43775 6103
rect 44453 6103 44511 6109
rect 44453 6100 44465 6103
rect 43763 6072 44465 6100
rect 43763 6069 43775 6072
rect 43717 6063 43775 6069
rect 44453 6069 44465 6072
rect 44499 6069 44511 6103
rect 44453 6063 44511 6069
rect 45462 6060 45468 6112
rect 45520 6060 45526 6112
rect 45646 6060 45652 6112
rect 45704 6100 45710 6112
rect 46477 6103 46535 6109
rect 46477 6100 46489 6103
rect 45704 6072 46489 6100
rect 45704 6060 45710 6072
rect 46477 6069 46489 6072
rect 46523 6100 46535 6103
rect 48866 6100 48872 6112
rect 46523 6072 48872 6100
rect 46523 6069 46535 6072
rect 46477 6063 46535 6069
rect 48866 6060 48872 6072
rect 48924 6100 48930 6112
rect 50338 6100 50344 6112
rect 48924 6072 50344 6100
rect 48924 6060 48930 6072
rect 50338 6060 50344 6072
rect 50396 6060 50402 6112
rect 50522 6060 50528 6112
rect 50580 6100 50586 6112
rect 50709 6103 50767 6109
rect 50709 6100 50721 6103
rect 50580 6072 50721 6100
rect 50580 6060 50586 6072
rect 50709 6069 50721 6072
rect 50755 6069 50767 6103
rect 52472 6100 52500 6276
rect 52546 6264 52552 6316
rect 52604 6304 52610 6316
rect 52733 6307 52791 6313
rect 52733 6304 52745 6307
rect 52604 6276 52745 6304
rect 52604 6264 52610 6276
rect 52733 6273 52745 6276
rect 52779 6273 52791 6307
rect 52733 6267 52791 6273
rect 54938 6264 54944 6316
rect 54996 6264 55002 6316
rect 55766 6264 55772 6316
rect 55824 6313 55830 6316
rect 55824 6307 55852 6313
rect 55840 6273 55852 6307
rect 55824 6267 55852 6273
rect 55824 6264 55830 6267
rect 56778 6264 56784 6316
rect 56836 6304 56842 6316
rect 57057 6307 57115 6313
rect 57057 6304 57069 6307
rect 56836 6276 57069 6304
rect 56836 6264 56842 6276
rect 57057 6273 57069 6276
rect 57103 6273 57115 6307
rect 57057 6267 57115 6273
rect 57701 6307 57759 6313
rect 57701 6273 57713 6307
rect 57747 6304 57759 6307
rect 57790 6304 57796 6316
rect 57747 6276 57796 6304
rect 57747 6273 57759 6276
rect 57701 6267 57759 6273
rect 57790 6264 57796 6276
rect 57848 6264 57854 6316
rect 54757 6239 54815 6245
rect 54757 6205 54769 6239
rect 54803 6205 54815 6239
rect 54757 6199 54815 6205
rect 52549 6171 52607 6177
rect 52549 6137 52561 6171
rect 52595 6168 52607 6171
rect 52730 6168 52736 6180
rect 52595 6140 52736 6168
rect 52595 6137 52607 6140
rect 52549 6131 52607 6137
rect 52730 6128 52736 6140
rect 52788 6128 52794 6180
rect 54772 6168 54800 6199
rect 55030 6196 55036 6248
rect 55088 6236 55094 6248
rect 55677 6239 55735 6245
rect 55677 6236 55689 6239
rect 55088 6208 55689 6236
rect 55088 6196 55094 6208
rect 55677 6205 55689 6208
rect 55723 6205 55735 6239
rect 55677 6199 55735 6205
rect 55953 6239 56011 6245
rect 55953 6205 55965 6239
rect 55999 6236 56011 6239
rect 56134 6236 56140 6248
rect 55999 6208 56140 6236
rect 55999 6205 56011 6208
rect 55953 6199 56011 6205
rect 56134 6196 56140 6208
rect 56192 6196 56198 6248
rect 56594 6236 56600 6248
rect 56520 6208 56600 6236
rect 55306 6168 55312 6180
rect 54772 6140 55312 6168
rect 55306 6128 55312 6140
rect 55364 6128 55370 6180
rect 55398 6128 55404 6180
rect 55456 6128 55462 6180
rect 54018 6100 54024 6112
rect 52472 6072 54024 6100
rect 50709 6063 50767 6069
rect 54018 6060 54024 6072
rect 54076 6060 54082 6112
rect 54113 6103 54171 6109
rect 54113 6069 54125 6103
rect 54159 6100 54171 6103
rect 55766 6100 55772 6112
rect 54159 6072 55772 6100
rect 54159 6069 54171 6072
rect 54113 6063 54171 6069
rect 55766 6060 55772 6072
rect 55824 6060 55830 6112
rect 55858 6060 55864 6112
rect 55916 6100 55922 6112
rect 56520 6100 56548 6208
rect 56594 6196 56600 6208
rect 56652 6196 56658 6248
rect 57146 6196 57152 6248
rect 57204 6196 57210 6248
rect 57238 6196 57244 6248
rect 57296 6196 57302 6248
rect 57885 6239 57943 6245
rect 57885 6205 57897 6239
rect 57931 6205 57943 6239
rect 57885 6199 57943 6205
rect 56689 6171 56747 6177
rect 56689 6137 56701 6171
rect 56735 6168 56747 6171
rect 57900 6168 57928 6199
rect 56735 6140 57928 6168
rect 56735 6137 56747 6140
rect 56689 6131 56747 6137
rect 55916 6072 56548 6100
rect 55916 6060 55922 6072
rect 56594 6060 56600 6112
rect 56652 6060 56658 6112
rect 57514 6060 57520 6112
rect 57572 6060 57578 6112
rect 58529 6103 58587 6109
rect 58529 6069 58541 6103
rect 58575 6100 58587 6103
rect 58575 6072 58940 6100
rect 58575 6069 58587 6072
rect 58529 6063 58587 6069
rect 1104 6010 58880 6032
rect 1104 5958 8172 6010
rect 8224 5958 8236 6010
rect 8288 5958 8300 6010
rect 8352 5958 8364 6010
rect 8416 5958 8428 6010
rect 8480 5958 22616 6010
rect 22668 5958 22680 6010
rect 22732 5958 22744 6010
rect 22796 5958 22808 6010
rect 22860 5958 22872 6010
rect 22924 5958 37060 6010
rect 37112 5958 37124 6010
rect 37176 5958 37188 6010
rect 37240 5958 37252 6010
rect 37304 5958 37316 6010
rect 37368 5958 51504 6010
rect 51556 5958 51568 6010
rect 51620 5958 51632 6010
rect 51684 5958 51696 6010
rect 51748 5958 51760 6010
rect 51812 5958 58880 6010
rect 1104 5936 58880 5958
rect 2498 5856 2504 5908
rect 2556 5856 2562 5908
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5261 5899 5319 5905
rect 5261 5896 5273 5899
rect 5224 5868 5273 5896
rect 5224 5856 5230 5868
rect 5261 5865 5273 5868
rect 5307 5865 5319 5899
rect 5261 5859 5319 5865
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 8076 5868 8493 5896
rect 8076 5856 8082 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 9582 5856 9588 5908
rect 9640 5856 9646 5908
rect 9674 5856 9680 5908
rect 9732 5856 9738 5908
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 11333 5899 11391 5905
rect 11333 5896 11345 5899
rect 10836 5868 11345 5896
rect 10836 5856 10842 5868
rect 11333 5865 11345 5868
rect 11379 5865 11391 5899
rect 11333 5859 11391 5865
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 11940 5868 12357 5896
rect 11940 5856 11946 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 12802 5856 12808 5908
rect 12860 5856 12866 5908
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 13538 5896 13544 5908
rect 13127 5868 13544 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 14734 5856 14740 5908
rect 14792 5856 14798 5908
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 17678 5896 17684 5908
rect 15160 5868 17684 5896
rect 15160 5856 15166 5868
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 17770 5856 17776 5908
rect 17828 5856 17834 5908
rect 22370 5856 22376 5908
rect 22428 5896 22434 5908
rect 22646 5896 22652 5908
rect 22428 5868 22652 5896
rect 22428 5856 22434 5868
rect 22646 5856 22652 5868
rect 22704 5896 22710 5908
rect 26142 5896 26148 5908
rect 22704 5868 26148 5896
rect 22704 5856 22710 5868
rect 26142 5856 26148 5868
rect 26200 5856 26206 5908
rect 28258 5856 28264 5908
rect 28316 5856 28322 5908
rect 29546 5856 29552 5908
rect 29604 5856 29610 5908
rect 30837 5899 30895 5905
rect 30837 5865 30849 5899
rect 30883 5896 30895 5899
rect 32858 5896 32864 5908
rect 30883 5868 31616 5896
rect 30883 5865 30895 5868
rect 30837 5859 30895 5865
rect 2516 5692 2544 5856
rect 3988 5760 4016 5856
rect 8570 5828 8576 5840
rect 4356 5800 8576 5828
rect 4356 5769 4384 5800
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 3804 5732 4016 5760
rect 4341 5763 4399 5769
rect 3804 5701 3832 5732
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 9692 5760 9720 5856
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 12621 5831 12679 5837
rect 12621 5828 12633 5831
rect 12216 5800 12633 5828
rect 12216 5788 12222 5800
rect 12621 5797 12633 5800
rect 12667 5797 12679 5831
rect 12621 5791 12679 5797
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 5224 5732 6316 5760
rect 9692 5732 11713 5760
rect 5224 5720 5230 5732
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 2516 5664 3801 5692
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 3878 5652 3884 5704
rect 3936 5692 3942 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3936 5664 3985 5692
rect 3936 5652 3942 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 5626 5692 5632 5704
rect 3973 5655 4031 5661
rect 5000 5664 5632 5692
rect 2590 5584 2596 5636
rect 2648 5624 2654 5636
rect 2685 5627 2743 5633
rect 2685 5624 2697 5627
rect 2648 5596 2697 5624
rect 2648 5584 2654 5596
rect 2685 5593 2697 5596
rect 2731 5593 2743 5627
rect 2685 5587 2743 5593
rect 2869 5627 2927 5633
rect 2869 5593 2881 5627
rect 2915 5624 2927 5627
rect 3326 5624 3332 5636
rect 2915 5596 3332 5624
rect 2915 5593 2927 5596
rect 2869 5587 2927 5593
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 3050 5516 3056 5568
rect 3108 5516 3114 5568
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 5000 5556 5028 5664
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 6288 5701 6316 5732
rect 11701 5729 11713 5732
rect 11747 5760 11759 5763
rect 12820 5760 12848 5856
rect 11747 5732 12848 5760
rect 11747 5729 11759 5732
rect 11701 5723 11759 5729
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 10686 5692 10692 5704
rect 6963 5664 10692 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 5077 5627 5135 5633
rect 5077 5593 5089 5627
rect 5123 5624 5135 5627
rect 5534 5624 5540 5636
rect 5123 5596 5540 5624
rect 5123 5593 5135 5596
rect 5077 5587 5135 5593
rect 5534 5584 5540 5596
rect 5592 5624 5598 5636
rect 5828 5624 5856 5655
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 13556 5692 13584 5856
rect 14108 5769 14136 5856
rect 14936 5828 14964 5856
rect 14936 5800 20300 5828
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15838 5760 15844 5772
rect 15519 5732 15844 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 16942 5760 16948 5772
rect 16316 5732 16948 5760
rect 16316 5692 16344 5732
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 19426 5720 19432 5772
rect 19484 5720 19490 5772
rect 19794 5720 19800 5772
rect 19852 5720 19858 5772
rect 19889 5763 19947 5769
rect 19889 5729 19901 5763
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 13556 5664 16344 5692
rect 16390 5652 16396 5704
rect 16448 5692 16454 5704
rect 16485 5695 16543 5701
rect 16485 5692 16497 5695
rect 16448 5664 16497 5692
rect 16448 5652 16454 5664
rect 16485 5661 16497 5664
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17828 5664 17877 5692
rect 17828 5652 17834 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18138 5692 18144 5704
rect 18095 5664 18144 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 19444 5692 19472 5720
rect 19904 5692 19932 5723
rect 18555 5664 19380 5692
rect 19444 5664 19932 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 5592 5596 5856 5624
rect 8205 5627 8263 5633
rect 5592 5584 5598 5596
rect 8205 5593 8217 5627
rect 8251 5624 8263 5627
rect 8846 5624 8852 5636
rect 8251 5596 8852 5624
rect 8251 5593 8263 5596
rect 8205 5587 8263 5593
rect 8846 5584 8852 5596
rect 8904 5624 8910 5636
rect 9306 5624 9312 5636
rect 8904 5596 9312 5624
rect 8904 5584 8910 5596
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 9766 5624 9772 5636
rect 9416 5596 9772 5624
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 4672 5528 5273 5556
rect 4672 5516 4678 5528
rect 5261 5525 5273 5528
rect 5307 5525 5319 5559
rect 5261 5519 5319 5525
rect 5445 5559 5503 5565
rect 5445 5525 5457 5559
rect 5491 5556 5503 5559
rect 6178 5556 6184 5568
rect 5491 5528 6184 5556
rect 5491 5525 5503 5528
rect 5445 5519 5503 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 7892 5528 9229 5556
rect 7892 5516 7898 5528
rect 9217 5525 9229 5528
rect 9263 5556 9275 5559
rect 9416 5556 9444 5596
rect 9766 5584 9772 5596
rect 9824 5624 9830 5636
rect 10134 5624 10140 5636
rect 9824 5596 10140 5624
rect 9824 5584 9830 5596
rect 10134 5584 10140 5596
rect 10192 5624 10198 5636
rect 15105 5627 15163 5633
rect 15105 5624 15117 5627
rect 10192 5596 15117 5624
rect 10192 5584 10198 5596
rect 15105 5593 15117 5596
rect 15151 5624 15163 5627
rect 15286 5624 15292 5636
rect 15151 5596 15292 5624
rect 15151 5593 15163 5596
rect 15105 5587 15163 5593
rect 15286 5584 15292 5596
rect 15344 5624 15350 5636
rect 15344 5596 15884 5624
rect 15344 5584 15350 5596
rect 9263 5528 9444 5556
rect 9953 5559 10011 5565
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9953 5525 9965 5559
rect 9999 5556 10011 5559
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 9999 5528 11069 5556
rect 9999 5525 10011 5528
rect 9953 5519 10011 5525
rect 11057 5525 11069 5528
rect 11103 5556 11115 5559
rect 12342 5556 12348 5568
rect 11103 5528 12348 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 12584 5528 13369 5556
rect 12584 5516 12590 5528
rect 13357 5525 13369 5528
rect 13403 5556 13415 5559
rect 14182 5556 14188 5568
rect 13403 5528 14188 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 14182 5516 14188 5528
rect 14240 5556 14246 5568
rect 15654 5556 15660 5568
rect 14240 5528 15660 5556
rect 14240 5516 14246 5528
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 15856 5565 15884 5596
rect 15930 5584 15936 5636
rect 15988 5624 15994 5636
rect 16666 5624 16672 5636
rect 15988 5596 16672 5624
rect 15988 5584 15994 5596
rect 16666 5584 16672 5596
rect 16724 5584 16730 5636
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16114 5556 16120 5568
rect 15887 5528 16120 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 17126 5516 17132 5568
rect 17184 5516 17190 5568
rect 18230 5516 18236 5568
rect 18288 5516 18294 5568
rect 19058 5516 19064 5568
rect 19116 5516 19122 5568
rect 19352 5565 19380 5664
rect 20272 5633 20300 5800
rect 22112 5800 22600 5828
rect 22112 5760 22140 5800
rect 22572 5769 22600 5800
rect 21744 5732 22140 5760
rect 22557 5763 22615 5769
rect 21744 5704 21772 5732
rect 22557 5729 22569 5763
rect 22603 5729 22615 5763
rect 22557 5723 22615 5729
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 23032 5732 24409 5760
rect 23032 5704 23060 5732
rect 24397 5729 24409 5732
rect 24443 5729 24455 5763
rect 24397 5723 24455 5729
rect 26234 5720 26240 5772
rect 26292 5720 26298 5772
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 27706 5760 27712 5772
rect 26476 5732 27712 5760
rect 26476 5720 26482 5732
rect 27706 5720 27712 5732
rect 27764 5720 27770 5772
rect 28276 5760 28304 5856
rect 28997 5763 29055 5769
rect 28997 5760 29009 5763
rect 28276 5732 29009 5760
rect 28997 5729 29009 5732
rect 29043 5729 29055 5763
rect 29564 5760 29592 5856
rect 29564 5732 29776 5760
rect 28997 5723 29055 5729
rect 21726 5652 21732 5704
rect 21784 5652 21790 5704
rect 22186 5692 22192 5704
rect 21836 5664 22192 5692
rect 20257 5627 20315 5633
rect 20257 5593 20269 5627
rect 20303 5624 20315 5627
rect 21836 5624 21864 5664
rect 22186 5652 22192 5664
rect 22244 5652 22250 5704
rect 23014 5652 23020 5704
rect 23072 5652 23078 5704
rect 23382 5652 23388 5704
rect 23440 5652 23446 5704
rect 23658 5652 23664 5704
rect 23716 5652 23722 5704
rect 26252 5692 26280 5720
rect 26160 5664 26280 5692
rect 20303 5596 21864 5624
rect 24664 5627 24722 5633
rect 20303 5593 20315 5596
rect 20257 5587 20315 5593
rect 24664 5593 24676 5627
rect 24710 5624 24722 5627
rect 25314 5624 25320 5636
rect 24710 5596 25320 5624
rect 24710 5593 24722 5596
rect 24664 5587 24722 5593
rect 25314 5584 25320 5596
rect 25372 5584 25378 5636
rect 19337 5559 19395 5565
rect 19337 5525 19349 5559
rect 19383 5525 19395 5559
rect 19337 5519 19395 5525
rect 19705 5559 19763 5565
rect 19705 5525 19717 5559
rect 19751 5556 19763 5559
rect 19794 5556 19800 5568
rect 19751 5528 19800 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21545 5559 21603 5565
rect 21545 5556 21557 5559
rect 20772 5528 21557 5556
rect 20772 5516 20778 5528
rect 21545 5525 21557 5528
rect 21591 5556 21603 5559
rect 21910 5556 21916 5568
rect 21591 5528 21916 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 21910 5516 21916 5528
rect 21968 5516 21974 5568
rect 22002 5516 22008 5568
rect 22060 5556 22066 5568
rect 22097 5559 22155 5565
rect 22097 5556 22109 5559
rect 22060 5528 22109 5556
rect 22060 5516 22066 5528
rect 22097 5525 22109 5528
rect 22143 5525 22155 5559
rect 22097 5519 22155 5525
rect 22370 5516 22376 5568
rect 22428 5556 22434 5568
rect 22465 5559 22523 5565
rect 22465 5556 22477 5559
rect 22428 5528 22477 5556
rect 22428 5516 22434 5528
rect 22465 5525 22477 5528
rect 22511 5525 22523 5559
rect 22465 5519 22523 5525
rect 23934 5516 23940 5568
rect 23992 5556 23998 5568
rect 24213 5559 24271 5565
rect 24213 5556 24225 5559
rect 23992 5528 24225 5556
rect 23992 5516 23998 5528
rect 24213 5525 24225 5528
rect 24259 5525 24271 5559
rect 24213 5519 24271 5525
rect 24394 5516 24400 5568
rect 24452 5556 24458 5568
rect 25777 5559 25835 5565
rect 25777 5556 25789 5559
rect 24452 5528 25789 5556
rect 24452 5516 24458 5528
rect 25777 5525 25789 5528
rect 25823 5525 25835 5559
rect 25777 5519 25835 5525
rect 25866 5516 25872 5568
rect 25924 5516 25930 5568
rect 26160 5556 26188 5664
rect 26326 5652 26332 5704
rect 26384 5692 26390 5704
rect 26697 5695 26755 5701
rect 26697 5692 26709 5695
rect 26384 5664 26709 5692
rect 26384 5652 26390 5664
rect 26697 5661 26709 5664
rect 26743 5661 26755 5695
rect 26697 5655 26755 5661
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5692 28963 5695
rect 29270 5692 29276 5704
rect 28951 5664 29276 5692
rect 28951 5661 28963 5664
rect 28905 5655 28963 5661
rect 29270 5652 29276 5664
rect 29328 5692 29334 5704
rect 29748 5701 29776 5732
rect 30650 5720 30656 5772
rect 30708 5760 30714 5772
rect 31389 5763 31447 5769
rect 31389 5760 31401 5763
rect 30708 5732 31156 5760
rect 30708 5720 30714 5732
rect 31128 5708 31156 5732
rect 31312 5732 31401 5760
rect 31312 5708 31340 5732
rect 31389 5729 31401 5732
rect 31435 5729 31447 5763
rect 31588 5760 31616 5868
rect 31864 5868 32864 5896
rect 31864 5760 31892 5868
rect 32858 5856 32864 5868
rect 32916 5856 32922 5908
rect 32950 5856 32956 5908
rect 33008 5896 33014 5908
rect 33321 5899 33379 5905
rect 33321 5896 33333 5899
rect 33008 5868 33333 5896
rect 33008 5856 33014 5868
rect 33321 5865 33333 5868
rect 33367 5865 33379 5899
rect 33321 5859 33379 5865
rect 34517 5899 34575 5905
rect 34517 5865 34529 5899
rect 34563 5896 34575 5899
rect 34606 5896 34612 5908
rect 34563 5868 34612 5896
rect 34563 5865 34575 5868
rect 34517 5859 34575 5865
rect 34606 5856 34612 5868
rect 34664 5856 34670 5908
rect 35802 5856 35808 5908
rect 35860 5896 35866 5908
rect 38105 5899 38163 5905
rect 38105 5896 38117 5899
rect 35860 5868 38117 5896
rect 35860 5856 35866 5868
rect 38105 5865 38117 5868
rect 38151 5865 38163 5899
rect 38105 5859 38163 5865
rect 38562 5856 38568 5908
rect 38620 5896 38626 5908
rect 38749 5899 38807 5905
rect 38749 5896 38761 5899
rect 38620 5868 38761 5896
rect 38620 5856 38626 5868
rect 38749 5865 38761 5868
rect 38795 5865 38807 5899
rect 40218 5896 40224 5908
rect 38749 5859 38807 5865
rect 39224 5868 40224 5896
rect 31588 5732 31892 5760
rect 31389 5723 31447 5729
rect 32214 5720 32220 5772
rect 32272 5760 32278 5772
rect 32677 5763 32735 5769
rect 32677 5760 32689 5763
rect 32272 5732 32689 5760
rect 32272 5720 32278 5732
rect 32677 5729 32689 5732
rect 32723 5729 32735 5763
rect 34624 5760 34652 5856
rect 37277 5831 37335 5837
rect 37277 5797 37289 5831
rect 37323 5828 37335 5831
rect 37323 5800 37504 5828
rect 37323 5797 37335 5800
rect 37277 5791 37335 5797
rect 35897 5763 35955 5769
rect 35897 5760 35909 5763
rect 34624 5732 35909 5760
rect 32677 5723 32735 5729
rect 35897 5729 35909 5732
rect 35943 5729 35955 5763
rect 35897 5723 35955 5729
rect 29733 5695 29791 5701
rect 29328 5664 29684 5692
rect 29328 5652 29334 5664
rect 26237 5627 26295 5633
rect 26237 5593 26249 5627
rect 26283 5624 26295 5627
rect 27341 5627 27399 5633
rect 27341 5624 27353 5627
rect 26283 5596 27353 5624
rect 26283 5593 26295 5596
rect 26237 5587 26295 5593
rect 27341 5593 27353 5596
rect 27387 5593 27399 5627
rect 27341 5587 27399 5593
rect 28813 5627 28871 5633
rect 28813 5593 28825 5627
rect 28859 5624 28871 5627
rect 29546 5624 29552 5636
rect 28859 5596 29552 5624
rect 28859 5593 28871 5596
rect 28813 5587 28871 5593
rect 29546 5584 29552 5596
rect 29604 5584 29610 5636
rect 26329 5559 26387 5565
rect 26329 5556 26341 5559
rect 26160 5528 26341 5556
rect 26329 5525 26341 5528
rect 26375 5525 26387 5559
rect 26329 5519 26387 5525
rect 28442 5516 28448 5568
rect 28500 5516 28506 5568
rect 29656 5556 29684 5664
rect 29733 5661 29745 5695
rect 29779 5661 29791 5695
rect 31128 5680 31340 5708
rect 37476 5704 37504 5800
rect 39224 5769 39252 5868
rect 40218 5856 40224 5868
rect 40276 5856 40282 5908
rect 44910 5856 44916 5908
rect 44968 5896 44974 5908
rect 45005 5899 45063 5905
rect 45005 5896 45017 5899
rect 44968 5868 45017 5896
rect 44968 5856 44974 5868
rect 45005 5865 45017 5868
rect 45051 5865 45063 5899
rect 45005 5859 45063 5865
rect 45646 5856 45652 5908
rect 45704 5856 45710 5908
rect 46845 5899 46903 5905
rect 46845 5865 46857 5899
rect 46891 5896 46903 5899
rect 46934 5896 46940 5908
rect 46891 5868 46940 5896
rect 46891 5865 46903 5868
rect 46845 5859 46903 5865
rect 46934 5856 46940 5868
rect 46992 5856 46998 5908
rect 49602 5856 49608 5908
rect 49660 5856 49666 5908
rect 54021 5899 54079 5905
rect 54021 5865 54033 5899
rect 54067 5896 54079 5899
rect 54202 5896 54208 5908
rect 54067 5868 54208 5896
rect 54067 5865 54079 5868
rect 54021 5859 54079 5865
rect 54202 5856 54208 5868
rect 54260 5896 54266 5908
rect 55030 5896 55036 5908
rect 54260 5868 55036 5896
rect 54260 5856 54266 5868
rect 55030 5856 55036 5868
rect 55088 5856 55094 5908
rect 55306 5856 55312 5908
rect 55364 5896 55370 5908
rect 57054 5896 57060 5908
rect 55364 5868 57060 5896
rect 55364 5856 55370 5868
rect 57054 5856 57060 5868
rect 57112 5896 57118 5908
rect 57333 5899 57391 5905
rect 57333 5896 57345 5899
rect 57112 5868 57345 5896
rect 57112 5856 57118 5868
rect 57333 5865 57345 5868
rect 57379 5865 57391 5899
rect 57333 5859 57391 5865
rect 57422 5856 57428 5908
rect 57480 5856 57486 5908
rect 58253 5899 58311 5905
rect 58253 5865 58265 5899
rect 58299 5896 58311 5899
rect 58342 5896 58348 5908
rect 58299 5868 58348 5896
rect 58299 5865 58311 5868
rect 58253 5859 58311 5865
rect 58342 5856 58348 5868
rect 58400 5856 58406 5908
rect 40236 5828 40264 5856
rect 41141 5831 41199 5837
rect 40236 5800 40724 5828
rect 39209 5763 39267 5769
rect 39209 5729 39221 5763
rect 39255 5729 39267 5763
rect 39209 5723 39267 5729
rect 39390 5720 39396 5772
rect 39448 5720 39454 5772
rect 40586 5760 40592 5772
rect 39776 5732 40592 5760
rect 29733 5655 29791 5661
rect 31846 5652 31852 5704
rect 31904 5652 31910 5704
rect 33594 5652 33600 5704
rect 33652 5652 33658 5704
rect 34698 5652 34704 5704
rect 34756 5652 34762 5704
rect 36906 5652 36912 5704
rect 36964 5692 36970 5704
rect 37369 5695 37427 5701
rect 37369 5692 37381 5695
rect 36964 5664 37381 5692
rect 36964 5652 36970 5664
rect 37369 5661 37381 5664
rect 37415 5661 37427 5695
rect 37369 5655 37427 5661
rect 37458 5652 37464 5704
rect 37516 5652 37522 5704
rect 38289 5695 38347 5701
rect 38289 5661 38301 5695
rect 38335 5692 38347 5695
rect 39776 5692 39804 5732
rect 40586 5720 40592 5732
rect 40644 5720 40650 5772
rect 40696 5760 40724 5800
rect 41141 5797 41153 5831
rect 41187 5828 41199 5831
rect 41187 5800 42012 5828
rect 41187 5797 41199 5800
rect 41141 5791 41199 5797
rect 41601 5763 41659 5769
rect 41601 5760 41613 5763
rect 40696 5732 41613 5760
rect 41601 5729 41613 5732
rect 41647 5729 41659 5763
rect 41601 5723 41659 5729
rect 41785 5763 41843 5769
rect 41785 5729 41797 5763
rect 41831 5760 41843 5763
rect 41874 5760 41880 5772
rect 41831 5732 41880 5760
rect 41831 5729 41843 5732
rect 41785 5723 41843 5729
rect 41874 5720 41880 5732
rect 41932 5720 41938 5772
rect 41984 5769 42012 5800
rect 45664 5769 45692 5856
rect 41969 5763 42027 5769
rect 41969 5729 41981 5763
rect 42015 5729 42027 5763
rect 41969 5723 42027 5729
rect 45649 5763 45707 5769
rect 45649 5729 45661 5763
rect 45695 5729 45707 5763
rect 46952 5760 46980 5856
rect 50157 5831 50215 5837
rect 50157 5797 50169 5831
rect 50203 5828 50215 5831
rect 58912 5828 58940 6072
rect 50203 5800 51074 5828
rect 50203 5797 50215 5800
rect 50157 5791 50215 5797
rect 47213 5763 47271 5769
rect 47213 5760 47225 5763
rect 46952 5732 47225 5760
rect 45649 5723 45707 5729
rect 47213 5729 47225 5732
rect 47259 5729 47271 5763
rect 47213 5723 47271 5729
rect 50338 5720 50344 5772
rect 50396 5760 50402 5772
rect 50709 5763 50767 5769
rect 50709 5760 50721 5763
rect 50396 5732 50721 5760
rect 50396 5720 50402 5732
rect 50709 5729 50721 5732
rect 50755 5729 50767 5763
rect 51046 5760 51074 5800
rect 57348 5800 58940 5828
rect 51721 5763 51779 5769
rect 51721 5760 51733 5763
rect 51046 5732 51733 5760
rect 50709 5723 50767 5729
rect 51721 5729 51733 5732
rect 51767 5729 51779 5763
rect 51721 5723 51779 5729
rect 52546 5720 52552 5772
rect 52604 5760 52610 5772
rect 52641 5763 52699 5769
rect 52641 5760 52653 5763
rect 52604 5732 52653 5760
rect 52604 5720 52610 5732
rect 52641 5729 52653 5732
rect 52687 5729 52699 5763
rect 55953 5763 56011 5769
rect 55953 5760 55965 5763
rect 52641 5723 52699 5729
rect 53760 5732 55965 5760
rect 38335 5664 39804 5692
rect 38335 5661 38347 5664
rect 38289 5655 38347 5661
rect 39850 5652 39856 5704
rect 39908 5652 39914 5704
rect 39942 5652 39948 5704
rect 40000 5692 40006 5704
rect 40000 5664 40632 5692
rect 40000 5652 40006 5664
rect 30558 5584 30564 5636
rect 30616 5624 30622 5636
rect 30742 5624 30748 5636
rect 30616 5596 30748 5624
rect 30616 5584 30622 5596
rect 30742 5584 30748 5596
rect 30800 5584 30806 5636
rect 31294 5584 31300 5636
rect 31352 5584 31358 5636
rect 31478 5584 31484 5636
rect 31536 5624 31542 5636
rect 32309 5627 32367 5633
rect 32309 5624 32321 5627
rect 31536 5596 32321 5624
rect 31536 5584 31542 5596
rect 32309 5593 32321 5596
rect 32355 5624 32367 5627
rect 32953 5627 33011 5633
rect 32953 5624 32965 5627
rect 32355 5596 32965 5624
rect 32355 5593 32367 5596
rect 32309 5587 32367 5593
rect 32953 5593 32965 5596
rect 32999 5593 33011 5627
rect 32953 5587 33011 5593
rect 34606 5584 34612 5636
rect 34664 5624 34670 5636
rect 35526 5624 35532 5636
rect 34664 5596 35532 5624
rect 34664 5584 34670 5596
rect 35526 5584 35532 5596
rect 35584 5584 35590 5636
rect 36164 5627 36222 5633
rect 36164 5593 36176 5627
rect 36210 5624 36222 5627
rect 38013 5627 38071 5633
rect 38013 5624 38025 5627
rect 36210 5596 38025 5624
rect 36210 5593 36222 5596
rect 36164 5587 36222 5593
rect 38013 5593 38025 5596
rect 38059 5593 38071 5627
rect 38013 5587 38071 5593
rect 39117 5627 39175 5633
rect 39117 5593 39129 5627
rect 39163 5624 39175 5627
rect 40497 5627 40555 5633
rect 40497 5624 40509 5627
rect 39163 5596 40509 5624
rect 39163 5593 39175 5596
rect 39117 5587 39175 5593
rect 40497 5593 40509 5596
rect 40543 5593 40555 5627
rect 40604 5624 40632 5664
rect 40678 5652 40684 5704
rect 40736 5692 40742 5704
rect 42889 5695 42947 5701
rect 42889 5692 42901 5695
rect 40736 5664 42901 5692
rect 40736 5652 40742 5664
rect 42889 5661 42901 5664
rect 42935 5661 42947 5695
rect 42889 5655 42947 5661
rect 43257 5695 43315 5701
rect 43257 5661 43269 5695
rect 43303 5692 43315 5695
rect 43346 5692 43352 5704
rect 43303 5664 43352 5692
rect 43303 5661 43315 5664
rect 43257 5655 43315 5661
rect 43346 5652 43352 5664
rect 43404 5652 43410 5704
rect 43990 5652 43996 5704
rect 44048 5652 44054 5704
rect 44174 5652 44180 5704
rect 44232 5692 44238 5704
rect 45370 5692 45376 5704
rect 44232 5664 45376 5692
rect 44232 5652 44238 5664
rect 45370 5652 45376 5664
rect 45428 5652 45434 5704
rect 45830 5652 45836 5704
rect 45888 5652 45894 5704
rect 48682 5652 48688 5704
rect 48740 5652 48746 5704
rect 50154 5652 50160 5704
rect 50212 5692 50218 5704
rect 50525 5695 50583 5701
rect 50525 5692 50537 5695
rect 50212 5664 50537 5692
rect 50212 5652 50218 5664
rect 50525 5661 50537 5664
rect 50571 5661 50583 5695
rect 50525 5655 50583 5661
rect 50982 5652 50988 5704
rect 51040 5652 51046 5704
rect 52656 5692 52684 5723
rect 53760 5692 53788 5732
rect 55953 5729 55965 5732
rect 55999 5729 56011 5763
rect 55953 5723 56011 5729
rect 52656 5664 53788 5692
rect 53926 5652 53932 5704
rect 53984 5692 53990 5704
rect 54113 5695 54171 5701
rect 54113 5692 54125 5695
rect 53984 5664 54125 5692
rect 53984 5652 53990 5664
rect 54113 5661 54125 5664
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 55122 5652 55128 5704
rect 55180 5652 55186 5704
rect 55490 5652 55496 5704
rect 55548 5652 55554 5704
rect 55677 5695 55735 5701
rect 55677 5661 55689 5695
rect 55723 5692 55735 5695
rect 55858 5692 55864 5704
rect 55723 5664 55864 5692
rect 55723 5661 55735 5664
rect 55677 5655 55735 5661
rect 55858 5652 55864 5664
rect 55916 5652 55922 5704
rect 56220 5695 56278 5701
rect 56220 5661 56232 5695
rect 56266 5692 56278 5695
rect 57348 5692 57376 5800
rect 57514 5720 57520 5772
rect 57572 5720 57578 5772
rect 57974 5720 57980 5772
rect 58032 5720 58038 5772
rect 56266 5664 57376 5692
rect 56266 5661 56278 5664
rect 56220 5655 56278 5661
rect 41414 5624 41420 5636
rect 40604 5596 41420 5624
rect 40497 5587 40555 5593
rect 41414 5584 41420 5596
rect 41472 5584 41478 5636
rect 41509 5627 41567 5633
rect 41509 5593 41521 5627
rect 41555 5624 41567 5627
rect 43070 5624 43076 5636
rect 41555 5596 43076 5624
rect 41555 5593 41567 5596
rect 41509 5587 41567 5593
rect 43070 5584 43076 5596
rect 43128 5584 43134 5636
rect 47480 5627 47538 5633
rect 43916 5596 47440 5624
rect 43916 5568 43944 5596
rect 31110 5556 31116 5568
rect 29656 5528 31116 5556
rect 31110 5516 31116 5528
rect 31168 5516 31174 5568
rect 31202 5516 31208 5568
rect 31260 5516 31266 5568
rect 34146 5516 34152 5568
rect 34204 5516 34210 5568
rect 36262 5516 36268 5568
rect 36320 5556 36326 5568
rect 38657 5559 38715 5565
rect 38657 5556 38669 5559
rect 36320 5528 38669 5556
rect 36320 5516 36326 5528
rect 38657 5525 38669 5528
rect 38703 5556 38715 5559
rect 40126 5556 40132 5568
rect 38703 5528 40132 5556
rect 38703 5525 38715 5528
rect 38657 5519 38715 5525
rect 40126 5516 40132 5528
rect 40184 5516 40190 5568
rect 40770 5516 40776 5568
rect 40828 5516 40834 5568
rect 41966 5516 41972 5568
rect 42024 5556 42030 5568
rect 42613 5559 42671 5565
rect 42613 5556 42625 5559
rect 42024 5528 42625 5556
rect 42024 5516 42030 5528
rect 42613 5525 42625 5528
rect 42659 5525 42671 5559
rect 42613 5519 42671 5525
rect 43806 5516 43812 5568
rect 43864 5516 43870 5568
rect 43898 5516 43904 5568
rect 43956 5516 43962 5568
rect 44082 5516 44088 5568
rect 44140 5556 44146 5568
rect 44637 5559 44695 5565
rect 44637 5556 44649 5559
rect 44140 5528 44649 5556
rect 44140 5516 44146 5528
rect 44637 5525 44649 5528
rect 44683 5525 44695 5559
rect 44637 5519 44695 5525
rect 45465 5559 45523 5565
rect 45465 5525 45477 5559
rect 45511 5556 45523 5559
rect 46477 5559 46535 5565
rect 46477 5556 46489 5559
rect 45511 5528 46489 5556
rect 45511 5525 45523 5528
rect 45465 5519 45523 5525
rect 46477 5525 46489 5528
rect 46523 5525 46535 5559
rect 47412 5556 47440 5596
rect 47480 5593 47492 5627
rect 47526 5624 47538 5627
rect 49329 5627 49387 5633
rect 49329 5624 49341 5627
rect 47526 5596 49341 5624
rect 47526 5593 47538 5596
rect 47480 5587 47538 5593
rect 49329 5593 49341 5596
rect 49375 5593 49387 5627
rect 49329 5587 49387 5593
rect 52908 5627 52966 5633
rect 52908 5593 52920 5627
rect 52954 5624 52966 5627
rect 54757 5627 54815 5633
rect 54757 5624 54769 5627
rect 52954 5596 54769 5624
rect 52954 5593 52966 5596
rect 52908 5587 52966 5593
rect 54757 5593 54769 5596
rect 54803 5593 54815 5627
rect 54757 5587 54815 5593
rect 55030 5584 55036 5636
rect 55088 5624 55094 5636
rect 57532 5624 57560 5720
rect 57698 5652 57704 5704
rect 57756 5692 57762 5704
rect 57793 5695 57851 5701
rect 57793 5692 57805 5695
rect 57756 5664 57805 5692
rect 57756 5652 57762 5664
rect 57793 5661 57805 5664
rect 57839 5661 57851 5695
rect 57793 5655 57851 5661
rect 57882 5652 57888 5704
rect 57940 5692 57946 5704
rect 58437 5695 58495 5701
rect 58437 5692 58449 5695
rect 57940 5664 58449 5692
rect 57940 5652 57946 5664
rect 58437 5661 58449 5664
rect 58483 5661 58495 5695
rect 58437 5655 58495 5661
rect 55088 5596 57560 5624
rect 55088 5584 55094 5596
rect 48498 5556 48504 5568
rect 47412 5528 48504 5556
rect 46477 5519 46535 5525
rect 48498 5516 48504 5528
rect 48556 5516 48562 5568
rect 48593 5559 48651 5565
rect 48593 5525 48605 5559
rect 48639 5556 48651 5559
rect 49418 5556 49424 5568
rect 48639 5528 49424 5556
rect 48639 5525 48651 5528
rect 48593 5519 48651 5525
rect 49418 5516 49424 5528
rect 49476 5516 49482 5568
rect 50617 5559 50675 5565
rect 50617 5525 50629 5559
rect 50663 5556 50675 5559
rect 51629 5559 51687 5565
rect 51629 5556 51641 5559
rect 50663 5528 51641 5556
rect 50663 5525 50675 5528
rect 50617 5519 50675 5525
rect 51629 5525 51641 5528
rect 51675 5525 51687 5559
rect 51629 5519 51687 5525
rect 52362 5516 52368 5568
rect 52420 5516 52426 5568
rect 54938 5516 54944 5568
rect 54996 5516 55002 5568
rect 55861 5559 55919 5565
rect 55861 5525 55873 5559
rect 55907 5556 55919 5559
rect 56502 5556 56508 5568
rect 55907 5528 56508 5556
rect 55907 5525 55919 5528
rect 55861 5519 55919 5525
rect 56502 5516 56508 5528
rect 56560 5516 56566 5568
rect 56778 5516 56784 5568
rect 56836 5556 56842 5568
rect 57885 5559 57943 5565
rect 57885 5556 57897 5559
rect 56836 5528 57897 5556
rect 56836 5516 56842 5528
rect 57885 5525 57897 5528
rect 57931 5525 57943 5559
rect 57885 5519 57943 5525
rect 1104 5466 59040 5488
rect 1104 5414 15394 5466
rect 15446 5414 15458 5466
rect 15510 5414 15522 5466
rect 15574 5414 15586 5466
rect 15638 5414 15650 5466
rect 15702 5414 29838 5466
rect 29890 5414 29902 5466
rect 29954 5414 29966 5466
rect 30018 5414 30030 5466
rect 30082 5414 30094 5466
rect 30146 5414 44282 5466
rect 44334 5414 44346 5466
rect 44398 5414 44410 5466
rect 44462 5414 44474 5466
rect 44526 5414 44538 5466
rect 44590 5414 58726 5466
rect 58778 5414 58790 5466
rect 58842 5414 58854 5466
rect 58906 5414 58918 5466
rect 58970 5414 58982 5466
rect 59034 5414 59040 5466
rect 1104 5392 59040 5414
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 3384 5324 4537 5352
rect 3384 5312 3390 5324
rect 4525 5321 4537 5324
rect 4571 5321 4583 5355
rect 4525 5315 4583 5321
rect 5460 5324 6684 5352
rect 5460 5296 5488 5324
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 3660 5256 3801 5284
rect 3660 5244 3666 5256
rect 3789 5253 3801 5256
rect 3835 5284 3847 5287
rect 3835 5256 3924 5284
rect 3835 5253 3847 5256
rect 3789 5247 3847 5253
rect 3896 5225 3924 5256
rect 5442 5244 5448 5296
rect 5500 5244 5506 5296
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 5684 5256 6561 5284
rect 5684 5244 5690 5256
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 5166 5216 5172 5228
rect 3927 5188 5172 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 5166 5176 5172 5188
rect 5224 5216 5230 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 5224 5188 5365 5216
rect 5224 5176 5230 5188
rect 5353 5185 5365 5188
rect 5399 5216 5411 5219
rect 5718 5216 5724 5228
rect 5399 5188 5724 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5718 5176 5724 5188
rect 5776 5216 5782 5228
rect 6656 5225 6684 5324
rect 7834 5312 7840 5364
rect 7892 5312 7898 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 10502 5352 10508 5364
rect 10275 5324 10508 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 10502 5312 10508 5324
rect 10560 5352 10566 5364
rect 11698 5352 11704 5364
rect 10560 5324 11704 5352
rect 10560 5312 10566 5324
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 13078 5352 13084 5364
rect 12400 5324 13084 5352
rect 12400 5312 12406 5324
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 14461 5355 14519 5361
rect 14461 5352 14473 5355
rect 13872 5324 14473 5352
rect 13872 5312 13878 5324
rect 14461 5321 14473 5324
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 14737 5355 14795 5361
rect 14737 5321 14749 5355
rect 14783 5321 14795 5355
rect 14737 5315 14795 5321
rect 15565 5355 15623 5361
rect 15565 5321 15577 5355
rect 15611 5352 15623 5355
rect 15746 5352 15752 5364
rect 15611 5324 15752 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 12066 5284 12072 5296
rect 7024 5256 12072 5284
rect 7024 5225 7052 5256
rect 12066 5244 12072 5256
rect 12124 5284 12130 5296
rect 14369 5287 14427 5293
rect 12124 5256 12434 5284
rect 12124 5244 12130 5256
rect 6641 5219 6699 5225
rect 5776 5188 5948 5216
rect 5776 5176 5782 5188
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 2133 5151 2191 5157
rect 2133 5148 2145 5151
rect 1820 5120 2145 5148
rect 1820 5108 1826 5120
rect 2133 5117 2145 5120
rect 2179 5117 2191 5151
rect 2133 5111 2191 5117
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2866 5148 2872 5160
rect 2455 5120 2872 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 5132 5120 5273 5148
rect 5132 5108 5138 5120
rect 5261 5117 5273 5120
rect 5307 5148 5319 5151
rect 5442 5148 5448 5160
rect 5307 5120 5448 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5117 5871 5151
rect 5920 5148 5948 5188
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 7892 5188 9689 5216
rect 7892 5176 7898 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 9677 5179 9735 5185
rect 10336 5188 11529 5216
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 5920 5120 7113 5148
rect 5813 5111 5871 5117
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 5626 5080 5632 5092
rect 3936 5052 5632 5080
rect 3936 5040 3942 5052
rect 5626 5040 5632 5052
rect 5684 5080 5690 5092
rect 5828 5080 5856 5111
rect 8018 5108 8024 5160
rect 8076 5108 8082 5160
rect 8846 5108 8852 5160
rect 8904 5108 8910 5160
rect 9030 5108 9036 5160
rect 9088 5148 9094 5160
rect 10336 5148 10364 5188
rect 11517 5185 11529 5188
rect 11563 5216 11575 5219
rect 11698 5216 11704 5228
rect 11563 5188 11704 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12406 5216 12434 5256
rect 14369 5253 14381 5287
rect 14415 5284 14427 5287
rect 14752 5284 14780 5315
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 19518 5352 19524 5364
rect 17972 5324 19524 5352
rect 14415 5256 14780 5284
rect 16485 5287 16543 5293
rect 14415 5253 14427 5256
rect 14369 5247 14427 5253
rect 16485 5253 16497 5287
rect 16531 5284 16543 5287
rect 17678 5284 17684 5296
rect 16531 5256 17684 5284
rect 16531 5253 16543 5256
rect 16485 5247 16543 5253
rect 17678 5244 17684 5256
rect 17736 5244 17742 5296
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12406 5188 12541 5216
rect 12529 5185 12541 5188
rect 12575 5216 12587 5219
rect 13722 5216 13728 5228
rect 12575 5188 13728 5216
rect 12575 5185 12587 5188
rect 12529 5179 12587 5185
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 14918 5176 14924 5228
rect 14976 5176 14982 5228
rect 15194 5176 15200 5228
rect 15252 5176 15258 5228
rect 15746 5176 15752 5228
rect 15804 5176 15810 5228
rect 16850 5176 16856 5228
rect 16908 5176 16914 5228
rect 17972 5214 18000 5324
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 19702 5312 19708 5364
rect 19760 5312 19766 5364
rect 21450 5352 21456 5364
rect 19812 5324 21456 5352
rect 18414 5284 18420 5296
rect 18340 5256 18420 5284
rect 18340 5225 18368 5256
rect 18414 5244 18420 5256
rect 18472 5244 18478 5296
rect 18592 5287 18650 5293
rect 18592 5253 18604 5287
rect 18638 5284 18650 5287
rect 19058 5284 19064 5296
rect 18638 5256 19064 5284
rect 18638 5253 18650 5256
rect 18592 5247 18650 5253
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 19812 5225 19840 5324
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 22278 5312 22284 5364
rect 22336 5312 22342 5364
rect 23658 5312 23664 5364
rect 23716 5352 23722 5364
rect 24121 5355 24179 5361
rect 24121 5352 24133 5355
rect 23716 5324 24133 5352
rect 23716 5312 23722 5324
rect 24121 5321 24133 5324
rect 24167 5321 24179 5355
rect 24121 5315 24179 5321
rect 21910 5244 21916 5296
rect 21968 5284 21974 5296
rect 22922 5284 22928 5296
rect 21968 5256 22928 5284
rect 21968 5244 21974 5256
rect 18069 5217 18127 5223
rect 18069 5214 18081 5217
rect 17972 5186 18081 5214
rect 18069 5183 18081 5186
rect 18115 5183 18127 5217
rect 18069 5177 18127 5183
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5185 18383 5219
rect 19797 5219 19855 5225
rect 18325 5179 18383 5185
rect 18432 5188 19748 5216
rect 9088 5120 10364 5148
rect 9088 5108 9094 5120
rect 10778 5108 10784 5160
rect 10836 5108 10842 5160
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 11020 5120 12173 5148
rect 11020 5108 11026 5120
rect 12161 5117 12173 5120
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 13078 5108 13084 5160
rect 13136 5148 13142 5160
rect 14185 5151 14243 5157
rect 14185 5148 14197 5151
rect 13136 5120 14197 5148
rect 13136 5108 13142 5120
rect 14185 5117 14197 5120
rect 14231 5148 14243 5151
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14231 5120 15025 5148
rect 14231 5117 14243 5120
rect 14185 5111 14243 5117
rect 15013 5117 15025 5120
rect 15059 5148 15071 5151
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 15059 5120 17417 5148
rect 15059 5117 15071 5120
rect 15013 5111 15071 5117
rect 17405 5117 17417 5120
rect 17451 5148 17463 5151
rect 17770 5148 17776 5160
rect 17451 5120 17776 5148
rect 17451 5117 17463 5120
rect 17405 5111 17463 5117
rect 17770 5108 17776 5120
rect 17828 5148 17834 5160
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 17828 5120 17877 5148
rect 17828 5108 17834 5120
rect 17865 5117 17877 5120
rect 17911 5117 17923 5151
rect 18432 5148 18460 5188
rect 17865 5111 17923 5117
rect 18340 5120 18460 5148
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 5684 5052 5856 5080
rect 6012 5052 10517 5080
rect 5684 5040 5690 5052
rect 6012 5024 6040 5052
rect 10505 5049 10517 5052
rect 10551 5080 10563 5083
rect 11146 5080 11152 5092
rect 10551 5052 11152 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 11790 5080 11796 5092
rect 11256 5052 11796 5080
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5500 4984 5733 5012
rect 5500 4972 5506 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 6089 5015 6147 5021
rect 6089 4981 6101 5015
rect 6135 5012 6147 5015
rect 7558 5012 7564 5024
rect 6135 4984 7564 5012
rect 6135 4981 6147 4984
rect 6089 4975 6147 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 7984 4984 8585 5012
rect 7984 4972 7990 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 8573 4975 8631 4981
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 8720 4984 9413 5012
rect 8720 4972 8726 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 11256 5012 11284 5052
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 13449 5083 13507 5089
rect 13449 5049 13461 5083
rect 13495 5080 13507 5083
rect 14734 5080 14740 5092
rect 13495 5052 14740 5080
rect 13495 5049 13507 5052
rect 13449 5043 13507 5049
rect 14734 5040 14740 5052
rect 14792 5080 14798 5092
rect 18046 5080 18052 5092
rect 14792 5052 18052 5080
rect 14792 5040 14798 5052
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 18340 5080 18368 5120
rect 18156 5052 18368 5080
rect 19720 5080 19748 5188
rect 19797 5185 19809 5219
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 20990 5176 20996 5228
rect 21048 5176 21054 5228
rect 22756 5225 22784 5256
rect 22922 5244 22928 5256
rect 22980 5244 22986 5296
rect 21637 5219 21695 5225
rect 21637 5185 21649 5219
rect 21683 5216 21695 5219
rect 22189 5219 22247 5225
rect 22189 5216 22201 5219
rect 21683 5188 22201 5216
rect 21683 5185 21695 5188
rect 21637 5179 21695 5185
rect 22189 5185 22201 5188
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 23008 5219 23066 5225
rect 23008 5185 23020 5219
rect 23054 5216 23066 5219
rect 23566 5216 23572 5228
rect 23054 5188 23572 5216
rect 23054 5185 23066 5188
rect 23008 5179 23066 5185
rect 23566 5176 23572 5188
rect 23624 5176 23630 5228
rect 24136 5216 24164 5315
rect 26602 5312 26608 5364
rect 26660 5352 26666 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26660 5324 27353 5352
rect 26660 5312 26666 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 28902 5312 28908 5364
rect 28960 5312 28966 5364
rect 28997 5355 29055 5361
rect 28997 5321 29009 5355
rect 29043 5352 29055 5355
rect 29086 5352 29092 5364
rect 29043 5324 29092 5352
rect 29043 5321 29055 5324
rect 28997 5315 29055 5321
rect 29086 5312 29092 5324
rect 29144 5312 29150 5364
rect 29546 5312 29552 5364
rect 29604 5352 29610 5364
rect 30193 5355 30251 5361
rect 30193 5352 30205 5355
rect 29604 5324 30205 5352
rect 29604 5312 29610 5324
rect 30193 5321 30205 5324
rect 30239 5321 30251 5355
rect 30193 5315 30251 5321
rect 30650 5312 30656 5364
rect 30708 5352 30714 5364
rect 30929 5355 30987 5361
rect 30929 5352 30941 5355
rect 30708 5324 30941 5352
rect 30708 5312 30714 5324
rect 30929 5321 30941 5324
rect 30975 5321 30987 5355
rect 30929 5315 30987 5321
rect 31110 5312 31116 5364
rect 31168 5352 31174 5364
rect 31297 5355 31355 5361
rect 31297 5352 31309 5355
rect 31168 5324 31309 5352
rect 31168 5312 31174 5324
rect 31297 5321 31309 5324
rect 31343 5321 31355 5355
rect 37458 5352 37464 5364
rect 31297 5315 31355 5321
rect 35084 5324 37464 5352
rect 26789 5287 26847 5293
rect 26789 5253 26801 5287
rect 26835 5284 26847 5287
rect 27062 5284 27068 5296
rect 26835 5256 27068 5284
rect 26835 5253 26847 5256
rect 26789 5247 26847 5253
rect 27062 5244 27068 5256
rect 27120 5284 27126 5296
rect 32030 5284 32036 5296
rect 27120 5256 32036 5284
rect 27120 5244 27126 5256
rect 24136 5188 24716 5216
rect 19978 5108 19984 5160
rect 20036 5108 20042 5160
rect 20717 5151 20775 5157
rect 20717 5148 20729 5151
rect 20548 5120 20729 5148
rect 20254 5080 20260 5092
rect 19720 5052 20260 5080
rect 9815 4984 11284 5012
rect 11333 5015 11391 5021
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 11882 5012 11888 5024
rect 11379 4984 11888 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 14458 5012 14464 5024
rect 13863 4984 14464 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 14458 4972 14464 4984
rect 14516 5012 14522 5024
rect 15102 5012 15108 5024
rect 14516 4984 15108 5012
rect 14516 4972 14522 4984
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 15378 4972 15384 5024
rect 15436 4972 15442 5024
rect 16022 4972 16028 5024
rect 16080 4972 16086 5024
rect 16945 5015 17003 5021
rect 16945 4981 16957 5015
rect 16991 5012 17003 5015
rect 17034 5012 17040 5024
rect 16991 4984 17040 5012
rect 16991 4981 17003 4984
rect 16945 4975 17003 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 17773 5015 17831 5021
rect 17773 4981 17785 5015
rect 17819 5012 17831 5015
rect 18156 5012 18184 5052
rect 20254 5040 20260 5052
rect 20312 5080 20318 5092
rect 20441 5083 20499 5089
rect 20441 5080 20453 5083
rect 20312 5052 20453 5080
rect 20312 5040 20318 5052
rect 20441 5049 20453 5052
rect 20487 5049 20499 5083
rect 20441 5043 20499 5049
rect 17819 4984 18184 5012
rect 18233 5015 18291 5021
rect 17819 4981 17831 4984
rect 17773 4975 17831 4981
rect 18233 4981 18245 5015
rect 18279 5012 18291 5015
rect 19334 5012 19340 5024
rect 18279 4984 19340 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 19702 4972 19708 5024
rect 19760 5012 19766 5024
rect 20548 5012 20576 5120
rect 20717 5117 20729 5120
rect 20763 5117 20775 5151
rect 20717 5111 20775 5117
rect 20806 5108 20812 5160
rect 20864 5157 20870 5160
rect 20864 5151 20892 5157
rect 20880 5117 20892 5151
rect 20864 5111 20892 5117
rect 20864 5108 20870 5111
rect 21542 5108 21548 5160
rect 21600 5148 21606 5160
rect 22373 5151 22431 5157
rect 21600 5120 22094 5148
rect 21600 5108 21606 5120
rect 22066 5080 22094 5120
rect 22373 5117 22385 5151
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 22388 5080 22416 5111
rect 24394 5108 24400 5160
rect 24452 5108 24458 5160
rect 24581 5151 24639 5157
rect 24581 5117 24593 5151
rect 24627 5117 24639 5151
rect 24688 5148 24716 5188
rect 25590 5176 25596 5228
rect 25648 5176 25654 5228
rect 25317 5151 25375 5157
rect 25317 5148 25329 5151
rect 24688 5120 25329 5148
rect 24581 5111 24639 5117
rect 25317 5117 25329 5120
rect 25363 5117 25375 5151
rect 25317 5111 25375 5117
rect 22066 5052 22416 5080
rect 19760 4984 20576 5012
rect 19760 4972 19766 4984
rect 21818 4972 21824 5024
rect 21876 4972 21882 5024
rect 24596 5012 24624 5111
rect 25406 5108 25412 5160
rect 25464 5157 25470 5160
rect 27540 5157 27568 5256
rect 32030 5244 32036 5256
rect 32088 5284 32094 5296
rect 32309 5287 32367 5293
rect 32309 5284 32321 5287
rect 32088 5256 32321 5284
rect 32088 5244 32094 5256
rect 32309 5253 32321 5256
rect 32355 5253 32367 5287
rect 32309 5247 32367 5253
rect 33312 5287 33370 5293
rect 33312 5253 33324 5287
rect 33358 5284 33370 5287
rect 34146 5284 34152 5296
rect 33358 5256 34152 5284
rect 33358 5253 33370 5256
rect 33312 5247 33370 5253
rect 34146 5244 34152 5256
rect 34204 5244 34210 5296
rect 28353 5219 28411 5225
rect 28353 5185 28365 5219
rect 28399 5216 28411 5219
rect 28442 5216 28448 5228
rect 28399 5188 28448 5216
rect 28399 5185 28411 5188
rect 28353 5179 28411 5185
rect 28442 5176 28448 5188
rect 28500 5176 28506 5228
rect 29181 5219 29239 5225
rect 29181 5185 29193 5219
rect 29227 5216 29239 5219
rect 29270 5216 29276 5228
rect 29227 5188 29276 5216
rect 29227 5185 29239 5188
rect 29181 5179 29239 5185
rect 29270 5176 29276 5188
rect 29328 5176 29334 5228
rect 29638 5176 29644 5228
rect 29696 5176 29702 5228
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5216 30527 5219
rect 31018 5216 31024 5228
rect 30515 5188 31024 5216
rect 30515 5185 30527 5188
rect 30469 5179 30527 5185
rect 31018 5176 31024 5188
rect 31076 5176 31082 5228
rect 31205 5219 31263 5225
rect 31205 5185 31217 5219
rect 31251 5216 31263 5219
rect 31570 5216 31576 5228
rect 31251 5188 31576 5216
rect 31251 5185 31263 5188
rect 31205 5179 31263 5185
rect 31570 5176 31576 5188
rect 31628 5176 31634 5228
rect 33042 5176 33048 5228
rect 33100 5176 33106 5228
rect 34790 5176 34796 5228
rect 34848 5176 34854 5228
rect 35084 5225 35112 5324
rect 37458 5312 37464 5324
rect 37516 5312 37522 5364
rect 37550 5312 37556 5364
rect 37608 5312 37614 5364
rect 39301 5355 39359 5361
rect 39301 5321 39313 5355
rect 39347 5352 39359 5355
rect 39850 5352 39856 5364
rect 39347 5324 39856 5352
rect 39347 5321 39359 5324
rect 39301 5315 39359 5321
rect 39850 5312 39856 5324
rect 39908 5352 39914 5364
rect 40402 5352 40408 5364
rect 39908 5324 40408 5352
rect 39908 5312 39914 5324
rect 40402 5312 40408 5324
rect 40460 5312 40466 5364
rect 41690 5312 41696 5364
rect 41748 5352 41754 5364
rect 41785 5355 41843 5361
rect 41785 5352 41797 5355
rect 41748 5324 41797 5352
rect 41748 5312 41754 5324
rect 41785 5321 41797 5324
rect 41831 5321 41843 5355
rect 41785 5315 41843 5321
rect 44910 5312 44916 5364
rect 44968 5352 44974 5364
rect 45554 5352 45560 5364
rect 44968 5324 45560 5352
rect 44968 5312 44974 5324
rect 45554 5312 45560 5324
rect 45612 5312 45618 5364
rect 45646 5312 45652 5364
rect 45704 5352 45710 5364
rect 45830 5352 45836 5364
rect 45704 5324 45836 5352
rect 45704 5312 45710 5324
rect 45830 5312 45836 5324
rect 45888 5312 45894 5364
rect 46109 5355 46167 5361
rect 46109 5321 46121 5355
rect 46155 5352 46167 5355
rect 46842 5352 46848 5364
rect 46155 5324 46848 5352
rect 46155 5321 46167 5324
rect 46109 5315 46167 5321
rect 46842 5312 46848 5324
rect 46900 5312 46906 5364
rect 48133 5355 48191 5361
rect 48133 5321 48145 5355
rect 48179 5352 48191 5355
rect 48406 5352 48412 5364
rect 48179 5324 48412 5352
rect 48179 5321 48191 5324
rect 48133 5315 48191 5321
rect 48406 5312 48412 5324
rect 48464 5312 48470 5364
rect 50982 5352 50988 5364
rect 48516 5324 50988 5352
rect 35069 5219 35127 5225
rect 35069 5185 35081 5219
rect 35115 5185 35127 5219
rect 35069 5179 35127 5185
rect 35253 5219 35311 5225
rect 35253 5185 35265 5219
rect 35299 5216 35311 5219
rect 35434 5216 35440 5228
rect 35299 5188 35440 5216
rect 35299 5185 35311 5188
rect 35253 5179 35311 5185
rect 35434 5176 35440 5188
rect 35492 5176 35498 5228
rect 35986 5176 35992 5228
rect 36044 5176 36050 5228
rect 36262 5176 36268 5228
rect 36320 5176 36326 5228
rect 37568 5216 37596 5312
rect 38188 5287 38246 5293
rect 38188 5253 38200 5287
rect 38234 5284 38246 5287
rect 39114 5284 39120 5296
rect 38234 5256 39120 5284
rect 38234 5253 38246 5256
rect 38188 5247 38246 5253
rect 39114 5244 39120 5256
rect 39172 5244 39178 5296
rect 42518 5244 42524 5296
rect 42576 5284 42582 5296
rect 42972 5287 43030 5293
rect 42576 5256 42840 5284
rect 42576 5244 42582 5256
rect 37645 5219 37703 5225
rect 37645 5216 37657 5219
rect 37568 5188 37657 5216
rect 37645 5185 37657 5188
rect 37691 5185 37703 5219
rect 37645 5179 37703 5185
rect 40310 5176 40316 5228
rect 40368 5176 40374 5228
rect 40402 5176 40408 5228
rect 40460 5225 40466 5228
rect 40460 5219 40488 5225
rect 40476 5185 40488 5219
rect 40460 5179 40488 5185
rect 41233 5219 41291 5225
rect 41233 5185 41245 5219
rect 41279 5216 41291 5219
rect 41693 5219 41751 5225
rect 41693 5216 41705 5219
rect 41279 5188 41705 5216
rect 41279 5185 41291 5188
rect 41233 5179 41291 5185
rect 41693 5185 41705 5188
rect 41739 5185 41751 5219
rect 41693 5179 41751 5185
rect 40460 5176 40466 5179
rect 25464 5151 25492 5157
rect 25480 5117 25492 5151
rect 25464 5111 25492 5117
rect 26237 5151 26295 5157
rect 26237 5117 26249 5151
rect 26283 5148 26295 5151
rect 27433 5151 27491 5157
rect 27433 5148 27445 5151
rect 26283 5120 27445 5148
rect 26283 5117 26295 5120
rect 26237 5111 26295 5117
rect 27433 5117 27445 5120
rect 27479 5117 27491 5151
rect 27433 5111 27491 5117
rect 27525 5151 27583 5157
rect 27525 5117 27537 5151
rect 27571 5117 27583 5151
rect 27525 5111 27583 5117
rect 25464 5108 25470 5111
rect 29730 5108 29736 5160
rect 29788 5148 29794 5160
rect 30285 5151 30343 5157
rect 30285 5148 30297 5151
rect 29788 5120 30297 5148
rect 29788 5108 29794 5120
rect 30285 5117 30297 5120
rect 30331 5148 30343 5151
rect 34609 5151 34667 5157
rect 30331 5120 31800 5148
rect 30331 5117 30343 5120
rect 30285 5111 30343 5117
rect 24762 5040 24768 5092
rect 24820 5080 24826 5092
rect 25041 5083 25099 5089
rect 25041 5080 25053 5083
rect 24820 5052 25053 5080
rect 24820 5040 24826 5052
rect 25041 5049 25053 5052
rect 25087 5049 25099 5083
rect 25041 5043 25099 5049
rect 26142 5040 26148 5092
rect 26200 5080 26206 5092
rect 31772 5089 31800 5120
rect 34609 5117 34621 5151
rect 34655 5148 34667 5151
rect 34698 5148 34704 5160
rect 34655 5120 34704 5148
rect 34655 5117 34667 5120
rect 34609 5111 34667 5117
rect 34698 5108 34704 5120
rect 34756 5108 34762 5160
rect 36106 5151 36164 5157
rect 36106 5148 36118 5151
rect 35360 5120 36118 5148
rect 26973 5083 27031 5089
rect 26973 5080 26985 5083
rect 26200 5052 26985 5080
rect 26200 5040 26206 5052
rect 26973 5049 26985 5052
rect 27019 5049 27031 5083
rect 26973 5043 27031 5049
rect 31757 5083 31815 5089
rect 31757 5049 31769 5083
rect 31803 5080 31815 5083
rect 35360 5080 35388 5120
rect 36106 5117 36118 5120
rect 36152 5117 36164 5151
rect 36106 5111 36164 5117
rect 36446 5108 36452 5160
rect 36504 5148 36510 5160
rect 37461 5151 37519 5157
rect 37461 5148 37473 5151
rect 36504 5120 37473 5148
rect 36504 5108 36510 5120
rect 36740 5092 36768 5120
rect 37461 5117 37473 5120
rect 37507 5117 37519 5151
rect 37461 5111 37519 5117
rect 37550 5108 37556 5160
rect 37608 5148 37614 5160
rect 37921 5151 37979 5157
rect 37921 5148 37933 5151
rect 37608 5120 37933 5148
rect 37608 5108 37614 5120
rect 37921 5117 37933 5120
rect 37967 5117 37979 5151
rect 37921 5111 37979 5117
rect 39390 5108 39396 5160
rect 39448 5108 39454 5160
rect 39574 5108 39580 5160
rect 39632 5108 39638 5160
rect 40126 5108 40132 5160
rect 40184 5148 40190 5160
rect 40589 5151 40647 5157
rect 40589 5148 40601 5151
rect 40184 5120 40601 5148
rect 40184 5108 40190 5120
rect 40589 5117 40601 5120
rect 40635 5117 40647 5151
rect 40589 5111 40647 5117
rect 41414 5108 41420 5160
rect 41472 5148 41478 5160
rect 41969 5151 42027 5157
rect 41969 5148 41981 5151
rect 41472 5120 41981 5148
rect 41472 5108 41478 5120
rect 41969 5117 41981 5120
rect 42015 5148 42027 5151
rect 42536 5148 42564 5244
rect 42702 5176 42708 5228
rect 42760 5176 42766 5228
rect 42812 5216 42840 5256
rect 42972 5253 42984 5287
rect 43018 5284 43030 5287
rect 43806 5284 43812 5296
rect 43018 5256 43812 5284
rect 43018 5253 43030 5256
rect 42972 5247 43030 5253
rect 43806 5244 43812 5256
rect 43864 5244 43870 5296
rect 44536 5287 44594 5293
rect 44536 5253 44548 5287
rect 44582 5284 44594 5287
rect 45462 5284 45468 5296
rect 44582 5256 45468 5284
rect 44582 5253 44594 5256
rect 44536 5247 44594 5253
rect 45462 5244 45468 5256
rect 45520 5244 45526 5296
rect 48041 5219 48099 5225
rect 42812 5188 46428 5216
rect 42015 5120 42564 5148
rect 44269 5151 44327 5157
rect 42015 5117 42027 5120
rect 41969 5111 42027 5117
rect 44269 5117 44281 5151
rect 44315 5117 44327 5151
rect 44269 5111 44327 5117
rect 31803 5052 32812 5080
rect 31803 5049 31815 5052
rect 31757 5043 31815 5049
rect 26326 5012 26332 5024
rect 24596 4984 26332 5012
rect 26326 4972 26332 4984
rect 26384 4972 26390 5024
rect 28166 4972 28172 5024
rect 28224 4972 28230 5024
rect 29638 4972 29644 5024
rect 29696 5012 29702 5024
rect 30282 5012 30288 5024
rect 29696 4984 30288 5012
rect 29696 4972 29702 4984
rect 30282 4972 30288 4984
rect 30340 4972 30346 5024
rect 30650 4972 30656 5024
rect 30708 4972 30714 5024
rect 32674 4972 32680 5024
rect 32732 4972 32738 5024
rect 32784 5012 32812 5052
rect 34440 5052 35388 5080
rect 34146 5012 34152 5024
rect 32784 4984 34152 5012
rect 34146 4972 34152 4984
rect 34204 4972 34210 5024
rect 34330 4972 34336 5024
rect 34388 5012 34394 5024
rect 34440 5021 34468 5052
rect 35618 5040 35624 5092
rect 35676 5080 35682 5092
rect 35713 5083 35771 5089
rect 35713 5080 35725 5083
rect 35676 5052 35725 5080
rect 35676 5040 35682 5052
rect 35713 5049 35725 5052
rect 35759 5049 35771 5083
rect 35713 5043 35771 5049
rect 36722 5040 36728 5092
rect 36780 5040 36786 5092
rect 37642 5080 37648 5092
rect 36832 5052 37648 5080
rect 34425 5015 34483 5021
rect 34425 5012 34437 5015
rect 34388 4984 34437 5012
rect 34388 4972 34394 4984
rect 34425 4981 34437 4984
rect 34471 4981 34483 5015
rect 34425 4975 34483 4981
rect 34977 5015 35035 5021
rect 34977 4981 34989 5015
rect 35023 5012 35035 5015
rect 36832 5012 36860 5052
rect 37642 5040 37648 5052
rect 37700 5040 37706 5092
rect 40037 5083 40095 5089
rect 40037 5049 40049 5083
rect 40083 5049 40095 5083
rect 40037 5043 40095 5049
rect 35023 4984 36860 5012
rect 35023 4981 35035 4984
rect 34977 4975 35035 4981
rect 36906 4972 36912 5024
rect 36964 4972 36970 5024
rect 37826 4972 37832 5024
rect 37884 4972 37890 5024
rect 40052 5012 40080 5043
rect 40678 5012 40684 5024
rect 40052 4984 40684 5012
rect 40678 4972 40684 4984
rect 40736 4972 40742 5024
rect 41325 5015 41383 5021
rect 41325 4981 41337 5015
rect 41371 5012 41383 5015
rect 41414 5012 41420 5024
rect 41371 4984 41420 5012
rect 41371 4981 41383 4984
rect 41325 4975 41383 4981
rect 41414 4972 41420 4984
rect 41472 4972 41478 5024
rect 43990 4972 43996 5024
rect 44048 5012 44054 5024
rect 44085 5015 44143 5021
rect 44085 5012 44097 5015
rect 44048 4984 44097 5012
rect 44048 4972 44054 4984
rect 44085 4981 44097 4984
rect 44131 4981 44143 5015
rect 44284 5012 44312 5111
rect 46198 5108 46204 5160
rect 46256 5108 46262 5160
rect 46400 5157 46428 5188
rect 48041 5185 48053 5219
rect 48087 5185 48099 5219
rect 48041 5179 48099 5185
rect 46385 5151 46443 5157
rect 46385 5117 46397 5151
rect 46431 5117 46443 5151
rect 46385 5111 46443 5117
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 46891 5120 47716 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 46400 5080 46428 5111
rect 47118 5080 47124 5092
rect 46400 5052 47124 5080
rect 47118 5040 47124 5052
rect 47176 5040 47182 5092
rect 47688 5089 47716 5120
rect 47673 5083 47731 5089
rect 47673 5049 47685 5083
rect 47719 5049 47731 5083
rect 48056 5080 48084 5179
rect 48222 5108 48228 5160
rect 48280 5108 48286 5160
rect 48516 5157 48544 5324
rect 50982 5312 50988 5324
rect 51040 5352 51046 5364
rect 51813 5355 51871 5361
rect 51813 5352 51825 5355
rect 51040 5324 51825 5352
rect 51040 5312 51046 5324
rect 51813 5321 51825 5324
rect 51859 5321 51871 5355
rect 51813 5315 51871 5321
rect 53742 5312 53748 5364
rect 53800 5312 53806 5364
rect 54110 5312 54116 5364
rect 54168 5352 54174 5364
rect 54757 5355 54815 5361
rect 54757 5352 54769 5355
rect 54168 5324 54769 5352
rect 54168 5312 54174 5324
rect 54757 5321 54769 5324
rect 54803 5321 54815 5355
rect 54757 5315 54815 5321
rect 57146 5312 57152 5364
rect 57204 5352 57210 5364
rect 57701 5355 57759 5361
rect 57701 5352 57713 5355
rect 57204 5324 57713 5352
rect 57204 5312 57210 5324
rect 57701 5321 57713 5324
rect 57747 5321 57759 5355
rect 57701 5315 57759 5321
rect 57882 5312 57888 5364
rect 57940 5312 57946 5364
rect 58526 5312 58532 5364
rect 58584 5312 58590 5364
rect 52086 5244 52092 5296
rect 52144 5284 52150 5296
rect 53285 5287 53343 5293
rect 53285 5284 53297 5287
rect 52144 5256 53297 5284
rect 52144 5244 52150 5256
rect 53285 5253 53297 5256
rect 53331 5284 53343 5287
rect 55493 5287 55551 5293
rect 53331 5256 55444 5284
rect 53331 5253 53343 5256
rect 53285 5247 53343 5253
rect 49418 5176 49424 5228
rect 49476 5176 49482 5228
rect 49694 5176 49700 5228
rect 49752 5176 49758 5228
rect 50433 5219 50491 5225
rect 50433 5185 50445 5219
rect 50479 5216 50491 5219
rect 50522 5216 50528 5228
rect 50479 5188 50528 5216
rect 50479 5185 50491 5188
rect 50433 5179 50491 5185
rect 50522 5176 50528 5188
rect 50580 5176 50586 5228
rect 50700 5219 50758 5225
rect 50700 5185 50712 5219
rect 50746 5216 50758 5219
rect 52362 5216 52368 5228
rect 50746 5188 52368 5216
rect 50746 5185 50758 5188
rect 50700 5179 50758 5185
rect 52362 5176 52368 5188
rect 52420 5176 52426 5228
rect 54021 5219 54079 5225
rect 54021 5185 54033 5219
rect 54067 5216 54079 5219
rect 54478 5216 54484 5228
rect 54067 5188 54484 5216
rect 54067 5185 54079 5188
rect 54021 5179 54079 5185
rect 54478 5176 54484 5188
rect 54536 5176 54542 5228
rect 55416 5216 55444 5256
rect 55493 5253 55505 5287
rect 55539 5284 55551 5287
rect 57900 5284 57928 5312
rect 55539 5256 57928 5284
rect 55539 5253 55551 5256
rect 55493 5247 55551 5253
rect 56686 5216 56692 5228
rect 55416 5188 56692 5216
rect 56686 5176 56692 5188
rect 56744 5216 56750 5228
rect 56744 5188 56824 5216
rect 56744 5176 56750 5188
rect 48501 5151 48559 5157
rect 48501 5117 48513 5151
rect 48547 5117 48559 5151
rect 48501 5111 48559 5117
rect 48685 5151 48743 5157
rect 48685 5117 48697 5151
rect 48731 5117 48743 5151
rect 48685 5111 48743 5117
rect 48590 5080 48596 5092
rect 48056 5052 48596 5080
rect 47673 5043 47731 5049
rect 48590 5040 48596 5052
rect 48648 5040 48654 5092
rect 48700 5080 48728 5111
rect 48774 5108 48780 5160
rect 48832 5148 48838 5160
rect 49538 5151 49596 5157
rect 49538 5148 49550 5151
rect 48832 5120 49550 5148
rect 48832 5108 48838 5120
rect 49538 5117 49550 5120
rect 49584 5117 49596 5151
rect 49538 5111 49596 5117
rect 52270 5108 52276 5160
rect 52328 5148 52334 5160
rect 52549 5151 52607 5157
rect 52549 5148 52561 5151
rect 52328 5120 52561 5148
rect 52328 5108 52334 5120
rect 52549 5117 52561 5120
rect 52595 5148 52607 5151
rect 53650 5148 53656 5160
rect 52595 5120 53656 5148
rect 52595 5117 52607 5120
rect 52549 5111 52607 5117
rect 53650 5108 53656 5120
rect 53708 5108 53714 5160
rect 54202 5108 54208 5160
rect 54260 5108 54266 5160
rect 54941 5151 54999 5157
rect 54941 5117 54953 5151
rect 54987 5117 54999 5151
rect 54941 5111 54999 5117
rect 48700 5052 49096 5080
rect 45186 5012 45192 5024
rect 44284 4984 45192 5012
rect 44085 4975 44143 4981
rect 45186 4972 45192 4984
rect 45244 4972 45250 5024
rect 45741 5015 45799 5021
rect 45741 4981 45753 5015
rect 45787 5012 45799 5015
rect 47026 5012 47032 5024
rect 45787 4984 47032 5012
rect 45787 4981 45799 4984
rect 45741 4975 45799 4981
rect 47026 4972 47032 4984
rect 47084 4972 47090 5024
rect 47210 4972 47216 5024
rect 47268 5012 47274 5024
rect 47397 5015 47455 5021
rect 47397 5012 47409 5015
rect 47268 4984 47409 5012
rect 47268 4972 47274 4984
rect 47397 4981 47409 4984
rect 47443 4981 47455 5015
rect 49068 5012 49096 5052
rect 49142 5040 49148 5092
rect 49200 5040 49206 5092
rect 54956 5080 54984 5111
rect 55674 5108 55680 5160
rect 55732 5108 55738 5160
rect 56318 5108 56324 5160
rect 56376 5108 56382 5160
rect 56686 5080 56692 5092
rect 52932 5052 54892 5080
rect 54956 5052 56692 5080
rect 52932 5024 52960 5052
rect 49786 5012 49792 5024
rect 49068 4984 49792 5012
rect 47397 4975 47455 4981
rect 49786 4972 49792 4984
rect 49844 4972 49850 5024
rect 50338 4972 50344 5024
rect 50396 4972 50402 5024
rect 51074 4972 51080 5024
rect 51132 5012 51138 5024
rect 52086 5012 52092 5024
rect 51132 4984 52092 5012
rect 51132 4972 51138 4984
rect 52086 4972 52092 4984
rect 52144 4972 52150 5024
rect 52914 4972 52920 5024
rect 52972 4972 52978 5024
rect 53834 4972 53840 5024
rect 53892 4972 53898 5024
rect 54864 5012 54892 5052
rect 56686 5040 56692 5052
rect 56744 5040 56750 5092
rect 56796 5080 56824 5188
rect 57054 5176 57060 5228
rect 57112 5176 57118 5228
rect 57422 5176 57428 5228
rect 57480 5216 57486 5228
rect 57885 5219 57943 5225
rect 57885 5216 57897 5219
rect 57480 5188 57897 5216
rect 57480 5176 57486 5188
rect 57885 5185 57897 5188
rect 57931 5185 57943 5219
rect 57885 5179 57943 5185
rect 57054 5080 57060 5092
rect 56796 5052 57060 5080
rect 57054 5040 57060 5052
rect 57112 5040 57118 5092
rect 55582 5012 55588 5024
rect 54864 4984 55588 5012
rect 55582 4972 55588 4984
rect 55640 4972 55646 5024
rect 56226 4972 56232 5024
rect 56284 4972 56290 5024
rect 56962 4972 56968 5024
rect 57020 4972 57026 5024
rect 1104 4922 58880 4944
rect 1104 4870 8172 4922
rect 8224 4870 8236 4922
rect 8288 4870 8300 4922
rect 8352 4870 8364 4922
rect 8416 4870 8428 4922
rect 8480 4870 22616 4922
rect 22668 4870 22680 4922
rect 22732 4870 22744 4922
rect 22796 4870 22808 4922
rect 22860 4870 22872 4922
rect 22924 4870 37060 4922
rect 37112 4870 37124 4922
rect 37176 4870 37188 4922
rect 37240 4870 37252 4922
rect 37304 4870 37316 4922
rect 37368 4870 51504 4922
rect 51556 4870 51568 4922
rect 51620 4870 51632 4922
rect 51684 4870 51696 4922
rect 51748 4870 51760 4922
rect 51812 4870 58880 4922
rect 1104 4848 58880 4870
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 2222 4808 2228 4820
rect 2179 4780 2228 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 2222 4768 2228 4780
rect 2280 4808 2286 4820
rect 2685 4811 2743 4817
rect 2685 4808 2697 4811
rect 2280 4780 2697 4808
rect 2280 4768 2286 4780
rect 2685 4777 2697 4780
rect 2731 4777 2743 4811
rect 2685 4771 2743 4777
rect 2866 4768 2872 4820
rect 2924 4768 2930 4820
rect 3418 4768 3424 4820
rect 3476 4808 3482 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3476 4780 3985 4808
rect 3476 4768 3482 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 3973 4771 4031 4777
rect 5994 4768 6000 4820
rect 6052 4768 6058 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7708 4780 7849 4808
rect 7708 4768 7714 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 2590 4740 2596 4752
rect 2056 4712 2596 4740
rect 2056 4613 2084 4712
rect 2590 4700 2596 4712
rect 2648 4740 2654 4752
rect 4157 4743 4215 4749
rect 4157 4740 4169 4743
rect 2648 4712 4169 4740
rect 2648 4700 2654 4712
rect 4157 4709 4169 4712
rect 4203 4709 4215 4743
rect 4157 4703 4215 4709
rect 4522 4700 4528 4752
rect 4580 4740 4586 4752
rect 5442 4740 5448 4752
rect 4580 4712 5448 4740
rect 4580 4700 4586 4712
rect 5442 4700 5448 4712
rect 5500 4740 5506 4752
rect 5537 4743 5595 4749
rect 5537 4740 5549 4743
rect 5500 4712 5549 4740
rect 5500 4700 5506 4712
rect 5537 4709 5549 4712
rect 5583 4709 5595 4743
rect 5537 4703 5595 4709
rect 3326 4672 3332 4684
rect 2240 4644 3332 4672
rect 2240 4613 2268 4644
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5169 4675 5227 4681
rect 5169 4672 5181 4675
rect 5132 4644 5181 4672
rect 5132 4632 5138 4644
rect 5169 4641 5181 4644
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 2590 4604 2596 4616
rect 2372 4576 2596 4604
rect 2372 4564 2378 4576
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 2866 4564 2872 4616
rect 2924 4604 2930 4616
rect 3145 4607 3203 4613
rect 3145 4604 3157 4607
rect 2924 4576 3157 4604
rect 2924 4564 2930 4576
rect 3145 4573 3157 4576
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3467 4576 4016 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 2685 4539 2743 4545
rect 2685 4505 2697 4539
rect 2731 4536 2743 4539
rect 3050 4536 3056 4548
rect 2731 4508 3056 4536
rect 2731 4505 2743 4508
rect 2685 4499 2743 4505
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 3160 4536 3188 4567
rect 3988 4548 4016 4576
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 3160 4508 3801 4536
rect 3789 4505 3801 4508
rect 3835 4505 3847 4539
rect 3789 4499 3847 4505
rect 3970 4496 3976 4548
rect 4028 4545 4034 4548
rect 4028 4539 4047 4545
rect 4035 4505 4047 4539
rect 5184 4536 5212 4635
rect 5552 4604 5580 4703
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 6270 4740 6276 4752
rect 5684 4712 6276 4740
rect 5684 4700 5690 4712
rect 6270 4700 6276 4712
rect 6328 4749 6334 4752
rect 6328 4743 6377 4749
rect 6328 4709 6331 4743
rect 6365 4709 6377 4743
rect 6328 4703 6377 4709
rect 6457 4743 6515 4749
rect 6457 4709 6469 4743
rect 6503 4709 6515 4743
rect 7852 4740 7880 4771
rect 8018 4768 8024 4820
rect 8076 4768 8082 4820
rect 17494 4808 17500 4820
rect 8496 4780 8708 4808
rect 8496 4740 8524 4780
rect 7852 4712 8524 4740
rect 6457 4703 6515 4709
rect 6328 4700 6334 4703
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 6472 4672 6500 4703
rect 5776 4644 6500 4672
rect 6549 4675 6607 4681
rect 5776 4632 5782 4644
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5552 4576 6193 4604
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6564 4536 6592 4635
rect 8478 4632 8484 4684
rect 8536 4632 8542 4684
rect 8680 4681 8708 4780
rect 15948 4780 17500 4808
rect 10226 4700 10232 4752
rect 10284 4700 10290 4752
rect 10505 4743 10563 4749
rect 10505 4709 10517 4743
rect 10551 4740 10563 4743
rect 10551 4712 12480 4740
rect 10551 4709 10563 4712
rect 10505 4703 10563 4709
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8711 4644 9321 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 10870 4632 10876 4684
rect 10928 4632 10934 4684
rect 10962 4632 10968 4684
rect 11020 4632 11026 4684
rect 12452 4681 12480 4712
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11103 4644 11713 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 11701 4641 11713 4644
rect 11747 4672 11759 4675
rect 12437 4675 12495 4681
rect 11747 4644 11928 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 9122 4604 9128 4616
rect 7616 4576 9128 4604
rect 7616 4564 7622 4576
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10686 4604 10692 4616
rect 10459 4576 10692 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10888 4604 10916 4632
rect 11072 4604 11100 4635
rect 10888 4576 11100 4604
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11204 4576 11345 4604
rect 11204 4564 11210 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 5184 4508 6592 4536
rect 4028 4499 4047 4505
rect 4028 4496 4034 4499
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8018 4536 8024 4548
rect 7800 4508 8024 4536
rect 7800 4496 7806 4508
rect 8018 4496 8024 4508
rect 8076 4536 8082 4548
rect 8389 4539 8447 4545
rect 8389 4536 8401 4539
rect 8076 4508 8401 4536
rect 8076 4496 8082 4508
rect 8389 4505 8401 4508
rect 8435 4536 8447 4539
rect 10873 4539 10931 4545
rect 10873 4536 10885 4539
rect 8435 4508 10885 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 10873 4505 10885 4508
rect 10919 4536 10931 4539
rect 11606 4536 11612 4548
rect 10919 4508 11612 4536
rect 10919 4505 10931 4508
rect 10873 4499 10931 4505
rect 11606 4496 11612 4508
rect 11664 4536 11670 4548
rect 11808 4536 11836 4564
rect 11664 4508 11836 4536
rect 11900 4536 11928 4644
rect 12437 4641 12449 4675
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 14826 4632 14832 4684
rect 14884 4672 14890 4684
rect 15948 4681 15976 4780
rect 17494 4768 17500 4780
rect 17552 4808 17558 4820
rect 18414 4808 18420 4820
rect 17552 4780 18420 4808
rect 17552 4768 17558 4780
rect 18414 4768 18420 4780
rect 18472 4808 18478 4820
rect 18472 4780 19288 4808
rect 18472 4768 18478 4780
rect 19260 4681 19288 4780
rect 19978 4768 19984 4820
rect 20036 4808 20042 4820
rect 21910 4808 21916 4820
rect 20036 4780 21916 4808
rect 20036 4768 20042 4780
rect 21910 4768 21916 4780
rect 21968 4808 21974 4820
rect 22281 4811 22339 4817
rect 22281 4808 22293 4811
rect 21968 4780 22293 4808
rect 21968 4768 21974 4780
rect 22281 4777 22293 4780
rect 22327 4777 22339 4811
rect 22281 4771 22339 4777
rect 26326 4768 26332 4820
rect 26384 4808 26390 4820
rect 26789 4811 26847 4817
rect 26789 4808 26801 4811
rect 26384 4780 26801 4808
rect 26384 4768 26390 4780
rect 26789 4777 26801 4780
rect 26835 4777 26847 4811
rect 29730 4808 29736 4820
rect 26789 4771 26847 4777
rect 27540 4780 29736 4808
rect 23032 4712 25452 4740
rect 23032 4684 23060 4712
rect 15933 4675 15991 4681
rect 15933 4672 15945 4675
rect 14884 4644 15945 4672
rect 14884 4632 14890 4644
rect 15933 4641 15945 4644
rect 15979 4641 15991 4675
rect 15933 4635 15991 4641
rect 19245 4675 19303 4681
rect 19245 4641 19257 4675
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 14090 4604 14096 4616
rect 13403 4576 14096 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 15010 4564 15016 4616
rect 15068 4564 15074 4616
rect 16200 4607 16258 4613
rect 16200 4573 16212 4607
rect 16246 4604 16258 4607
rect 17126 4604 17132 4616
rect 16246 4576 17132 4604
rect 16246 4573 16258 4576
rect 16200 4567 16258 4573
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17328 4576 17417 4604
rect 16022 4536 16028 4548
rect 11900 4508 16028 4536
rect 11664 4496 11670 4508
rect 16022 4496 16028 4508
rect 16080 4536 16086 4548
rect 17218 4536 17224 4548
rect 16080 4508 17224 4536
rect 16080 4496 16086 4508
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 2958 4428 2964 4480
rect 3016 4428 3022 4480
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 4709 4471 4767 4477
rect 4709 4437 4721 4471
rect 4755 4468 4767 4471
rect 4798 4468 4804 4480
rect 4755 4440 4804 4468
rect 4755 4437 4767 4440
rect 4709 4431 4767 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5077 4471 5135 4477
rect 5077 4437 5089 4471
rect 5123 4468 5135 4471
rect 5902 4468 5908 4480
rect 5123 4440 5908 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6825 4471 6883 4477
rect 6825 4437 6837 4471
rect 6871 4468 6883 4471
rect 11238 4468 11244 4480
rect 6871 4440 11244 4468
rect 6871 4437 6883 4440
rect 6825 4431 6883 4437
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 11848 4440 13093 4468
rect 11848 4428 11854 4440
rect 13081 4437 13093 4440
rect 13127 4437 13139 4471
rect 13081 4431 13139 4437
rect 13906 4428 13912 4480
rect 13964 4428 13970 4480
rect 14826 4428 14832 4480
rect 14884 4428 14890 4480
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 15252 4440 15577 4468
rect 15252 4428 15258 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 15565 4431 15623 4437
rect 15838 4428 15844 4480
rect 15896 4468 15902 4480
rect 17328 4477 17356 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17678 4564 17684 4616
rect 17736 4604 17742 4616
rect 18046 4604 18052 4616
rect 17736 4576 18052 4604
rect 17736 4564 17742 4576
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4573 18567 4607
rect 19260 4604 19288 4635
rect 23014 4632 23020 4684
rect 23072 4632 23078 4684
rect 23934 4632 23940 4684
rect 23992 4632 23998 4684
rect 24118 4632 24124 4684
rect 24176 4672 24182 4684
rect 24394 4672 24400 4684
rect 24176 4644 24400 4672
rect 24176 4632 24182 4644
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 25038 4632 25044 4684
rect 25096 4632 25102 4684
rect 25424 4681 25452 4712
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4641 25191 4675
rect 25133 4635 25191 4641
rect 25409 4675 25467 4681
rect 25409 4641 25421 4675
rect 25455 4641 25467 4675
rect 25409 4635 25467 4641
rect 20714 4604 20720 4616
rect 19260 4576 20720 4604
rect 18509 4567 18567 4573
rect 18524 4536 18552 4567
rect 20714 4564 20720 4576
rect 20772 4604 20778 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20772 4576 20913 4604
rect 20772 4564 20778 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 22002 4564 22008 4616
rect 22060 4604 22066 4616
rect 22373 4607 22431 4613
rect 22373 4604 22385 4607
rect 22060 4576 22385 4604
rect 22060 4564 22066 4576
rect 22373 4573 22385 4576
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 23385 4607 23443 4613
rect 23385 4573 23397 4607
rect 23431 4604 23443 4607
rect 25148 4604 25176 4635
rect 23431 4576 25176 4604
rect 25424 4604 25452 4635
rect 26234 4604 26240 4616
rect 25424 4576 26240 4604
rect 23431 4573 23443 4576
rect 23385 4567 23443 4573
rect 19512 4539 19570 4545
rect 18524 4508 19472 4536
rect 17313 4471 17371 4477
rect 17313 4468 17325 4471
rect 15896 4440 17325 4468
rect 15896 4428 15902 4440
rect 17313 4437 17325 4440
rect 17359 4437 17371 4471
rect 17313 4431 17371 4437
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17828 4440 18061 4468
rect 17828 4428 17834 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18049 4431 18107 4437
rect 19058 4428 19064 4480
rect 19116 4428 19122 4480
rect 19444 4468 19472 4508
rect 19512 4505 19524 4539
rect 19558 4536 19570 4539
rect 19978 4536 19984 4548
rect 19558 4508 19984 4536
rect 19558 4505 19570 4508
rect 19512 4499 19570 4505
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 21168 4539 21226 4545
rect 21168 4505 21180 4539
rect 21214 4536 21226 4539
rect 23017 4539 23075 4545
rect 23017 4536 23029 4539
rect 21214 4508 23029 4536
rect 21214 4505 21226 4508
rect 21168 4499 21226 4505
rect 23017 4505 23029 4508
rect 23063 4505 23075 4539
rect 23017 4499 23075 4505
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24762 4536 24768 4548
rect 23891 4508 24768 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24762 4496 24768 4508
rect 24820 4536 24826 4548
rect 25148 4536 25176 4576
rect 26234 4564 26240 4576
rect 26292 4564 26298 4616
rect 25498 4536 25504 4548
rect 24820 4508 24992 4536
rect 25148 4508 25504 4536
rect 24820 4496 24826 4508
rect 20625 4471 20683 4477
rect 20625 4468 20637 4471
rect 19444 4440 20637 4468
rect 20625 4437 20637 4440
rect 20671 4468 20683 4471
rect 20806 4468 20812 4480
rect 20671 4440 20812 4468
rect 20671 4437 20683 4440
rect 20625 4431 20683 4437
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 23474 4428 23480 4480
rect 23532 4428 23538 4480
rect 24578 4428 24584 4480
rect 24636 4428 24642 4480
rect 24964 4477 24992 4508
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 25676 4539 25734 4545
rect 25676 4505 25688 4539
rect 25722 4536 25734 4539
rect 26418 4536 26424 4548
rect 25722 4508 26424 4536
rect 25722 4505 25734 4508
rect 25676 4499 25734 4505
rect 26418 4496 26424 4508
rect 26476 4496 26482 4548
rect 24949 4471 25007 4477
rect 24949 4437 24961 4471
rect 24995 4468 25007 4471
rect 26326 4468 26332 4480
rect 24995 4440 26332 4468
rect 24995 4437 25007 4440
rect 24949 4431 25007 4437
rect 26326 4428 26332 4440
rect 26384 4428 26390 4480
rect 26602 4428 26608 4480
rect 26660 4468 26666 4480
rect 27157 4471 27215 4477
rect 27157 4468 27169 4471
rect 26660 4440 27169 4468
rect 26660 4428 26666 4440
rect 27157 4437 27169 4440
rect 27203 4468 27215 4471
rect 27540 4468 27568 4780
rect 29730 4768 29736 4780
rect 29788 4768 29794 4820
rect 33226 4808 33232 4820
rect 31726 4780 33232 4808
rect 27614 4700 27620 4752
rect 27672 4740 27678 4752
rect 28077 4743 28135 4749
rect 28077 4740 28089 4743
rect 27672 4712 28089 4740
rect 27672 4700 27678 4712
rect 28077 4709 28089 4712
rect 28123 4709 28135 4743
rect 28077 4703 28135 4709
rect 31202 4700 31208 4752
rect 31260 4700 31266 4752
rect 27706 4632 27712 4684
rect 27764 4672 27770 4684
rect 31726 4672 31754 4780
rect 33226 4768 33232 4780
rect 33284 4768 33290 4820
rect 33594 4768 33600 4820
rect 33652 4768 33658 4820
rect 34698 4768 34704 4820
rect 34756 4808 34762 4820
rect 34756 4780 35940 4808
rect 34756 4768 34762 4780
rect 32030 4700 32036 4752
rect 32088 4700 32094 4752
rect 34606 4740 34612 4752
rect 34256 4712 34612 4740
rect 27764 4644 31754 4672
rect 31849 4675 31907 4681
rect 27764 4632 27770 4644
rect 31849 4641 31861 4675
rect 31895 4641 31907 4675
rect 31849 4635 31907 4641
rect 27617 4607 27675 4613
rect 27617 4573 27629 4607
rect 27663 4604 27675 4607
rect 27724 4604 27752 4632
rect 27663 4576 27752 4604
rect 27663 4573 27675 4576
rect 27617 4567 27675 4573
rect 27982 4564 27988 4616
rect 28040 4604 28046 4616
rect 28261 4607 28319 4613
rect 28261 4604 28273 4607
rect 28040 4576 28273 4604
rect 28040 4564 28046 4576
rect 28261 4573 28273 4576
rect 28307 4573 28319 4607
rect 28261 4567 28319 4573
rect 28813 4607 28871 4613
rect 28813 4573 28825 4607
rect 28859 4604 28871 4607
rect 29178 4604 29184 4616
rect 28859 4576 29184 4604
rect 28859 4573 28871 4576
rect 28813 4567 28871 4573
rect 29178 4564 29184 4576
rect 29236 4564 29242 4616
rect 29546 4564 29552 4616
rect 29604 4604 29610 4616
rect 29733 4607 29791 4613
rect 29733 4604 29745 4607
rect 29604 4576 29745 4604
rect 29604 4564 29610 4576
rect 29733 4573 29745 4576
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 30558 4564 30564 4616
rect 30616 4604 30622 4616
rect 31386 4604 31392 4616
rect 30616 4576 31392 4604
rect 30616 4564 30622 4576
rect 31386 4564 31392 4576
rect 31444 4564 31450 4616
rect 31478 4536 31484 4548
rect 28644 4508 31484 4536
rect 28644 4477 28672 4508
rect 31478 4496 31484 4508
rect 31536 4496 31542 4548
rect 31573 4539 31631 4545
rect 31573 4505 31585 4539
rect 31619 4536 31631 4539
rect 31754 4536 31760 4548
rect 31619 4508 31760 4536
rect 31619 4505 31631 4508
rect 31573 4499 31631 4505
rect 31754 4496 31760 4508
rect 31812 4496 31818 4548
rect 31864 4536 31892 4635
rect 32048 4613 32076 4700
rect 34054 4632 34060 4684
rect 34112 4632 34118 4684
rect 34256 4681 34284 4712
rect 34606 4700 34612 4712
rect 34664 4700 34670 4752
rect 35912 4740 35940 4780
rect 35986 4768 35992 4820
rect 36044 4808 36050 4820
rect 36081 4811 36139 4817
rect 36081 4808 36093 4811
rect 36044 4780 36093 4808
rect 36044 4768 36050 4780
rect 36081 4777 36093 4780
rect 36127 4777 36139 4811
rect 36906 4808 36912 4820
rect 36081 4771 36139 4777
rect 36648 4780 36912 4808
rect 36446 4740 36452 4752
rect 35912 4712 36452 4740
rect 36446 4700 36452 4712
rect 36504 4700 36510 4752
rect 34241 4675 34299 4681
rect 34241 4641 34253 4675
rect 34287 4641 34299 4675
rect 34241 4635 34299 4641
rect 34422 4632 34428 4684
rect 34480 4672 34486 4684
rect 36648 4681 36676 4780
rect 36906 4768 36912 4780
rect 36964 4768 36970 4820
rect 37108 4780 39344 4808
rect 36814 4700 36820 4752
rect 36872 4740 36878 4752
rect 37001 4743 37059 4749
rect 37001 4740 37013 4743
rect 36872 4712 37013 4740
rect 36872 4700 36878 4712
rect 37001 4709 37013 4712
rect 37047 4709 37059 4743
rect 37001 4703 37059 4709
rect 34701 4675 34759 4681
rect 34701 4672 34713 4675
rect 34480 4644 34713 4672
rect 34480 4632 34486 4644
rect 34701 4641 34713 4644
rect 34747 4641 34759 4675
rect 34701 4635 34759 4641
rect 36633 4675 36691 4681
rect 36633 4641 36645 4675
rect 36679 4641 36691 4675
rect 36633 4635 36691 4641
rect 36725 4675 36783 4681
rect 36725 4641 36737 4675
rect 36771 4672 36783 4675
rect 37108 4672 37136 4780
rect 38286 4700 38292 4752
rect 38344 4700 38350 4752
rect 36771 4644 37136 4672
rect 36771 4641 36783 4644
rect 36725 4635 36783 4641
rect 32033 4607 32091 4613
rect 32033 4573 32045 4607
rect 32079 4573 32091 4607
rect 32033 4567 32091 4573
rect 32674 4564 32680 4616
rect 32732 4604 32738 4616
rect 32861 4607 32919 4613
rect 32861 4604 32873 4607
rect 32732 4576 32873 4604
rect 32732 4564 32738 4576
rect 32861 4573 32873 4576
rect 32907 4604 32919 4607
rect 34716 4604 34744 4635
rect 35802 4604 35808 4616
rect 32907 4576 34652 4604
rect 34716 4576 35808 4604
rect 32907 4573 32919 4576
rect 32861 4567 32919 4573
rect 32692 4536 32720 4564
rect 31864 4508 32720 4536
rect 33318 4496 33324 4548
rect 33376 4496 33382 4548
rect 34624 4536 34652 4576
rect 35802 4564 35808 4576
rect 35860 4564 35866 4616
rect 36538 4564 36544 4616
rect 36596 4564 36602 4616
rect 34968 4539 35026 4545
rect 34624 4508 34928 4536
rect 27893 4471 27951 4477
rect 27893 4468 27905 4471
rect 27203 4440 27905 4468
rect 27203 4437 27215 4440
rect 27157 4431 27215 4437
rect 27893 4437 27905 4440
rect 27939 4437 27951 4471
rect 27893 4431 27951 4437
rect 28629 4471 28687 4477
rect 28629 4437 28641 4471
rect 28675 4437 28687 4471
rect 28629 4431 28687 4437
rect 29362 4428 29368 4480
rect 29420 4428 29426 4480
rect 30282 4428 30288 4480
rect 30340 4468 30346 4480
rect 30377 4471 30435 4477
rect 30377 4468 30389 4471
rect 30340 4440 30389 4468
rect 30340 4428 30346 4440
rect 30377 4437 30389 4440
rect 30423 4437 30435 4471
rect 30377 4431 30435 4437
rect 31110 4428 31116 4480
rect 31168 4428 31174 4480
rect 31665 4471 31723 4477
rect 31665 4437 31677 4471
rect 31711 4468 31723 4471
rect 31938 4468 31944 4480
rect 31711 4440 31944 4468
rect 31711 4437 31723 4440
rect 31665 4431 31723 4437
rect 31938 4428 31944 4440
rect 31996 4428 32002 4480
rect 33410 4428 33416 4480
rect 33468 4428 33474 4480
rect 33962 4428 33968 4480
rect 34020 4428 34026 4480
rect 34900 4468 34928 4508
rect 34968 4505 34980 4539
rect 35014 4536 35026 4539
rect 35894 4536 35900 4548
rect 35014 4508 35900 4536
rect 35014 4505 35026 4508
rect 34968 4499 35026 4505
rect 35894 4496 35900 4508
rect 35952 4496 35958 4548
rect 36740 4536 36768 4635
rect 37274 4632 37280 4684
rect 37332 4672 37338 4684
rect 37645 4675 37703 4681
rect 37645 4672 37657 4675
rect 37332 4644 37657 4672
rect 37332 4632 37338 4644
rect 37645 4641 37657 4644
rect 37691 4672 37703 4675
rect 38304 4672 38332 4700
rect 37691 4644 38332 4672
rect 39316 4672 39344 4780
rect 39574 4768 39580 4820
rect 39632 4768 39638 4820
rect 39669 4811 39727 4817
rect 39669 4777 39681 4811
rect 39715 4808 39727 4811
rect 40034 4808 40040 4820
rect 39715 4780 40040 4808
rect 39715 4777 39727 4780
rect 39669 4771 39727 4777
rect 40034 4768 40040 4780
rect 40092 4808 40098 4820
rect 40310 4808 40316 4820
rect 40092 4780 40316 4808
rect 40092 4768 40098 4780
rect 40310 4768 40316 4780
rect 40368 4768 40374 4820
rect 42337 4811 42395 4817
rect 42337 4808 42349 4811
rect 40512 4780 42349 4808
rect 39592 4740 39620 4768
rect 40512 4740 40540 4780
rect 42337 4777 42349 4780
rect 42383 4777 42395 4811
rect 42337 4771 42395 4777
rect 39592 4712 40540 4740
rect 39942 4672 39948 4684
rect 39316 4644 39948 4672
rect 37691 4641 37703 4644
rect 37645 4635 37703 4641
rect 39942 4632 39948 4644
rect 40000 4632 40006 4684
rect 40494 4632 40500 4684
rect 40552 4632 40558 4684
rect 40770 4672 40776 4684
rect 40696 4644 40776 4672
rect 36814 4564 36820 4616
rect 36872 4604 36878 4616
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 36872 4576 37841 4604
rect 36872 4564 36878 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 38010 4564 38016 4616
rect 38068 4564 38074 4616
rect 38289 4607 38347 4613
rect 38289 4573 38301 4607
rect 38335 4604 38347 4607
rect 40696 4604 40724 4644
rect 40770 4632 40776 4644
rect 40828 4672 40834 4684
rect 40957 4675 41015 4681
rect 40957 4672 40969 4675
rect 40828 4644 40969 4672
rect 40828 4632 40834 4644
rect 40957 4641 40969 4644
rect 41003 4672 41015 4675
rect 42352 4672 42380 4771
rect 43070 4768 43076 4820
rect 43128 4768 43134 4820
rect 43346 4768 43352 4820
rect 43404 4768 43410 4820
rect 43990 4768 43996 4820
rect 44048 4808 44054 4820
rect 44048 4780 45784 4808
rect 44048 4768 44054 4780
rect 44177 4743 44235 4749
rect 44177 4709 44189 4743
rect 44223 4709 44235 4743
rect 44177 4703 44235 4709
rect 44545 4743 44603 4749
rect 44545 4709 44557 4743
rect 44591 4740 44603 4743
rect 44910 4740 44916 4752
rect 44591 4712 44916 4740
rect 44591 4709 44603 4712
rect 44545 4703 44603 4709
rect 42429 4675 42487 4681
rect 42429 4672 42441 4675
rect 41003 4644 41092 4672
rect 42352 4644 42441 4672
rect 41003 4641 41015 4644
rect 40957 4635 41015 4641
rect 38335 4576 40724 4604
rect 38335 4573 38347 4576
rect 38289 4567 38347 4573
rect 36004 4508 36768 4536
rect 36004 4468 36032 4508
rect 37550 4496 37556 4548
rect 37608 4536 37614 4548
rect 38304 4536 38332 4567
rect 40862 4564 40868 4616
rect 40920 4564 40926 4616
rect 41064 4604 41092 4644
rect 42429 4641 42441 4644
rect 42475 4641 42487 4675
rect 42429 4635 42487 4641
rect 43898 4632 43904 4684
rect 43956 4632 43962 4684
rect 44082 4632 44088 4684
rect 44140 4632 44146 4684
rect 44192 4672 44220 4703
rect 44910 4700 44916 4712
rect 44968 4700 44974 4752
rect 45462 4740 45468 4752
rect 45020 4712 45468 4740
rect 44634 4672 44640 4684
rect 44192 4644 44640 4672
rect 44634 4632 44640 4644
rect 44692 4632 44698 4684
rect 45020 4681 45048 4712
rect 45462 4700 45468 4712
rect 45520 4700 45526 4752
rect 45005 4675 45063 4681
rect 45005 4641 45017 4675
rect 45051 4641 45063 4675
rect 45005 4635 45063 4641
rect 45189 4675 45247 4681
rect 45189 4641 45201 4675
rect 45235 4672 45247 4675
rect 45554 4672 45560 4684
rect 45235 4644 45560 4672
rect 45235 4641 45247 4644
rect 45189 4635 45247 4641
rect 45554 4632 45560 4644
rect 45612 4632 45618 4684
rect 45646 4632 45652 4684
rect 45704 4632 45710 4684
rect 45756 4672 45784 4780
rect 46198 4768 46204 4820
rect 46256 4808 46262 4820
rect 46845 4811 46903 4817
rect 46845 4808 46857 4811
rect 46256 4780 46857 4808
rect 46256 4768 46262 4780
rect 46845 4777 46857 4780
rect 46891 4777 46903 4811
rect 46845 4771 46903 4777
rect 48317 4811 48375 4817
rect 48317 4777 48329 4811
rect 48363 4777 48375 4811
rect 48317 4771 48375 4777
rect 48409 4811 48467 4817
rect 48409 4777 48421 4811
rect 48455 4808 48467 4811
rect 48682 4808 48688 4820
rect 48455 4780 48688 4808
rect 48455 4777 48467 4780
rect 48409 4771 48467 4777
rect 48222 4700 48228 4752
rect 48280 4740 48286 4752
rect 48332 4740 48360 4771
rect 48682 4768 48688 4780
rect 48740 4768 48746 4820
rect 48774 4768 48780 4820
rect 48832 4768 48838 4820
rect 50062 4808 50068 4820
rect 48976 4780 50068 4808
rect 48792 4740 48820 4768
rect 48280 4712 48820 4740
rect 48280 4700 48286 4712
rect 45925 4675 45983 4681
rect 45925 4672 45937 4675
rect 45756 4644 45937 4672
rect 45925 4641 45937 4644
rect 45971 4641 45983 4675
rect 45925 4635 45983 4641
rect 46201 4675 46259 4681
rect 46201 4641 46213 4675
rect 46247 4672 46259 4675
rect 46382 4672 46388 4684
rect 46247 4644 46388 4672
rect 46247 4641 46259 4644
rect 46201 4635 46259 4641
rect 46382 4632 46388 4644
rect 46440 4632 46446 4684
rect 46934 4632 46940 4684
rect 46992 4632 46998 4684
rect 48498 4632 48504 4684
rect 48556 4672 48562 4684
rect 48976 4681 49004 4780
rect 50062 4768 50068 4780
rect 50120 4768 50126 4820
rect 50338 4768 50344 4820
rect 50396 4768 50402 4820
rect 51813 4811 51871 4817
rect 51813 4777 51825 4811
rect 51859 4808 51871 4811
rect 52270 4808 52276 4820
rect 51859 4780 52276 4808
rect 51859 4777 51871 4780
rect 51813 4771 51871 4777
rect 52270 4768 52276 4780
rect 52328 4768 52334 4820
rect 54018 4768 54024 4820
rect 54076 4808 54082 4820
rect 54941 4811 54999 4817
rect 54941 4808 54953 4811
rect 54076 4780 54953 4808
rect 54076 4768 54082 4780
rect 54941 4777 54953 4780
rect 54987 4777 54999 4811
rect 54941 4771 54999 4777
rect 56318 4768 56324 4820
rect 56376 4768 56382 4820
rect 56502 4768 56508 4820
rect 56560 4808 56566 4820
rect 56560 4780 57192 4808
rect 56560 4768 56566 4780
rect 48961 4675 49019 4681
rect 48961 4672 48973 4675
rect 48556 4644 48973 4672
rect 48556 4632 48562 4644
rect 48961 4641 48973 4644
rect 49007 4641 49019 4675
rect 48961 4635 49019 4641
rect 49329 4675 49387 4681
rect 49329 4641 49341 4675
rect 49375 4672 49387 4675
rect 49418 4672 49424 4684
rect 49375 4644 49424 4672
rect 49375 4641 49387 4644
rect 49329 4635 49387 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 50356 4672 50384 4768
rect 52549 4743 52607 4749
rect 52549 4709 52561 4743
rect 52595 4740 52607 4743
rect 52595 4712 53420 4740
rect 52595 4709 52607 4712
rect 52549 4703 52607 4709
rect 50617 4675 50675 4681
rect 50617 4672 50629 4675
rect 50356 4644 50629 4672
rect 50617 4641 50629 4644
rect 50663 4641 50675 4675
rect 50617 4635 50675 4641
rect 50801 4675 50859 4681
rect 50801 4641 50813 4675
rect 50847 4672 50859 4675
rect 52914 4672 52920 4684
rect 50847 4644 52920 4672
rect 50847 4641 50859 4644
rect 50801 4635 50859 4641
rect 42702 4604 42708 4616
rect 41064 4576 42708 4604
rect 42702 4564 42708 4576
rect 42760 4564 42766 4616
rect 43809 4607 43867 4613
rect 43809 4573 43821 4607
rect 43855 4604 43867 4607
rect 44100 4604 44128 4632
rect 43855 4576 44128 4604
rect 43855 4573 43867 4576
rect 43809 4567 43867 4573
rect 44174 4564 44180 4616
rect 44232 4564 44238 4616
rect 44361 4607 44419 4613
rect 44361 4573 44373 4607
rect 44407 4573 44419 4607
rect 44361 4567 44419 4573
rect 44729 4607 44787 4613
rect 44729 4573 44741 4607
rect 44775 4604 44787 4607
rect 45370 4604 45376 4616
rect 44775 4576 45376 4604
rect 44775 4573 44787 4576
rect 44729 4567 44787 4573
rect 37608 4508 38332 4536
rect 38556 4539 38614 4545
rect 37608 4496 37614 4508
rect 38556 4505 38568 4539
rect 38602 4536 38614 4539
rect 39206 4536 39212 4548
rect 38602 4508 39212 4536
rect 38602 4505 38614 4508
rect 38556 4499 38614 4505
rect 39206 4496 39212 4508
rect 39264 4496 39270 4548
rect 40218 4496 40224 4548
rect 40276 4496 40282 4548
rect 41224 4539 41282 4545
rect 41224 4505 41236 4539
rect 41270 4536 41282 4539
rect 41966 4536 41972 4548
rect 41270 4508 41972 4536
rect 41270 4505 41282 4508
rect 41224 4499 41282 4505
rect 41966 4496 41972 4508
rect 42024 4496 42030 4548
rect 42058 4496 42064 4548
rect 42116 4536 42122 4548
rect 43717 4539 43775 4545
rect 42116 4508 42288 4536
rect 42116 4496 42122 4508
rect 34900 4440 36032 4468
rect 36078 4428 36084 4480
rect 36136 4468 36142 4480
rect 36173 4471 36231 4477
rect 36173 4468 36185 4471
rect 36136 4440 36185 4468
rect 36136 4428 36142 4440
rect 36173 4437 36185 4440
rect 36219 4437 36231 4471
rect 36173 4431 36231 4437
rect 36262 4428 36268 4480
rect 36320 4468 36326 4480
rect 37369 4471 37427 4477
rect 37369 4468 37381 4471
rect 36320 4440 37381 4468
rect 36320 4428 36326 4440
rect 37369 4437 37381 4440
rect 37415 4437 37427 4471
rect 37369 4431 37427 4437
rect 37458 4428 37464 4480
rect 37516 4428 37522 4480
rect 38194 4428 38200 4480
rect 38252 4428 38258 4480
rect 39850 4428 39856 4480
rect 39908 4428 39914 4480
rect 40310 4428 40316 4480
rect 40368 4428 40374 4480
rect 40681 4471 40739 4477
rect 40681 4437 40693 4471
rect 40727 4468 40739 4471
rect 41874 4468 41880 4480
rect 40727 4440 41880 4468
rect 40727 4437 40739 4440
rect 40681 4431 40739 4437
rect 41874 4428 41880 4440
rect 41932 4428 41938 4480
rect 42260 4468 42288 4508
rect 43717 4505 43729 4539
rect 43763 4536 43775 4539
rect 44192 4536 44220 4564
rect 43763 4508 44220 4536
rect 44376 4536 44404 4567
rect 45370 4564 45376 4576
rect 45428 4564 45434 4616
rect 46014 4564 46020 4616
rect 46072 4613 46078 4616
rect 47210 4613 47216 4616
rect 46072 4607 46100 4613
rect 46088 4573 46100 4607
rect 47204 4604 47216 4613
rect 47171 4576 47216 4604
rect 46072 4567 46100 4573
rect 47204 4567 47216 4576
rect 46072 4564 46078 4567
rect 47210 4564 47216 4567
rect 47268 4564 47274 4616
rect 48406 4564 48412 4616
rect 48464 4604 48470 4616
rect 48777 4607 48835 4613
rect 48777 4604 48789 4607
rect 48464 4576 48789 4604
rect 48464 4564 48470 4576
rect 48777 4573 48789 4576
rect 48823 4604 48835 4607
rect 49234 4604 49240 4616
rect 48823 4576 49240 4604
rect 48823 4573 48835 4576
rect 48777 4567 48835 4573
rect 49234 4564 49240 4576
rect 49292 4564 49298 4616
rect 50816 4604 50844 4635
rect 52914 4632 52920 4644
rect 52972 4632 52978 4684
rect 53098 4632 53104 4684
rect 53156 4632 53162 4684
rect 53392 4681 53420 4712
rect 55692 4712 56263 4740
rect 53377 4675 53435 4681
rect 53377 4641 53389 4675
rect 53423 4641 53435 4675
rect 55692 4672 55720 4712
rect 53377 4635 53435 4641
rect 53944 4644 55720 4672
rect 49344 4576 50844 4604
rect 44376 4508 45232 4536
rect 43763 4505 43775 4508
rect 43717 4499 43775 4505
rect 43622 4468 43628 4480
rect 42260 4440 43628 4468
rect 43622 4428 43628 4440
rect 43680 4428 43686 4480
rect 45204 4468 45232 4508
rect 47118 4496 47124 4548
rect 47176 4536 47182 4548
rect 49344 4536 49372 4576
rect 51442 4564 51448 4616
rect 51500 4564 51506 4616
rect 53282 4604 53288 4616
rect 52932 4576 53288 4604
rect 47176 4508 49372 4536
rect 50525 4539 50583 4545
rect 47176 4496 47182 4508
rect 50525 4505 50537 4539
rect 50571 4536 50583 4539
rect 50706 4536 50712 4548
rect 50571 4508 50712 4536
rect 50571 4505 50583 4508
rect 50525 4499 50583 4505
rect 50706 4496 50712 4508
rect 50764 4496 50770 4548
rect 52932 4545 52960 4576
rect 53282 4564 53288 4576
rect 53340 4604 53346 4616
rect 53944 4604 53972 4644
rect 53340 4576 53972 4604
rect 53340 4564 53346 4576
rect 54018 4564 54024 4616
rect 54076 4564 54082 4616
rect 54110 4564 54116 4616
rect 54168 4564 54174 4616
rect 55692 4613 55720 4644
rect 55953 4675 56011 4681
rect 55953 4641 55965 4675
rect 55999 4641 56011 4675
rect 56235 4672 56263 4712
rect 56778 4672 56784 4684
rect 56235 4644 56784 4672
rect 55953 4635 56011 4641
rect 55125 4607 55183 4613
rect 55125 4573 55137 4607
rect 55171 4573 55183 4607
rect 55125 4567 55183 4573
rect 55677 4607 55735 4613
rect 55677 4573 55689 4607
rect 55723 4573 55735 4607
rect 55968 4604 55996 4635
rect 56778 4632 56784 4644
rect 56836 4632 56842 4684
rect 56965 4675 57023 4681
rect 56965 4641 56977 4675
rect 57011 4672 57023 4675
rect 57054 4672 57060 4684
rect 57011 4644 57060 4672
rect 57011 4641 57023 4644
rect 56965 4635 57023 4641
rect 57054 4632 57060 4644
rect 57112 4632 57118 4684
rect 56042 4604 56048 4616
rect 55968 4576 56048 4604
rect 55677 4567 55735 4573
rect 52917 4539 52975 4545
rect 52917 4505 52929 4539
rect 52963 4505 52975 4539
rect 52917 4499 52975 4505
rect 53009 4539 53067 4545
rect 53009 4505 53021 4539
rect 53055 4536 53067 4539
rect 54757 4539 54815 4545
rect 54757 4536 54769 4539
rect 53055 4508 54769 4536
rect 53055 4505 53067 4508
rect 53009 4499 53067 4505
rect 54757 4505 54769 4508
rect 54803 4505 54815 4539
rect 55140 4536 55168 4567
rect 56042 4564 56048 4576
rect 56100 4564 56106 4616
rect 56226 4564 56232 4616
rect 56284 4604 56290 4616
rect 57164 4613 57192 4780
rect 56689 4607 56747 4613
rect 56689 4604 56701 4607
rect 56284 4576 56701 4604
rect 56284 4564 56290 4576
rect 56689 4573 56701 4576
rect 56735 4573 56747 4607
rect 56689 4567 56747 4573
rect 57149 4607 57207 4613
rect 57149 4573 57161 4607
rect 57195 4573 57207 4607
rect 57149 4567 57207 4573
rect 58345 4539 58403 4545
rect 55140 4508 55996 4536
rect 54757 4499 54815 4505
rect 45646 4468 45652 4480
rect 45204 4440 45652 4468
rect 45646 4428 45652 4440
rect 45704 4428 45710 4480
rect 48869 4471 48927 4477
rect 48869 4437 48881 4471
rect 48915 4468 48927 4471
rect 49881 4471 49939 4477
rect 49881 4468 49893 4471
rect 48915 4440 49893 4468
rect 48915 4437 48927 4440
rect 48869 4431 48927 4437
rect 49881 4437 49893 4440
rect 49927 4437 49939 4471
rect 49881 4431 49939 4437
rect 50154 4428 50160 4480
rect 50212 4428 50218 4480
rect 51258 4428 51264 4480
rect 51316 4428 51322 4480
rect 52086 4428 52092 4480
rect 52144 4428 52150 4480
rect 55306 4428 55312 4480
rect 55364 4428 55370 4480
rect 55766 4428 55772 4480
rect 55824 4428 55830 4480
rect 55968 4468 55996 4508
rect 58345 4505 58357 4539
rect 58391 4536 58403 4539
rect 59078 4536 59084 4548
rect 58391 4508 59084 4536
rect 58391 4505 58403 4508
rect 58345 4499 58403 4505
rect 59078 4496 59084 4508
rect 59136 4496 59142 4548
rect 58526 4468 58532 4480
rect 55968 4440 58532 4468
rect 58526 4428 58532 4440
rect 58584 4428 58590 4480
rect 1104 4378 59040 4400
rect 1104 4326 15394 4378
rect 15446 4326 15458 4378
rect 15510 4326 15522 4378
rect 15574 4326 15586 4378
rect 15638 4326 15650 4378
rect 15702 4326 29838 4378
rect 29890 4326 29902 4378
rect 29954 4326 29966 4378
rect 30018 4326 30030 4378
rect 30082 4326 30094 4378
rect 30146 4326 44282 4378
rect 44334 4326 44346 4378
rect 44398 4326 44410 4378
rect 44462 4326 44474 4378
rect 44526 4326 44538 4378
rect 44590 4326 58726 4378
rect 58778 4326 58790 4378
rect 58842 4326 58854 4378
rect 58906 4326 58918 4378
rect 58970 4326 58982 4378
rect 59034 4326 59040 4378
rect 1104 4304 59040 4326
rect 3970 4224 3976 4276
rect 4028 4224 4034 4276
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7834 4264 7840 4276
rect 7055 4236 7840 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8904 4236 8953 4264
rect 8904 4224 8910 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 8941 4227 8999 4233
rect 2682 4156 2688 4208
rect 2740 4196 2746 4208
rect 3878 4196 3884 4208
rect 2740 4168 3884 4196
rect 2740 4156 2746 4168
rect 3878 4156 3884 4168
rect 3936 4156 3942 4208
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2958 4128 2964 4140
rect 2455 4100 2964 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3142 4128 3148 4140
rect 3099 4100 3148 4128
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3988 4128 4016 4224
rect 6362 4156 6368 4208
rect 6420 4156 6426 4208
rect 7926 4156 7932 4208
rect 7984 4156 7990 4208
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 3988 4100 4445 4128
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4614 4088 4620 4140
rect 4672 4088 4678 4140
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6236 4100 6868 4128
rect 6236 4088 6242 4100
rect 3160 4060 3188 4088
rect 6840 4072 6868 4100
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 7064 4100 7205 4128
rect 7064 4088 7070 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7828 4131 7886 4137
rect 7828 4097 7840 4131
rect 7874 4128 7886 4131
rect 7944 4128 7972 4156
rect 7874 4100 7972 4128
rect 8956 4128 8984 4227
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 9732 4236 10824 4264
rect 9732 4224 9738 4236
rect 10796 4208 10824 4236
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14332 4236 14749 4264
rect 14332 4224 14338 4236
rect 14737 4233 14749 4236
rect 14783 4233 14795 4267
rect 14737 4227 14795 4233
rect 15194 4224 15200 4276
rect 15252 4224 15258 4276
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16209 4267 16267 4273
rect 16209 4264 16221 4267
rect 15804 4236 16221 4264
rect 15804 4224 15810 4236
rect 16209 4233 16221 4236
rect 16255 4233 16267 4267
rect 17865 4267 17923 4273
rect 17865 4264 17877 4267
rect 16209 4227 16267 4233
rect 17788 4236 17877 4264
rect 10778 4156 10784 4208
rect 10836 4156 10842 4208
rect 11532 4168 13308 4196
rect 8956 4100 9352 4128
rect 7874 4097 7886 4100
rect 7828 4091 7886 4097
rect 4341 4063 4399 4069
rect 3160 4032 3924 4060
rect 3896 4001 3924 4032
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4387 4032 4752 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 3237 3995 3295 4001
rect 3237 3992 3249 3995
rect 2884 3964 3249 3992
rect 2884 3936 2912 3964
rect 3237 3961 3249 3964
rect 3283 3961 3295 3995
rect 3237 3955 3295 3961
rect 3881 3995 3939 4001
rect 3881 3961 3893 3995
rect 3927 3961 3939 3995
rect 3881 3955 3939 3961
rect 4724 3936 4752 4032
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6328 4032 6745 4060
rect 6328 4020 6334 4032
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 6822 4020 6828 4072
rect 6880 4020 6886 4072
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7432 4032 7573 4060
rect 7432 4020 7438 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4029 9275 4063
rect 9324 4060 9352 4100
rect 11330 4088 11336 4140
rect 11388 4088 11394 4140
rect 11422 4088 11428 4140
rect 11480 4128 11486 4140
rect 11532 4137 11560 4168
rect 13280 4140 13308 4168
rect 14826 4156 14832 4208
rect 14884 4156 14890 4208
rect 15105 4199 15163 4205
rect 15105 4165 15117 4199
rect 15151 4196 15163 4199
rect 15151 4168 17080 4196
rect 15151 4165 15163 4168
rect 15105 4159 15163 4165
rect 11790 4137 11796 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11480 4100 11529 4128
rect 11480 4088 11486 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11784 4128 11796 4137
rect 11751 4100 11796 4128
rect 11517 4091 11575 4097
rect 11784 4091 11796 4100
rect 11790 4088 11796 4091
rect 11848 4088 11854 4140
rect 13170 4088 13176 4140
rect 13228 4088 13234 4140
rect 13262 4088 13268 4140
rect 13320 4088 13326 4140
rect 13532 4131 13590 4137
rect 13532 4097 13544 4131
rect 13578 4128 13590 4131
rect 14844 4128 14872 4156
rect 13578 4100 14872 4128
rect 13578 4097 13590 4100
rect 13532 4091 13590 4097
rect 10134 4069 10140 4072
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9324 4032 9965 4060
rect 9217 4023 9275 4029
rect 9953 4029 9965 4032
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 10091 4063 10140 4069
rect 10091 4029 10103 4063
rect 10137 4029 10140 4063
rect 10091 4023 10140 4029
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 6549 3995 6607 4001
rect 5123 3964 6040 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 6012 3936 6040 3964
rect 6549 3961 6561 3995
rect 6595 3992 6607 3995
rect 9232 3992 9260 4023
rect 10134 4020 10140 4023
rect 10192 4020 10198 4072
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10410 4060 10416 4072
rect 10275 4032 10416 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10410 4020 10416 4032
rect 10468 4020 10474 4072
rect 11054 4020 11060 4072
rect 11112 4020 11118 4072
rect 14458 4020 14464 4072
rect 14516 4020 14522 4072
rect 14550 4020 14556 4072
rect 14608 4060 14614 4072
rect 15120 4060 15148 4159
rect 17052 4140 17080 4168
rect 17402 4156 17408 4208
rect 17460 4196 17466 4208
rect 17788 4196 17816 4236
rect 17865 4233 17877 4236
rect 17911 4233 17923 4267
rect 17865 4227 17923 4233
rect 19058 4224 19064 4276
rect 19116 4264 19122 4276
rect 19521 4267 19579 4273
rect 19521 4264 19533 4267
rect 19116 4236 19533 4264
rect 19116 4224 19122 4236
rect 19521 4233 19533 4236
rect 19567 4233 19579 4267
rect 21542 4264 21548 4276
rect 19521 4227 19579 4233
rect 19628 4236 21548 4264
rect 19628 4196 19656 4236
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 21818 4224 21824 4276
rect 21876 4224 21882 4276
rect 23106 4264 23112 4276
rect 22848 4236 23112 4264
rect 21836 4196 21864 4224
rect 17460 4168 17816 4196
rect 18064 4168 19656 4196
rect 20824 4168 21864 4196
rect 17460 4156 17466 4168
rect 14608 4032 15148 4060
rect 15212 4100 16344 4128
rect 14608 4020 14614 4032
rect 9582 3992 9588 4004
rect 6595 3964 7604 3992
rect 9232 3964 9588 3992
rect 6595 3961 6607 3964
rect 6549 3955 6607 3961
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 4154 3924 4160 3936
rect 3007 3896 4160 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4706 3884 4712 3936
rect 4764 3884 4770 3936
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 5902 3924 5908 3936
rect 5859 3896 5908 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 5994 3884 6000 3936
rect 6052 3884 6058 3936
rect 6178 3884 6184 3936
rect 6236 3924 6242 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6236 3896 6377 3924
rect 6236 3884 6242 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6638 3884 6644 3936
rect 6696 3884 6702 3936
rect 7576 3924 7604 3964
rect 9582 3952 9588 3964
rect 9640 3952 9646 4004
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 9766 3992 9772 4004
rect 9723 3964 9772 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 11072 3992 11100 4020
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 11072 3964 11161 3992
rect 11149 3961 11161 3964
rect 11195 3961 11207 3995
rect 11149 3955 11207 3961
rect 10226 3924 10232 3936
rect 7576 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10870 3884 10876 3936
rect 10928 3884 10934 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 11756 3896 12909 3924
rect 11756 3884 11762 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 14476 3924 14504 4020
rect 14645 3995 14703 4001
rect 14645 3961 14657 3995
rect 14691 3992 14703 3995
rect 15010 3992 15016 4004
rect 14691 3964 15016 3992
rect 14691 3961 14703 3964
rect 14645 3955 14703 3961
rect 15010 3952 15016 3964
rect 15068 3992 15074 4004
rect 15212 3992 15240 4100
rect 16316 4072 16344 4100
rect 16482 4088 16488 4140
rect 16540 4088 16546 4140
rect 17034 4088 17040 4140
rect 17092 4088 17098 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17770 4128 17776 4140
rect 17175 4100 17776 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 18064 4072 18092 4168
rect 18138 4088 18144 4140
rect 18196 4088 18202 4140
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4128 19671 4131
rect 19794 4128 19800 4140
rect 19659 4100 19800 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 19794 4088 19800 4100
rect 19852 4128 19858 4140
rect 20257 4131 20315 4137
rect 19852 4100 20208 4128
rect 19852 4088 19858 4100
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 15068 3964 15240 3992
rect 15068 3952 15074 3964
rect 15304 3924 15332 4023
rect 15378 4020 15384 4072
rect 15436 4060 15442 4072
rect 15565 4063 15623 4069
rect 15565 4060 15577 4063
rect 15436 4032 15577 4060
rect 15436 4020 15442 4032
rect 15565 4029 15577 4032
rect 15611 4029 15623 4063
rect 15565 4023 15623 4029
rect 16298 4020 16304 4072
rect 16356 4020 16362 4072
rect 17218 4020 17224 4072
rect 17276 4020 17282 4072
rect 17310 4020 17316 4072
rect 17368 4060 17374 4072
rect 17957 4063 18015 4069
rect 17957 4060 17969 4063
rect 17368 4032 17969 4060
rect 17368 4020 17374 4032
rect 17957 4029 17969 4032
rect 18003 4029 18015 4063
rect 17957 4023 18015 4029
rect 18046 4020 18052 4072
rect 18104 4020 18110 4072
rect 17497 3995 17555 4001
rect 17497 3961 17509 3995
rect 17543 3992 17555 3995
rect 18156 3992 18184 4088
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18340 4032 18429 4060
rect 18340 4004 18368 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19705 4063 19763 4069
rect 19705 4060 19717 4063
rect 19484 4032 19717 4060
rect 19484 4020 19490 4032
rect 19705 4029 19717 4032
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 20070 4020 20076 4072
rect 20128 4020 20134 4072
rect 20180 4060 20208 4100
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 20824 4128 20852 4168
rect 20303 4100 20852 4128
rect 20901 4131 20959 4137
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 20901 4097 20913 4131
rect 20947 4128 20959 4131
rect 21545 4131 21603 4137
rect 20947 4100 21211 4128
rect 20947 4097 20959 4100
rect 20901 4091 20959 4097
rect 20916 4060 20944 4091
rect 20180 4032 20944 4060
rect 20990 4020 20996 4072
rect 21048 4020 21054 4072
rect 21082 4020 21088 4072
rect 21140 4020 21146 4072
rect 21183 4060 21211 4100
rect 21545 4097 21557 4131
rect 21591 4128 21603 4131
rect 22094 4128 22100 4140
rect 21591 4100 22100 4128
rect 21591 4097 21603 4100
rect 21545 4091 21603 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22370 4088 22376 4140
rect 22428 4128 22434 4140
rect 22848 4137 22876 4236
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 23566 4224 23572 4276
rect 23624 4264 23630 4276
rect 23937 4267 23995 4273
rect 23937 4264 23949 4267
rect 23624 4236 23949 4264
rect 23624 4224 23630 4236
rect 23937 4233 23949 4236
rect 23983 4233 23995 4267
rect 23937 4227 23995 4233
rect 26418 4224 26424 4276
rect 26476 4224 26482 4276
rect 29457 4267 29515 4273
rect 29457 4233 29469 4267
rect 29503 4264 29515 4267
rect 29546 4264 29552 4276
rect 29503 4236 29552 4264
rect 29503 4233 29515 4236
rect 29457 4227 29515 4233
rect 29546 4224 29552 4236
rect 29604 4224 29610 4276
rect 29730 4224 29736 4276
rect 29788 4224 29794 4276
rect 30558 4264 30564 4276
rect 30300 4236 30564 4264
rect 23124 4196 23152 4224
rect 25682 4196 25688 4208
rect 23124 4168 25688 4196
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 22428 4100 22477 4128
rect 22428 4088 22434 4100
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22833 4131 22891 4137
rect 22833 4097 22845 4131
rect 22879 4097 22891 4131
rect 22833 4091 22891 4097
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 23385 4131 23443 4137
rect 23385 4097 23397 4131
rect 23431 4128 23443 4131
rect 23474 4128 23480 4140
rect 23431 4100 23480 4128
rect 23431 4097 23443 4100
rect 23385 4091 23443 4097
rect 21726 4060 21732 4072
rect 21183 4032 21732 4060
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 21910 4020 21916 4072
rect 21968 4020 21974 4072
rect 23032 4060 23060 4091
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 24228 4137 24256 4168
rect 25682 4156 25688 4168
rect 25740 4196 25746 4208
rect 26602 4196 26608 4208
rect 25740 4168 26608 4196
rect 25740 4156 25746 4168
rect 26602 4156 26608 4168
rect 26660 4156 26666 4208
rect 27338 4156 27344 4208
rect 27396 4156 27402 4208
rect 29362 4156 29368 4208
rect 29420 4156 29426 4208
rect 24213 4131 24271 4137
rect 24213 4097 24225 4131
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 24397 4131 24455 4137
rect 24397 4097 24409 4131
rect 24443 4097 24455 4131
rect 24397 4091 24455 4097
rect 23566 4060 23572 4072
rect 23032 4032 23572 4060
rect 23566 4020 23572 4032
rect 23624 4020 23630 4072
rect 24412 4060 24440 4091
rect 24578 4088 24584 4140
rect 24636 4128 24642 4140
rect 24673 4131 24731 4137
rect 24673 4128 24685 4131
rect 24636 4100 24685 4128
rect 24636 4088 24642 4100
rect 24673 4097 24685 4100
rect 24719 4097 24731 4131
rect 24673 4091 24731 4097
rect 25314 4088 25320 4140
rect 25372 4088 25378 4140
rect 25590 4088 25596 4140
rect 25648 4088 25654 4140
rect 25866 4088 25872 4140
rect 25924 4088 25930 4140
rect 26789 4131 26847 4137
rect 26789 4128 26801 4131
rect 26252 4100 26801 4128
rect 26142 4060 26148 4072
rect 24412 4032 26148 4060
rect 26142 4020 26148 4032
rect 26200 4020 26206 4072
rect 17543 3964 18184 3992
rect 17543 3961 17555 3964
rect 17497 3955 17555 3961
rect 18322 3952 18328 4004
rect 18380 3952 18386 4004
rect 20441 3995 20499 4001
rect 20441 3961 20453 3995
rect 20487 3992 20499 3995
rect 22186 3992 22192 4004
rect 20487 3964 22192 3992
rect 20487 3961 20499 3964
rect 20441 3955 20499 3961
rect 22186 3952 22192 3964
rect 22244 3952 22250 4004
rect 23382 3952 23388 4004
rect 23440 3992 23446 4004
rect 26252 3992 26280 4100
rect 26789 4097 26801 4100
rect 26835 4097 26847 4131
rect 26789 4091 26847 4097
rect 27157 4131 27215 4137
rect 27157 4097 27169 4131
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 27172 4060 27200 4091
rect 27246 4088 27252 4140
rect 27304 4128 27310 4140
rect 27617 4131 27675 4137
rect 27617 4128 27629 4131
rect 27304 4100 27629 4128
rect 27304 4088 27310 4100
rect 27617 4097 27629 4100
rect 27663 4097 27675 4131
rect 27617 4091 27675 4097
rect 28344 4131 28402 4137
rect 28344 4097 28356 4131
rect 28390 4128 28402 4131
rect 29380 4128 29408 4156
rect 28390 4100 29408 4128
rect 28390 4097 28402 4100
rect 28344 4091 28402 4097
rect 26384 4032 27200 4060
rect 26384 4020 26390 4032
rect 27430 4020 27436 4072
rect 27488 4020 27494 4072
rect 28077 4063 28135 4069
rect 28077 4029 28089 4063
rect 28123 4029 28135 4063
rect 29564 4060 29592 4224
rect 29748 4196 29776 4224
rect 30300 4196 30328 4236
rect 30558 4224 30564 4236
rect 30616 4224 30622 4276
rect 31938 4224 31944 4276
rect 31996 4224 32002 4276
rect 34054 4224 34060 4276
rect 34112 4264 34118 4276
rect 34885 4267 34943 4273
rect 34885 4264 34897 4267
rect 34112 4236 34897 4264
rect 34112 4224 34118 4236
rect 34885 4233 34897 4236
rect 34931 4233 34943 4267
rect 34885 4227 34943 4233
rect 29656 4168 29776 4196
rect 30116 4168 30328 4196
rect 34900 4196 34928 4227
rect 35894 4224 35900 4276
rect 35952 4264 35958 4276
rect 35989 4267 36047 4273
rect 35989 4264 36001 4267
rect 35952 4236 36001 4264
rect 35952 4224 35958 4236
rect 35989 4233 36001 4236
rect 36035 4233 36047 4267
rect 35989 4227 36047 4233
rect 36814 4224 36820 4276
rect 36872 4224 36878 4276
rect 37458 4224 37464 4276
rect 37516 4264 37522 4276
rect 38013 4267 38071 4273
rect 38013 4264 38025 4267
rect 37516 4236 38025 4264
rect 37516 4224 37522 4236
rect 38013 4233 38025 4236
rect 38059 4233 38071 4267
rect 38013 4227 38071 4233
rect 39206 4224 39212 4276
rect 39264 4264 39270 4276
rect 39853 4267 39911 4273
rect 39853 4264 39865 4267
rect 39264 4236 39865 4264
rect 39264 4224 39270 4236
rect 39853 4233 39865 4236
rect 39899 4233 39911 4267
rect 39853 4227 39911 4233
rect 40310 4224 40316 4276
rect 40368 4264 40374 4276
rect 40681 4267 40739 4273
rect 40681 4264 40693 4267
rect 40368 4236 40693 4264
rect 40368 4224 40374 4236
rect 40681 4233 40693 4236
rect 40727 4233 40739 4267
rect 42058 4264 42064 4276
rect 40681 4227 40739 4233
rect 41800 4236 42064 4264
rect 36262 4196 36268 4208
rect 34900 4168 36268 4196
rect 29656 4137 29684 4168
rect 29641 4131 29699 4137
rect 29641 4097 29653 4131
rect 29687 4097 29699 4131
rect 29641 4091 29699 4097
rect 29730 4088 29736 4140
rect 29788 4088 29794 4140
rect 30116 4137 30144 4168
rect 36262 4156 36268 4168
rect 36320 4156 36326 4208
rect 36832 4196 36860 4224
rect 41800 4205 41828 4236
rect 42058 4224 42064 4236
rect 42116 4224 42122 4276
rect 43622 4224 43628 4276
rect 43680 4224 43686 4276
rect 45186 4224 45192 4276
rect 45244 4224 45250 4276
rect 45741 4267 45799 4273
rect 45741 4233 45753 4267
rect 45787 4233 45799 4267
rect 45741 4227 45799 4233
rect 41785 4199 41843 4205
rect 36832 4168 41276 4196
rect 30101 4131 30159 4137
rect 30101 4097 30113 4131
rect 30147 4097 30159 4131
rect 30101 4091 30159 4097
rect 30208 4098 30411 4126
rect 30208 4060 30236 4098
rect 29564 4032 30236 4060
rect 30285 4063 30343 4069
rect 28077 4023 28135 4029
rect 30285 4029 30297 4063
rect 30331 4029 30343 4063
rect 30383 4060 30411 4098
rect 31294 4088 31300 4140
rect 31352 4088 31358 4140
rect 32214 4088 32220 4140
rect 32272 4088 32278 4140
rect 33226 4088 33232 4140
rect 33284 4088 33290 4140
rect 34977 4131 35035 4137
rect 34977 4097 34989 4131
rect 35023 4128 35035 4131
rect 35023 4100 35848 4128
rect 35023 4097 35035 4100
rect 34977 4091 35035 4097
rect 31202 4069 31208 4072
rect 31021 4063 31079 4069
rect 31021 4060 31033 4063
rect 30383 4032 31033 4060
rect 30285 4023 30343 4029
rect 31021 4029 31033 4032
rect 31067 4029 31079 4063
rect 31021 4023 31079 4029
rect 31159 4063 31208 4069
rect 31159 4029 31171 4063
rect 31205 4029 31208 4063
rect 31159 4023 31208 4029
rect 23440 3964 26280 3992
rect 23440 3952 23446 3964
rect 26510 3952 26516 4004
rect 26568 3992 26574 4004
rect 26605 3995 26663 4001
rect 26605 3992 26617 3995
rect 26568 3964 26617 3992
rect 26568 3952 26574 3964
rect 26605 3961 26617 3964
rect 26651 3961 26663 3995
rect 26605 3955 26663 3961
rect 27062 3952 27068 4004
rect 27120 3992 27126 4004
rect 27890 3992 27896 4004
rect 27120 3964 27896 3992
rect 27120 3952 27126 3964
rect 27890 3952 27896 3964
rect 27948 3992 27954 4004
rect 28092 3992 28120 4023
rect 27948 3964 28120 3992
rect 27948 3952 27954 3964
rect 14476 3896 15332 3924
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 15620 3896 16313 3924
rect 15620 3884 15626 3896
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 16301 3887 16359 3893
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16448 3896 16681 3924
rect 16448 3884 16454 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 17736 3896 18981 3924
rect 17736 3884 17742 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 19150 3884 19156 3936
rect 19208 3884 19214 3936
rect 20530 3884 20536 3936
rect 20588 3884 20594 3936
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 21634 3924 21640 3936
rect 21407 3896 21640 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 21634 3884 21640 3896
rect 21692 3884 21698 3936
rect 23201 3927 23259 3933
rect 23201 3893 23213 3927
rect 23247 3924 23259 3927
rect 23750 3924 23756 3936
rect 23247 3896 23756 3924
rect 23247 3893 23259 3896
rect 23201 3887 23259 3893
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 24581 3927 24639 3933
rect 24581 3893 24593 3927
rect 24627 3924 24639 3927
rect 25130 3924 25136 3936
rect 24627 3896 25136 3924
rect 24627 3893 24639 3896
rect 24581 3887 24639 3893
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 25409 3927 25467 3933
rect 25409 3893 25421 3927
rect 25455 3924 25467 3927
rect 25774 3924 25780 3936
rect 25455 3896 25780 3924
rect 25455 3893 25467 3896
rect 25409 3887 25467 3893
rect 25774 3884 25780 3896
rect 25832 3884 25838 3936
rect 26970 3884 26976 3936
rect 27028 3884 27034 3936
rect 27338 3884 27344 3936
rect 27396 3884 27402 3936
rect 27798 3884 27804 3936
rect 27856 3884 27862 3936
rect 29546 3884 29552 3936
rect 29604 3924 29610 3936
rect 29917 3927 29975 3933
rect 29917 3924 29929 3927
rect 29604 3896 29929 3924
rect 29604 3884 29610 3896
rect 29917 3893 29929 3896
rect 29963 3893 29975 3927
rect 30300 3924 30328 4023
rect 31202 4020 31208 4023
rect 31260 4020 31266 4072
rect 31478 4020 31484 4072
rect 31536 4060 31542 4072
rect 31846 4060 31852 4072
rect 31536 4032 31852 4060
rect 31536 4020 31542 4032
rect 31846 4020 31852 4032
rect 31904 4060 31910 4072
rect 32950 4060 32956 4072
rect 31904 4032 32956 4060
rect 31904 4020 31910 4032
rect 32950 4020 32956 4032
rect 33008 4020 33014 4072
rect 34057 4063 34115 4069
rect 34057 4029 34069 4063
rect 34103 4060 34115 4063
rect 34422 4060 34428 4072
rect 34103 4032 34428 4060
rect 34103 4029 34115 4032
rect 34057 4023 34115 4029
rect 34422 4020 34428 4032
rect 34480 4020 34486 4072
rect 35066 4020 35072 4072
rect 35124 4020 35130 4072
rect 35345 4063 35403 4069
rect 35345 4029 35357 4063
rect 35391 4029 35403 4063
rect 35345 4023 35403 4029
rect 30742 3952 30748 4004
rect 30800 3952 30806 4004
rect 34517 3995 34575 4001
rect 34517 3961 34529 3995
rect 34563 3992 34575 3995
rect 35360 3992 35388 4023
rect 35526 4020 35532 4072
rect 35584 4020 35590 4072
rect 35820 4060 35848 4100
rect 35986 4088 35992 4140
rect 36044 4128 36050 4140
rect 36081 4131 36139 4137
rect 36081 4128 36093 4131
rect 36044 4100 36093 4128
rect 36044 4088 36050 4100
rect 36081 4097 36093 4100
rect 36127 4097 36139 4131
rect 36081 4091 36139 4097
rect 37093 4131 37151 4137
rect 37093 4097 37105 4131
rect 37139 4128 37151 4131
rect 38654 4128 38660 4140
rect 37139 4100 38660 4128
rect 37139 4097 37151 4100
rect 37093 4091 37151 4097
rect 38654 4088 38660 4100
rect 38712 4088 38718 4140
rect 39022 4088 39028 4140
rect 39080 4088 39086 4140
rect 39301 4131 39359 4137
rect 39301 4097 39313 4131
rect 39347 4128 39359 4131
rect 39850 4128 39856 4140
rect 39347 4100 39856 4128
rect 39347 4097 39359 4100
rect 39301 4091 39359 4097
rect 39850 4088 39856 4100
rect 39908 4088 39914 4140
rect 40034 4088 40040 4140
rect 40092 4088 40098 4140
rect 40880 4137 40908 4168
rect 40865 4131 40923 4137
rect 40865 4097 40877 4131
rect 40911 4097 40923 4131
rect 40865 4091 40923 4097
rect 40957 4131 41015 4137
rect 40957 4097 40969 4131
rect 41003 4097 41015 4131
rect 40957 4091 41015 4097
rect 36725 4063 36783 4069
rect 36725 4060 36737 4063
rect 35820 4032 36737 4060
rect 36725 4029 36737 4032
rect 36771 4029 36783 4063
rect 36725 4023 36783 4029
rect 37366 4020 37372 4072
rect 37424 4020 37430 4072
rect 38105 4063 38163 4069
rect 38105 4029 38117 4063
rect 38151 4029 38163 4063
rect 39758 4060 39764 4072
rect 38105 4023 38163 4029
rect 38856 4032 39764 4060
rect 34563 3964 35388 3992
rect 35544 3992 35572 4020
rect 38120 3992 38148 4023
rect 38856 4001 38884 4032
rect 39758 4020 39764 4032
rect 39816 4020 39822 4072
rect 35544 3964 38148 3992
rect 38841 3995 38899 4001
rect 34563 3961 34575 3964
rect 34517 3955 34575 3961
rect 38841 3961 38853 3995
rect 38887 3961 38899 3995
rect 38841 3955 38899 3961
rect 39482 3952 39488 4004
rect 39540 3992 39546 4004
rect 40972 3992 41000 4091
rect 41248 4069 41276 4168
rect 41785 4165 41797 4199
rect 41831 4165 41843 4199
rect 41785 4159 41843 4165
rect 41874 4156 41880 4208
rect 41932 4196 41938 4208
rect 41932 4168 42104 4196
rect 41932 4156 41938 4168
rect 41414 4088 41420 4140
rect 41472 4088 41478 4140
rect 42076 4137 42104 4168
rect 42334 4156 42340 4208
rect 42392 4196 42398 4208
rect 42429 4199 42487 4205
rect 42429 4196 42441 4199
rect 42392 4168 42441 4196
rect 42392 4156 42398 4168
rect 42429 4165 42441 4168
rect 42475 4165 42487 4199
rect 42429 4159 42487 4165
rect 43254 4156 43260 4208
rect 43312 4196 43318 4208
rect 43901 4199 43959 4205
rect 43901 4196 43913 4199
rect 43312 4168 43913 4196
rect 43312 4156 43318 4168
rect 43901 4165 43913 4168
rect 43947 4165 43959 4199
rect 45756 4196 45784 4227
rect 48590 4224 48596 4276
rect 48648 4264 48654 4276
rect 48869 4267 48927 4273
rect 48869 4264 48881 4267
rect 48648 4236 48881 4264
rect 48648 4224 48654 4236
rect 48869 4233 48881 4236
rect 48915 4233 48927 4267
rect 48869 4227 48927 4233
rect 49234 4224 49240 4276
rect 49292 4264 49298 4276
rect 49418 4264 49424 4276
rect 49292 4236 49424 4264
rect 49292 4224 49298 4236
rect 49418 4224 49424 4236
rect 49476 4224 49482 4276
rect 53742 4224 53748 4276
rect 53800 4224 53806 4276
rect 55674 4264 55680 4276
rect 54680 4236 55680 4264
rect 45830 4196 45836 4208
rect 45756 4168 45836 4196
rect 43901 4159 43959 4165
rect 45830 4156 45836 4168
rect 45888 4156 45894 4208
rect 46109 4199 46167 4205
rect 46109 4165 46121 4199
rect 46155 4196 46167 4199
rect 47213 4199 47271 4205
rect 47213 4196 47225 4199
rect 46155 4168 47225 4196
rect 46155 4165 46167 4168
rect 46109 4159 46167 4165
rect 47213 4165 47225 4168
rect 47259 4165 47271 4199
rect 47213 4159 47271 4165
rect 49329 4199 49387 4205
rect 49329 4165 49341 4199
rect 49375 4196 49387 4199
rect 51169 4199 51227 4205
rect 51169 4196 51181 4199
rect 49375 4168 51181 4196
rect 49375 4165 49387 4168
rect 49329 4159 49387 4165
rect 51169 4165 51181 4168
rect 51215 4165 51227 4199
rect 53760 4196 53788 4224
rect 51169 4159 51227 4165
rect 52748 4168 53788 4196
rect 52748 4140 52776 4168
rect 54018 4156 54024 4208
rect 54076 4156 54082 4208
rect 42061 4131 42119 4137
rect 42061 4097 42073 4131
rect 42107 4097 42119 4131
rect 42061 4091 42119 4097
rect 43073 4131 43131 4137
rect 43073 4097 43085 4131
rect 43119 4128 43131 4131
rect 43162 4128 43168 4140
rect 43119 4100 43168 4128
rect 43119 4097 43131 4100
rect 43073 4091 43131 4097
rect 43162 4088 43168 4100
rect 43220 4088 43226 4140
rect 43530 4088 43536 4140
rect 43588 4088 43594 4140
rect 43809 4131 43867 4137
rect 43809 4097 43821 4131
rect 43855 4097 43867 4131
rect 43809 4091 43867 4097
rect 41233 4063 41291 4069
rect 41233 4029 41245 4063
rect 41279 4060 41291 4063
rect 41322 4060 41328 4072
rect 41279 4032 41328 4060
rect 41279 4029 41291 4032
rect 41233 4023 41291 4029
rect 41322 4020 41328 4032
rect 41380 4020 41386 4072
rect 41969 4063 42027 4069
rect 41969 4029 41981 4063
rect 42015 4029 42027 4063
rect 41969 4023 42027 4029
rect 42076 4032 42748 4060
rect 39540 3964 41000 3992
rect 39540 3952 39546 3964
rect 41984 3936 42012 4023
rect 33134 3924 33140 3936
rect 30300 3896 33140 3924
rect 29917 3887 29975 3893
rect 33134 3884 33140 3896
rect 33192 3924 33198 3936
rect 33594 3924 33600 3936
rect 33192 3896 33600 3924
rect 33192 3884 33198 3896
rect 33594 3884 33600 3896
rect 33652 3884 33658 3936
rect 35250 3884 35256 3936
rect 35308 3924 35314 3936
rect 36909 3927 36967 3933
rect 36909 3924 36921 3927
rect 35308 3896 36921 3924
rect 35308 3884 35314 3896
rect 36909 3893 36921 3896
rect 36955 3893 36967 3927
rect 36909 3887 36967 3893
rect 37734 3884 37740 3936
rect 37792 3924 37798 3936
rect 38749 3927 38807 3933
rect 38749 3924 38761 3927
rect 37792 3896 38761 3924
rect 37792 3884 37798 3896
rect 38749 3893 38761 3896
rect 38795 3893 38807 3927
rect 38749 3887 38807 3893
rect 40034 3884 40040 3936
rect 40092 3924 40098 3936
rect 41141 3927 41199 3933
rect 41141 3924 41153 3927
rect 40092 3896 41153 3924
rect 40092 3884 40098 3896
rect 41141 3893 41153 3896
rect 41187 3893 41199 3927
rect 41141 3887 41199 3893
rect 41598 3884 41604 3936
rect 41656 3884 41662 3936
rect 41966 3884 41972 3936
rect 42024 3884 42030 3936
rect 42076 3933 42104 4032
rect 42245 3995 42303 4001
rect 42245 3961 42257 3995
rect 42291 3992 42303 3995
rect 42613 3995 42671 4001
rect 42613 3992 42625 3995
rect 42291 3964 42625 3992
rect 42291 3961 42303 3964
rect 42245 3955 42303 3961
rect 42613 3961 42625 3964
rect 42659 3961 42671 3995
rect 42720 3992 42748 4032
rect 42794 4020 42800 4072
rect 42852 4020 42858 4072
rect 42886 4020 42892 4072
rect 42944 4020 42950 4072
rect 42978 4020 42984 4072
rect 43036 4060 43042 4072
rect 43824 4060 43852 4091
rect 45554 4088 45560 4140
rect 45612 4128 45618 4140
rect 46474 4128 46480 4140
rect 45612 4100 46480 4128
rect 45612 4088 45618 4100
rect 46474 4088 46480 4100
rect 46532 4128 46538 4140
rect 46569 4131 46627 4137
rect 46569 4128 46581 4131
rect 46532 4100 46581 4128
rect 46532 4088 46538 4100
rect 46569 4097 46581 4100
rect 46615 4097 46627 4131
rect 46569 4091 46627 4097
rect 47854 4088 47860 4140
rect 47912 4088 47918 4140
rect 48222 4088 48228 4140
rect 48280 4088 48286 4140
rect 52730 4088 52736 4140
rect 52788 4088 52794 4140
rect 53000 4131 53058 4137
rect 53000 4097 53012 4131
rect 53046 4128 53058 4131
rect 54036 4128 54064 4156
rect 54680 4137 54708 4236
rect 55674 4224 55680 4236
rect 55732 4264 55738 4276
rect 55732 4236 56272 4264
rect 55732 4224 55738 4236
rect 53046 4100 54064 4128
rect 54389 4131 54447 4137
rect 53046 4097 53058 4100
rect 53000 4091 53058 4097
rect 54389 4097 54401 4131
rect 54435 4097 54447 4131
rect 54389 4091 54447 4097
rect 54665 4131 54723 4137
rect 54665 4097 54677 4131
rect 54711 4097 54723 4131
rect 54665 4091 54723 4097
rect 43036 4032 43852 4060
rect 43036 4020 43042 4032
rect 44082 4020 44088 4072
rect 44140 4060 44146 4072
rect 46014 4060 46020 4072
rect 44140 4032 46020 4060
rect 44140 4020 44146 4032
rect 46014 4020 46020 4032
rect 46072 4020 46078 4072
rect 46201 4063 46259 4069
rect 46201 4029 46213 4063
rect 46247 4029 46259 4063
rect 46201 4023 46259 4029
rect 46293 4063 46351 4069
rect 46293 4029 46305 4063
rect 46339 4060 46351 4063
rect 49326 4060 49332 4072
rect 46339 4032 49332 4060
rect 46339 4029 46351 4032
rect 46293 4023 46351 4029
rect 44818 3992 44824 4004
rect 42720 3964 44824 3992
rect 42613 3955 42671 3961
rect 44818 3952 44824 3964
rect 44876 3952 44882 4004
rect 45278 3952 45284 4004
rect 45336 3992 45342 4004
rect 46216 3992 46244 4023
rect 45336 3964 46244 3992
rect 45336 3952 45342 3964
rect 42061 3927 42119 3933
rect 42061 3893 42073 3927
rect 42107 3893 42119 3927
rect 42061 3887 42119 3893
rect 42426 3884 42432 3936
rect 42484 3884 42490 3936
rect 42705 3927 42763 3933
rect 42705 3893 42717 3927
rect 42751 3924 42763 3927
rect 43070 3924 43076 3936
rect 42751 3896 43076 3924
rect 42751 3893 42763 3896
rect 42705 3887 42763 3893
rect 43070 3884 43076 3896
rect 43128 3884 43134 3936
rect 43254 3884 43260 3936
rect 43312 3884 43318 3936
rect 43346 3884 43352 3936
rect 43404 3884 43410 3936
rect 43714 3884 43720 3936
rect 43772 3924 43778 3936
rect 46308 3924 46336 4023
rect 49326 4020 49332 4032
rect 49384 4060 49390 4072
rect 49513 4063 49571 4069
rect 49513 4060 49525 4063
rect 49384 4032 49525 4060
rect 49384 4020 49390 4032
rect 49513 4029 49525 4032
rect 49559 4029 49571 4063
rect 49513 4023 49571 4029
rect 49789 4063 49847 4069
rect 49789 4029 49801 4063
rect 49835 4029 49847 4063
rect 49789 4023 49847 4029
rect 48961 3995 49019 4001
rect 48961 3961 48973 3995
rect 49007 3992 49019 3995
rect 49804 3992 49832 4023
rect 49878 4020 49884 4072
rect 49936 4060 49942 4072
rect 50525 4063 50583 4069
rect 50525 4060 50537 4063
rect 49936 4032 50537 4060
rect 49936 4020 49942 4032
rect 50525 4029 50537 4032
rect 50571 4029 50583 4063
rect 50525 4023 50583 4029
rect 51629 4063 51687 4069
rect 51629 4029 51641 4063
rect 51675 4060 51687 4063
rect 51994 4060 52000 4072
rect 51675 4032 52000 4060
rect 51675 4029 51687 4032
rect 51629 4023 51687 4029
rect 51994 4020 52000 4032
rect 52052 4020 52058 4072
rect 54404 4060 54432 4091
rect 53760 4032 54432 4060
rect 54481 4063 54539 4069
rect 49007 3964 49832 3992
rect 49007 3961 49019 3964
rect 48961 3955 49019 3961
rect 43772 3896 46336 3924
rect 43772 3884 43778 3896
rect 47670 3884 47676 3936
rect 47728 3884 47734 3936
rect 49510 3884 49516 3936
rect 49568 3924 49574 3936
rect 50433 3927 50491 3933
rect 50433 3924 50445 3927
rect 49568 3896 50445 3924
rect 49568 3884 49574 3896
rect 50433 3893 50445 3896
rect 50479 3893 50491 3927
rect 50433 3887 50491 3893
rect 52546 3884 52552 3936
rect 52604 3884 52610 3936
rect 53098 3884 53104 3936
rect 53156 3924 53162 3936
rect 53760 3924 53788 4032
rect 54481 4029 54493 4063
rect 54527 4060 54539 4063
rect 54570 4060 54576 4072
rect 54527 4032 54576 4060
rect 54527 4029 54539 4032
rect 54481 4023 54539 4029
rect 54570 4020 54576 4032
rect 54628 4020 54634 4072
rect 55401 4063 55459 4069
rect 55401 4060 55413 4063
rect 54772 4032 55413 4060
rect 54110 3952 54116 4004
rect 54168 3992 54174 4004
rect 54772 3992 54800 4032
rect 55401 4029 55413 4032
rect 55447 4029 55459 4063
rect 55401 4023 55459 4029
rect 55490 4020 55496 4072
rect 55548 4069 55554 4072
rect 55548 4063 55576 4069
rect 55564 4029 55576 4063
rect 55548 4023 55576 4029
rect 55677 4063 55735 4069
rect 55677 4029 55689 4063
rect 55723 4060 55735 4063
rect 55723 4032 56180 4060
rect 55723 4029 55735 4032
rect 55677 4023 55735 4029
rect 55548 4020 55554 4023
rect 56152 4004 56180 4032
rect 54168 3964 54800 3992
rect 54168 3952 54174 3964
rect 54846 3952 54852 4004
rect 54904 3992 54910 4004
rect 55125 3995 55183 4001
rect 55125 3992 55137 3995
rect 54904 3964 55137 3992
rect 54904 3952 54910 3964
rect 55125 3961 55137 3964
rect 55171 3961 55183 3995
rect 55125 3955 55183 3961
rect 56134 3952 56140 4004
rect 56192 3952 56198 4004
rect 56244 3992 56272 4236
rect 56594 4224 56600 4276
rect 56652 4264 56658 4276
rect 56781 4267 56839 4273
rect 56781 4264 56793 4267
rect 56652 4236 56793 4264
rect 56652 4224 56658 4236
rect 56781 4233 56793 4236
rect 56827 4233 56839 4267
rect 56781 4227 56839 4233
rect 56410 4088 56416 4140
rect 56468 4128 56474 4140
rect 57425 4131 57483 4137
rect 57425 4128 57437 4131
rect 56468 4100 57008 4128
rect 56468 4088 56474 4100
rect 56980 4069 57008 4100
rect 57164 4100 57437 4128
rect 57164 4072 57192 4100
rect 57425 4097 57437 4100
rect 57471 4097 57483 4131
rect 57425 4091 57483 4097
rect 57882 4088 57888 4140
rect 57940 4088 57946 4140
rect 56321 4063 56379 4069
rect 56321 4029 56333 4063
rect 56367 4060 56379 4063
rect 56873 4063 56931 4069
rect 56873 4060 56885 4063
rect 56367 4032 56885 4060
rect 56367 4029 56379 4032
rect 56321 4023 56379 4029
rect 56873 4029 56885 4032
rect 56919 4029 56931 4063
rect 56873 4023 56931 4029
rect 56965 4063 57023 4069
rect 56965 4029 56977 4063
rect 57011 4029 57023 4063
rect 56965 4023 57023 4029
rect 57146 4020 57152 4072
rect 57204 4020 57210 4072
rect 57238 4020 57244 4072
rect 57296 4020 57302 4072
rect 56244 3964 58296 3992
rect 58268 3936 58296 3964
rect 53156 3896 53788 3924
rect 53156 3884 53162 3896
rect 54202 3884 54208 3936
rect 54260 3884 54266 3936
rect 54294 3884 54300 3936
rect 54352 3924 54358 3936
rect 55490 3924 55496 3936
rect 54352 3896 55496 3924
rect 54352 3884 54358 3896
rect 55490 3884 55496 3896
rect 55548 3884 55554 3936
rect 55582 3884 55588 3936
rect 55640 3924 55646 3936
rect 56318 3924 56324 3936
rect 55640 3896 56324 3924
rect 55640 3884 55646 3896
rect 56318 3884 56324 3896
rect 56376 3884 56382 3936
rect 56410 3884 56416 3936
rect 56468 3884 56474 3936
rect 56594 3884 56600 3936
rect 56652 3924 56658 3936
rect 57238 3924 57244 3936
rect 56652 3896 57244 3924
rect 56652 3884 56658 3896
rect 57238 3884 57244 3896
rect 57296 3884 57302 3936
rect 57606 3884 57612 3936
rect 57664 3884 57670 3936
rect 58250 3884 58256 3936
rect 58308 3884 58314 3936
rect 58529 3927 58587 3933
rect 58529 3893 58541 3927
rect 58575 3924 58587 3927
rect 58575 3896 58940 3924
rect 58575 3893 58587 3896
rect 58529 3887 58587 3893
rect 1104 3834 58880 3856
rect 1104 3782 8172 3834
rect 8224 3782 8236 3834
rect 8288 3782 8300 3834
rect 8352 3782 8364 3834
rect 8416 3782 8428 3834
rect 8480 3782 22616 3834
rect 22668 3782 22680 3834
rect 22732 3782 22744 3834
rect 22796 3782 22808 3834
rect 22860 3782 22872 3834
rect 22924 3782 37060 3834
rect 37112 3782 37124 3834
rect 37176 3782 37188 3834
rect 37240 3782 37252 3834
rect 37304 3782 37316 3834
rect 37368 3782 51504 3834
rect 51556 3782 51568 3834
rect 51620 3782 51632 3834
rect 51684 3782 51696 3834
rect 51748 3782 51760 3834
rect 51812 3782 58880 3834
rect 1104 3760 58880 3782
rect 3142 3680 3148 3732
rect 3200 3680 3206 3732
rect 5442 3680 5448 3732
rect 5500 3680 5506 3732
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6638 3720 6644 3732
rect 6595 3692 6644 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 8938 3720 8944 3732
rect 6880 3692 8944 3720
rect 6880 3680 6886 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 10134 3680 10140 3732
rect 10192 3680 10198 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11977 3723 12035 3729
rect 11977 3720 11989 3723
rect 10836 3692 11989 3720
rect 10836 3680 10842 3692
rect 11977 3689 11989 3692
rect 12023 3689 12035 3723
rect 11977 3683 12035 3689
rect 12986 3680 12992 3732
rect 13044 3720 13050 3732
rect 14921 3723 14979 3729
rect 14921 3720 14933 3723
rect 13044 3692 14933 3720
rect 13044 3680 13050 3692
rect 14921 3689 14933 3692
rect 14967 3689 14979 3723
rect 14921 3683 14979 3689
rect 15856 3692 17264 3720
rect 3421 3655 3479 3661
rect 3421 3621 3433 3655
rect 3467 3621 3479 3655
rect 3421 3615 3479 3621
rect 1762 3544 1768 3596
rect 1820 3544 1826 3596
rect 3436 3584 3464 3615
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4157 3655 4215 3661
rect 4157 3652 4169 3655
rect 4028 3624 4169 3652
rect 4028 3612 4034 3624
rect 4157 3621 4169 3624
rect 4203 3652 4215 3655
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 4203 3624 4445 3652
rect 4203 3621 4215 3624
rect 4157 3615 4215 3621
rect 4433 3621 4445 3624
rect 4479 3621 4491 3655
rect 4433 3615 4491 3621
rect 4798 3612 4804 3664
rect 4856 3652 4862 3664
rect 5460 3652 5488 3680
rect 4856 3624 5488 3652
rect 8665 3655 8723 3661
rect 4856 3612 4862 3624
rect 5368 3593 5396 3624
rect 8665 3621 8677 3655
rect 8711 3652 8723 3655
rect 8754 3652 8760 3664
rect 8711 3624 8760 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 8754 3612 8760 3624
rect 8812 3652 8818 3664
rect 10152 3652 10180 3680
rect 8812 3624 10180 3652
rect 8812 3612 8818 3624
rect 14090 3612 14096 3664
rect 14148 3612 14154 3664
rect 14200 3624 14780 3652
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 3436 3556 5089 3584
rect 5077 3553 5089 3556
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3553 5411 3587
rect 5353 3547 5411 3553
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 6178 3584 6184 3596
rect 5491 3556 6184 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4246 3516 4252 3528
rect 3651 3488 4252 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4706 3516 4712 3528
rect 4356 3488 4712 3516
rect 2032 3451 2090 3457
rect 2032 3417 2044 3451
rect 2078 3448 2090 3451
rect 2774 3448 2780 3460
rect 2078 3420 2780 3448
rect 2078 3417 2090 3420
rect 2032 3411 2090 3417
rect 2774 3408 2780 3420
rect 2832 3408 2838 3460
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 3326 3448 3332 3460
rect 3108 3420 3332 3448
rect 3108 3408 3114 3420
rect 3326 3408 3332 3420
rect 3384 3448 3390 3460
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3384 3420 3893 3448
rect 3384 3408 3390 3420
rect 3881 3417 3893 3420
rect 3927 3448 3939 3451
rect 4356 3448 4384 3488
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 5460 3516 5488 3547
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 8496 3556 10609 3584
rect 4847 3488 5488 3516
rect 5813 3519 5871 3525
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 5994 3516 6000 3528
rect 5859 3488 6000 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6512 3488 6745 3516
rect 6512 3476 6518 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 7374 3516 7380 3528
rect 7331 3488 7380 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 4890 3448 4896 3460
rect 3927 3420 4384 3448
rect 4540 3420 4896 3448
rect 3927 3417 3939 3420
rect 3881 3411 3939 3417
rect 4341 3383 4399 3389
rect 4341 3349 4353 3383
rect 4387 3380 4399 3383
rect 4540 3380 4568 3420
rect 4890 3408 4896 3420
rect 4948 3448 4954 3460
rect 5537 3451 5595 3457
rect 5537 3448 5549 3451
rect 4948 3420 5549 3448
rect 4948 3408 4954 3420
rect 5537 3417 5549 3420
rect 5583 3417 5595 3451
rect 5537 3411 5595 3417
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6365 3451 6423 3457
rect 6365 3448 6377 3451
rect 5960 3420 6377 3448
rect 5960 3408 5966 3420
rect 6365 3417 6377 3420
rect 6411 3448 6423 3451
rect 6840 3448 6868 3476
rect 6411 3420 6868 3448
rect 7024 3448 7052 3479
rect 7374 3476 7380 3488
rect 7432 3516 7438 3528
rect 8496 3516 8524 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 14200 3584 14228 3624
rect 14752 3596 14780 3624
rect 10597 3547 10655 3553
rect 11624 3556 14228 3584
rect 7432 3488 8524 3516
rect 7432 3476 7438 3488
rect 8938 3476 8944 3528
rect 8996 3476 9002 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9088 3488 10241 3516
rect 9088 3476 9094 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 11624 3516 11652 3556
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14734 3544 14740 3596
rect 14792 3544 14798 3596
rect 15746 3584 15752 3596
rect 15212 3556 15752 3584
rect 10229 3479 10287 3485
rect 10796 3488 11652 3516
rect 7552 3451 7610 3457
rect 7024 3420 7512 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 4387 3352 4568 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 4614 3340 4620 3392
rect 4672 3340 4678 3392
rect 4709 3383 4767 3389
rect 4709 3349 4721 3383
rect 4755 3380 4767 3383
rect 4798 3380 4804 3392
rect 4755 3352 4804 3380
rect 4755 3349 4767 3352
rect 4709 3343 4767 3349
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 4982 3340 4988 3392
rect 5040 3340 5046 3392
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 7484 3380 7512 3420
rect 7552 3417 7564 3451
rect 7598 3448 7610 3451
rect 7742 3448 7748 3460
rect 7598 3420 7748 3448
rect 7598 3417 7610 3420
rect 7552 3411 7610 3417
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 9769 3451 9827 3457
rect 9769 3448 9781 3451
rect 9364 3420 9781 3448
rect 9364 3408 9370 3420
rect 9769 3417 9781 3420
rect 9815 3448 9827 3451
rect 10796 3448 10824 3488
rect 12066 3476 12072 3528
rect 12124 3476 12130 3528
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13403 3488 14688 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 9815 3420 10824 3448
rect 10864 3451 10922 3457
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 10864 3417 10876 3451
rect 10910 3448 10922 3451
rect 11330 3448 11336 3460
rect 10910 3420 11336 3448
rect 10910 3417 10922 3420
rect 10864 3411 10922 3417
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12584 3420 12909 3448
rect 12584 3408 12590 3420
rect 12897 3417 12909 3420
rect 12943 3417 12955 3451
rect 12897 3411 12955 3417
rect 13909 3451 13967 3457
rect 13909 3417 13921 3451
rect 13955 3448 13967 3451
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 13955 3420 14473 3448
rect 13955 3417 13967 3420
rect 13909 3411 13967 3417
rect 14461 3417 14473 3420
rect 14507 3417 14519 3451
rect 14461 3411 14519 3417
rect 14660 3392 14688 3488
rect 15102 3476 15108 3528
rect 15160 3476 15166 3528
rect 15212 3525 15240 3556
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 15470 3476 15476 3528
rect 15528 3476 15534 3528
rect 15562 3476 15568 3528
rect 15620 3476 15626 3528
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 15856 3516 15884 3692
rect 16114 3612 16120 3664
rect 16172 3612 16178 3664
rect 17236 3652 17264 3692
rect 17310 3680 17316 3732
rect 17368 3680 17374 3732
rect 18322 3720 18328 3732
rect 17420 3692 18328 3720
rect 17420 3652 17448 3692
rect 18322 3680 18328 3692
rect 18380 3720 18386 3732
rect 18785 3723 18843 3729
rect 18785 3720 18797 3723
rect 18380 3692 18797 3720
rect 18380 3680 18386 3692
rect 18785 3689 18797 3692
rect 18831 3689 18843 3723
rect 18785 3683 18843 3689
rect 19150 3680 19156 3732
rect 19208 3680 19214 3732
rect 19978 3680 19984 3732
rect 20036 3680 20042 3732
rect 20990 3680 20996 3732
rect 21048 3720 21054 3732
rect 22189 3723 22247 3729
rect 22189 3720 22201 3723
rect 21048 3692 22201 3720
rect 21048 3680 21054 3692
rect 22189 3689 22201 3692
rect 22235 3689 22247 3723
rect 22189 3683 22247 3689
rect 22278 3680 22284 3732
rect 22336 3680 22342 3732
rect 24302 3720 24308 3732
rect 22388 3692 24308 3720
rect 17236 3624 17448 3652
rect 16206 3544 16212 3596
rect 16264 3584 16270 3596
rect 16510 3587 16568 3593
rect 16510 3584 16522 3587
rect 16264 3556 16522 3584
rect 16264 3544 16270 3556
rect 16510 3553 16522 3556
rect 16556 3553 16568 3587
rect 16510 3547 16568 3553
rect 16666 3544 16672 3596
rect 16724 3544 16730 3596
rect 19168 3584 19196 3680
rect 21450 3612 21456 3664
rect 21508 3612 21514 3664
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 19168 3556 19349 3584
rect 19337 3553 19349 3556
rect 19383 3553 19395 3587
rect 21468 3584 21496 3612
rect 22388 3593 22416 3692
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 24394 3680 24400 3732
rect 24452 3720 24458 3732
rect 26602 3720 26608 3732
rect 24452 3692 26608 3720
rect 24452 3680 24458 3692
rect 26602 3680 26608 3692
rect 26660 3680 26666 3732
rect 26694 3680 26700 3732
rect 26752 3680 26758 3732
rect 27246 3720 27252 3732
rect 26804 3692 27252 3720
rect 22738 3612 22744 3664
rect 22796 3612 22802 3664
rect 24213 3655 24271 3661
rect 24213 3621 24225 3655
rect 24259 3652 24271 3655
rect 26804 3652 26832 3692
rect 27246 3680 27252 3692
rect 27304 3680 27310 3732
rect 29178 3680 29184 3732
rect 29236 3720 29242 3732
rect 29549 3723 29607 3729
rect 29549 3720 29561 3723
rect 29236 3692 29561 3720
rect 29236 3680 29242 3692
rect 29549 3689 29561 3692
rect 29595 3689 29607 3723
rect 31662 3720 31668 3732
rect 29549 3683 29607 3689
rect 30392 3692 31668 3720
rect 24259 3624 25360 3652
rect 24259 3621 24271 3624
rect 24213 3615 24271 3621
rect 25332 3596 25360 3624
rect 25424 3624 26832 3652
rect 21545 3587 21603 3593
rect 21545 3584 21557 3587
rect 21468 3556 21557 3584
rect 19337 3547 19395 3553
rect 21545 3553 21557 3556
rect 21591 3553 21603 3587
rect 21545 3547 21603 3553
rect 22373 3587 22431 3593
rect 22373 3553 22385 3587
rect 22419 3553 22431 3587
rect 22373 3547 22431 3553
rect 22830 3544 22836 3596
rect 22888 3544 22894 3596
rect 24762 3544 24768 3596
rect 24820 3584 24826 3596
rect 24857 3587 24915 3593
rect 24857 3584 24869 3587
rect 24820 3556 24869 3584
rect 24820 3544 24826 3556
rect 24857 3553 24869 3556
rect 24903 3553 24915 3587
rect 24857 3547 24915 3553
rect 25038 3544 25044 3596
rect 25096 3544 25102 3596
rect 25314 3544 25320 3596
rect 25372 3544 25378 3596
rect 15703 3488 15884 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16390 3476 16396 3528
rect 16448 3476 16454 3528
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3516 17463 3519
rect 17494 3516 17500 3528
rect 17451 3488 17500 3516
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 19610 3476 19616 3528
rect 19668 3476 19674 3528
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20714 3516 20720 3528
rect 20119 3488 20720 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 22066 3488 22569 3516
rect 14921 3451 14979 3457
rect 14921 3417 14933 3451
rect 14967 3448 14979 3451
rect 15580 3448 15608 3476
rect 14967 3420 15608 3448
rect 17672 3451 17730 3457
rect 14967 3417 14979 3420
rect 14921 3411 14979 3417
rect 17672 3417 17684 3451
rect 17718 3448 17730 3451
rect 17770 3448 17776 3460
rect 17718 3420 17776 3448
rect 17718 3417 17730 3420
rect 17672 3411 17730 3417
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 9858 3380 9864 3392
rect 7484 3352 9864 3380
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 14642 3340 14648 3392
rect 14700 3340 14706 3392
rect 15381 3383 15439 3389
rect 15381 3349 15393 3383
rect 15427 3380 15439 3383
rect 16298 3380 16304 3392
rect 15427 3352 16304 3380
rect 15427 3349 15439 3352
rect 15381 3343 15439 3349
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 19628 3380 19656 3476
rect 20340 3451 20398 3457
rect 20340 3417 20352 3451
rect 20386 3448 20398 3451
rect 21358 3448 21364 3460
rect 20386 3420 21364 3448
rect 20386 3417 20398 3420
rect 20340 3411 20398 3417
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 16724 3352 19656 3380
rect 16724 3340 16730 3352
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 22066 3380 22094 3488
rect 22557 3485 22569 3488
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 25424 3516 25452 3624
rect 25774 3544 25780 3596
rect 25832 3544 25838 3596
rect 26234 3544 26240 3596
rect 26292 3584 26298 3596
rect 27062 3584 27068 3596
rect 26292 3556 27068 3584
rect 26292 3544 26298 3556
rect 27062 3544 27068 3556
rect 27120 3544 27126 3596
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 29089 3587 29147 3593
rect 29089 3584 29101 3587
rect 28224 3556 29101 3584
rect 28224 3544 28230 3556
rect 29089 3553 29101 3556
rect 29135 3553 29147 3587
rect 30101 3587 30159 3593
rect 30101 3584 30113 3587
rect 29089 3547 29147 3553
rect 29196 3556 30113 3584
rect 22796 3488 25452 3516
rect 25792 3516 25820 3544
rect 26053 3519 26111 3525
rect 26053 3516 26065 3519
rect 25792 3488 26065 3516
rect 22796 3476 22802 3488
rect 26053 3485 26065 3488
rect 26099 3485 26111 3519
rect 26053 3479 26111 3485
rect 26418 3476 26424 3528
rect 26476 3476 26482 3528
rect 26878 3476 26884 3528
rect 26936 3476 26942 3528
rect 29196 3516 29224 3556
rect 30101 3553 30113 3556
rect 30147 3553 30159 3587
rect 30101 3547 30159 3553
rect 30282 3544 30288 3596
rect 30340 3544 30346 3596
rect 30392 3593 30420 3692
rect 31662 3680 31668 3692
rect 31720 3720 31726 3732
rect 31720 3692 32260 3720
rect 31720 3680 31726 3692
rect 31386 3612 31392 3664
rect 31444 3652 31450 3664
rect 31757 3655 31815 3661
rect 31757 3652 31769 3655
rect 31444 3624 31769 3652
rect 31444 3612 31450 3624
rect 31757 3621 31769 3624
rect 31803 3621 31815 3655
rect 31757 3615 31815 3621
rect 32232 3593 32260 3692
rect 33594 3680 33600 3732
rect 33652 3680 33658 3732
rect 33962 3680 33968 3732
rect 34020 3720 34026 3732
rect 34425 3723 34483 3729
rect 34425 3720 34437 3723
rect 34020 3692 34437 3720
rect 34020 3680 34026 3692
rect 34425 3689 34437 3692
rect 34471 3689 34483 3723
rect 34425 3683 34483 3689
rect 34701 3723 34759 3729
rect 34701 3689 34713 3723
rect 34747 3689 34759 3723
rect 34701 3683 34759 3689
rect 34716 3652 34744 3683
rect 35158 3680 35164 3732
rect 35216 3680 35222 3732
rect 35894 3680 35900 3732
rect 35952 3720 35958 3732
rect 37550 3720 37556 3732
rect 35952 3692 37556 3720
rect 35952 3680 35958 3692
rect 37550 3680 37556 3692
rect 37608 3680 37614 3732
rect 39022 3680 39028 3732
rect 39080 3720 39086 3732
rect 41325 3723 41383 3729
rect 41325 3720 41337 3723
rect 39080 3692 41337 3720
rect 39080 3680 39086 3692
rect 41325 3689 41337 3692
rect 41371 3689 41383 3723
rect 42702 3720 42708 3732
rect 41325 3683 41383 3689
rect 42352 3692 42708 3720
rect 33244 3624 34744 3652
rect 30377 3587 30435 3593
rect 30377 3553 30389 3587
rect 30423 3553 30435 3587
rect 32217 3587 32275 3593
rect 30377 3547 30435 3553
rect 31726 3556 32168 3584
rect 26988 3488 29224 3516
rect 30009 3519 30067 3525
rect 22281 3451 22339 3457
rect 22281 3417 22293 3451
rect 22327 3448 22339 3451
rect 23100 3451 23158 3457
rect 22327 3420 22692 3448
rect 22327 3417 22339 3420
rect 22281 3411 22339 3417
rect 21600 3352 22094 3380
rect 22664 3380 22692 3420
rect 23100 3417 23112 3451
rect 23146 3448 23158 3451
rect 24118 3448 24124 3460
rect 23146 3420 24124 3448
rect 23146 3417 23158 3420
rect 23100 3411 23158 3417
rect 24118 3408 24124 3420
rect 24176 3408 24182 3460
rect 24765 3451 24823 3457
rect 24765 3417 24777 3451
rect 24811 3448 24823 3451
rect 25869 3451 25927 3457
rect 25869 3448 25881 3451
rect 24811 3420 25881 3448
rect 24811 3417 24823 3420
rect 24765 3411 24823 3417
rect 25869 3417 25881 3420
rect 25915 3417 25927 3451
rect 25869 3411 25927 3417
rect 26237 3451 26295 3457
rect 26237 3417 26249 3451
rect 26283 3448 26295 3451
rect 26436 3448 26464 3476
rect 26283 3420 26464 3448
rect 26283 3417 26295 3420
rect 26237 3411 26295 3417
rect 26602 3408 26608 3460
rect 26660 3448 26666 3460
rect 26988 3448 27016 3488
rect 30009 3485 30021 3519
rect 30055 3516 30067 3519
rect 30300 3516 30328 3544
rect 30055 3488 30328 3516
rect 30392 3488 31340 3516
rect 30055 3485 30067 3488
rect 30009 3479 30067 3485
rect 26660 3420 27016 3448
rect 27332 3451 27390 3457
rect 26660 3408 26666 3420
rect 27332 3417 27344 3451
rect 27378 3448 27390 3451
rect 28350 3448 28356 3460
rect 27378 3420 28356 3448
rect 27378 3417 27390 3420
rect 27332 3411 27390 3417
rect 28350 3408 28356 3420
rect 28408 3408 28414 3460
rect 30392 3448 30420 3488
rect 31312 3460 31340 3488
rect 28460 3420 30420 3448
rect 30644 3451 30702 3457
rect 28460 3392 28488 3420
rect 30644 3417 30656 3451
rect 30690 3448 30702 3451
rect 31202 3448 31208 3460
rect 30690 3420 31208 3448
rect 30690 3417 30702 3420
rect 30644 3411 30702 3417
rect 31202 3408 31208 3420
rect 31260 3408 31266 3460
rect 31294 3408 31300 3460
rect 31352 3408 31358 3460
rect 24026 3380 24032 3392
rect 22664 3352 24032 3380
rect 21600 3340 21606 3352
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 24394 3340 24400 3392
rect 24452 3340 24458 3392
rect 25038 3340 25044 3392
rect 25096 3380 25102 3392
rect 28166 3380 28172 3392
rect 25096 3352 28172 3380
rect 25096 3340 25102 3352
rect 28166 3340 28172 3352
rect 28224 3340 28230 3392
rect 28442 3340 28448 3392
rect 28500 3340 28506 3392
rect 28534 3340 28540 3392
rect 28592 3340 28598 3392
rect 28902 3340 28908 3392
rect 28960 3340 28966 3392
rect 28997 3383 29055 3389
rect 28997 3349 29009 3383
rect 29043 3380 29055 3383
rect 29086 3380 29092 3392
rect 29043 3352 29092 3380
rect 29043 3349 29055 3352
rect 28997 3343 29055 3349
rect 29086 3340 29092 3352
rect 29144 3380 29150 3392
rect 29917 3383 29975 3389
rect 29917 3380 29929 3383
rect 29144 3352 29929 3380
rect 29144 3340 29150 3352
rect 29917 3349 29929 3352
rect 29963 3380 29975 3383
rect 30742 3380 30748 3392
rect 29963 3352 30748 3380
rect 29963 3349 29975 3352
rect 29917 3343 29975 3349
rect 30742 3340 30748 3352
rect 30800 3340 30806 3392
rect 30834 3340 30840 3392
rect 30892 3380 30898 3392
rect 31726 3380 31754 3556
rect 32030 3476 32036 3528
rect 32088 3476 32094 3528
rect 32140 3516 32168 3556
rect 32217 3553 32229 3587
rect 32263 3553 32275 3587
rect 32217 3547 32275 3553
rect 33244 3516 33272 3624
rect 33873 3587 33931 3593
rect 33873 3553 33885 3587
rect 33919 3584 33931 3587
rect 34330 3584 34336 3596
rect 33919 3556 34336 3584
rect 33919 3553 33931 3556
rect 33873 3547 33931 3553
rect 34330 3544 34336 3556
rect 34388 3544 34394 3596
rect 35912 3593 35940 3680
rect 35253 3587 35311 3593
rect 35253 3584 35265 3587
rect 34808 3556 35265 3584
rect 34808 3528 34836 3556
rect 35253 3553 35265 3556
rect 35299 3553 35311 3587
rect 35253 3547 35311 3553
rect 35897 3587 35955 3593
rect 35897 3553 35909 3587
rect 35943 3553 35955 3587
rect 37568 3584 37596 3680
rect 39390 3612 39396 3664
rect 39448 3652 39454 3664
rect 39669 3655 39727 3661
rect 39669 3652 39681 3655
rect 39448 3624 39681 3652
rect 39448 3612 39454 3624
rect 39669 3621 39681 3624
rect 39715 3652 39727 3655
rect 39715 3624 41460 3652
rect 39715 3621 39727 3624
rect 39669 3615 39727 3621
rect 38289 3587 38347 3593
rect 38289 3584 38301 3587
rect 35897 3547 35955 3553
rect 37292 3556 37504 3584
rect 37568 3556 38301 3584
rect 32140 3488 33272 3516
rect 34790 3476 34796 3528
rect 34848 3476 34854 3528
rect 34882 3476 34888 3528
rect 34940 3476 34946 3528
rect 34974 3476 34980 3528
rect 35032 3476 35038 3528
rect 35437 3519 35495 3525
rect 35437 3485 35449 3519
rect 35483 3516 35495 3519
rect 35986 3516 35992 3528
rect 35483 3488 35992 3516
rect 35483 3485 35495 3488
rect 35437 3479 35495 3485
rect 35986 3476 35992 3488
rect 36044 3476 36050 3528
rect 37292 3516 37320 3556
rect 36096 3488 37320 3516
rect 32484 3451 32542 3457
rect 32484 3417 32496 3451
rect 32530 3448 32542 3451
rect 34238 3448 34244 3460
rect 32530 3420 34244 3448
rect 32530 3417 32542 3420
rect 32484 3411 32542 3417
rect 34238 3408 34244 3420
rect 34296 3408 34302 3460
rect 34701 3451 34759 3457
rect 34701 3417 34713 3451
rect 34747 3448 34759 3451
rect 36096 3448 36124 3488
rect 37366 3476 37372 3528
rect 37424 3476 37430 3528
rect 37476 3516 37504 3556
rect 38289 3553 38301 3556
rect 38335 3553 38347 3587
rect 38289 3547 38347 3553
rect 40497 3587 40555 3593
rect 40497 3553 40509 3587
rect 40543 3584 40555 3587
rect 40954 3584 40960 3596
rect 40543 3556 40960 3584
rect 40543 3553 40555 3556
rect 40497 3547 40555 3553
rect 40954 3544 40960 3556
rect 41012 3544 41018 3596
rect 41432 3593 41460 3624
rect 41417 3587 41475 3593
rect 41417 3553 41429 3587
rect 41463 3553 41475 3587
rect 41417 3547 41475 3553
rect 42242 3544 42248 3596
rect 42300 3544 42306 3596
rect 42352 3593 42380 3692
rect 42702 3680 42708 3692
rect 42760 3680 42766 3732
rect 43070 3680 43076 3732
rect 43128 3720 43134 3732
rect 44637 3723 44695 3729
rect 43128 3692 44588 3720
rect 43128 3680 43134 3692
rect 43717 3655 43775 3661
rect 43717 3621 43729 3655
rect 43763 3652 43775 3655
rect 44082 3652 44088 3664
rect 43763 3624 44088 3652
rect 43763 3621 43775 3624
rect 43717 3615 43775 3621
rect 44082 3612 44088 3624
rect 44140 3612 44146 3664
rect 42337 3587 42395 3593
rect 42337 3553 42349 3587
rect 42383 3553 42395 3587
rect 42337 3547 42395 3553
rect 44174 3544 44180 3596
rect 44232 3584 44238 3596
rect 44269 3587 44327 3593
rect 44269 3584 44281 3587
rect 44232 3556 44281 3584
rect 44232 3544 44238 3556
rect 44269 3553 44281 3556
rect 44315 3553 44327 3587
rect 44269 3547 44327 3553
rect 44450 3544 44456 3596
rect 44508 3544 44514 3596
rect 38930 3516 38936 3528
rect 37476 3488 38936 3516
rect 38930 3476 38936 3488
rect 38988 3476 38994 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 39316 3488 40693 3516
rect 34747 3420 36124 3448
rect 36164 3451 36222 3457
rect 34747 3417 34759 3420
rect 34701 3411 34759 3417
rect 36164 3417 36176 3451
rect 36210 3448 36222 3451
rect 38013 3451 38071 3457
rect 38013 3448 38025 3451
rect 36210 3420 38025 3448
rect 36210 3417 36222 3420
rect 36164 3411 36222 3417
rect 38013 3417 38025 3420
rect 38059 3417 38071 3451
rect 38013 3411 38071 3417
rect 38556 3451 38614 3457
rect 38556 3417 38568 3451
rect 38602 3448 38614 3451
rect 39206 3448 39212 3460
rect 38602 3420 39212 3448
rect 38602 3417 38614 3420
rect 38556 3411 38614 3417
rect 39206 3408 39212 3420
rect 39264 3408 39270 3460
rect 30892 3352 31754 3380
rect 31849 3383 31907 3389
rect 30892 3340 30898 3352
rect 31849 3349 31861 3383
rect 31895 3380 31907 3383
rect 33502 3380 33508 3392
rect 31895 3352 33508 3380
rect 31895 3349 31907 3352
rect 31849 3343 31907 3349
rect 33502 3340 33508 3352
rect 33560 3340 33566 3392
rect 35618 3340 35624 3392
rect 35676 3340 35682 3392
rect 35710 3340 35716 3392
rect 35768 3380 35774 3392
rect 37277 3383 37335 3389
rect 37277 3380 37289 3383
rect 35768 3352 37289 3380
rect 35768 3340 35774 3352
rect 37277 3349 37289 3352
rect 37323 3349 37335 3383
rect 37277 3343 37335 3349
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39316 3380 39344 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 42260 3516 42288 3544
rect 43346 3516 43352 3528
rect 42260 3488 43352 3516
rect 40681 3479 40739 3485
rect 43346 3476 43352 3488
rect 43404 3476 43410 3528
rect 40218 3408 40224 3460
rect 40276 3408 40282 3460
rect 40313 3451 40371 3457
rect 40313 3417 40325 3451
rect 40359 3448 40371 3451
rect 42061 3451 42119 3457
rect 42061 3448 42073 3451
rect 40359 3420 42073 3448
rect 40359 3417 40371 3420
rect 40313 3411 40371 3417
rect 42061 3417 42073 3420
rect 42107 3417 42119 3451
rect 42061 3411 42119 3417
rect 42604 3451 42662 3457
rect 42604 3417 42616 3451
rect 42650 3448 42662 3451
rect 43898 3448 43904 3460
rect 42650 3420 43904 3448
rect 42650 3417 42662 3420
rect 42604 3411 42662 3417
rect 43898 3408 43904 3420
rect 43956 3408 43962 3460
rect 38436 3352 39344 3380
rect 38436 3340 38442 3352
rect 39850 3340 39856 3392
rect 39908 3340 39914 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 43714 3380 43720 3392
rect 41932 3352 43720 3380
rect 41932 3340 41938 3352
rect 43714 3340 43720 3352
rect 43772 3340 43778 3392
rect 43806 3340 43812 3392
rect 43864 3340 43870 3392
rect 44174 3340 44180 3392
rect 44232 3340 44238 3392
rect 44560 3380 44588 3692
rect 44637 3689 44649 3723
rect 44683 3720 44695 3723
rect 44818 3720 44824 3732
rect 44683 3692 44824 3720
rect 44683 3689 44695 3692
rect 44637 3683 44695 3689
rect 44818 3680 44824 3692
rect 44876 3680 44882 3732
rect 45830 3680 45836 3732
rect 45888 3720 45894 3732
rect 45888 3692 46244 3720
rect 45888 3680 45894 3692
rect 46216 3584 46244 3692
rect 46474 3680 46480 3732
rect 46532 3680 46538 3732
rect 47394 3680 47400 3732
rect 47452 3680 47458 3732
rect 47762 3680 47768 3732
rect 47820 3680 47826 3732
rect 49418 3680 49424 3732
rect 49476 3680 49482 3732
rect 49786 3680 49792 3732
rect 49844 3680 49850 3732
rect 50706 3680 50712 3732
rect 50764 3720 50770 3732
rect 50764 3692 52868 3720
rect 50764 3680 50770 3692
rect 47670 3612 47676 3664
rect 47728 3612 47734 3664
rect 46569 3587 46627 3593
rect 46569 3584 46581 3587
rect 46216 3556 46581 3584
rect 46569 3553 46581 3556
rect 46615 3553 46627 3587
rect 46569 3547 46627 3553
rect 47578 3544 47584 3596
rect 47636 3544 47642 3596
rect 44818 3476 44824 3528
rect 44876 3476 44882 3528
rect 45097 3519 45155 3525
rect 45097 3485 45109 3519
rect 45143 3516 45155 3519
rect 45186 3516 45192 3528
rect 45143 3488 45192 3516
rect 45143 3485 45155 3488
rect 45097 3479 45155 3485
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 47681 3525 47709 3612
rect 47780 3584 47808 3680
rect 49436 3652 49464 3680
rect 50433 3655 50491 3661
rect 50433 3652 50445 3655
rect 49436 3624 50445 3652
rect 50433 3621 50445 3624
rect 50479 3621 50491 3655
rect 50433 3615 50491 3621
rect 47780 3556 48176 3584
rect 47673 3519 47731 3525
rect 47673 3485 47685 3519
rect 47719 3485 47731 3519
rect 47673 3479 47731 3485
rect 48038 3476 48044 3528
rect 48096 3476 48102 3528
rect 48148 3525 48176 3556
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 52730 3584 52736 3596
rect 50580 3556 51396 3584
rect 50580 3544 50586 3556
rect 48133 3519 48191 3525
rect 48133 3485 48145 3519
rect 48179 3485 48191 3519
rect 48133 3479 48191 3485
rect 48409 3519 48467 3525
rect 48409 3485 48421 3519
rect 48455 3516 48467 3519
rect 50540 3516 50568 3544
rect 48455 3488 50568 3516
rect 48455 3485 48467 3488
rect 48409 3479 48467 3485
rect 50982 3476 50988 3528
rect 51040 3476 51046 3528
rect 51368 3525 51396 3556
rect 52656 3556 52736 3584
rect 51077 3519 51135 3525
rect 51077 3485 51089 3519
rect 51123 3485 51135 3519
rect 51077 3479 51135 3485
rect 51353 3519 51411 3525
rect 51353 3485 51365 3519
rect 51399 3516 51411 3519
rect 52656 3516 52684 3556
rect 52730 3544 52736 3556
rect 52788 3544 52794 3596
rect 52840 3584 52868 3692
rect 54202 3680 54208 3732
rect 54260 3680 54266 3732
rect 54941 3723 54999 3729
rect 54941 3689 54953 3723
rect 54987 3720 54999 3723
rect 58345 3723 58403 3729
rect 58345 3720 58357 3723
rect 54987 3692 58357 3720
rect 54987 3689 54999 3692
rect 54941 3683 54999 3689
rect 58345 3689 58357 3692
rect 58391 3689 58403 3723
rect 58345 3683 58403 3689
rect 53760 3624 54156 3652
rect 53760 3593 53788 3624
rect 54128 3596 54156 3624
rect 53377 3587 53435 3593
rect 53377 3584 53389 3587
rect 52840 3556 53389 3584
rect 53377 3553 53389 3556
rect 53423 3553 53435 3587
rect 53377 3547 53435 3553
rect 53745 3587 53803 3593
rect 53745 3553 53757 3587
rect 53791 3553 53803 3587
rect 53745 3547 53803 3553
rect 53760 3516 53788 3547
rect 53834 3544 53840 3596
rect 53892 3544 53898 3596
rect 54110 3544 54116 3596
rect 54168 3544 54174 3596
rect 54220 3584 54248 3680
rect 58250 3612 58256 3664
rect 58308 3612 58314 3664
rect 54220 3556 54616 3584
rect 51399 3488 52684 3516
rect 52748 3488 53788 3516
rect 53852 3516 53880 3544
rect 54588 3525 54616 3556
rect 56870 3544 56876 3596
rect 56928 3544 56934 3596
rect 54481 3519 54539 3525
rect 54481 3516 54493 3519
rect 53852 3488 54493 3516
rect 51399 3485 51411 3488
rect 51353 3479 51411 3485
rect 45364 3451 45422 3457
rect 45364 3417 45376 3451
rect 45410 3448 45422 3451
rect 47213 3451 47271 3457
rect 47213 3448 47225 3451
rect 45410 3420 47225 3448
rect 45410 3417 45422 3420
rect 45364 3411 45422 3417
rect 47213 3417 47225 3420
rect 47259 3417 47271 3451
rect 47213 3411 47271 3417
rect 47397 3451 47455 3457
rect 47397 3417 47409 3451
rect 47443 3448 47455 3451
rect 48676 3451 48734 3457
rect 47443 3420 48636 3448
rect 47443 3417 47455 3420
rect 47397 3411 47455 3417
rect 47857 3383 47915 3389
rect 47857 3380 47869 3383
rect 44560 3352 47869 3380
rect 47857 3349 47869 3352
rect 47903 3349 47915 3383
rect 47857 3343 47915 3349
rect 48314 3340 48320 3392
rect 48372 3340 48378 3392
rect 48608 3380 48636 3420
rect 48676 3417 48688 3451
rect 48722 3448 48734 3451
rect 49510 3448 49516 3460
rect 48722 3420 49516 3448
rect 48722 3417 48734 3420
rect 48676 3411 48734 3417
rect 49510 3408 49516 3420
rect 49568 3408 49574 3460
rect 50246 3408 50252 3460
rect 50304 3408 50310 3460
rect 50430 3408 50436 3460
rect 50488 3448 50494 3460
rect 51092 3448 51120 3479
rect 50488 3420 51120 3448
rect 51620 3451 51678 3457
rect 50488 3408 50494 3420
rect 51620 3417 51632 3451
rect 51666 3448 51678 3451
rect 52546 3448 52552 3460
rect 51666 3420 52552 3448
rect 51666 3417 51678 3420
rect 51620 3411 51678 3417
rect 52546 3408 52552 3420
rect 52604 3408 52610 3460
rect 49694 3380 49700 3392
rect 48608 3352 49700 3380
rect 49694 3340 49700 3352
rect 49752 3340 49758 3392
rect 51258 3340 51264 3392
rect 51316 3340 51322 3392
rect 52748 3389 52776 3488
rect 54481 3485 54493 3488
rect 54527 3485 54539 3519
rect 54481 3479 54539 3485
rect 54573 3519 54631 3525
rect 54573 3485 54585 3519
rect 54619 3485 54631 3519
rect 54573 3479 54631 3485
rect 54941 3519 54999 3525
rect 54941 3485 54953 3519
rect 54987 3516 54999 3519
rect 55030 3516 55036 3528
rect 54987 3488 55036 3516
rect 54987 3485 54999 3488
rect 54941 3479 54999 3485
rect 55030 3476 55036 3488
rect 55088 3476 55094 3528
rect 55306 3476 55312 3528
rect 55364 3516 55370 3528
rect 56888 3516 56916 3544
rect 55364 3488 56916 3516
rect 55364 3476 55370 3488
rect 56962 3476 56968 3528
rect 57020 3516 57026 3528
rect 57129 3519 57187 3525
rect 57129 3516 57141 3519
rect 57020 3488 57141 3516
rect 57020 3476 57026 3488
rect 57129 3485 57141 3488
rect 57175 3485 57187 3519
rect 57129 3479 57187 3485
rect 57422 3476 57428 3528
rect 57480 3516 57486 3528
rect 58529 3519 58587 3525
rect 58529 3516 58541 3519
rect 57480 3488 58541 3516
rect 57480 3476 57486 3488
rect 58529 3485 58541 3488
rect 58575 3485 58587 3519
rect 58529 3479 58587 3485
rect 53193 3451 53251 3457
rect 53193 3417 53205 3451
rect 53239 3448 53251 3451
rect 54297 3451 54355 3457
rect 54297 3448 54309 3451
rect 53239 3420 54309 3448
rect 53239 3417 53251 3420
rect 53193 3411 53251 3417
rect 54297 3417 54309 3420
rect 54343 3417 54355 3451
rect 55576 3451 55634 3457
rect 54297 3411 54355 3417
rect 54588 3420 55536 3448
rect 54588 3392 54616 3420
rect 52733 3383 52791 3389
rect 52733 3349 52745 3383
rect 52779 3349 52791 3383
rect 52733 3343 52791 3349
rect 52822 3340 52828 3392
rect 52880 3340 52886 3392
rect 53282 3340 53288 3392
rect 53340 3340 53346 3392
rect 54570 3340 54576 3392
rect 54628 3340 54634 3392
rect 55122 3340 55128 3392
rect 55180 3340 55186 3392
rect 55508 3380 55536 3420
rect 55576 3417 55588 3451
rect 55622 3448 55634 3451
rect 58912 3448 58940 3896
rect 55622 3420 58940 3448
rect 55622 3417 55634 3420
rect 55576 3411 55634 3417
rect 56689 3383 56747 3389
rect 56689 3380 56701 3383
rect 55508 3352 56701 3380
rect 56689 3349 56701 3352
rect 56735 3349 56747 3383
rect 56689 3343 56747 3349
rect 1104 3290 59040 3312
rect 1104 3238 15394 3290
rect 15446 3238 15458 3290
rect 15510 3238 15522 3290
rect 15574 3238 15586 3290
rect 15638 3238 15650 3290
rect 15702 3238 29838 3290
rect 29890 3238 29902 3290
rect 29954 3238 29966 3290
rect 30018 3238 30030 3290
rect 30082 3238 30094 3290
rect 30146 3238 44282 3290
rect 44334 3238 44346 3290
rect 44398 3238 44410 3290
rect 44462 3238 44474 3290
rect 44526 3238 44538 3290
rect 44590 3238 58726 3290
rect 58778 3238 58790 3290
rect 58842 3238 58854 3290
rect 58906 3238 58918 3290
rect 58970 3238 58982 3290
rect 59034 3238 59040 3290
rect 1104 3216 59040 3238
rect 2774 3136 2780 3188
rect 2832 3136 2838 3188
rect 4525 3179 4583 3185
rect 3068 3148 3280 3176
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 3068 3108 3096 3148
rect 2648 3080 3096 3108
rect 3252 3108 3280 3148
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4614 3176 4620 3188
rect 4571 3148 4620 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 4764 3148 6193 3176
rect 4764 3136 4770 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7742 3136 7748 3188
rect 7800 3136 7806 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 8076 3148 8309 3176
rect 8076 3136 8082 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 8297 3139 8355 3145
rect 9214 3136 9220 3188
rect 9272 3136 9278 3188
rect 9858 3136 9864 3188
rect 9916 3136 9922 3188
rect 10321 3179 10379 3185
rect 10321 3145 10333 3179
rect 10367 3176 10379 3179
rect 10870 3176 10876 3188
rect 10367 3148 10876 3176
rect 10367 3145 10379 3148
rect 10321 3139 10379 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11330 3136 11336 3188
rect 11388 3136 11394 3188
rect 11514 3136 11520 3188
rect 11572 3136 11578 3188
rect 11606 3136 11612 3188
rect 11664 3136 11670 3188
rect 11882 3136 11888 3188
rect 11940 3136 11946 3188
rect 14642 3136 14648 3188
rect 14700 3176 14706 3188
rect 16114 3176 16120 3188
rect 14700 3148 16120 3176
rect 14700 3136 14706 3148
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 16209 3179 16267 3185
rect 16209 3145 16221 3179
rect 16255 3176 16267 3179
rect 16850 3176 16856 3188
rect 16255 3148 16856 3176
rect 16255 3145 16267 3148
rect 16209 3139 16267 3145
rect 16850 3136 16856 3148
rect 16908 3136 16914 3188
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 17678 3176 17684 3188
rect 17451 3148 17684 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 17828 3148 18889 3176
rect 17828 3136 17834 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 18877 3139 18935 3145
rect 20530 3136 20536 3188
rect 20588 3136 20594 3188
rect 21358 3136 21364 3188
rect 21416 3136 21422 3188
rect 21453 3179 21511 3185
rect 21453 3145 21465 3179
rect 21499 3176 21511 3179
rect 21542 3176 21548 3188
rect 21499 3148 21548 3176
rect 21499 3145 21511 3148
rect 21453 3139 21511 3145
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 21634 3136 21640 3188
rect 21692 3136 21698 3188
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 22005 3179 22063 3185
rect 22005 3176 22017 3179
rect 21784 3148 22017 3176
rect 21784 3136 21790 3148
rect 22005 3145 22017 3148
rect 22051 3145 22063 3179
rect 22005 3139 22063 3145
rect 22649 3179 22707 3185
rect 22649 3145 22661 3179
rect 22695 3176 22707 3179
rect 23106 3176 23112 3188
rect 22695 3148 23112 3176
rect 22695 3145 22707 3148
rect 22649 3139 22707 3145
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 23382 3136 23388 3188
rect 23440 3136 23446 3188
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 24394 3136 24400 3188
rect 24452 3136 24458 3188
rect 26789 3179 26847 3185
rect 26789 3145 26801 3179
rect 26835 3176 26847 3179
rect 26878 3176 26884 3188
rect 26835 3148 26884 3176
rect 26835 3145 26847 3148
rect 26789 3139 26847 3145
rect 26878 3136 26884 3148
rect 26936 3136 26942 3188
rect 28350 3136 28356 3188
rect 28408 3136 28414 3188
rect 28534 3136 28540 3188
rect 28592 3136 28598 3188
rect 28902 3136 28908 3188
rect 28960 3176 28966 3188
rect 29089 3179 29147 3185
rect 29089 3176 29101 3179
rect 28960 3148 29101 3176
rect 28960 3136 28966 3148
rect 29089 3145 29101 3148
rect 29135 3145 29147 3179
rect 29089 3139 29147 3145
rect 29546 3136 29552 3188
rect 29604 3136 29610 3188
rect 30653 3179 30711 3185
rect 30653 3145 30665 3179
rect 30699 3176 30711 3179
rect 30834 3176 30840 3188
rect 30699 3148 30840 3176
rect 30699 3145 30711 3148
rect 30653 3139 30711 3145
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 30929 3179 30987 3185
rect 30929 3145 30941 3179
rect 30975 3145 30987 3179
rect 30929 3139 30987 3145
rect 9232 3108 9260 3136
rect 10229 3111 10287 3117
rect 3252 3080 4752 3108
rect 9232 3080 9628 3108
rect 2648 3068 2654 3080
rect 2866 3000 2872 3052
rect 2924 3000 2930 3052
rect 3050 3000 3056 3052
rect 3108 3000 3114 3052
rect 3513 3043 3571 3049
rect 3160 3012 3464 3040
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 2240 2904 2268 2935
rect 3160 2904 3188 3012
rect 3237 2975 3295 2981
rect 3237 2941 3249 2975
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 2240 2876 3188 2904
rect 3252 2836 3280 2935
rect 3436 2904 3464 3012
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3528 2972 3556 3003
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 3970 3040 3976 3052
rect 3896 3012 3976 3040
rect 3896 2981 3924 3012
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4724 3049 4752 3080
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5408 3012 5733 3040
rect 5408 3000 5414 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5902 3000 5908 3052
rect 5960 3000 5966 3052
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 8251 3012 9321 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3528 2944 3893 2972
rect 3881 2941 3893 2944
rect 3927 2941 3939 2975
rect 3881 2935 3939 2941
rect 4798 2932 4804 2984
rect 4856 2932 4862 2984
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 5920 2972 5948 3000
rect 5583 2944 5948 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 4338 2904 4344 2916
rect 3436 2876 4344 2904
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 6012 2904 6040 3003
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 9600 3049 9628 3080
rect 10229 3077 10241 3111
rect 10275 3108 10287 3111
rect 11532 3108 11560 3136
rect 10275 3080 11560 3108
rect 11624 3108 11652 3136
rect 11977 3111 12035 3117
rect 11977 3108 11989 3111
rect 11624 3080 11989 3108
rect 10275 3077 10287 3080
rect 10229 3071 10287 3077
rect 11977 3077 11989 3080
rect 12023 3077 12035 3111
rect 11977 3071 12035 3077
rect 13532 3111 13590 3117
rect 13532 3077 13544 3111
rect 13578 3108 13590 3111
rect 13906 3108 13912 3120
rect 13578 3080 13912 3108
rect 13578 3077 13590 3080
rect 13532 3071 13590 3077
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 20162 3108 20168 3120
rect 18064 3080 20168 3108
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 13262 3000 13268 3052
rect 13320 3000 13326 3052
rect 14734 3000 14740 3052
rect 14792 3000 14798 3052
rect 16390 3000 16396 3052
rect 16448 3000 16454 3052
rect 16666 3000 16672 3052
rect 16724 3000 16730 3052
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 18064 3049 18092 3080
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17092 3012 17509 3040
rect 17092 3000 17098 3012
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 18196 3012 19165 3040
rect 18196 3000 18202 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 20548 3040 20576 3136
rect 21652 3108 21680 3136
rect 21913 3111 21971 3117
rect 21913 3108 21925 3111
rect 21652 3080 21925 3108
rect 21913 3077 21925 3080
rect 21959 3077 21971 3111
rect 24412 3108 24440 3136
rect 21913 3071 21971 3077
rect 23584 3080 24440 3108
rect 26053 3111 26111 3117
rect 20717 3043 20775 3049
rect 20717 3040 20729 3043
rect 19475 3012 20116 3040
rect 20548 3012 20729 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 6457 2975 6515 2981
rect 6457 2941 6469 2975
rect 6503 2972 6515 2975
rect 7006 2972 7012 2984
rect 6503 2944 7012 2972
rect 6503 2941 6515 2944
rect 6457 2935 6515 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 8481 2975 8539 2981
rect 7239 2944 7880 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7852 2913 7880 2944
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 4448 2876 6040 2904
rect 7837 2907 7895 2913
rect 3602 2836 3608 2848
rect 3252 2808 3608 2836
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 4448 2836 4476 2876
rect 7837 2873 7849 2907
rect 7883 2873 7895 2907
rect 8496 2904 8524 2935
rect 8754 2932 8760 2984
rect 8812 2932 8818 2984
rect 9306 2904 9312 2916
rect 8496 2876 9312 2904
rect 7837 2867 7895 2873
rect 9306 2864 9312 2876
rect 9364 2864 9370 2916
rect 3752 2808 4476 2836
rect 3752 2796 3758 2808
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 5445 2839 5503 2845
rect 5445 2836 5457 2839
rect 4764 2808 5457 2836
rect 4764 2796 4770 2808
rect 5445 2805 5457 2808
rect 5491 2805 5503 2839
rect 5445 2799 5503 2805
rect 5902 2796 5908 2848
rect 5960 2796 5966 2848
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 9508 2836 9536 3000
rect 10502 2932 10508 2984
rect 10560 2932 10566 2984
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2972 10839 2975
rect 12161 2975 12219 2981
rect 10827 2944 11560 2972
rect 10827 2941 10839 2944
rect 10781 2935 10839 2941
rect 11532 2913 11560 2944
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 12526 2972 12532 2984
rect 12207 2944 12532 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 12621 2975 12679 2981
rect 12621 2941 12633 2975
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 11517 2907 11575 2913
rect 11517 2873 11529 2907
rect 11563 2873 11575 2907
rect 12636 2904 12664 2935
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 14332 2944 15209 2972
rect 14332 2932 14338 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 13262 2904 13268 2916
rect 12636 2876 13268 2904
rect 11517 2867 11575 2873
rect 13262 2864 13268 2876
rect 13320 2864 13326 2916
rect 14918 2864 14924 2916
rect 14976 2864 14982 2916
rect 16684 2913 16712 3000
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17589 2975 17647 2981
rect 17589 2972 17601 2975
rect 16816 2944 17601 2972
rect 16816 2932 16822 2944
rect 17589 2941 17601 2944
rect 17635 2941 17647 2975
rect 17589 2935 17647 2941
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 19705 2975 19763 2981
rect 19705 2941 19717 2975
rect 19751 2941 19763 2975
rect 20088 2972 20116 3012
rect 20717 3009 20729 3012
rect 20763 3009 20775 3043
rect 20717 3003 20775 3009
rect 20898 3000 20904 3052
rect 20956 3000 20962 3052
rect 21358 3000 21364 3052
rect 21416 3040 21422 3052
rect 23584 3049 23612 3080
rect 26053 3077 26065 3111
rect 26099 3108 26111 3111
rect 27706 3108 27712 3120
rect 26099 3080 27712 3108
rect 26099 3077 26111 3080
rect 26053 3071 26111 3077
rect 27706 3068 27712 3080
rect 27764 3068 27770 3120
rect 21637 3043 21695 3049
rect 21637 3040 21649 3043
rect 21416 3012 21649 3040
rect 21416 3000 21422 3012
rect 21637 3009 21649 3012
rect 21683 3009 21695 3043
rect 21637 3003 21695 3009
rect 23569 3043 23627 3049
rect 23569 3009 23581 3043
rect 23615 3009 23627 3043
rect 23569 3003 23627 3009
rect 23750 3000 23756 3052
rect 23808 3040 23814 3052
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 23808 3012 24225 3040
rect 23808 3000 23814 3012
rect 24213 3009 24225 3012
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 25682 3000 25688 3052
rect 25740 3000 25746 3052
rect 25866 3000 25872 3052
rect 25924 3000 25930 3052
rect 27801 3043 27859 3049
rect 27801 3009 27813 3043
rect 27847 3040 27859 3043
rect 28552 3040 28580 3136
rect 27847 3012 28580 3040
rect 29365 3043 29423 3049
rect 27847 3009 27859 3012
rect 27801 3003 27859 3009
rect 29365 3009 29377 3043
rect 29411 3040 29423 3043
rect 29564 3040 29592 3136
rect 30944 3108 30972 3139
rect 31110 3136 31116 3188
rect 31168 3176 31174 3188
rect 31389 3179 31447 3185
rect 31389 3176 31401 3179
rect 31168 3148 31401 3176
rect 31168 3136 31174 3148
rect 31389 3145 31401 3148
rect 31435 3145 31447 3179
rect 31389 3139 31447 3145
rect 31478 3136 31484 3188
rect 31536 3176 31542 3188
rect 31846 3176 31852 3188
rect 31536 3148 31852 3176
rect 31536 3136 31542 3148
rect 31846 3136 31852 3148
rect 31904 3136 31910 3188
rect 32306 3136 32312 3188
rect 32364 3136 32370 3188
rect 32508 3148 33916 3176
rect 32508 3108 32536 3148
rect 30944 3080 32536 3108
rect 32677 3111 32735 3117
rect 32677 3077 32689 3111
rect 32723 3108 32735 3111
rect 33781 3111 33839 3117
rect 33781 3108 33793 3111
rect 32723 3080 33793 3108
rect 32723 3077 32735 3080
rect 32677 3071 32735 3077
rect 33781 3077 33793 3080
rect 33827 3077 33839 3111
rect 33781 3071 33839 3077
rect 29411 3012 29592 3040
rect 30837 3043 30895 3049
rect 29411 3009 29423 3012
rect 29365 3003 29423 3009
rect 30837 3009 30849 3043
rect 30883 3009 30895 3043
rect 30837 3003 30895 3009
rect 20916 2972 20944 3000
rect 20088 2944 20944 2972
rect 22833 2975 22891 2981
rect 19705 2935 19763 2941
rect 22833 2941 22845 2975
rect 22879 2941 22891 2975
rect 22833 2935 22891 2941
rect 16669 2907 16727 2913
rect 16669 2873 16681 2907
rect 16715 2873 16727 2907
rect 16669 2867 16727 2873
rect 17037 2907 17095 2913
rect 17037 2873 17049 2907
rect 17083 2904 17095 2907
rect 18248 2904 18276 2935
rect 17083 2876 18276 2904
rect 17083 2873 17095 2876
rect 17037 2867 17095 2873
rect 18506 2864 18512 2916
rect 18564 2864 18570 2916
rect 18966 2864 18972 2916
rect 19024 2864 19030 2916
rect 19150 2864 19156 2916
rect 19208 2904 19214 2916
rect 19720 2904 19748 2935
rect 19208 2876 19748 2904
rect 22848 2904 22876 2935
rect 24118 2932 24124 2984
rect 24176 2972 24182 2984
rect 24673 2975 24731 2981
rect 24673 2972 24685 2975
rect 24176 2944 24685 2972
rect 24176 2932 24182 2944
rect 24673 2941 24685 2944
rect 24719 2941 24731 2975
rect 24673 2935 24731 2941
rect 26237 2975 26295 2981
rect 26237 2941 26249 2975
rect 26283 2972 26295 2975
rect 26878 2972 26884 2984
rect 26283 2944 26884 2972
rect 26283 2941 26295 2944
rect 26237 2935 26295 2941
rect 26878 2932 26884 2944
rect 26936 2932 26942 2984
rect 27065 2975 27123 2981
rect 27065 2941 27077 2975
rect 27111 2972 27123 2975
rect 28350 2972 28356 2984
rect 27111 2944 28356 2972
rect 27111 2941 27123 2944
rect 27065 2935 27123 2941
rect 28350 2932 28356 2944
rect 28408 2932 28414 2984
rect 28442 2932 28448 2984
rect 28500 2932 28506 2984
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 29144 2944 29653 2972
rect 29144 2932 29150 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 27617 2907 27675 2913
rect 22848 2876 23520 2904
rect 19208 2864 19214 2876
rect 6880 2808 9536 2836
rect 6880 2796 6886 2808
rect 9766 2796 9772 2848
rect 9824 2796 9830 2848
rect 13173 2839 13231 2845
rect 13173 2805 13185 2839
rect 13219 2836 13231 2839
rect 14936 2836 14964 2864
rect 13219 2808 14964 2836
rect 17865 2839 17923 2845
rect 13219 2805 13231 2808
rect 13173 2799 13231 2805
rect 17865 2805 17877 2839
rect 17911 2836 17923 2839
rect 18524 2836 18552 2864
rect 23492 2848 23520 2876
rect 27617 2873 27629 2907
rect 27663 2904 27675 2907
rect 29270 2904 29276 2916
rect 27663 2876 29276 2904
rect 27663 2873 27675 2876
rect 27617 2867 27675 2873
rect 29270 2864 29276 2876
rect 29328 2864 29334 2916
rect 30852 2904 30880 3003
rect 30926 3000 30932 3052
rect 30984 3040 30990 3052
rect 31297 3043 31355 3049
rect 31297 3040 31309 3043
rect 30984 3012 31309 3040
rect 30984 3000 30990 3012
rect 31297 3009 31309 3012
rect 31343 3040 31355 3043
rect 31343 3012 31616 3040
rect 31343 3009 31355 3012
rect 31297 3003 31355 3009
rect 31478 2932 31484 2984
rect 31536 2932 31542 2984
rect 31588 2972 31616 3012
rect 31662 3000 31668 3052
rect 31720 3040 31726 3052
rect 33888 3049 33916 3148
rect 34238 3136 34244 3188
rect 34296 3176 34302 3188
rect 35253 3179 35311 3185
rect 35253 3176 35265 3179
rect 34296 3148 35265 3176
rect 34296 3136 34302 3148
rect 35253 3145 35265 3148
rect 35299 3145 35311 3179
rect 35253 3139 35311 3145
rect 36173 3179 36231 3185
rect 36173 3145 36185 3179
rect 36219 3176 36231 3179
rect 37366 3176 37372 3188
rect 36219 3148 37372 3176
rect 36219 3145 36231 3148
rect 36173 3139 36231 3145
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 37458 3136 37464 3188
rect 37516 3176 37522 3188
rect 37516 3148 37964 3176
rect 37516 3136 37522 3148
rect 36262 3068 36268 3120
rect 36320 3068 36326 3120
rect 36541 3111 36599 3117
rect 36541 3077 36553 3111
rect 36587 3108 36599 3111
rect 37734 3108 37740 3120
rect 36587 3080 37740 3108
rect 36587 3077 36599 3080
rect 36541 3071 36599 3077
rect 37734 3068 37740 3080
rect 37792 3068 37798 3120
rect 31941 3043 31999 3049
rect 31941 3040 31953 3043
rect 31720 3012 31953 3040
rect 31720 3000 31726 3012
rect 31941 3009 31953 3012
rect 31987 3009 31999 3043
rect 31941 3003 31999 3009
rect 33873 3043 33931 3049
rect 33873 3009 33885 3043
rect 33919 3009 33931 3043
rect 33873 3003 33931 3009
rect 34054 3000 34060 3052
rect 34112 3040 34118 3052
rect 34517 3043 34575 3049
rect 34517 3040 34529 3043
rect 34112 3012 34529 3040
rect 34112 3000 34118 3012
rect 34517 3009 34529 3012
rect 34563 3009 34575 3043
rect 34517 3003 34575 3009
rect 34606 3000 34612 3052
rect 34664 3000 34670 3052
rect 36170 3040 36176 3052
rect 35452 3012 36176 3040
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 31588 2944 32781 2972
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 32769 2935 32827 2941
rect 32858 2932 32864 2984
rect 32916 2972 32922 2984
rect 32916 2944 33088 2972
rect 32916 2932 32922 2944
rect 32950 2904 32956 2916
rect 30852 2876 32956 2904
rect 32950 2864 32956 2876
rect 33008 2864 33014 2916
rect 33060 2904 33088 2944
rect 33134 2932 33140 2984
rect 33192 2932 33198 2984
rect 35342 2932 35348 2984
rect 35400 2932 35406 2984
rect 33060 2876 33364 2904
rect 17911 2808 18552 2836
rect 17911 2805 17923 2808
rect 17865 2799 17923 2805
rect 23474 2796 23480 2848
rect 23532 2796 23538 2848
rect 31754 2796 31760 2848
rect 31812 2796 31818 2848
rect 33336 2836 33364 2876
rect 33502 2864 33508 2916
rect 33560 2904 33566 2916
rect 35452 2904 35480 3012
rect 36170 3000 36176 3012
rect 36228 3000 36234 3052
rect 36280 3040 36308 3068
rect 36633 3043 36691 3049
rect 36633 3040 36645 3043
rect 36280 3012 36645 3040
rect 36633 3009 36645 3012
rect 36679 3009 36691 3043
rect 36633 3003 36691 3009
rect 37553 3043 37611 3049
rect 37553 3009 37565 3043
rect 37599 3040 37611 3043
rect 37826 3040 37832 3052
rect 37599 3012 37832 3040
rect 37599 3009 37611 3012
rect 37553 3003 37611 3009
rect 37826 3000 37832 3012
rect 37884 3000 37890 3052
rect 37936 3040 37964 3148
rect 38930 3136 38936 3188
rect 38988 3136 38994 3188
rect 39206 3136 39212 3188
rect 39264 3136 39270 3188
rect 39850 3136 39856 3188
rect 39908 3136 39914 3188
rect 40586 3136 40592 3188
rect 40644 3136 40650 3188
rect 41598 3176 41604 3188
rect 41386 3148 41604 3176
rect 39117 3043 39175 3049
rect 39117 3040 39129 3043
rect 37936 3012 39129 3040
rect 39117 3009 39129 3012
rect 39163 3009 39175 3043
rect 39117 3003 39175 3009
rect 36725 2975 36783 2981
rect 36725 2941 36737 2975
rect 36771 2941 36783 2975
rect 36725 2935 36783 2941
rect 36630 2904 36636 2916
rect 33560 2876 35480 2904
rect 35636 2876 36636 2904
rect 33560 2864 33566 2876
rect 34422 2836 34428 2848
rect 33336 2808 34428 2836
rect 34422 2796 34428 2808
rect 34480 2836 34486 2848
rect 35636 2836 35664 2876
rect 36630 2864 36636 2876
rect 36688 2904 36694 2916
rect 36740 2904 36768 2935
rect 37642 2932 37648 2984
rect 37700 2972 37706 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37700 2944 37933 2972
rect 37700 2932 37706 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 39224 2972 39252 3136
rect 39301 3043 39359 3049
rect 39301 3009 39313 3043
rect 39347 3040 39359 3043
rect 39868 3040 39896 3136
rect 39942 3068 39948 3120
rect 40000 3068 40006 3120
rect 39347 3012 39896 3040
rect 39960 3040 39988 3068
rect 40957 3043 41015 3049
rect 39960 3012 40172 3040
rect 39347 3009 39359 3012
rect 39301 3003 39359 3009
rect 39853 2975 39911 2981
rect 39853 2972 39865 2975
rect 39224 2944 39865 2972
rect 37921 2935 37979 2941
rect 39853 2941 39865 2944
rect 39899 2941 39911 2975
rect 39853 2935 39911 2941
rect 39945 2975 40003 2981
rect 39945 2941 39957 2975
rect 39991 2941 40003 2975
rect 39945 2935 40003 2941
rect 36688 2876 36768 2904
rect 36688 2864 36694 2876
rect 36814 2864 36820 2916
rect 36872 2904 36878 2916
rect 36872 2876 37780 2904
rect 36872 2864 36878 2876
rect 34480 2808 35664 2836
rect 34480 2796 34486 2808
rect 35986 2796 35992 2848
rect 36044 2796 36050 2848
rect 36262 2796 36268 2848
rect 36320 2836 36326 2848
rect 37458 2836 37464 2848
rect 36320 2808 37464 2836
rect 36320 2796 36326 2808
rect 37458 2796 37464 2808
rect 37516 2796 37522 2848
rect 37752 2836 37780 2876
rect 39960 2836 39988 2935
rect 40144 2904 40172 3012
rect 40957 3009 40969 3043
rect 41003 3040 41015 3043
rect 41386 3040 41414 3148
rect 41598 3136 41604 3148
rect 41656 3136 41662 3188
rect 43073 3179 43131 3185
rect 43073 3145 43085 3179
rect 43119 3176 43131 3179
rect 43530 3176 43536 3188
rect 43119 3148 43536 3176
rect 43119 3145 43131 3148
rect 43073 3139 43131 3145
rect 43530 3136 43536 3148
rect 43588 3136 43594 3188
rect 43806 3136 43812 3188
rect 43864 3136 43870 3188
rect 43898 3136 43904 3188
rect 43956 3136 43962 3188
rect 45554 3136 45560 3188
rect 45612 3176 45618 3188
rect 46201 3179 46259 3185
rect 46201 3176 46213 3179
rect 45612 3148 46213 3176
rect 45612 3136 45618 3148
rect 46201 3145 46213 3148
rect 46247 3145 46259 3179
rect 46201 3139 46259 3145
rect 47026 3136 47032 3188
rect 47084 3136 47090 3188
rect 47854 3136 47860 3188
rect 47912 3176 47918 3188
rect 48225 3179 48283 3185
rect 48225 3176 48237 3179
rect 47912 3148 48237 3176
rect 47912 3136 47918 3148
rect 48225 3145 48237 3148
rect 48271 3145 48283 3179
rect 51074 3176 51080 3188
rect 48225 3139 48283 3145
rect 48332 3148 51080 3176
rect 41003 3012 41414 3040
rect 43349 3043 43407 3049
rect 41003 3009 41015 3012
rect 40957 3003 41015 3009
rect 43349 3009 43361 3043
rect 43395 3040 43407 3043
rect 43824 3040 43852 3136
rect 45094 3108 45100 3120
rect 44284 3080 45100 3108
rect 44284 3049 44312 3080
rect 45094 3068 45100 3080
rect 45152 3068 45158 3120
rect 45278 3068 45284 3120
rect 45336 3108 45342 3120
rect 46661 3111 46719 3117
rect 46661 3108 46673 3111
rect 45336 3080 46673 3108
rect 45336 3068 45342 3080
rect 46661 3077 46673 3080
rect 46707 3077 46719 3111
rect 46661 3071 46719 3077
rect 43395 3012 43852 3040
rect 44269 3043 44327 3049
rect 43395 3009 43407 3012
rect 43349 3003 43407 3009
rect 44269 3009 44281 3043
rect 44315 3009 44327 3043
rect 44818 3040 44824 3052
rect 44269 3003 44327 3009
rect 44652 3012 44824 3040
rect 40678 2932 40684 2984
rect 40736 2972 40742 2984
rect 41233 2975 41291 2981
rect 41233 2972 41245 2975
rect 40736 2944 41245 2972
rect 40736 2932 40742 2944
rect 41233 2941 41245 2944
rect 41279 2941 41291 2975
rect 41233 2935 41291 2941
rect 41782 2932 41788 2984
rect 41840 2972 41846 2984
rect 42429 2975 42487 2981
rect 42429 2972 42441 2975
rect 41840 2944 42441 2972
rect 41840 2932 41846 2944
rect 42429 2941 42441 2944
rect 42475 2941 42487 2975
rect 42429 2935 42487 2941
rect 43990 2932 43996 2984
rect 44048 2972 44054 2984
rect 44545 2975 44603 2981
rect 44545 2972 44557 2975
rect 44048 2944 44557 2972
rect 44048 2932 44054 2944
rect 44545 2941 44557 2944
rect 44591 2941 44603 2975
rect 44545 2935 44603 2941
rect 44652 2904 44680 3012
rect 44818 3000 44824 3012
rect 44876 3000 44882 3052
rect 46382 3000 46388 3052
rect 46440 3000 46446 3052
rect 46474 3000 46480 3052
rect 46532 3000 46538 3052
rect 46750 3000 46756 3052
rect 46808 3000 46814 3052
rect 46937 3043 46995 3049
rect 46937 3009 46949 3043
rect 46983 3040 46995 3043
rect 47044 3040 47072 3136
rect 48038 3068 48044 3120
rect 48096 3108 48102 3120
rect 48332 3108 48360 3148
rect 51046 3136 51080 3148
rect 51132 3136 51138 3188
rect 52546 3136 52552 3188
rect 52604 3136 52610 3188
rect 52822 3136 52828 3188
rect 52880 3136 52886 3188
rect 54386 3136 54392 3188
rect 54444 3136 54450 3188
rect 54570 3136 54576 3188
rect 54628 3136 54634 3188
rect 55766 3136 55772 3188
rect 55824 3176 55830 3188
rect 56137 3179 56195 3185
rect 56137 3176 56149 3179
rect 55824 3148 56149 3176
rect 55824 3136 55830 3148
rect 56137 3145 56149 3148
rect 56183 3145 56195 3179
rect 56137 3139 56195 3145
rect 56318 3136 56324 3188
rect 56376 3176 56382 3188
rect 57422 3176 57428 3188
rect 56376 3148 57428 3176
rect 56376 3136 56382 3148
rect 57422 3136 57428 3148
rect 57480 3136 57486 3188
rect 57606 3136 57612 3188
rect 57664 3136 57670 3188
rect 57974 3136 57980 3188
rect 58032 3176 58038 3188
rect 58529 3179 58587 3185
rect 58529 3176 58541 3179
rect 58032 3148 58541 3176
rect 58032 3136 58038 3148
rect 58529 3145 58541 3148
rect 58575 3145 58587 3179
rect 58529 3139 58587 3145
rect 50154 3108 50160 3120
rect 48096 3080 48360 3108
rect 48096 3068 48102 3080
rect 46983 3012 47072 3040
rect 46983 3009 46995 3012
rect 46937 3003 46995 3009
rect 47118 3000 47124 3052
rect 47176 3000 47182 3052
rect 48332 3049 48360 3080
rect 48516 3080 50160 3108
rect 48516 3049 48544 3080
rect 50154 3068 50160 3080
rect 50212 3068 50218 3120
rect 47397 3043 47455 3049
rect 47397 3009 47409 3043
rect 47443 3040 47455 3043
rect 48317 3043 48375 3049
rect 47443 3012 47716 3040
rect 47443 3009 47455 3012
rect 47397 3003 47455 3009
rect 45094 2932 45100 2984
rect 45152 2972 45158 2984
rect 45557 2975 45615 2981
rect 45557 2972 45569 2975
rect 45152 2944 45569 2972
rect 45152 2932 45158 2944
rect 45557 2941 45569 2944
rect 45603 2941 45615 2975
rect 45557 2935 45615 2941
rect 46842 2932 46848 2984
rect 46900 2972 46906 2984
rect 47581 2975 47639 2981
rect 47581 2972 47593 2975
rect 46900 2944 47593 2972
rect 46900 2932 46906 2944
rect 47581 2941 47593 2944
rect 47627 2941 47639 2975
rect 47581 2935 47639 2941
rect 40144 2876 44680 2904
rect 44726 2864 44732 2916
rect 44784 2904 44790 2916
rect 47688 2904 47716 3012
rect 48317 3009 48329 3043
rect 48363 3009 48375 3043
rect 48317 3003 48375 3009
rect 48501 3043 48559 3049
rect 48501 3009 48513 3043
rect 48547 3009 48559 3043
rect 48961 3043 49019 3049
rect 48961 3040 48973 3043
rect 48501 3003 48559 3009
rect 48608 3012 48973 3040
rect 47854 2932 47860 2984
rect 47912 2972 47918 2984
rect 48608 2972 48636 3012
rect 48961 3009 48973 3012
rect 49007 3009 49019 3043
rect 48961 3003 49019 3009
rect 49053 3043 49111 3049
rect 49053 3009 49065 3043
rect 49099 3009 49111 3043
rect 49053 3003 49111 3009
rect 47912 2944 48636 2972
rect 48685 2975 48743 2981
rect 47912 2932 47918 2944
rect 48685 2941 48697 2975
rect 48731 2972 48743 2975
rect 49068 2972 49096 3003
rect 48731 2944 49096 2972
rect 48731 2941 48743 2944
rect 48685 2935 48743 2941
rect 49234 2932 49240 2984
rect 49292 2972 49298 2984
rect 49513 2975 49571 2981
rect 49513 2972 49525 2975
rect 49292 2944 49525 2972
rect 49292 2932 49298 2944
rect 49513 2941 49525 2944
rect 49559 2941 49571 2975
rect 49513 2935 49571 2941
rect 50062 2932 50068 2984
rect 50120 2972 50126 2984
rect 50525 2975 50583 2981
rect 50525 2972 50537 2975
rect 50120 2944 50537 2972
rect 50120 2932 50126 2944
rect 50525 2941 50537 2944
rect 50571 2941 50583 2975
rect 51046 2972 51074 3136
rect 51629 3043 51687 3049
rect 51629 3009 51641 3043
rect 51675 3040 51687 3043
rect 52454 3040 52460 3052
rect 51675 3012 52460 3040
rect 51675 3009 51687 3012
rect 51629 3003 51687 3009
rect 52454 3000 52460 3012
rect 52512 3000 52518 3052
rect 51445 2975 51503 2981
rect 51445 2972 51457 2975
rect 51046 2944 51457 2972
rect 50525 2935 50583 2941
rect 51445 2941 51457 2944
rect 51491 2941 51503 2975
rect 51445 2935 51503 2941
rect 48777 2907 48835 2913
rect 48777 2904 48789 2907
rect 44784 2876 47716 2904
rect 48286 2876 48789 2904
rect 44784 2864 44790 2876
rect 37752 2808 39988 2836
rect 41138 2796 41144 2848
rect 41196 2836 41202 2848
rect 41874 2836 41880 2848
rect 41196 2808 41880 2836
rect 41196 2796 41202 2808
rect 41874 2796 41880 2808
rect 41932 2796 41938 2848
rect 41966 2796 41972 2848
rect 42024 2836 42030 2848
rect 47213 2839 47271 2845
rect 47213 2836 47225 2839
rect 42024 2808 47225 2836
rect 42024 2796 42030 2808
rect 47213 2805 47225 2808
rect 47259 2805 47271 2839
rect 47213 2799 47271 2805
rect 47670 2796 47676 2848
rect 47728 2836 47734 2848
rect 48286 2836 48314 2876
rect 48777 2873 48789 2876
rect 48823 2873 48835 2907
rect 51460 2904 51488 2935
rect 51902 2932 51908 2984
rect 51960 2932 51966 2984
rect 52564 2972 52592 3136
rect 52840 3049 52868 3136
rect 54404 3108 54432 3136
rect 53760 3080 54432 3108
rect 52825 3043 52883 3049
rect 52825 3009 52837 3043
rect 52871 3009 52883 3043
rect 52825 3003 52883 3009
rect 53650 3000 53656 3052
rect 53708 3000 53714 3052
rect 53760 3049 53788 3080
rect 53745 3043 53803 3049
rect 53745 3009 53757 3043
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 53929 3043 53987 3049
rect 53929 3009 53941 3043
rect 53975 3040 53987 3043
rect 54021 3043 54079 3049
rect 54021 3040 54033 3043
rect 53975 3012 54033 3040
rect 53975 3009 53987 3012
rect 53929 3003 53987 3009
rect 54021 3009 54033 3012
rect 54067 3009 54079 3043
rect 54588 3040 54616 3136
rect 55493 3043 55551 3049
rect 55493 3040 55505 3043
rect 54588 3012 55505 3040
rect 54021 3003 54079 3009
rect 55493 3009 55505 3012
rect 55539 3009 55551 3043
rect 55493 3003 55551 3009
rect 56505 3043 56563 3049
rect 56505 3009 56517 3043
rect 56551 3040 56563 3043
rect 57624 3040 57652 3136
rect 56551 3012 57652 3040
rect 56551 3009 56563 3012
rect 56505 3003 56563 3009
rect 53377 2975 53435 2981
rect 53377 2972 53389 2975
rect 52564 2944 53389 2972
rect 53377 2941 53389 2944
rect 53423 2941 53435 2975
rect 53377 2935 53435 2941
rect 53668 2904 53696 3000
rect 54202 2932 54208 2984
rect 54260 2972 54266 2984
rect 54481 2975 54539 2981
rect 54481 2972 54493 2975
rect 54260 2944 54493 2972
rect 54260 2932 54266 2944
rect 54481 2941 54493 2944
rect 54527 2941 54539 2975
rect 54481 2935 54539 2941
rect 57238 2932 57244 2984
rect 57296 2932 57302 2984
rect 57885 2975 57943 2981
rect 57885 2941 57897 2975
rect 57931 2941 57943 2975
rect 57885 2935 57943 2941
rect 51460 2876 53696 2904
rect 48777 2867 48835 2873
rect 55030 2864 55036 2916
rect 55088 2904 55094 2916
rect 57900 2904 57928 2935
rect 55088 2876 57928 2904
rect 55088 2864 55094 2876
rect 47728 2808 48314 2836
rect 47728 2796 47734 2808
rect 51166 2796 51172 2848
rect 51224 2796 51230 2848
rect 51813 2839 51871 2845
rect 51813 2805 51825 2839
rect 51859 2836 51871 2839
rect 52454 2836 52460 2848
rect 51859 2808 52460 2836
rect 51859 2805 51871 2808
rect 51813 2799 51871 2805
rect 52454 2796 52460 2808
rect 52512 2796 52518 2848
rect 52549 2839 52607 2845
rect 52549 2805 52561 2839
rect 52595 2836 52607 2839
rect 55398 2836 55404 2848
rect 52595 2808 55404 2836
rect 52595 2805 52607 2808
rect 52549 2799 52607 2805
rect 55398 2796 55404 2808
rect 55456 2796 55462 2848
rect 1104 2746 58880 2768
rect 1104 2694 8172 2746
rect 8224 2694 8236 2746
rect 8288 2694 8300 2746
rect 8352 2694 8364 2746
rect 8416 2694 8428 2746
rect 8480 2694 22616 2746
rect 22668 2694 22680 2746
rect 22732 2694 22744 2746
rect 22796 2694 22808 2746
rect 22860 2694 22872 2746
rect 22924 2694 37060 2746
rect 37112 2694 37124 2746
rect 37176 2694 37188 2746
rect 37240 2694 37252 2746
rect 37304 2694 37316 2746
rect 37368 2694 51504 2746
rect 51556 2694 51568 2746
rect 51620 2694 51632 2746
rect 51684 2694 51696 2746
rect 51748 2694 51760 2746
rect 51812 2694 58880 2746
rect 1104 2672 58880 2694
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 4157 2635 4215 2641
rect 4157 2632 4169 2635
rect 3660 2604 4169 2632
rect 3660 2592 3666 2604
rect 4157 2601 4169 2604
rect 4203 2601 4215 2635
rect 4157 2595 4215 2601
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2682 2564 2688 2576
rect 1995 2536 2688 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2682 2524 2688 2536
rect 2740 2564 2746 2576
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 2740 2536 3801 2564
rect 2740 2524 2746 2536
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 4172 2564 4200 2595
rect 4338 2592 4344 2644
rect 4396 2592 4402 2644
rect 4982 2592 4988 2644
rect 5040 2592 5046 2644
rect 6362 2592 6368 2644
rect 6420 2592 6426 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 9030 2632 9036 2644
rect 7331 2604 9036 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 11146 2632 11152 2644
rect 9815 2604 11152 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 13909 2635 13967 2641
rect 13909 2601 13921 2635
rect 13955 2632 13967 2635
rect 14734 2632 14740 2644
rect 13955 2604 14740 2632
rect 13955 2601 13967 2604
rect 13909 2595 13967 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 15013 2635 15071 2641
rect 15013 2601 15025 2635
rect 15059 2632 15071 2635
rect 16390 2632 16396 2644
rect 15059 2604 16396 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 16850 2592 16856 2644
rect 16908 2632 16914 2644
rect 17497 2635 17555 2641
rect 17497 2632 17509 2635
rect 16908 2604 17509 2632
rect 16908 2592 16914 2604
rect 17497 2601 17509 2604
rect 17543 2601 17555 2635
rect 17497 2595 17555 2601
rect 20162 2592 20168 2644
rect 20220 2592 20226 2644
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22465 2635 22523 2641
rect 22465 2632 22477 2635
rect 22152 2604 22477 2632
rect 22152 2592 22158 2604
rect 22465 2601 22477 2604
rect 22511 2601 22523 2635
rect 22465 2595 22523 2601
rect 24026 2592 24032 2644
rect 24084 2592 24090 2644
rect 24394 2592 24400 2644
rect 24452 2592 24458 2644
rect 25317 2635 25375 2641
rect 25317 2601 25329 2635
rect 25363 2632 25375 2635
rect 25590 2632 25596 2644
rect 25363 2604 25596 2632
rect 25363 2601 25375 2604
rect 25317 2595 25375 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 27062 2592 27068 2644
rect 27120 2592 27126 2644
rect 27430 2592 27436 2644
rect 27488 2592 27494 2644
rect 28994 2592 29000 2644
rect 29052 2632 29058 2644
rect 29089 2635 29147 2641
rect 29089 2632 29101 2635
rect 29052 2604 29101 2632
rect 29052 2592 29058 2604
rect 29089 2601 29101 2604
rect 29135 2601 29147 2635
rect 29089 2595 29147 2601
rect 31570 2592 31576 2644
rect 31628 2632 31634 2644
rect 32217 2635 32275 2641
rect 32217 2632 32229 2635
rect 31628 2604 32229 2632
rect 31628 2592 31634 2604
rect 32217 2601 32229 2604
rect 32263 2601 32275 2635
rect 32217 2595 32275 2601
rect 34425 2635 34483 2641
rect 34425 2601 34437 2635
rect 34471 2632 34483 2635
rect 34790 2632 34796 2644
rect 34471 2604 34796 2632
rect 34471 2601 34483 2604
rect 34425 2595 34483 2601
rect 34790 2592 34796 2604
rect 34848 2592 34854 2644
rect 34974 2592 34980 2644
rect 35032 2632 35038 2644
rect 36909 2635 36967 2641
rect 36909 2632 36921 2635
rect 35032 2604 36921 2632
rect 35032 2592 35038 2604
rect 36909 2601 36921 2604
rect 36955 2601 36967 2635
rect 36909 2595 36967 2601
rect 38654 2592 38660 2644
rect 38712 2632 38718 2644
rect 39393 2635 39451 2641
rect 39393 2632 39405 2635
rect 38712 2604 39405 2632
rect 38712 2592 38718 2604
rect 39393 2601 39405 2604
rect 39439 2601 39451 2635
rect 39393 2595 39451 2601
rect 39482 2592 39488 2644
rect 39540 2592 39546 2644
rect 41506 2592 41512 2644
rect 41564 2632 41570 2644
rect 42061 2635 42119 2641
rect 42061 2632 42073 2635
rect 41564 2604 42073 2632
rect 41564 2592 41570 2604
rect 42061 2601 42073 2604
rect 42107 2601 42119 2635
rect 42061 2595 42119 2601
rect 44174 2592 44180 2644
rect 44232 2632 44238 2644
rect 44637 2635 44695 2641
rect 44637 2632 44649 2635
rect 44232 2604 44649 2632
rect 44232 2592 44238 2604
rect 44637 2601 44649 2604
rect 44683 2601 44695 2635
rect 44637 2595 44695 2601
rect 45554 2592 45560 2644
rect 45612 2632 45618 2644
rect 45649 2635 45707 2641
rect 45649 2632 45661 2635
rect 45612 2604 45661 2632
rect 45612 2592 45618 2604
rect 45649 2601 45661 2604
rect 45695 2601 45707 2635
rect 45649 2595 45707 2601
rect 47213 2635 47271 2641
rect 47213 2601 47225 2635
rect 47259 2632 47271 2635
rect 47394 2632 47400 2644
rect 47259 2604 47400 2632
rect 47259 2601 47271 2604
rect 47213 2595 47271 2601
rect 47394 2592 47400 2604
rect 47452 2592 47458 2644
rect 49694 2592 49700 2644
rect 49752 2632 49758 2644
rect 49789 2635 49847 2641
rect 49789 2632 49801 2635
rect 49752 2604 49801 2632
rect 49752 2592 49758 2604
rect 49789 2601 49801 2604
rect 49835 2601 49847 2635
rect 49789 2595 49847 2601
rect 50246 2592 50252 2644
rect 50304 2592 50310 2644
rect 52457 2635 52515 2641
rect 52457 2601 52469 2635
rect 52503 2632 52515 2635
rect 52730 2632 52736 2644
rect 52503 2604 52736 2632
rect 52503 2601 52515 2604
rect 52457 2595 52515 2601
rect 52730 2592 52736 2604
rect 52788 2592 52794 2644
rect 53282 2592 53288 2644
rect 53340 2592 53346 2644
rect 54481 2635 54539 2641
rect 54481 2601 54493 2635
rect 54527 2632 54539 2635
rect 55306 2632 55312 2644
rect 54527 2604 55312 2632
rect 54527 2601 54539 2604
rect 54481 2595 54539 2601
rect 55306 2592 55312 2604
rect 55364 2592 55370 2644
rect 56410 2592 56416 2644
rect 56468 2592 56474 2644
rect 58526 2592 58532 2644
rect 58584 2592 58590 2644
rect 4522 2564 4528 2576
rect 4172 2536 4528 2564
rect 3789 2527 3847 2533
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 2038 2456 2044 2508
rect 2096 2496 2102 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2096 2468 2789 2496
rect 2096 2456 2102 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 5000 2496 5028 2592
rect 14093 2567 14151 2573
rect 14093 2533 14105 2567
rect 14139 2564 14151 2567
rect 15746 2564 15752 2576
rect 14139 2536 15752 2564
rect 14139 2533 14151 2536
rect 14093 2527 14151 2533
rect 15746 2524 15752 2536
rect 15804 2524 15810 2576
rect 19245 2567 19303 2573
rect 19245 2533 19257 2567
rect 19291 2564 19303 2567
rect 22278 2564 22284 2576
rect 19291 2536 22284 2564
rect 19291 2533 19303 2536
rect 19245 2527 19303 2533
rect 22278 2524 22284 2536
rect 22336 2524 22342 2576
rect 35986 2564 35992 2576
rect 27172 2536 31800 2564
rect 2777 2459 2835 2465
rect 3528 2468 5028 2496
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 3528 2428 3556 2468
rect 5534 2456 5540 2508
rect 5592 2456 5598 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6779 2468 7512 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 2363 2400 3556 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5902 2428 5908 2440
rect 5031 2400 5908 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6595 2400 6914 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 1670 2320 1676 2372
rect 1728 2320 1734 2372
rect 4154 2320 4160 2372
rect 4212 2320 4218 2372
rect 5258 2360 5264 2372
rect 4540 2332 5264 2360
rect 4540 2301 4568 2332
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 6886 2360 6914 2400
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7248 2400 7389 2428
rect 7248 2388 7254 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7484 2428 7512 2468
rect 7558 2456 7564 2508
rect 7616 2496 7622 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7616 2468 7849 2496
rect 7616 2456 7622 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 10008 2468 10333 2496
rect 10008 2456 10014 2468
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11664 2468 12204 2496
rect 11664 2456 11670 2468
rect 8754 2428 8760 2440
rect 7484 2400 8760 2428
rect 7377 2391 7435 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 8386 2360 8392 2372
rect 6886 2332 8392 2360
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 9232 2360 9260 2391
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9824 2400 9873 2428
rect 9824 2388 9830 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11790 2388 11796 2440
rect 11848 2388 11854 2440
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 12023 2400 12081 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12176 2428 12204 2468
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12400 2468 12541 2496
rect 12400 2456 12406 2468
rect 12529 2465 12541 2468
rect 12575 2465 12587 2499
rect 12529 2459 12587 2465
rect 15838 2456 15844 2508
rect 15896 2456 15902 2508
rect 17862 2456 17868 2508
rect 17920 2496 17926 2508
rect 18049 2499 18107 2505
rect 18049 2496 18061 2499
rect 17920 2468 18061 2496
rect 17920 2456 17926 2468
rect 18049 2465 18061 2468
rect 18095 2465 18107 2499
rect 18049 2459 18107 2465
rect 19352 2468 20300 2496
rect 19352 2440 19380 2468
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 12176 2400 13553 2428
rect 12069 2391 12127 2397
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 13998 2428 14004 2440
rect 13771 2400 14004 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14507 2400 15056 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 11146 2360 11152 2372
rect 9232 2332 11152 2360
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 14292 2360 14320 2391
rect 14734 2360 14740 2372
rect 14292 2332 14740 2360
rect 14734 2320 14740 2332
rect 14792 2320 14798 2372
rect 15028 2360 15056 2400
rect 15194 2388 15200 2440
rect 15252 2388 15258 2440
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 18230 2428 18236 2440
rect 17819 2400 18236 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 16574 2360 16580 2372
rect 15028 2332 16580 2360
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 16960 2360 16988 2391
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 19334 2388 19340 2440
rect 19392 2388 19398 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 20070 2428 20076 2440
rect 19659 2400 20076 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20272 2437 20300 2468
rect 20806 2456 20812 2508
rect 20864 2456 20870 2508
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 25866 2456 25872 2508
rect 25924 2456 25930 2508
rect 27172 2505 27200 2536
rect 31772 2508 31800 2536
rect 32416 2536 35992 2564
rect 27157 2499 27215 2505
rect 27157 2465 27169 2499
rect 27203 2465 27215 2499
rect 27157 2459 27215 2465
rect 27430 2456 27436 2508
rect 27488 2496 27494 2508
rect 27985 2499 28043 2505
rect 27985 2496 27997 2499
rect 27488 2468 27997 2496
rect 27488 2456 27494 2468
rect 27985 2465 27997 2468
rect 28031 2465 28043 2499
rect 30469 2499 30527 2505
rect 30469 2496 30481 2499
rect 27985 2459 28043 2465
rect 29288 2468 30481 2496
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 21910 2388 21916 2440
rect 21968 2388 21974 2440
rect 22186 2388 22192 2440
rect 22244 2428 22250 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22244 2400 22569 2428
rect 22244 2388 22250 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 23382 2388 23388 2440
rect 23440 2428 23446 2440
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 23440 2400 24225 2428
rect 23440 2388 23446 2400
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 24765 2431 24823 2437
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 25222 2428 25228 2440
rect 24811 2400 25228 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25314 2388 25320 2440
rect 25372 2428 25378 2440
rect 25409 2431 25467 2437
rect 25409 2428 25421 2431
rect 25372 2400 25421 2428
rect 25372 2388 25378 2400
rect 25409 2397 25421 2400
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 27249 2431 27307 2437
rect 27249 2397 27261 2431
rect 27295 2428 27307 2431
rect 27522 2428 27528 2440
rect 27295 2400 27528 2428
rect 27295 2397 27307 2400
rect 27249 2391 27307 2397
rect 27522 2388 27528 2400
rect 27580 2388 27586 2440
rect 27706 2388 27712 2440
rect 27764 2388 27770 2440
rect 29288 2437 29316 2468
rect 30469 2465 30481 2468
rect 30515 2465 30527 2499
rect 30469 2459 30527 2465
rect 30742 2456 30748 2508
rect 30800 2496 30806 2508
rect 31021 2499 31079 2505
rect 31021 2496 31033 2499
rect 30800 2468 31033 2496
rect 30800 2456 30806 2468
rect 31021 2465 31033 2468
rect 31067 2465 31079 2499
rect 31021 2459 31079 2465
rect 31754 2456 31760 2508
rect 31812 2456 31818 2508
rect 29273 2431 29331 2437
rect 29273 2397 29285 2431
rect 29319 2397 29331 2431
rect 29273 2391 29331 2397
rect 29730 2388 29736 2440
rect 29788 2388 29794 2440
rect 29917 2431 29975 2437
rect 29917 2397 29929 2431
rect 29963 2428 29975 2431
rect 30190 2428 30196 2440
rect 29963 2400 30196 2428
rect 29963 2397 29975 2400
rect 29917 2391 29975 2397
rect 30190 2388 30196 2400
rect 30248 2388 30254 2440
rect 30650 2388 30656 2440
rect 30708 2388 30714 2440
rect 32416 2437 32444 2536
rect 35986 2524 35992 2536
rect 36044 2524 36050 2576
rect 53300 2564 53328 2592
rect 54941 2567 54999 2573
rect 54941 2564 54953 2567
rect 53300 2536 54953 2564
rect 54941 2533 54953 2536
rect 54987 2533 54999 2567
rect 54941 2527 54999 2533
rect 32674 2456 32680 2508
rect 32732 2496 32738 2508
rect 32953 2499 33011 2505
rect 32953 2496 32965 2499
rect 32732 2468 32965 2496
rect 32732 2456 32738 2468
rect 32953 2465 32965 2468
rect 32999 2465 33011 2499
rect 35618 2496 35624 2508
rect 32953 2459 33011 2465
rect 34900 2468 35624 2496
rect 32401 2431 32459 2437
rect 32401 2397 32413 2431
rect 32447 2397 32459 2431
rect 32401 2391 32459 2397
rect 32585 2431 32643 2437
rect 32585 2397 32597 2431
rect 32631 2397 32643 2431
rect 32585 2391 32643 2397
rect 18598 2360 18604 2372
rect 16960 2332 18604 2360
rect 18598 2320 18604 2332
rect 18656 2320 18662 2372
rect 26973 2363 27031 2369
rect 26973 2329 26985 2363
rect 27019 2360 27031 2363
rect 27019 2332 29592 2360
rect 27019 2329 27031 2332
rect 26973 2323 27031 2329
rect 29564 2301 29592 2332
rect 4525 2295 4583 2301
rect 4525 2261 4537 2295
rect 4571 2261 4583 2295
rect 4525 2255 4583 2261
rect 29549 2295 29607 2301
rect 29549 2261 29561 2295
rect 29595 2261 29607 2295
rect 32600 2292 32628 2391
rect 34146 2388 34152 2440
rect 34204 2388 34210 2440
rect 34900 2437 34928 2468
rect 35618 2456 35624 2468
rect 35676 2456 35682 2508
rect 35710 2456 35716 2508
rect 35768 2496 35774 2508
rect 37737 2499 37795 2505
rect 37737 2496 37749 2499
rect 35768 2468 37749 2496
rect 35768 2456 35774 2468
rect 37737 2465 37749 2468
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 38746 2456 38752 2508
rect 38804 2456 38810 2508
rect 39022 2456 39028 2508
rect 39080 2496 39086 2508
rect 40313 2499 40371 2505
rect 40313 2496 40325 2499
rect 39080 2468 40325 2496
rect 39080 2456 39086 2468
rect 40313 2465 40325 2468
rect 40359 2465 40371 2499
rect 40313 2459 40371 2465
rect 42610 2456 42616 2508
rect 42668 2496 42674 2508
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 42668 2468 42901 2496
rect 42668 2456 42674 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 44082 2456 44088 2508
rect 44140 2456 44146 2508
rect 45646 2456 45652 2508
rect 45704 2496 45710 2508
rect 46201 2499 46259 2505
rect 46201 2496 46213 2499
rect 45704 2468 46213 2496
rect 45704 2456 45710 2468
rect 46201 2465 46213 2468
rect 46247 2465 46259 2499
rect 46201 2459 46259 2465
rect 47486 2456 47492 2508
rect 47544 2496 47550 2508
rect 48041 2499 48099 2505
rect 48041 2496 48053 2499
rect 47544 2468 48053 2496
rect 47544 2456 47550 2468
rect 48041 2465 48053 2468
rect 48087 2465 48099 2499
rect 48041 2459 48099 2465
rect 50614 2456 50620 2508
rect 50672 2496 50678 2508
rect 51261 2499 51319 2505
rect 51261 2496 51273 2499
rect 50672 2468 51273 2496
rect 50672 2456 50678 2468
rect 51261 2465 51273 2468
rect 51307 2465 51319 2499
rect 51261 2459 51319 2465
rect 52362 2456 52368 2508
rect 52420 2496 52426 2508
rect 53193 2499 53251 2505
rect 53193 2496 53205 2499
rect 52420 2468 53205 2496
rect 52420 2456 52426 2468
rect 53193 2465 53205 2468
rect 53239 2465 53251 2499
rect 53193 2459 53251 2465
rect 55582 2456 55588 2508
rect 55640 2496 55646 2508
rect 56137 2499 56195 2505
rect 56137 2496 56149 2499
rect 55640 2468 56149 2496
rect 55640 2456 55646 2468
rect 56137 2465 56149 2468
rect 56183 2465 56195 2499
rect 56428 2496 56456 2592
rect 56428 2468 57376 2496
rect 56137 2459 56195 2465
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 36170 2388 36176 2440
rect 36228 2388 36234 2440
rect 37093 2431 37151 2437
rect 37093 2397 37105 2431
rect 37139 2397 37151 2431
rect 37093 2391 37151 2397
rect 37277 2431 37335 2437
rect 37277 2397 37289 2431
rect 37323 2428 37335 2431
rect 37550 2428 37556 2440
rect 37323 2400 37556 2428
rect 37323 2397 37335 2400
rect 37277 2391 37335 2397
rect 34422 2320 34428 2372
rect 34480 2360 34486 2372
rect 35621 2363 35679 2369
rect 35621 2360 35633 2363
rect 34480 2332 35633 2360
rect 34480 2320 34486 2332
rect 35621 2329 35633 2332
rect 35667 2329 35679 2363
rect 37108 2360 37136 2391
rect 37550 2388 37556 2400
rect 37608 2388 37614 2440
rect 39669 2431 39727 2437
rect 39669 2397 39681 2431
rect 39715 2397 39727 2431
rect 39669 2391 39727 2397
rect 39945 2431 40003 2437
rect 39945 2397 39957 2431
rect 39991 2428 40003 2431
rect 40034 2428 40040 2440
rect 39991 2400 40040 2428
rect 39991 2397 40003 2400
rect 39945 2391 40003 2397
rect 35621 2323 35679 2329
rect 35728 2332 37136 2360
rect 34054 2292 34060 2304
rect 32600 2264 34060 2292
rect 29549 2255 29607 2261
rect 34054 2252 34060 2264
rect 34112 2252 34118 2304
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35728 2292 35756 2332
rect 38010 2320 38016 2372
rect 38068 2360 38074 2372
rect 39684 2360 39712 2391
rect 40034 2388 40040 2400
rect 40092 2388 40098 2440
rect 40126 2388 40132 2440
rect 40184 2428 40190 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 40184 2400 41337 2428
rect 40184 2388 40190 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 41969 2431 42027 2437
rect 41969 2397 41981 2431
rect 42015 2428 42027 2431
rect 42245 2431 42303 2437
rect 42245 2428 42257 2431
rect 42015 2400 42257 2428
rect 42015 2397 42027 2400
rect 41969 2391 42027 2397
rect 42245 2397 42257 2400
rect 42291 2397 42303 2431
rect 42245 2391 42303 2397
rect 42521 2431 42579 2437
rect 42521 2397 42533 2431
rect 42567 2428 42579 2431
rect 43254 2428 43260 2440
rect 42567 2400 43260 2428
rect 42567 2397 42579 2400
rect 42521 2391 42579 2397
rect 43254 2388 43260 2400
rect 43312 2388 43318 2440
rect 45005 2431 45063 2437
rect 45005 2397 45017 2431
rect 45051 2397 45063 2431
rect 45005 2391 45063 2397
rect 45925 2431 45983 2437
rect 45925 2397 45937 2431
rect 45971 2428 45983 2431
rect 47118 2428 47124 2440
rect 45971 2400 47124 2428
rect 45971 2397 45983 2400
rect 45925 2391 45983 2397
rect 38068 2332 39712 2360
rect 38068 2320 38074 2332
rect 43898 2320 43904 2372
rect 43956 2360 43962 2372
rect 45020 2360 45048 2391
rect 47118 2388 47124 2400
rect 47176 2388 47182 2440
rect 47397 2431 47455 2437
rect 47397 2397 47409 2431
rect 47443 2397 47455 2431
rect 47397 2391 47455 2397
rect 47765 2431 47823 2437
rect 47765 2397 47777 2431
rect 47811 2428 47823 2431
rect 48314 2428 48320 2440
rect 47811 2400 48320 2428
rect 47811 2397 47823 2400
rect 47765 2391 47823 2397
rect 43956 2332 45048 2360
rect 43956 2320 43962 2332
rect 46198 2320 46204 2372
rect 46256 2360 46262 2372
rect 47412 2360 47440 2391
rect 48314 2388 48320 2400
rect 48372 2388 48378 2440
rect 48406 2388 48412 2440
rect 48464 2428 48470 2440
rect 49053 2431 49111 2437
rect 49053 2428 49065 2431
rect 48464 2400 49065 2428
rect 48464 2388 48470 2400
rect 49053 2397 49065 2400
rect 49099 2397 49111 2431
rect 49053 2391 49111 2397
rect 49694 2388 49700 2440
rect 49752 2428 49758 2440
rect 49973 2431 50031 2437
rect 49973 2428 49985 2431
rect 49752 2400 49985 2428
rect 49752 2388 49758 2400
rect 49973 2397 49985 2400
rect 50019 2397 50031 2431
rect 49973 2391 50031 2397
rect 50433 2431 50491 2437
rect 50433 2397 50445 2431
rect 50479 2397 50491 2431
rect 50433 2391 50491 2397
rect 50893 2431 50951 2437
rect 50893 2397 50905 2431
rect 50939 2428 50951 2431
rect 51074 2428 51080 2440
rect 50939 2400 51080 2428
rect 50939 2397 50951 2400
rect 50893 2391 50951 2397
rect 50448 2360 50476 2391
rect 51074 2388 51080 2400
rect 51132 2388 51138 2440
rect 51166 2388 51172 2440
rect 51224 2428 51230 2440
rect 52273 2431 52331 2437
rect 52273 2428 52285 2431
rect 51224 2400 52285 2428
rect 51224 2388 51230 2400
rect 52273 2397 52285 2400
rect 52319 2397 52331 2431
rect 52273 2391 52331 2397
rect 52454 2388 52460 2440
rect 52512 2428 52518 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52512 2400 52745 2428
rect 52512 2388 52518 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 54757 2431 54815 2437
rect 54757 2397 54769 2431
rect 54803 2428 54815 2431
rect 54938 2428 54944 2440
rect 54803 2400 54944 2428
rect 54803 2397 54815 2400
rect 54757 2391 54815 2397
rect 54938 2388 54944 2400
rect 54996 2388 55002 2440
rect 55398 2388 55404 2440
rect 55456 2388 55462 2440
rect 55861 2431 55919 2437
rect 55861 2397 55873 2431
rect 55907 2397 55919 2431
rect 55861 2391 55919 2397
rect 46256 2332 47440 2360
rect 49712 2332 50476 2360
rect 55876 2360 55904 2391
rect 57146 2388 57152 2440
rect 57204 2388 57210 2440
rect 57348 2437 57376 2468
rect 57882 2456 57888 2508
rect 57940 2456 57946 2508
rect 57333 2431 57391 2437
rect 57333 2397 57345 2431
rect 57379 2397 57391 2431
rect 57333 2391 57391 2397
rect 57517 2363 57575 2369
rect 57517 2360 57529 2363
rect 55876 2332 57529 2360
rect 46256 2320 46262 2332
rect 34848 2264 35756 2292
rect 34848 2252 34854 2264
rect 35802 2252 35808 2304
rect 35860 2292 35866 2304
rect 49712 2301 49740 2332
rect 57517 2329 57529 2332
rect 57563 2329 57575 2363
rect 57517 2323 57575 2329
rect 36817 2295 36875 2301
rect 36817 2292 36829 2295
rect 35860 2264 36829 2292
rect 35860 2252 35866 2264
rect 36817 2261 36829 2264
rect 36863 2261 36875 2295
rect 36817 2255 36875 2261
rect 49697 2295 49755 2301
rect 49697 2261 49709 2295
rect 49743 2261 49755 2295
rect 49697 2255 49755 2261
rect 53190 2252 53196 2304
rect 53248 2292 53254 2304
rect 55585 2295 55643 2301
rect 55585 2292 55597 2295
rect 53248 2264 55597 2292
rect 53248 2252 53254 2264
rect 55585 2261 55597 2264
rect 55631 2261 55643 2295
rect 55585 2255 55643 2261
rect 1104 2202 59040 2224
rect 1104 2150 15394 2202
rect 15446 2150 15458 2202
rect 15510 2150 15522 2202
rect 15574 2150 15586 2202
rect 15638 2150 15650 2202
rect 15702 2150 29838 2202
rect 29890 2150 29902 2202
rect 29954 2150 29966 2202
rect 30018 2150 30030 2202
rect 30082 2150 30094 2202
rect 30146 2150 44282 2202
rect 44334 2150 44346 2202
rect 44398 2150 44410 2202
rect 44462 2150 44474 2202
rect 44526 2150 44538 2202
rect 44590 2150 58726 2202
rect 58778 2150 58790 2202
rect 58842 2150 58854 2202
rect 58906 2150 58918 2202
rect 58970 2150 58982 2202
rect 59034 2150 59040 2202
rect 1104 2128 59040 2150
rect 32030 2048 32036 2100
rect 32088 2048 32094 2100
rect 34054 2048 34060 2100
rect 34112 2088 34118 2100
rect 38194 2088 38200 2100
rect 34112 2060 38200 2088
rect 34112 2048 34118 2060
rect 38194 2048 38200 2060
rect 38252 2048 38258 2100
rect 32048 2020 32076 2048
rect 35802 2020 35808 2032
rect 32048 1992 35808 2020
rect 35802 1980 35808 1992
rect 35860 1980 35866 2032
rect 31846 1504 31852 1556
rect 31904 1544 31910 1556
rect 35342 1544 35348 1556
rect 31904 1516 35348 1544
rect 31904 1504 31910 1516
rect 35342 1504 35348 1516
rect 35400 1504 35406 1556
<< via1 >>
rect 8172 27718 8224 27770
rect 8236 27718 8288 27770
rect 8300 27718 8352 27770
rect 8364 27718 8416 27770
rect 8428 27718 8480 27770
rect 22616 27718 22668 27770
rect 22680 27718 22732 27770
rect 22744 27718 22796 27770
rect 22808 27718 22860 27770
rect 22872 27718 22924 27770
rect 37060 27718 37112 27770
rect 37124 27718 37176 27770
rect 37188 27718 37240 27770
rect 37252 27718 37304 27770
rect 37316 27718 37368 27770
rect 51504 27718 51556 27770
rect 51568 27718 51620 27770
rect 51632 27718 51684 27770
rect 51696 27718 51748 27770
rect 51760 27718 51812 27770
rect 15394 27174 15446 27226
rect 15458 27174 15510 27226
rect 15522 27174 15574 27226
rect 15586 27174 15638 27226
rect 15650 27174 15702 27226
rect 29838 27174 29890 27226
rect 29902 27174 29954 27226
rect 29966 27174 30018 27226
rect 30030 27174 30082 27226
rect 30094 27174 30146 27226
rect 44282 27174 44334 27226
rect 44346 27174 44398 27226
rect 44410 27174 44462 27226
rect 44474 27174 44526 27226
rect 44538 27174 44590 27226
rect 58726 27174 58778 27226
rect 58790 27174 58842 27226
rect 58854 27174 58906 27226
rect 58918 27174 58970 27226
rect 58982 27174 59034 27226
rect 8172 26630 8224 26682
rect 8236 26630 8288 26682
rect 8300 26630 8352 26682
rect 8364 26630 8416 26682
rect 8428 26630 8480 26682
rect 22616 26630 22668 26682
rect 22680 26630 22732 26682
rect 22744 26630 22796 26682
rect 22808 26630 22860 26682
rect 22872 26630 22924 26682
rect 37060 26630 37112 26682
rect 37124 26630 37176 26682
rect 37188 26630 37240 26682
rect 37252 26630 37304 26682
rect 37316 26630 37368 26682
rect 51504 26630 51556 26682
rect 51568 26630 51620 26682
rect 51632 26630 51684 26682
rect 51696 26630 51748 26682
rect 51760 26630 51812 26682
rect 15394 26086 15446 26138
rect 15458 26086 15510 26138
rect 15522 26086 15574 26138
rect 15586 26086 15638 26138
rect 15650 26086 15702 26138
rect 29838 26086 29890 26138
rect 29902 26086 29954 26138
rect 29966 26086 30018 26138
rect 30030 26086 30082 26138
rect 30094 26086 30146 26138
rect 44282 26086 44334 26138
rect 44346 26086 44398 26138
rect 44410 26086 44462 26138
rect 44474 26086 44526 26138
rect 44538 26086 44590 26138
rect 58726 26086 58778 26138
rect 58790 26086 58842 26138
rect 58854 26086 58906 26138
rect 58918 26086 58970 26138
rect 58982 26086 59034 26138
rect 8172 25542 8224 25594
rect 8236 25542 8288 25594
rect 8300 25542 8352 25594
rect 8364 25542 8416 25594
rect 8428 25542 8480 25594
rect 22616 25542 22668 25594
rect 22680 25542 22732 25594
rect 22744 25542 22796 25594
rect 22808 25542 22860 25594
rect 22872 25542 22924 25594
rect 37060 25542 37112 25594
rect 37124 25542 37176 25594
rect 37188 25542 37240 25594
rect 37252 25542 37304 25594
rect 37316 25542 37368 25594
rect 51504 25542 51556 25594
rect 51568 25542 51620 25594
rect 51632 25542 51684 25594
rect 51696 25542 51748 25594
rect 51760 25542 51812 25594
rect 15394 24998 15446 25050
rect 15458 24998 15510 25050
rect 15522 24998 15574 25050
rect 15586 24998 15638 25050
rect 15650 24998 15702 25050
rect 29838 24998 29890 25050
rect 29902 24998 29954 25050
rect 29966 24998 30018 25050
rect 30030 24998 30082 25050
rect 30094 24998 30146 25050
rect 44282 24998 44334 25050
rect 44346 24998 44398 25050
rect 44410 24998 44462 25050
rect 44474 24998 44526 25050
rect 44538 24998 44590 25050
rect 58726 24998 58778 25050
rect 58790 24998 58842 25050
rect 58854 24998 58906 25050
rect 58918 24998 58970 25050
rect 58982 24998 59034 25050
rect 8172 24454 8224 24506
rect 8236 24454 8288 24506
rect 8300 24454 8352 24506
rect 8364 24454 8416 24506
rect 8428 24454 8480 24506
rect 22616 24454 22668 24506
rect 22680 24454 22732 24506
rect 22744 24454 22796 24506
rect 22808 24454 22860 24506
rect 22872 24454 22924 24506
rect 37060 24454 37112 24506
rect 37124 24454 37176 24506
rect 37188 24454 37240 24506
rect 37252 24454 37304 24506
rect 37316 24454 37368 24506
rect 51504 24454 51556 24506
rect 51568 24454 51620 24506
rect 51632 24454 51684 24506
rect 51696 24454 51748 24506
rect 51760 24454 51812 24506
rect 15394 23910 15446 23962
rect 15458 23910 15510 23962
rect 15522 23910 15574 23962
rect 15586 23910 15638 23962
rect 15650 23910 15702 23962
rect 29838 23910 29890 23962
rect 29902 23910 29954 23962
rect 29966 23910 30018 23962
rect 30030 23910 30082 23962
rect 30094 23910 30146 23962
rect 44282 23910 44334 23962
rect 44346 23910 44398 23962
rect 44410 23910 44462 23962
rect 44474 23910 44526 23962
rect 44538 23910 44590 23962
rect 58726 23910 58778 23962
rect 58790 23910 58842 23962
rect 58854 23910 58906 23962
rect 58918 23910 58970 23962
rect 58982 23910 59034 23962
rect 8172 23366 8224 23418
rect 8236 23366 8288 23418
rect 8300 23366 8352 23418
rect 8364 23366 8416 23418
rect 8428 23366 8480 23418
rect 22616 23366 22668 23418
rect 22680 23366 22732 23418
rect 22744 23366 22796 23418
rect 22808 23366 22860 23418
rect 22872 23366 22924 23418
rect 37060 23366 37112 23418
rect 37124 23366 37176 23418
rect 37188 23366 37240 23418
rect 37252 23366 37304 23418
rect 37316 23366 37368 23418
rect 51504 23366 51556 23418
rect 51568 23366 51620 23418
rect 51632 23366 51684 23418
rect 51696 23366 51748 23418
rect 51760 23366 51812 23418
rect 38844 23103 38896 23112
rect 38844 23069 38853 23103
rect 38853 23069 38887 23103
rect 38887 23069 38896 23103
rect 38844 23060 38896 23069
rect 47860 23103 47912 23112
rect 47860 23069 47869 23103
rect 47869 23069 47903 23103
rect 47903 23069 47912 23103
rect 47860 23060 47912 23069
rect 39396 22967 39448 22976
rect 39396 22933 39405 22967
rect 39405 22933 39439 22967
rect 39439 22933 39448 22967
rect 39396 22924 39448 22933
rect 40040 22967 40092 22976
rect 40040 22933 40049 22967
rect 40049 22933 40083 22967
rect 40083 22933 40092 22967
rect 40040 22924 40092 22933
rect 48504 22967 48556 22976
rect 48504 22933 48513 22967
rect 48513 22933 48547 22967
rect 48547 22933 48556 22967
rect 48504 22924 48556 22933
rect 15394 22822 15446 22874
rect 15458 22822 15510 22874
rect 15522 22822 15574 22874
rect 15586 22822 15638 22874
rect 15650 22822 15702 22874
rect 29838 22822 29890 22874
rect 29902 22822 29954 22874
rect 29966 22822 30018 22874
rect 30030 22822 30082 22874
rect 30094 22822 30146 22874
rect 44282 22822 44334 22874
rect 44346 22822 44398 22874
rect 44410 22822 44462 22874
rect 44474 22822 44526 22874
rect 44538 22822 44590 22874
rect 58726 22822 58778 22874
rect 58790 22822 58842 22874
rect 58854 22822 58906 22874
rect 58918 22822 58970 22874
rect 58982 22822 59034 22874
rect 48504 22720 48556 22772
rect 40040 22652 40092 22704
rect 47584 22652 47636 22704
rect 38292 22627 38344 22636
rect 38292 22593 38301 22627
rect 38301 22593 38335 22627
rect 38335 22593 38344 22627
rect 38292 22584 38344 22593
rect 39396 22584 39448 22636
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 24308 22423 24360 22432
rect 24308 22389 24317 22423
rect 24317 22389 24351 22423
rect 24351 22389 24360 22423
rect 24308 22380 24360 22389
rect 24676 22423 24728 22432
rect 24676 22389 24685 22423
rect 24685 22389 24719 22423
rect 24719 22389 24728 22423
rect 24676 22380 24728 22389
rect 25412 22423 25464 22432
rect 25412 22389 25421 22423
rect 25421 22389 25455 22423
rect 25455 22389 25464 22423
rect 25412 22380 25464 22389
rect 37924 22380 37976 22432
rect 38568 22380 38620 22432
rect 38660 22380 38712 22432
rect 40408 22423 40460 22432
rect 40408 22389 40417 22423
rect 40417 22389 40451 22423
rect 40451 22389 40460 22423
rect 40408 22380 40460 22389
rect 50712 22559 50764 22568
rect 50712 22525 50721 22559
rect 50721 22525 50755 22559
rect 50755 22525 50764 22559
rect 50712 22516 50764 22525
rect 51356 22559 51408 22568
rect 51356 22525 51365 22559
rect 51365 22525 51399 22559
rect 51399 22525 51408 22559
rect 51356 22516 51408 22525
rect 52920 22559 52972 22568
rect 52920 22525 52929 22559
rect 52929 22525 52963 22559
rect 52963 22525 52972 22559
rect 52920 22516 52972 22525
rect 55312 22516 55364 22568
rect 55956 22516 56008 22568
rect 48504 22380 48556 22432
rect 49700 22423 49752 22432
rect 49700 22389 49709 22423
rect 49709 22389 49743 22423
rect 49743 22389 49752 22423
rect 49700 22380 49752 22389
rect 50804 22380 50856 22432
rect 52000 22423 52052 22432
rect 52000 22389 52009 22423
rect 52009 22389 52043 22423
rect 52043 22389 52052 22423
rect 52000 22380 52052 22389
rect 52368 22423 52420 22432
rect 52368 22389 52377 22423
rect 52377 22389 52411 22423
rect 52411 22389 52420 22423
rect 52368 22380 52420 22389
rect 53564 22423 53616 22432
rect 53564 22389 53573 22423
rect 53573 22389 53607 22423
rect 53607 22389 53616 22423
rect 53564 22380 53616 22389
rect 54852 22380 54904 22432
rect 55772 22380 55824 22432
rect 56692 22423 56744 22432
rect 56692 22389 56701 22423
rect 56701 22389 56735 22423
rect 56735 22389 56744 22423
rect 56692 22380 56744 22389
rect 8172 22278 8224 22330
rect 8236 22278 8288 22330
rect 8300 22278 8352 22330
rect 8364 22278 8416 22330
rect 8428 22278 8480 22330
rect 22616 22278 22668 22330
rect 22680 22278 22732 22330
rect 22744 22278 22796 22330
rect 22808 22278 22860 22330
rect 22872 22278 22924 22330
rect 37060 22278 37112 22330
rect 37124 22278 37176 22330
rect 37188 22278 37240 22330
rect 37252 22278 37304 22330
rect 37316 22278 37368 22330
rect 51504 22278 51556 22330
rect 51568 22278 51620 22330
rect 51632 22278 51684 22330
rect 51696 22278 51748 22330
rect 51760 22278 51812 22330
rect 47860 22176 47912 22228
rect 55312 22219 55364 22228
rect 55312 22185 55321 22219
rect 55321 22185 55355 22219
rect 55355 22185 55364 22219
rect 55312 22176 55364 22185
rect 38568 22108 38620 22160
rect 24308 22040 24360 22092
rect 40776 22108 40828 22160
rect 48228 22108 48280 22160
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 25412 21972 25464 22024
rect 14832 21947 14884 21956
rect 5356 21836 5408 21888
rect 7564 21836 7616 21888
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 14832 21913 14841 21947
rect 14841 21913 14875 21947
rect 14875 21913 14884 21947
rect 14832 21904 14884 21913
rect 11336 21836 11388 21845
rect 23020 21879 23072 21888
rect 23020 21845 23029 21879
rect 23029 21845 23063 21879
rect 23063 21845 23072 21879
rect 23020 21836 23072 21845
rect 24216 21879 24268 21888
rect 24216 21845 24225 21879
rect 24225 21845 24259 21879
rect 24259 21845 24268 21879
rect 24216 21836 24268 21845
rect 24400 21836 24452 21888
rect 38292 21972 38344 22024
rect 49700 22040 49752 22092
rect 55772 22083 55824 22092
rect 55772 22049 55781 22083
rect 55781 22049 55815 22083
rect 55815 22049 55824 22083
rect 55772 22040 55824 22049
rect 55864 22040 55916 22092
rect 48504 21972 48556 22024
rect 52368 21972 52420 22024
rect 52460 21972 52512 22024
rect 56692 22108 56744 22160
rect 26516 21879 26568 21888
rect 26516 21845 26525 21879
rect 26525 21845 26559 21879
rect 26559 21845 26568 21879
rect 26516 21836 26568 21845
rect 38752 21836 38804 21888
rect 50804 21904 50856 21956
rect 39212 21836 39264 21888
rect 39396 21879 39448 21888
rect 39396 21845 39405 21879
rect 39405 21845 39439 21879
rect 39439 21845 39448 21879
rect 39396 21836 39448 21845
rect 47308 21836 47360 21888
rect 51356 21836 51408 21888
rect 52184 21836 52236 21888
rect 52736 21836 52788 21888
rect 58532 21904 58584 21956
rect 54484 21879 54536 21888
rect 54484 21845 54493 21879
rect 54493 21845 54527 21879
rect 54527 21845 54536 21879
rect 54484 21836 54536 21845
rect 54760 21879 54812 21888
rect 54760 21845 54769 21879
rect 54769 21845 54803 21879
rect 54803 21845 54812 21879
rect 54760 21836 54812 21845
rect 57796 21836 57848 21888
rect 57980 21879 58032 21888
rect 57980 21845 57989 21879
rect 57989 21845 58023 21879
rect 58023 21845 58032 21879
rect 57980 21836 58032 21845
rect 15394 21734 15446 21786
rect 15458 21734 15510 21786
rect 15522 21734 15574 21786
rect 15586 21734 15638 21786
rect 15650 21734 15702 21786
rect 29838 21734 29890 21786
rect 29902 21734 29954 21786
rect 29966 21734 30018 21786
rect 30030 21734 30082 21786
rect 30094 21734 30146 21786
rect 44282 21734 44334 21786
rect 44346 21734 44398 21786
rect 44410 21734 44462 21786
rect 44474 21734 44526 21786
rect 44538 21734 44590 21786
rect 58726 21734 58778 21786
rect 58790 21734 58842 21786
rect 58854 21734 58906 21786
rect 58918 21734 58970 21786
rect 58982 21734 59034 21786
rect 4436 21675 4488 21684
rect 4436 21641 4445 21675
rect 4445 21641 4479 21675
rect 4479 21641 4488 21675
rect 4436 21632 4488 21641
rect 5816 21632 5868 21684
rect 9864 21632 9916 21684
rect 10508 21675 10560 21684
rect 10508 21641 10517 21675
rect 10517 21641 10551 21675
rect 10551 21641 10560 21675
rect 10508 21632 10560 21641
rect 24216 21632 24268 21684
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 26516 21632 26568 21684
rect 38844 21675 38896 21684
rect 38844 21641 38853 21675
rect 38853 21641 38887 21675
rect 38887 21641 38896 21675
rect 38844 21632 38896 21641
rect 39396 21632 39448 21684
rect 40408 21632 40460 21684
rect 50712 21675 50764 21684
rect 50712 21641 50721 21675
rect 50721 21641 50755 21675
rect 50755 21641 50764 21675
rect 50712 21632 50764 21641
rect 52000 21632 52052 21684
rect 54484 21632 54536 21684
rect 54760 21632 54812 21684
rect 55956 21632 56008 21684
rect 56508 21632 56560 21684
rect 57980 21632 58032 21684
rect 58532 21675 58584 21684
rect 58532 21641 58541 21675
rect 58541 21641 58575 21675
rect 58575 21641 58584 21675
rect 58532 21632 58584 21641
rect 8760 21496 8812 21548
rect 10416 21496 10468 21548
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 5356 21428 5408 21480
rect 5448 21428 5500 21480
rect 6276 21428 6328 21480
rect 7840 21428 7892 21480
rect 8668 21428 8720 21480
rect 9404 21428 9456 21480
rect 10968 21428 11020 21480
rect 11336 21564 11388 21616
rect 18972 21564 19024 21616
rect 23020 21564 23072 21616
rect 7564 21360 7616 21412
rect 13912 21471 13964 21480
rect 13912 21437 13921 21471
rect 13921 21437 13955 21471
rect 13955 21437 13964 21471
rect 13912 21428 13964 21437
rect 15200 21471 15252 21480
rect 15200 21437 15209 21471
rect 15209 21437 15243 21471
rect 15243 21437 15252 21471
rect 15200 21428 15252 21437
rect 18696 21471 18748 21480
rect 18696 21437 18705 21471
rect 18705 21437 18739 21471
rect 18739 21437 18748 21471
rect 18696 21428 18748 21437
rect 3700 21335 3752 21344
rect 3700 21301 3709 21335
rect 3709 21301 3743 21335
rect 3743 21301 3752 21335
rect 3700 21292 3752 21301
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 7104 21335 7156 21344
rect 7104 21301 7113 21335
rect 7113 21301 7147 21335
rect 7147 21301 7156 21335
rect 7104 21292 7156 21301
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 9680 21292 9732 21344
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 9772 21292 9824 21301
rect 9864 21292 9916 21344
rect 14740 21360 14792 21412
rect 14464 21335 14516 21344
rect 14464 21301 14473 21335
rect 14473 21301 14507 21335
rect 14507 21301 14516 21335
rect 14464 21292 14516 21301
rect 14648 21292 14700 21344
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 19340 21335 19392 21344
rect 19340 21301 19349 21335
rect 19349 21301 19383 21335
rect 19383 21301 19392 21335
rect 19340 21292 19392 21301
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 23020 21335 23072 21344
rect 23020 21301 23029 21335
rect 23029 21301 23063 21335
rect 23063 21301 23072 21335
rect 23020 21292 23072 21301
rect 27896 21564 27948 21616
rect 52368 21564 52420 21616
rect 23940 21471 23992 21480
rect 23940 21437 23949 21471
rect 23949 21437 23983 21471
rect 23983 21437 23992 21471
rect 23940 21428 23992 21437
rect 26792 21496 26844 21548
rect 38752 21496 38804 21548
rect 38936 21496 38988 21548
rect 39212 21539 39264 21548
rect 39212 21505 39221 21539
rect 39221 21505 39255 21539
rect 39255 21505 39264 21539
rect 39212 21496 39264 21505
rect 24860 21428 24912 21480
rect 26056 21471 26108 21480
rect 26056 21437 26065 21471
rect 26065 21437 26099 21471
rect 26099 21437 26108 21471
rect 26056 21428 26108 21437
rect 30196 21471 30248 21480
rect 30196 21437 30205 21471
rect 30205 21437 30239 21471
rect 30239 21437 30248 21471
rect 30196 21428 30248 21437
rect 52092 21496 52144 21548
rect 52460 21496 52512 21548
rect 53564 21496 53616 21548
rect 54852 21564 54904 21616
rect 56048 21539 56100 21548
rect 56048 21505 56057 21539
rect 56057 21505 56091 21539
rect 56091 21505 56100 21539
rect 56048 21496 56100 21505
rect 56876 21496 56928 21548
rect 39304 21428 39356 21480
rect 30012 21360 30064 21412
rect 35348 21360 35400 21412
rect 39028 21360 39080 21412
rect 42708 21471 42760 21480
rect 42708 21437 42717 21471
rect 42717 21437 42751 21471
rect 42751 21437 42760 21471
rect 42708 21428 42760 21437
rect 46664 21471 46716 21480
rect 46664 21437 46673 21471
rect 46673 21437 46707 21471
rect 46707 21437 46716 21471
rect 46664 21428 46716 21437
rect 51356 21471 51408 21480
rect 51356 21437 51365 21471
rect 51365 21437 51399 21471
rect 51399 21437 51408 21471
rect 51356 21428 51408 21437
rect 52276 21471 52328 21480
rect 42248 21403 42300 21412
rect 42248 21369 42257 21403
rect 42257 21369 42291 21403
rect 42291 21369 42300 21403
rect 52276 21437 52285 21471
rect 52285 21437 52319 21471
rect 52319 21437 52328 21471
rect 52276 21428 52328 21437
rect 42248 21360 42300 21369
rect 24032 21292 24084 21344
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 25780 21335 25832 21344
rect 25780 21301 25789 21335
rect 25789 21301 25823 21335
rect 25823 21301 25832 21335
rect 25780 21292 25832 21301
rect 26608 21335 26660 21344
rect 26608 21301 26617 21335
rect 26617 21301 26651 21335
rect 26651 21301 26660 21335
rect 26608 21292 26660 21301
rect 30840 21335 30892 21344
rect 30840 21301 30849 21335
rect 30849 21301 30883 21335
rect 30883 21301 30892 21335
rect 30840 21292 30892 21301
rect 38384 21335 38436 21344
rect 38384 21301 38393 21335
rect 38393 21301 38427 21335
rect 38427 21301 38436 21335
rect 38384 21292 38436 21301
rect 39212 21292 39264 21344
rect 41880 21335 41932 21344
rect 41880 21301 41889 21335
rect 41889 21301 41923 21335
rect 41923 21301 41932 21335
rect 41880 21292 41932 21301
rect 43260 21335 43312 21344
rect 43260 21301 43269 21335
rect 43269 21301 43303 21335
rect 43303 21301 43312 21335
rect 43260 21292 43312 21301
rect 43904 21292 43956 21344
rect 46112 21292 46164 21344
rect 46480 21335 46532 21344
rect 46480 21301 46489 21335
rect 46489 21301 46523 21335
rect 46523 21301 46532 21335
rect 46480 21292 46532 21301
rect 47216 21335 47268 21344
rect 47216 21301 47225 21335
rect 47225 21301 47259 21335
rect 47259 21301 47268 21335
rect 47216 21292 47268 21301
rect 47860 21335 47912 21344
rect 47860 21301 47869 21335
rect 47869 21301 47903 21335
rect 47903 21301 47912 21335
rect 47860 21292 47912 21301
rect 48228 21292 48280 21344
rect 51264 21292 51316 21344
rect 52644 21292 52696 21344
rect 53748 21292 53800 21344
rect 56508 21292 56560 21344
rect 57520 21335 57572 21344
rect 57520 21301 57529 21335
rect 57529 21301 57563 21335
rect 57563 21301 57572 21335
rect 57520 21292 57572 21301
rect 8172 21190 8224 21242
rect 8236 21190 8288 21242
rect 8300 21190 8352 21242
rect 8364 21190 8416 21242
rect 8428 21190 8480 21242
rect 22616 21190 22668 21242
rect 22680 21190 22732 21242
rect 22744 21190 22796 21242
rect 22808 21190 22860 21242
rect 22872 21190 22924 21242
rect 37060 21190 37112 21242
rect 37124 21190 37176 21242
rect 37188 21190 37240 21242
rect 37252 21190 37304 21242
rect 37316 21190 37368 21242
rect 51504 21190 51556 21242
rect 51568 21190 51620 21242
rect 51632 21190 51684 21242
rect 51696 21190 51748 21242
rect 51760 21190 51812 21242
rect 4436 21088 4488 21140
rect 6184 21088 6236 21140
rect 6276 21131 6328 21140
rect 6276 21097 6285 21131
rect 6285 21097 6319 21131
rect 6319 21097 6328 21131
rect 6276 21088 6328 21097
rect 7104 21088 7156 21140
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 5356 20884 5408 20936
rect 2872 20748 2924 20800
rect 3240 20791 3292 20800
rect 3240 20757 3249 20791
rect 3249 20757 3283 20791
rect 3283 20757 3292 20791
rect 3240 20748 3292 20757
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 4160 20748 4212 20800
rect 4528 20791 4580 20800
rect 4528 20757 4537 20791
rect 4537 20757 4571 20791
rect 4571 20757 4580 20791
rect 4528 20748 4580 20757
rect 7564 21088 7616 21140
rect 8760 21131 8812 21140
rect 8760 21097 8769 21131
rect 8769 21097 8803 21131
rect 8803 21097 8812 21131
rect 8760 21088 8812 21097
rect 8944 21088 8996 21140
rect 9772 21088 9824 21140
rect 9864 21088 9916 21140
rect 14464 21088 14516 21140
rect 14832 21088 14884 21140
rect 15200 21088 15252 21140
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 9680 20884 9732 20936
rect 7840 20816 7892 20868
rect 8668 20816 8720 20868
rect 5448 20748 5500 20800
rect 6644 20791 6696 20800
rect 6644 20757 6653 20791
rect 6653 20757 6687 20791
rect 6687 20757 6696 20791
rect 6644 20748 6696 20757
rect 11060 20816 11112 20868
rect 16488 20884 16540 20936
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 22192 20952 22244 21004
rect 24308 21088 24360 21140
rect 23664 21020 23716 21072
rect 25320 21088 25372 21140
rect 25780 21088 25832 21140
rect 26056 21088 26108 21140
rect 30012 21131 30064 21140
rect 30012 21097 30021 21131
rect 30021 21097 30055 21131
rect 30055 21097 30064 21131
rect 30012 21088 30064 21097
rect 30196 21131 30248 21140
rect 30196 21097 30205 21131
rect 30205 21097 30239 21131
rect 30239 21097 30248 21131
rect 30196 21088 30248 21097
rect 24400 20995 24452 21004
rect 24400 20961 24409 20995
rect 24409 20961 24443 20995
rect 24443 20961 24452 20995
rect 24400 20952 24452 20961
rect 24952 20952 25004 21004
rect 26700 20952 26752 21004
rect 26792 20995 26844 21004
rect 26792 20961 26801 20995
rect 26801 20961 26835 20995
rect 26835 20961 26844 20995
rect 26792 20952 26844 20961
rect 38384 21088 38436 21140
rect 39488 21088 39540 21140
rect 39948 21088 40000 21140
rect 41420 21131 41472 21140
rect 41420 21097 41429 21131
rect 41429 21097 41463 21131
rect 41463 21097 41472 21131
rect 41420 21088 41472 21097
rect 42248 21088 42300 21140
rect 46664 21088 46716 21140
rect 31668 21020 31720 21072
rect 43904 21063 43956 21072
rect 43904 21029 43913 21063
rect 43913 21029 43947 21063
rect 43947 21029 43956 21063
rect 43904 21020 43956 21029
rect 46112 21020 46164 21072
rect 51080 21020 51132 21072
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 19892 20927 19944 20936
rect 19892 20893 19901 20927
rect 19901 20893 19935 20927
rect 19935 20893 19944 20927
rect 19892 20884 19944 20893
rect 20628 20927 20680 20936
rect 20628 20893 20637 20927
rect 20637 20893 20671 20927
rect 20671 20893 20680 20927
rect 20628 20884 20680 20893
rect 23020 20884 23072 20936
rect 23940 20884 23992 20936
rect 24308 20816 24360 20868
rect 9404 20748 9456 20800
rect 9864 20748 9916 20800
rect 10968 20748 11020 20800
rect 13728 20791 13780 20800
rect 13728 20757 13737 20791
rect 13737 20757 13771 20791
rect 13771 20757 13780 20791
rect 13728 20748 13780 20757
rect 13820 20748 13872 20800
rect 14924 20748 14976 20800
rect 16580 20791 16632 20800
rect 16580 20757 16589 20791
rect 16589 20757 16623 20791
rect 16623 20757 16632 20791
rect 16580 20748 16632 20757
rect 18788 20791 18840 20800
rect 18788 20757 18797 20791
rect 18797 20757 18831 20791
rect 18831 20757 18840 20791
rect 18788 20748 18840 20757
rect 18972 20748 19024 20800
rect 19800 20748 19852 20800
rect 20444 20748 20496 20800
rect 20536 20791 20588 20800
rect 20536 20757 20545 20791
rect 20545 20757 20579 20791
rect 20579 20757 20588 20791
rect 20536 20748 20588 20757
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 25320 20927 25372 20936
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25320 20884 25372 20893
rect 25412 20927 25464 20936
rect 25412 20893 25446 20927
rect 25446 20893 25464 20927
rect 25412 20884 25464 20893
rect 25596 20927 25648 20936
rect 25596 20893 25605 20927
rect 25605 20893 25639 20927
rect 25639 20893 25648 20927
rect 25596 20884 25648 20893
rect 46480 20952 46532 21004
rect 51356 20952 51408 21004
rect 27988 20927 28040 20936
rect 27988 20893 27997 20927
rect 27997 20893 28031 20927
rect 28031 20893 28040 20927
rect 27988 20884 28040 20893
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 31024 20927 31076 20936
rect 31024 20893 31033 20927
rect 31033 20893 31067 20927
rect 31067 20893 31076 20927
rect 31024 20884 31076 20893
rect 32864 20927 32916 20936
rect 32864 20893 32873 20927
rect 32873 20893 32907 20927
rect 32907 20893 32916 20927
rect 32864 20884 32916 20893
rect 33692 20927 33744 20936
rect 33692 20893 33701 20927
rect 33701 20893 33735 20927
rect 33735 20893 33744 20927
rect 33692 20884 33744 20893
rect 35348 20884 35400 20936
rect 35900 20884 35952 20936
rect 37556 20927 37608 20936
rect 37556 20893 37565 20927
rect 37565 20893 37599 20927
rect 37599 20893 37608 20927
rect 37556 20884 37608 20893
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 41788 20927 41840 20936
rect 41788 20893 41797 20927
rect 41797 20893 41831 20927
rect 41831 20893 41840 20927
rect 41788 20884 41840 20893
rect 41880 20884 41932 20936
rect 44732 20884 44784 20936
rect 45008 20927 45060 20936
rect 45008 20893 45017 20927
rect 45017 20893 45051 20927
rect 45051 20893 45060 20927
rect 45008 20884 45060 20893
rect 47676 20927 47728 20936
rect 47676 20893 47685 20927
rect 47685 20893 47719 20927
rect 47719 20893 47728 20927
rect 47676 20884 47728 20893
rect 49516 20884 49568 20936
rect 51264 20884 51316 20936
rect 54760 21088 54812 21140
rect 53748 21020 53800 21072
rect 52000 20952 52052 21004
rect 52184 20952 52236 21004
rect 52644 20995 52696 21004
rect 52644 20961 52653 20995
rect 52653 20961 52687 20995
rect 52687 20961 52696 20995
rect 52644 20952 52696 20961
rect 45376 20816 45428 20868
rect 47308 20816 47360 20868
rect 48688 20816 48740 20868
rect 25412 20748 25464 20800
rect 26148 20748 26200 20800
rect 28540 20791 28592 20800
rect 28540 20757 28549 20791
rect 28549 20757 28583 20791
rect 28583 20757 28592 20791
rect 28540 20748 28592 20757
rect 28908 20748 28960 20800
rect 30564 20791 30616 20800
rect 30564 20757 30573 20791
rect 30573 20757 30607 20791
rect 30607 20757 30616 20791
rect 30564 20748 30616 20757
rect 33416 20791 33468 20800
rect 33416 20757 33425 20791
rect 33425 20757 33459 20791
rect 33459 20757 33468 20791
rect 33416 20748 33468 20757
rect 34244 20791 34296 20800
rect 34244 20757 34253 20791
rect 34253 20757 34287 20791
rect 34287 20757 34296 20791
rect 34244 20748 34296 20757
rect 35808 20748 35860 20800
rect 36728 20791 36780 20800
rect 36728 20757 36737 20791
rect 36737 20757 36771 20791
rect 36771 20757 36780 20791
rect 36728 20748 36780 20757
rect 37464 20748 37516 20800
rect 38108 20791 38160 20800
rect 38108 20757 38117 20791
rect 38117 20757 38151 20791
rect 38151 20757 38160 20791
rect 38108 20748 38160 20757
rect 38844 20791 38896 20800
rect 38844 20757 38853 20791
rect 38853 20757 38887 20791
rect 38887 20757 38896 20791
rect 38844 20748 38896 20757
rect 39212 20791 39264 20800
rect 39212 20757 39221 20791
rect 39221 20757 39255 20791
rect 39255 20757 39264 20791
rect 39212 20748 39264 20757
rect 42340 20791 42392 20800
rect 42340 20757 42349 20791
rect 42349 20757 42383 20791
rect 42383 20757 42392 20791
rect 42340 20748 42392 20757
rect 44640 20791 44692 20800
rect 44640 20757 44649 20791
rect 44649 20757 44683 20791
rect 44683 20757 44692 20791
rect 44640 20748 44692 20757
rect 45652 20791 45704 20800
rect 45652 20757 45661 20791
rect 45661 20757 45695 20791
rect 45695 20757 45704 20791
rect 45652 20748 45704 20757
rect 48780 20748 48832 20800
rect 49700 20791 49752 20800
rect 49700 20757 49709 20791
rect 49709 20757 49743 20791
rect 49743 20757 49752 20791
rect 49700 20748 49752 20757
rect 50160 20748 50212 20800
rect 51080 20791 51132 20800
rect 51080 20757 51089 20791
rect 51089 20757 51123 20791
rect 51123 20757 51132 20791
rect 51080 20748 51132 20757
rect 52460 20927 52512 20936
rect 52460 20893 52494 20927
rect 52494 20893 52512 20927
rect 52460 20884 52512 20893
rect 53564 20884 53616 20936
rect 55588 20952 55640 21004
rect 57520 21088 57572 21140
rect 56048 20952 56100 21004
rect 56232 20952 56284 21004
rect 56416 20952 56468 21004
rect 56876 20995 56928 21004
rect 56876 20961 56885 20995
rect 56885 20961 56919 20995
rect 56919 20961 56928 20995
rect 56876 20952 56928 20961
rect 58164 20995 58216 21004
rect 58164 20961 58173 20995
rect 58173 20961 58207 20995
rect 58207 20961 58216 20995
rect 58164 20952 58216 20961
rect 53196 20816 53248 20868
rect 52736 20748 52788 20800
rect 53288 20791 53340 20800
rect 53288 20757 53297 20791
rect 53297 20757 53331 20791
rect 53331 20757 53340 20791
rect 53288 20748 53340 20757
rect 55036 20816 55088 20868
rect 55772 20748 55824 20800
rect 56600 20927 56652 20936
rect 56600 20893 56609 20927
rect 56609 20893 56643 20927
rect 56643 20893 56652 20927
rect 56600 20884 56652 20893
rect 57796 20816 57848 20868
rect 56968 20748 57020 20800
rect 57520 20791 57572 20800
rect 57520 20757 57529 20791
rect 57529 20757 57563 20791
rect 57563 20757 57572 20791
rect 57520 20748 57572 20757
rect 57612 20791 57664 20800
rect 57612 20757 57621 20791
rect 57621 20757 57655 20791
rect 57655 20757 57664 20791
rect 57612 20748 57664 20757
rect 57704 20748 57756 20800
rect 15394 20646 15446 20698
rect 15458 20646 15510 20698
rect 15522 20646 15574 20698
rect 15586 20646 15638 20698
rect 15650 20646 15702 20698
rect 29838 20646 29890 20698
rect 29902 20646 29954 20698
rect 29966 20646 30018 20698
rect 30030 20646 30082 20698
rect 30094 20646 30146 20698
rect 44282 20646 44334 20698
rect 44346 20646 44398 20698
rect 44410 20646 44462 20698
rect 44474 20646 44526 20698
rect 44538 20646 44590 20698
rect 58726 20646 58778 20698
rect 58790 20646 58842 20698
rect 58854 20646 58906 20698
rect 58918 20646 58970 20698
rect 58982 20646 59034 20698
rect 4068 20544 4120 20596
rect 4436 20544 4488 20596
rect 6644 20544 6696 20596
rect 7564 20587 7616 20596
rect 7564 20553 7573 20587
rect 7573 20553 7607 20587
rect 7607 20553 7616 20587
rect 7564 20544 7616 20553
rect 13912 20544 13964 20596
rect 2780 20476 2832 20528
rect 3700 20408 3752 20460
rect 3976 20408 4028 20460
rect 4160 20340 4212 20392
rect 4988 20451 5040 20460
rect 4988 20417 4997 20451
rect 4997 20417 5031 20451
rect 5031 20417 5040 20451
rect 4988 20408 5040 20417
rect 6736 20451 6788 20460
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 13728 20476 13780 20528
rect 19340 20544 19392 20596
rect 15844 20476 15896 20528
rect 8760 20408 8812 20460
rect 9864 20408 9916 20460
rect 10416 20451 10468 20460
rect 10416 20417 10425 20451
rect 10425 20417 10459 20451
rect 10459 20417 10468 20451
rect 10416 20408 10468 20417
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 14648 20408 14700 20460
rect 15108 20408 15160 20460
rect 19156 20408 19208 20460
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 7288 20340 7340 20392
rect 9680 20383 9732 20392
rect 9680 20349 9689 20383
rect 9689 20349 9723 20383
rect 9723 20349 9732 20383
rect 9680 20340 9732 20349
rect 4436 20272 4488 20324
rect 6644 20272 6696 20324
rect 9864 20272 9916 20324
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 6368 20247 6420 20256
rect 6368 20213 6377 20247
rect 6377 20213 6411 20247
rect 6411 20213 6420 20247
rect 6368 20204 6420 20213
rect 9036 20247 9088 20256
rect 9036 20213 9045 20247
rect 9045 20213 9079 20247
rect 9079 20213 9088 20247
rect 9036 20204 9088 20213
rect 11520 20340 11572 20392
rect 11520 20204 11572 20256
rect 13820 20340 13872 20392
rect 15016 20383 15068 20392
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 18972 20340 19024 20392
rect 19524 20544 19576 20596
rect 20444 20544 20496 20596
rect 22192 20587 22244 20596
rect 22192 20553 22201 20587
rect 22201 20553 22235 20587
rect 22235 20553 22244 20587
rect 22192 20544 22244 20553
rect 23940 20544 23992 20596
rect 24584 20544 24636 20596
rect 26700 20587 26752 20596
rect 26700 20553 26709 20587
rect 26709 20553 26743 20587
rect 26743 20553 26752 20587
rect 26700 20544 26752 20553
rect 27896 20587 27948 20596
rect 27896 20553 27905 20587
rect 27905 20553 27939 20587
rect 27939 20553 27948 20587
rect 27896 20544 27948 20553
rect 27988 20544 28040 20596
rect 28908 20544 28960 20596
rect 19616 20476 19668 20528
rect 20536 20408 20588 20460
rect 23848 20408 23900 20460
rect 26608 20408 26660 20460
rect 18144 20272 18196 20324
rect 12072 20204 12124 20256
rect 14280 20204 14332 20256
rect 16672 20204 16724 20256
rect 16856 20247 16908 20256
rect 16856 20213 16865 20247
rect 16865 20213 16899 20247
rect 16899 20213 16908 20247
rect 16856 20204 16908 20213
rect 17960 20247 18012 20256
rect 17960 20213 17969 20247
rect 17969 20213 18003 20247
rect 18003 20213 18012 20247
rect 17960 20204 18012 20213
rect 24032 20340 24084 20392
rect 30564 20544 30616 20596
rect 30748 20544 30800 20596
rect 31668 20544 31720 20596
rect 32864 20544 32916 20596
rect 34244 20544 34296 20596
rect 37556 20587 37608 20596
rect 37556 20553 37565 20587
rect 37565 20553 37599 20587
rect 37599 20553 37608 20587
rect 37556 20544 37608 20553
rect 38844 20544 38896 20596
rect 40776 20587 40828 20596
rect 40776 20553 40785 20587
rect 40785 20553 40819 20587
rect 40819 20553 40828 20587
rect 40776 20544 40828 20553
rect 41788 20544 41840 20596
rect 43260 20544 43312 20596
rect 29460 20476 29512 20528
rect 30840 20476 30892 20528
rect 30564 20408 30616 20460
rect 24860 20315 24912 20324
rect 24860 20281 24869 20315
rect 24869 20281 24903 20315
rect 24903 20281 24912 20315
rect 24860 20272 24912 20281
rect 29736 20340 29788 20392
rect 34152 20476 34204 20528
rect 37832 20476 37884 20528
rect 33968 20408 34020 20460
rect 33784 20383 33836 20392
rect 33784 20349 33793 20383
rect 33793 20349 33827 20383
rect 33827 20349 33836 20383
rect 33784 20340 33836 20349
rect 19340 20204 19392 20256
rect 20628 20204 20680 20256
rect 21180 20204 21232 20256
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 23756 20247 23808 20256
rect 23756 20213 23765 20247
rect 23765 20213 23799 20247
rect 23799 20213 23808 20247
rect 23756 20204 23808 20213
rect 24216 20204 24268 20256
rect 25320 20204 25372 20256
rect 34336 20272 34388 20324
rect 35992 20383 36044 20392
rect 35992 20349 36001 20383
rect 36001 20349 36035 20383
rect 36035 20349 36044 20383
rect 35992 20340 36044 20349
rect 37464 20340 37516 20392
rect 39304 20451 39356 20460
rect 39304 20417 39313 20451
rect 39313 20417 39347 20451
rect 39347 20417 39356 20451
rect 39304 20408 39356 20417
rect 39580 20451 39632 20460
rect 39580 20417 39589 20451
rect 39589 20417 39623 20451
rect 39623 20417 39632 20451
rect 39580 20408 39632 20417
rect 27344 20204 27396 20256
rect 28632 20204 28684 20256
rect 29552 20247 29604 20256
rect 29552 20213 29561 20247
rect 29561 20213 29595 20247
rect 29595 20213 29604 20247
rect 29552 20204 29604 20213
rect 30104 20204 30156 20256
rect 31024 20204 31076 20256
rect 31852 20247 31904 20256
rect 31852 20213 31861 20247
rect 31861 20213 31895 20247
rect 31895 20213 31904 20247
rect 31852 20204 31904 20213
rect 33324 20204 33376 20256
rect 35900 20247 35952 20256
rect 35900 20213 35909 20247
rect 35909 20213 35943 20247
rect 35943 20213 35952 20247
rect 35900 20204 35952 20213
rect 36912 20247 36964 20256
rect 36912 20213 36921 20247
rect 36921 20213 36955 20247
rect 36955 20213 36964 20247
rect 36912 20204 36964 20213
rect 38200 20340 38252 20392
rect 38292 20340 38344 20392
rect 38568 20383 38620 20392
rect 38568 20349 38577 20383
rect 38577 20349 38611 20383
rect 38611 20349 38620 20383
rect 38568 20340 38620 20349
rect 38660 20340 38712 20392
rect 39948 20340 40000 20392
rect 41420 20476 41472 20528
rect 42064 20476 42116 20528
rect 42340 20408 42392 20460
rect 43168 20408 43220 20460
rect 43904 20476 43956 20528
rect 45652 20476 45704 20528
rect 43076 20383 43128 20392
rect 43076 20349 43085 20383
rect 43085 20349 43119 20383
rect 43119 20349 43128 20383
rect 43076 20340 43128 20349
rect 44916 20383 44968 20392
rect 44916 20349 44925 20383
rect 44925 20349 44959 20383
rect 44959 20349 44968 20383
rect 44916 20340 44968 20349
rect 45468 20340 45520 20392
rect 48228 20544 48280 20596
rect 49516 20587 49568 20596
rect 49516 20553 49525 20587
rect 49525 20553 49559 20587
rect 49559 20553 49568 20587
rect 49516 20544 49568 20553
rect 52920 20544 52972 20596
rect 57704 20587 57756 20596
rect 57704 20553 57713 20587
rect 57713 20553 57747 20587
rect 57747 20553 57756 20587
rect 57704 20544 57756 20553
rect 58164 20544 58216 20596
rect 47216 20476 47268 20528
rect 46112 20408 46164 20460
rect 47584 20451 47636 20460
rect 47584 20417 47593 20451
rect 47593 20417 47627 20451
rect 47627 20417 47636 20451
rect 47584 20408 47636 20417
rect 47676 20408 47728 20460
rect 39028 20315 39080 20324
rect 39028 20281 39037 20315
rect 39037 20281 39071 20315
rect 39071 20281 39080 20315
rect 39028 20272 39080 20281
rect 38844 20204 38896 20256
rect 40224 20247 40276 20256
rect 40224 20213 40233 20247
rect 40233 20213 40267 20247
rect 40267 20213 40276 20247
rect 40224 20204 40276 20213
rect 40776 20204 40828 20256
rect 56416 20408 56468 20460
rect 42708 20204 42760 20256
rect 43628 20204 43680 20256
rect 44732 20247 44784 20256
rect 44732 20213 44741 20247
rect 44741 20213 44775 20247
rect 44775 20213 44784 20247
rect 44732 20204 44784 20213
rect 45100 20204 45152 20256
rect 48596 20383 48648 20392
rect 48596 20349 48630 20383
rect 48630 20349 48648 20383
rect 48596 20340 48648 20349
rect 48780 20383 48832 20392
rect 48780 20349 48789 20383
rect 48789 20349 48823 20383
rect 48823 20349 48832 20383
rect 48780 20340 48832 20349
rect 49976 20383 50028 20392
rect 49976 20349 49985 20383
rect 49985 20349 50019 20383
rect 50019 20349 50028 20383
rect 49976 20340 50028 20349
rect 50160 20383 50212 20392
rect 50160 20349 50169 20383
rect 50169 20349 50203 20383
rect 50203 20349 50212 20383
rect 50160 20340 50212 20349
rect 47860 20272 47912 20324
rect 48320 20272 48372 20324
rect 50436 20383 50488 20392
rect 50436 20349 50445 20383
rect 50445 20349 50479 20383
rect 50479 20349 50488 20383
rect 50436 20340 50488 20349
rect 51264 20340 51316 20392
rect 53196 20383 53248 20392
rect 53196 20349 53205 20383
rect 53205 20349 53239 20383
rect 53239 20349 53248 20383
rect 53196 20340 53248 20349
rect 53748 20383 53800 20392
rect 53748 20349 53757 20383
rect 53757 20349 53791 20383
rect 53791 20349 53800 20383
rect 53748 20340 53800 20349
rect 54852 20340 54904 20392
rect 55220 20383 55272 20392
rect 55220 20349 55229 20383
rect 55229 20349 55263 20383
rect 55263 20349 55272 20383
rect 55220 20340 55272 20349
rect 55588 20383 55640 20392
rect 55588 20349 55597 20383
rect 55597 20349 55631 20383
rect 55631 20349 55640 20383
rect 55588 20340 55640 20349
rect 56968 20408 57020 20460
rect 57612 20408 57664 20460
rect 49332 20204 49384 20256
rect 50068 20204 50120 20256
rect 52000 20247 52052 20256
rect 52000 20213 52009 20247
rect 52009 20213 52043 20247
rect 52043 20213 52052 20247
rect 52000 20204 52052 20213
rect 54668 20247 54720 20256
rect 54668 20213 54677 20247
rect 54677 20213 54711 20247
rect 54711 20213 54720 20247
rect 54668 20204 54720 20213
rect 8172 20102 8224 20154
rect 8236 20102 8288 20154
rect 8300 20102 8352 20154
rect 8364 20102 8416 20154
rect 8428 20102 8480 20154
rect 22616 20102 22668 20154
rect 22680 20102 22732 20154
rect 22744 20102 22796 20154
rect 22808 20102 22860 20154
rect 22872 20102 22924 20154
rect 37060 20102 37112 20154
rect 37124 20102 37176 20154
rect 37188 20102 37240 20154
rect 37252 20102 37304 20154
rect 37316 20102 37368 20154
rect 51504 20102 51556 20154
rect 51568 20102 51620 20154
rect 51632 20102 51684 20154
rect 51696 20102 51748 20154
rect 51760 20102 51812 20154
rect 3148 20000 3200 20052
rect 4988 20000 5040 20052
rect 6368 20000 6420 20052
rect 6644 20043 6696 20052
rect 6644 20009 6653 20043
rect 6653 20009 6687 20043
rect 6687 20009 6696 20043
rect 6644 20000 6696 20009
rect 7564 20000 7616 20052
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 9036 20000 9088 20052
rect 9680 20000 9732 20052
rect 12348 20000 12400 20052
rect 3516 19932 3568 19984
rect 2780 19796 2832 19848
rect 4528 19796 4580 19848
rect 5356 19796 5408 19848
rect 2872 19728 2924 19780
rect 4712 19728 4764 19780
rect 6092 19796 6144 19848
rect 9680 19864 9732 19916
rect 12072 19864 12124 19916
rect 13820 20000 13872 20052
rect 14924 20000 14976 20052
rect 14096 19932 14148 19984
rect 14280 19907 14332 19916
rect 14280 19873 14289 19907
rect 14289 19873 14323 19907
rect 14323 19873 14332 19907
rect 14280 19864 14332 19873
rect 11336 19728 11388 19780
rect 13636 19728 13688 19780
rect 4344 19660 4396 19712
rect 4988 19660 5040 19712
rect 5264 19660 5316 19712
rect 8760 19660 8812 19712
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 13820 19660 13872 19712
rect 18696 20000 18748 20052
rect 20168 20000 20220 20052
rect 18604 19932 18656 19984
rect 16856 19907 16908 19916
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15476 19839 15528 19848
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 16580 19839 16632 19848
rect 16580 19805 16589 19839
rect 16589 19805 16623 19839
rect 16623 19805 16632 19839
rect 16580 19796 16632 19805
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 19800 19864 19852 19916
rect 20444 19907 20496 19916
rect 20444 19873 20453 19907
rect 20453 19873 20487 19907
rect 20487 19873 20496 19907
rect 20444 19864 20496 19873
rect 19340 19796 19392 19848
rect 16488 19728 16540 19780
rect 17960 19728 18012 19780
rect 16120 19703 16172 19712
rect 16120 19669 16129 19703
rect 16129 19669 16163 19703
rect 16163 19669 16172 19703
rect 16120 19660 16172 19669
rect 16212 19703 16264 19712
rect 16212 19669 16221 19703
rect 16221 19669 16255 19703
rect 16255 19669 16264 19703
rect 16212 19660 16264 19669
rect 19616 19796 19668 19848
rect 20168 19839 20220 19848
rect 20168 19805 20177 19839
rect 20177 19805 20211 19839
rect 20211 19805 20220 19839
rect 20168 19796 20220 19805
rect 21180 19796 21232 19848
rect 21640 20000 21692 20052
rect 23756 20000 23808 20052
rect 23848 20043 23900 20052
rect 23848 20009 23857 20043
rect 23857 20009 23891 20043
rect 23891 20009 23900 20043
rect 23848 20000 23900 20009
rect 28816 20043 28868 20052
rect 28816 20009 28825 20043
rect 28825 20009 28859 20043
rect 28859 20009 28868 20043
rect 28816 20000 28868 20009
rect 21640 19864 21692 19916
rect 25780 19796 25832 19848
rect 27344 19839 27396 19848
rect 27344 19805 27353 19839
rect 27353 19805 27387 19839
rect 27387 19805 27396 19839
rect 27344 19796 27396 19805
rect 29736 19932 29788 19984
rect 30104 19864 30156 19916
rect 30196 19907 30248 19916
rect 30196 19873 30205 19907
rect 30205 19873 30239 19907
rect 30239 19873 30248 19907
rect 30196 19864 30248 19873
rect 31852 20000 31904 20052
rect 33324 20000 33376 20052
rect 33784 20000 33836 20052
rect 30564 19907 30616 19916
rect 30564 19873 30598 19907
rect 30598 19873 30616 19907
rect 30564 19864 30616 19873
rect 30748 19907 30800 19916
rect 30748 19873 30757 19907
rect 30757 19873 30791 19907
rect 30791 19873 30800 19907
rect 30748 19864 30800 19873
rect 30932 19864 30984 19916
rect 28540 19796 28592 19848
rect 33600 19932 33652 19984
rect 34152 19907 34204 19916
rect 34152 19873 34161 19907
rect 34161 19873 34195 19907
rect 34195 19873 34204 19907
rect 34152 19864 34204 19873
rect 21088 19703 21140 19712
rect 21088 19669 21097 19703
rect 21097 19669 21131 19703
rect 21131 19669 21140 19703
rect 21088 19660 21140 19669
rect 21640 19703 21692 19712
rect 21640 19669 21649 19703
rect 21649 19669 21683 19703
rect 21683 19669 21692 19703
rect 21640 19660 21692 19669
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 24216 19703 24268 19712
rect 24216 19669 24225 19703
rect 24225 19669 24259 19703
rect 24259 19669 24268 19703
rect 24216 19660 24268 19669
rect 29000 19660 29052 19712
rect 34336 19728 34388 19780
rect 31208 19660 31260 19712
rect 33876 19703 33928 19712
rect 33876 19669 33885 19703
rect 33885 19669 33919 19703
rect 33919 19669 33928 19703
rect 33876 19660 33928 19669
rect 33968 19703 34020 19712
rect 33968 19669 33977 19703
rect 33977 19669 34011 19703
rect 34011 19669 34020 19703
rect 33968 19660 34020 19669
rect 34428 19660 34480 19712
rect 34704 19839 34756 19848
rect 34704 19805 34713 19839
rect 34713 19805 34747 19839
rect 34747 19805 34756 19839
rect 34704 19796 34756 19805
rect 35900 20000 35952 20052
rect 38292 20000 38344 20052
rect 40040 20000 40092 20052
rect 35348 19907 35400 19916
rect 35348 19873 35357 19907
rect 35357 19873 35391 19907
rect 35391 19873 35400 19907
rect 35348 19864 35400 19873
rect 38200 19864 38252 19916
rect 39028 19864 39080 19916
rect 35624 19839 35676 19848
rect 35624 19805 35633 19839
rect 35633 19805 35667 19839
rect 35667 19805 35676 19839
rect 35624 19796 35676 19805
rect 35900 19839 35952 19848
rect 35900 19805 35909 19839
rect 35909 19805 35943 19839
rect 35943 19805 35952 19839
rect 35900 19796 35952 19805
rect 36912 19796 36964 19848
rect 42616 19864 42668 19916
rect 44732 20000 44784 20052
rect 44916 20000 44968 20052
rect 43260 19864 43312 19916
rect 44088 19864 44140 19916
rect 44640 19864 44692 19916
rect 45468 19864 45520 19916
rect 46940 19864 46992 19916
rect 48504 20000 48556 20052
rect 49700 20000 49752 20052
rect 52000 20000 52052 20052
rect 54668 20000 54720 20052
rect 55036 20043 55088 20052
rect 55036 20009 55045 20043
rect 55045 20009 55079 20043
rect 55079 20009 55088 20043
rect 55036 20000 55088 20009
rect 57060 20000 57112 20052
rect 36544 19703 36596 19712
rect 36544 19669 36553 19703
rect 36553 19669 36587 19703
rect 36587 19669 36596 19703
rect 36544 19660 36596 19669
rect 38108 19728 38160 19780
rect 39948 19728 40000 19780
rect 41052 19728 41104 19780
rect 37464 19660 37516 19712
rect 38844 19660 38896 19712
rect 39304 19703 39356 19712
rect 39304 19669 39313 19703
rect 39313 19669 39347 19703
rect 39347 19669 39356 19703
rect 39304 19660 39356 19669
rect 39580 19660 39632 19712
rect 41512 19703 41564 19712
rect 41512 19669 41521 19703
rect 41521 19669 41555 19703
rect 41555 19669 41564 19703
rect 41512 19660 41564 19669
rect 41788 19660 41840 19712
rect 42064 19660 42116 19712
rect 43628 19839 43680 19848
rect 43628 19805 43637 19839
rect 43637 19805 43671 19839
rect 43671 19805 43680 19839
rect 43628 19796 43680 19805
rect 47308 19796 47360 19848
rect 49608 19796 49660 19848
rect 47216 19728 47268 19780
rect 43996 19660 44048 19712
rect 44180 19660 44232 19712
rect 44916 19660 44968 19712
rect 45468 19703 45520 19712
rect 45468 19669 45477 19703
rect 45477 19669 45511 19703
rect 45511 19669 45520 19703
rect 45468 19660 45520 19669
rect 46112 19660 46164 19712
rect 49332 19728 49384 19780
rect 47400 19703 47452 19712
rect 47400 19669 47409 19703
rect 47409 19669 47443 19703
rect 47443 19669 47452 19703
rect 47400 19660 47452 19669
rect 47768 19703 47820 19712
rect 47768 19669 47777 19703
rect 47777 19669 47811 19703
rect 47811 19669 47820 19703
rect 47768 19660 47820 19669
rect 48596 19660 48648 19712
rect 50436 19728 50488 19780
rect 52460 19864 52512 19916
rect 56508 19796 56560 19848
rect 51356 19660 51408 19712
rect 53012 19703 53064 19712
rect 53012 19669 53021 19703
rect 53021 19669 53055 19703
rect 53055 19669 53064 19703
rect 53012 19660 53064 19669
rect 53932 19660 53984 19712
rect 55128 19660 55180 19712
rect 15394 19558 15446 19610
rect 15458 19558 15510 19610
rect 15522 19558 15574 19610
rect 15586 19558 15638 19610
rect 15650 19558 15702 19610
rect 29838 19558 29890 19610
rect 29902 19558 29954 19610
rect 29966 19558 30018 19610
rect 30030 19558 30082 19610
rect 30094 19558 30146 19610
rect 44282 19558 44334 19610
rect 44346 19558 44398 19610
rect 44410 19558 44462 19610
rect 44474 19558 44526 19610
rect 44538 19558 44590 19610
rect 58726 19558 58778 19610
rect 58790 19558 58842 19610
rect 58854 19558 58906 19610
rect 58918 19558 58970 19610
rect 58982 19558 59034 19610
rect 3332 19456 3384 19508
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 6736 19456 6788 19508
rect 7288 19499 7340 19508
rect 7288 19465 7297 19499
rect 7297 19465 7331 19499
rect 7331 19465 7340 19499
rect 7288 19456 7340 19465
rect 11336 19499 11388 19508
rect 11336 19465 11345 19499
rect 11345 19465 11379 19499
rect 11379 19465 11388 19499
rect 11336 19456 11388 19465
rect 16488 19499 16540 19508
rect 16488 19465 16497 19499
rect 16497 19465 16531 19499
rect 16531 19465 16540 19499
rect 16488 19456 16540 19465
rect 18236 19456 18288 19508
rect 21180 19499 21232 19508
rect 21180 19465 21189 19499
rect 21189 19465 21223 19499
rect 21223 19465 21232 19499
rect 21180 19456 21232 19465
rect 22652 19456 22704 19508
rect 27344 19456 27396 19508
rect 28632 19499 28684 19508
rect 28632 19465 28641 19499
rect 28641 19465 28675 19499
rect 28675 19465 28684 19499
rect 28632 19456 28684 19465
rect 29000 19456 29052 19508
rect 29552 19456 29604 19508
rect 31208 19499 31260 19508
rect 31208 19465 31217 19499
rect 31217 19465 31251 19499
rect 31251 19465 31260 19499
rect 31208 19456 31260 19465
rect 33692 19499 33744 19508
rect 33692 19465 33701 19499
rect 33701 19465 33735 19499
rect 33735 19465 33744 19499
rect 33692 19456 33744 19465
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 6644 19320 6696 19372
rect 13728 19388 13780 19440
rect 14924 19388 14976 19440
rect 15016 19431 15068 19440
rect 15016 19397 15025 19431
rect 15025 19397 15059 19431
rect 15059 19397 15068 19431
rect 15016 19388 15068 19397
rect 11796 19320 11848 19372
rect 16948 19320 17000 19372
rect 18788 19388 18840 19440
rect 17316 19320 17368 19372
rect 19064 19363 19116 19372
rect 19064 19329 19073 19363
rect 19073 19329 19107 19363
rect 19107 19329 19116 19363
rect 19064 19320 19116 19329
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 19616 19320 19668 19372
rect 30196 19388 30248 19440
rect 28816 19320 28868 19372
rect 29736 19320 29788 19372
rect 30840 19320 30892 19372
rect 34704 19456 34756 19508
rect 33416 19320 33468 19372
rect 35624 19388 35676 19440
rect 35992 19456 36044 19508
rect 36728 19456 36780 19508
rect 36912 19499 36964 19508
rect 36912 19465 36921 19499
rect 36921 19465 36955 19499
rect 36955 19465 36964 19499
rect 36912 19456 36964 19465
rect 39304 19456 39356 19508
rect 41788 19456 41840 19508
rect 42064 19456 42116 19508
rect 36268 19388 36320 19440
rect 34336 19363 34388 19372
rect 34336 19329 34345 19363
rect 34345 19329 34379 19363
rect 34379 19329 34388 19363
rect 34336 19320 34388 19329
rect 36176 19320 36228 19372
rect 38660 19320 38712 19372
rect 39948 19320 40000 19372
rect 41972 19320 42024 19372
rect 9864 19184 9916 19236
rect 11152 19252 11204 19304
rect 12164 19252 12216 19304
rect 12348 19295 12400 19304
rect 12348 19261 12357 19295
rect 12357 19261 12391 19295
rect 12391 19261 12400 19295
rect 12348 19252 12400 19261
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 9496 19116 9548 19168
rect 9680 19116 9732 19168
rect 12900 19184 12952 19236
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 13084 19116 13136 19168
rect 18604 19227 18656 19236
rect 18604 19193 18613 19227
rect 18613 19193 18647 19227
rect 18647 19193 18656 19227
rect 18604 19184 18656 19193
rect 17408 19116 17460 19168
rect 18696 19116 18748 19168
rect 19340 19252 19392 19304
rect 23480 19252 23532 19304
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 29276 19252 29328 19261
rect 29460 19252 29512 19304
rect 39580 19295 39632 19304
rect 21548 19159 21600 19168
rect 21548 19125 21557 19159
rect 21557 19125 21591 19159
rect 21591 19125 21600 19159
rect 21548 19116 21600 19125
rect 28724 19159 28776 19168
rect 28724 19125 28733 19159
rect 28733 19125 28767 19159
rect 28767 19125 28776 19159
rect 28724 19116 28776 19125
rect 31944 19159 31996 19168
rect 31944 19125 31953 19159
rect 31953 19125 31987 19159
rect 31987 19125 31996 19159
rect 31944 19116 31996 19125
rect 34520 19116 34572 19168
rect 39580 19261 39589 19295
rect 39589 19261 39623 19295
rect 39623 19261 39632 19295
rect 39580 19252 39632 19261
rect 42616 19320 42668 19372
rect 43168 19363 43220 19372
rect 43168 19329 43177 19363
rect 43177 19329 43211 19363
rect 43211 19329 43220 19363
rect 43168 19320 43220 19329
rect 43996 19456 44048 19508
rect 44548 19499 44600 19508
rect 44548 19465 44557 19499
rect 44557 19465 44591 19499
rect 44591 19465 44600 19499
rect 44548 19456 44600 19465
rect 45008 19456 45060 19508
rect 45100 19456 45152 19508
rect 45376 19456 45428 19508
rect 45468 19456 45520 19508
rect 46112 19456 46164 19508
rect 48504 19456 48556 19508
rect 51264 19456 51316 19508
rect 53012 19456 53064 19508
rect 56600 19456 56652 19508
rect 57520 19456 57572 19508
rect 44916 19320 44968 19372
rect 47216 19388 47268 19440
rect 47400 19320 47452 19372
rect 47768 19388 47820 19440
rect 48596 19320 48648 19372
rect 48688 19320 48740 19372
rect 52092 19320 52144 19372
rect 53012 19320 53064 19372
rect 53196 19320 53248 19372
rect 58164 19320 58216 19372
rect 44548 19252 44600 19304
rect 45192 19295 45244 19304
rect 45192 19261 45201 19295
rect 45201 19261 45235 19295
rect 45235 19261 45244 19295
rect 45192 19252 45244 19261
rect 38292 19159 38344 19168
rect 38292 19125 38301 19159
rect 38301 19125 38335 19159
rect 38335 19125 38344 19159
rect 38292 19116 38344 19125
rect 38384 19116 38436 19168
rect 39028 19159 39080 19168
rect 39028 19125 39037 19159
rect 39037 19125 39071 19159
rect 39071 19125 39080 19159
rect 39028 19116 39080 19125
rect 45192 19116 45244 19168
rect 48412 19184 48464 19236
rect 50528 19295 50580 19304
rect 50528 19261 50537 19295
rect 50537 19261 50571 19295
rect 50571 19261 50580 19295
rect 50528 19252 50580 19261
rect 46940 19116 46992 19168
rect 53932 19252 53984 19304
rect 54024 19295 54076 19304
rect 54024 19261 54033 19295
rect 54033 19261 54067 19295
rect 54067 19261 54076 19295
rect 54024 19252 54076 19261
rect 57428 19295 57480 19304
rect 57428 19261 57437 19295
rect 57437 19261 57471 19295
rect 57471 19261 57480 19295
rect 57428 19252 57480 19261
rect 51172 19159 51224 19168
rect 51172 19125 51181 19159
rect 51181 19125 51215 19159
rect 51215 19125 51224 19159
rect 51172 19116 51224 19125
rect 54576 19159 54628 19168
rect 54576 19125 54585 19159
rect 54585 19125 54619 19159
rect 54619 19125 54628 19159
rect 54576 19116 54628 19125
rect 56784 19159 56836 19168
rect 56784 19125 56793 19159
rect 56793 19125 56827 19159
rect 56827 19125 56836 19159
rect 56784 19116 56836 19125
rect 57888 19116 57940 19168
rect 8172 19014 8224 19066
rect 8236 19014 8288 19066
rect 8300 19014 8352 19066
rect 8364 19014 8416 19066
rect 8428 19014 8480 19066
rect 22616 19014 22668 19066
rect 22680 19014 22732 19066
rect 22744 19014 22796 19066
rect 22808 19014 22860 19066
rect 22872 19014 22924 19066
rect 37060 19014 37112 19066
rect 37124 19014 37176 19066
rect 37188 19014 37240 19066
rect 37252 19014 37304 19066
rect 37316 19014 37368 19066
rect 51504 19014 51556 19066
rect 51568 19014 51620 19066
rect 51632 19014 51684 19066
rect 51696 19014 51748 19066
rect 51760 19014 51812 19066
rect 12072 18955 12124 18964
rect 12072 18921 12081 18955
rect 12081 18921 12115 18955
rect 12115 18921 12124 18955
rect 12072 18912 12124 18921
rect 12900 18955 12952 18964
rect 12900 18921 12909 18955
rect 12909 18921 12943 18955
rect 12943 18921 12952 18955
rect 12900 18912 12952 18921
rect 13636 18955 13688 18964
rect 13636 18921 13645 18955
rect 13645 18921 13679 18955
rect 13679 18921 13688 18955
rect 13636 18912 13688 18921
rect 15016 18912 15068 18964
rect 16856 18912 16908 18964
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 18696 18912 18748 18964
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 19892 18955 19944 18964
rect 19892 18921 19901 18955
rect 19901 18921 19935 18955
rect 19935 18921 19944 18955
rect 19892 18912 19944 18921
rect 23480 18912 23532 18964
rect 24216 18912 24268 18964
rect 12164 18844 12216 18896
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 15292 18776 15344 18828
rect 16212 18776 16264 18828
rect 24768 18844 24820 18896
rect 28816 18955 28868 18964
rect 28816 18921 28825 18955
rect 28825 18921 28859 18955
rect 28859 18921 28868 18955
rect 28816 18912 28868 18921
rect 29276 18912 29328 18964
rect 30840 18912 30892 18964
rect 34336 18912 34388 18964
rect 36176 18955 36228 18964
rect 36176 18921 36185 18955
rect 36185 18921 36219 18955
rect 36219 18921 36228 18955
rect 36176 18912 36228 18921
rect 41052 18955 41104 18964
rect 41052 18921 41061 18955
rect 41061 18921 41095 18955
rect 41095 18921 41104 18955
rect 41052 18912 41104 18921
rect 41972 18955 42024 18964
rect 41972 18921 41981 18955
rect 41981 18921 42015 18955
rect 42015 18921 42024 18955
rect 41972 18912 42024 18921
rect 43168 18912 43220 18964
rect 45100 18912 45152 18964
rect 48504 18912 48556 18964
rect 50528 18912 50580 18964
rect 54024 18912 54076 18964
rect 57888 18955 57940 18964
rect 57888 18921 57897 18955
rect 57897 18921 57931 18955
rect 57931 18921 57940 18955
rect 57888 18912 57940 18921
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 4252 18751 4304 18760
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 18604 18708 18656 18760
rect 9036 18640 9088 18692
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 4804 18615 4856 18624
rect 4804 18581 4813 18615
rect 4813 18581 4847 18615
rect 4847 18581 4856 18615
rect 4804 18572 4856 18581
rect 5080 18572 5132 18624
rect 6184 18572 6236 18624
rect 8024 18572 8076 18624
rect 12716 18572 12768 18624
rect 19432 18572 19484 18624
rect 21272 18776 21324 18828
rect 27068 18776 27120 18828
rect 28724 18776 28776 18828
rect 30656 18776 30708 18828
rect 33876 18844 33928 18896
rect 33600 18776 33652 18828
rect 38660 18844 38712 18896
rect 43260 18844 43312 18896
rect 45928 18844 45980 18896
rect 55680 18844 55732 18896
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22787 18751
rect 22787 18717 22796 18751
rect 22744 18708 22796 18717
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 26608 18751 26660 18760
rect 26608 18717 26617 18751
rect 26617 18717 26651 18751
rect 26651 18717 26660 18751
rect 26608 18708 26660 18717
rect 31944 18708 31996 18760
rect 35900 18776 35952 18828
rect 36268 18819 36320 18828
rect 36268 18785 36277 18819
rect 36277 18785 36311 18819
rect 36311 18785 36320 18819
rect 36268 18776 36320 18785
rect 36912 18776 36964 18828
rect 38292 18776 38344 18828
rect 38568 18640 38620 18692
rect 20352 18572 20404 18624
rect 21640 18572 21692 18624
rect 23296 18615 23348 18624
rect 23296 18581 23305 18615
rect 23305 18581 23339 18615
rect 23339 18581 23348 18615
rect 23296 18572 23348 18581
rect 24124 18615 24176 18624
rect 24124 18581 24133 18615
rect 24133 18581 24167 18615
rect 24167 18581 24176 18615
rect 24124 18572 24176 18581
rect 26056 18572 26108 18624
rect 26240 18615 26292 18624
rect 26240 18581 26249 18615
rect 26249 18581 26283 18615
rect 26283 18581 26292 18615
rect 26240 18572 26292 18581
rect 27252 18615 27304 18624
rect 27252 18581 27261 18615
rect 27261 18581 27295 18615
rect 27295 18581 27304 18615
rect 27252 18572 27304 18581
rect 28080 18615 28132 18624
rect 28080 18581 28089 18615
rect 28089 18581 28123 18615
rect 28123 18581 28132 18615
rect 28080 18572 28132 18581
rect 29092 18615 29144 18624
rect 29092 18581 29101 18615
rect 29101 18581 29135 18615
rect 29135 18581 29144 18615
rect 29092 18572 29144 18581
rect 30380 18572 30432 18624
rect 34428 18572 34480 18624
rect 34888 18572 34940 18624
rect 38476 18615 38528 18624
rect 38476 18581 38485 18615
rect 38485 18581 38519 18615
rect 38519 18581 38528 18615
rect 38476 18572 38528 18581
rect 38844 18615 38896 18624
rect 38844 18581 38853 18615
rect 38853 18581 38887 18615
rect 38887 18581 38896 18615
rect 38844 18572 38896 18581
rect 38936 18615 38988 18624
rect 38936 18581 38945 18615
rect 38945 18581 38979 18615
rect 38979 18581 38988 18615
rect 38936 18572 38988 18581
rect 40040 18776 40092 18828
rect 41512 18776 41564 18828
rect 50712 18819 50764 18828
rect 50712 18785 50721 18819
rect 50721 18785 50755 18819
rect 50755 18785 50764 18819
rect 50712 18776 50764 18785
rect 47492 18751 47544 18760
rect 47492 18717 47501 18751
rect 47501 18717 47535 18751
rect 47535 18717 47544 18751
rect 47492 18708 47544 18717
rect 50988 18751 51040 18760
rect 50988 18717 50997 18751
rect 50997 18717 51031 18751
rect 51031 18717 51040 18751
rect 50988 18708 51040 18717
rect 52828 18751 52880 18760
rect 52828 18717 52837 18751
rect 52837 18717 52871 18751
rect 52871 18717 52880 18751
rect 52828 18708 52880 18717
rect 56048 18708 56100 18760
rect 56508 18751 56560 18760
rect 56508 18717 56517 18751
rect 56517 18717 56551 18751
rect 56551 18717 56560 18751
rect 56508 18708 56560 18717
rect 58532 18640 58584 18692
rect 41236 18572 41288 18624
rect 47124 18572 47176 18624
rect 49976 18572 50028 18624
rect 53472 18615 53524 18624
rect 53472 18581 53481 18615
rect 53481 18581 53515 18615
rect 53515 18581 53524 18615
rect 53472 18572 53524 18581
rect 54024 18615 54076 18624
rect 54024 18581 54033 18615
rect 54033 18581 54067 18615
rect 54067 18581 54076 18615
rect 54024 18572 54076 18581
rect 54852 18572 54904 18624
rect 56508 18572 56560 18624
rect 15394 18470 15446 18522
rect 15458 18470 15510 18522
rect 15522 18470 15574 18522
rect 15586 18470 15638 18522
rect 15650 18470 15702 18522
rect 29838 18470 29890 18522
rect 29902 18470 29954 18522
rect 29966 18470 30018 18522
rect 30030 18470 30082 18522
rect 30094 18470 30146 18522
rect 44282 18470 44334 18522
rect 44346 18470 44398 18522
rect 44410 18470 44462 18522
rect 44474 18470 44526 18522
rect 44538 18470 44590 18522
rect 58726 18470 58778 18522
rect 58790 18470 58842 18522
rect 58854 18470 58906 18522
rect 58918 18470 58970 18522
rect 58982 18470 59034 18522
rect 3608 18368 3660 18420
rect 4252 18368 4304 18420
rect 8944 18368 8996 18420
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 22744 18368 22796 18420
rect 24124 18368 24176 18420
rect 24860 18411 24912 18420
rect 24860 18377 24869 18411
rect 24869 18377 24903 18411
rect 24903 18377 24912 18411
rect 24860 18368 24912 18377
rect 25044 18368 25096 18420
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 7656 18300 7708 18352
rect 4344 18096 4396 18148
rect 5080 18207 5132 18216
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 6644 18207 6696 18216
rect 6644 18173 6653 18207
rect 6653 18173 6687 18207
rect 6687 18173 6696 18207
rect 6644 18164 6696 18173
rect 8576 18164 8628 18216
rect 27252 18368 27304 18420
rect 38476 18368 38528 18420
rect 38568 18411 38620 18420
rect 38568 18377 38577 18411
rect 38577 18377 38611 18411
rect 38611 18377 38620 18411
rect 38568 18368 38620 18377
rect 38936 18368 38988 18420
rect 48320 18368 48372 18420
rect 48688 18368 48740 18420
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 25320 18232 25372 18284
rect 29460 18232 29512 18284
rect 30380 18232 30432 18284
rect 47584 18300 47636 18352
rect 48780 18300 48832 18352
rect 49332 18300 49384 18352
rect 51172 18300 51224 18352
rect 54576 18300 54628 18352
rect 56508 18368 56560 18420
rect 57428 18368 57480 18420
rect 58532 18411 58584 18420
rect 58532 18377 58541 18411
rect 58541 18377 58575 18411
rect 58575 18377 58584 18411
rect 58532 18368 58584 18377
rect 38660 18275 38712 18284
rect 38660 18241 38669 18275
rect 38669 18241 38703 18275
rect 38703 18241 38712 18275
rect 38660 18232 38712 18241
rect 53564 18232 53616 18284
rect 9036 18207 9088 18216
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 11612 18207 11664 18216
rect 11612 18173 11621 18207
rect 11621 18173 11655 18207
rect 11655 18173 11664 18207
rect 11612 18164 11664 18173
rect 14188 18164 14240 18216
rect 19800 18164 19852 18216
rect 9956 18096 10008 18148
rect 23848 18207 23900 18216
rect 23848 18173 23857 18207
rect 23857 18173 23891 18207
rect 23891 18173 23900 18207
rect 23848 18164 23900 18173
rect 24032 18164 24084 18216
rect 2504 18028 2556 18080
rect 4436 18028 4488 18080
rect 6184 18028 6236 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7932 18028 7984 18080
rect 9404 18028 9456 18080
rect 10784 18028 10836 18080
rect 12900 18028 12952 18080
rect 13820 18028 13872 18080
rect 15292 18071 15344 18080
rect 15292 18037 15301 18071
rect 15301 18037 15335 18071
rect 15335 18037 15344 18071
rect 15292 18028 15344 18037
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 22468 18028 22520 18080
rect 25136 18096 25188 18148
rect 28632 18207 28684 18216
rect 28632 18173 28641 18207
rect 28641 18173 28675 18207
rect 28675 18173 28684 18207
rect 28632 18164 28684 18173
rect 29092 18164 29144 18216
rect 24492 18071 24544 18080
rect 24492 18037 24501 18071
rect 24501 18037 24535 18071
rect 24535 18037 24544 18071
rect 24492 18028 24544 18037
rect 24952 18028 25004 18080
rect 30196 18207 30248 18216
rect 30196 18173 30205 18207
rect 30205 18173 30239 18207
rect 30239 18173 30248 18207
rect 30196 18164 30248 18173
rect 33508 18164 33560 18216
rect 33968 18207 34020 18216
rect 33968 18173 33977 18207
rect 33977 18173 34011 18207
rect 34011 18173 34020 18207
rect 33968 18164 34020 18173
rect 47400 18164 47452 18216
rect 48320 18164 48372 18216
rect 49608 18207 49660 18216
rect 49608 18173 49617 18207
rect 49617 18173 49651 18207
rect 49651 18173 49660 18207
rect 49608 18164 49660 18173
rect 53104 18164 53156 18216
rect 55680 18275 55732 18284
rect 55680 18241 55689 18275
rect 55689 18241 55723 18275
rect 55723 18241 55732 18275
rect 55680 18232 55732 18241
rect 56508 18275 56560 18284
rect 56508 18241 56542 18275
rect 56542 18241 56560 18275
rect 56508 18232 56560 18241
rect 56140 18207 56192 18216
rect 41328 18096 41380 18148
rect 41512 18096 41564 18148
rect 27620 18071 27672 18080
rect 27620 18037 27629 18071
rect 27629 18037 27663 18071
rect 27663 18037 27672 18071
rect 27620 18028 27672 18037
rect 29276 18071 29328 18080
rect 29276 18037 29285 18071
rect 29285 18037 29319 18071
rect 29319 18037 29328 18071
rect 29276 18028 29328 18037
rect 30472 18028 30524 18080
rect 33140 18028 33192 18080
rect 34612 18071 34664 18080
rect 34612 18037 34621 18071
rect 34621 18037 34655 18071
rect 34655 18037 34664 18071
rect 34612 18028 34664 18037
rect 35440 18028 35492 18080
rect 35900 18028 35952 18080
rect 36912 18028 36964 18080
rect 39948 18028 40000 18080
rect 42064 18028 42116 18080
rect 47584 18028 47636 18080
rect 47676 18028 47728 18080
rect 48228 18071 48280 18080
rect 48228 18037 48237 18071
rect 48237 18037 48271 18071
rect 48271 18037 48280 18071
rect 48228 18028 48280 18037
rect 48504 18028 48556 18080
rect 50988 18071 51040 18080
rect 50988 18037 50997 18071
rect 50997 18037 51031 18071
rect 51031 18037 51040 18071
rect 50988 18028 51040 18037
rect 52736 18028 52788 18080
rect 53380 18071 53432 18080
rect 53380 18037 53389 18071
rect 53389 18037 53423 18071
rect 53423 18037 53432 18071
rect 53380 18028 53432 18037
rect 56140 18173 56149 18207
rect 56149 18173 56183 18207
rect 56183 18173 56192 18207
rect 56140 18164 56192 18173
rect 56416 18207 56468 18216
rect 56416 18173 56425 18207
rect 56425 18173 56459 18207
rect 56459 18173 56468 18207
rect 56416 18164 56468 18173
rect 56692 18207 56744 18216
rect 56692 18173 56701 18207
rect 56701 18173 56735 18207
rect 56735 18173 56744 18207
rect 56692 18164 56744 18173
rect 57888 18207 57940 18216
rect 57888 18173 57897 18207
rect 57897 18173 57931 18207
rect 57931 18173 57940 18207
rect 57888 18164 57940 18173
rect 57428 18028 57480 18080
rect 8172 17926 8224 17978
rect 8236 17926 8288 17978
rect 8300 17926 8352 17978
rect 8364 17926 8416 17978
rect 8428 17926 8480 17978
rect 22616 17926 22668 17978
rect 22680 17926 22732 17978
rect 22744 17926 22796 17978
rect 22808 17926 22860 17978
rect 22872 17926 22924 17978
rect 37060 17926 37112 17978
rect 37124 17926 37176 17978
rect 37188 17926 37240 17978
rect 37252 17926 37304 17978
rect 37316 17926 37368 17978
rect 51504 17926 51556 17978
rect 51568 17926 51620 17978
rect 51632 17926 51684 17978
rect 51696 17926 51748 17978
rect 51760 17926 51812 17978
rect 3056 17824 3108 17876
rect 4712 17824 4764 17876
rect 8576 17824 8628 17876
rect 9312 17824 9364 17876
rect 4436 17731 4488 17740
rect 4436 17697 4445 17731
rect 4445 17697 4479 17731
rect 4479 17697 4488 17731
rect 4436 17688 4488 17697
rect 5172 17688 5224 17740
rect 8576 17688 8628 17740
rect 9404 17688 9456 17740
rect 4160 17620 4212 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 4896 17620 4948 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 2504 17552 2556 17604
rect 2780 17552 2832 17604
rect 6828 17620 6880 17672
rect 20444 17824 20496 17876
rect 12900 17756 12952 17808
rect 19524 17756 19576 17808
rect 7288 17552 7340 17604
rect 7932 17552 7984 17604
rect 10508 17552 10560 17604
rect 20536 17731 20588 17740
rect 10784 17663 10836 17672
rect 10784 17629 10818 17663
rect 10818 17629 10836 17663
rect 10784 17620 10836 17629
rect 11060 17620 11112 17672
rect 11520 17620 11572 17672
rect 12900 17663 12952 17672
rect 12900 17629 12909 17663
rect 12909 17629 12943 17663
rect 12943 17629 12952 17663
rect 12900 17620 12952 17629
rect 14096 17620 14148 17672
rect 14740 17620 14792 17672
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 11336 17552 11388 17604
rect 20536 17697 20545 17731
rect 20545 17697 20579 17731
rect 20579 17697 20588 17731
rect 20536 17688 20588 17697
rect 23572 17799 23624 17808
rect 23572 17765 23581 17799
rect 23581 17765 23615 17799
rect 23615 17765 23624 17799
rect 25412 17824 25464 17876
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 26608 17824 26660 17876
rect 30196 17867 30248 17876
rect 30196 17833 30205 17867
rect 30205 17833 30239 17867
rect 30239 17833 30248 17867
rect 30196 17824 30248 17833
rect 38292 17824 38344 17876
rect 47400 17824 47452 17876
rect 23572 17756 23624 17765
rect 26148 17756 26200 17808
rect 24952 17688 25004 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 25136 17688 25188 17740
rect 20720 17620 20772 17672
rect 23296 17620 23348 17672
rect 24768 17620 24820 17672
rect 25412 17731 25464 17740
rect 25412 17697 25446 17731
rect 25446 17697 25464 17731
rect 25412 17688 25464 17697
rect 26332 17688 26384 17740
rect 25596 17663 25648 17672
rect 25596 17629 25605 17663
rect 25605 17629 25639 17663
rect 25639 17629 25648 17663
rect 25596 17620 25648 17629
rect 27620 17756 27672 17808
rect 26976 17731 27028 17740
rect 26976 17697 26985 17731
rect 26985 17697 27019 17731
rect 27019 17697 27028 17731
rect 26976 17688 27028 17697
rect 29276 17688 29328 17740
rect 33140 17688 33192 17740
rect 34244 17731 34296 17740
rect 27620 17663 27672 17672
rect 27620 17629 27629 17663
rect 27629 17629 27663 17663
rect 27663 17629 27672 17663
rect 27620 17620 27672 17629
rect 30380 17620 30432 17672
rect 31116 17663 31168 17672
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 5540 17484 5592 17536
rect 5632 17527 5684 17536
rect 5632 17493 5641 17527
rect 5641 17493 5675 17527
rect 5675 17493 5684 17527
rect 5632 17484 5684 17493
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 8760 17484 8812 17536
rect 10876 17484 10928 17536
rect 11428 17484 11480 17536
rect 11980 17527 12032 17536
rect 11980 17493 11989 17527
rect 11989 17493 12023 17527
rect 12023 17493 12032 17527
rect 11980 17484 12032 17493
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 13820 17527 13872 17536
rect 13820 17493 13829 17527
rect 13829 17493 13863 17527
rect 13863 17493 13872 17527
rect 13820 17484 13872 17493
rect 14188 17484 14240 17536
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 18144 17484 18196 17493
rect 20076 17484 20128 17536
rect 20352 17484 20404 17536
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 22192 17484 22244 17536
rect 23940 17484 23992 17536
rect 24124 17527 24176 17536
rect 24124 17493 24133 17527
rect 24133 17493 24167 17527
rect 24167 17493 24176 17527
rect 24124 17484 24176 17493
rect 24308 17484 24360 17536
rect 25596 17484 25648 17536
rect 27344 17527 27396 17536
rect 27344 17493 27353 17527
rect 27353 17493 27387 17527
rect 27387 17493 27396 17527
rect 27344 17484 27396 17493
rect 34244 17697 34253 17731
rect 34253 17697 34287 17731
rect 34287 17697 34296 17731
rect 40776 17731 40828 17740
rect 34244 17688 34296 17697
rect 40776 17697 40785 17731
rect 40785 17697 40819 17731
rect 40819 17697 40828 17731
rect 40776 17688 40828 17697
rect 43352 17688 43404 17740
rect 34520 17620 34572 17672
rect 38108 17620 38160 17672
rect 38936 17620 38988 17672
rect 40132 17663 40184 17672
rect 40132 17629 40141 17663
rect 40141 17629 40175 17663
rect 40175 17629 40184 17663
rect 40132 17620 40184 17629
rect 41512 17663 41564 17672
rect 41512 17629 41521 17663
rect 41521 17629 41555 17663
rect 41555 17629 41564 17663
rect 41512 17620 41564 17629
rect 44180 17620 44232 17672
rect 27712 17484 27764 17536
rect 27896 17484 27948 17536
rect 29368 17527 29420 17536
rect 29368 17493 29377 17527
rect 29377 17493 29411 17527
rect 29411 17493 29420 17527
rect 29368 17484 29420 17493
rect 32772 17527 32824 17536
rect 32772 17493 32781 17527
rect 32781 17493 32815 17527
rect 32815 17493 32824 17527
rect 32772 17484 32824 17493
rect 33140 17484 33192 17536
rect 35348 17527 35400 17536
rect 35348 17493 35357 17527
rect 35357 17493 35391 17527
rect 35391 17493 35400 17527
rect 35348 17484 35400 17493
rect 36636 17484 36688 17536
rect 36728 17484 36780 17536
rect 38200 17527 38252 17536
rect 38200 17493 38209 17527
rect 38209 17493 38243 17527
rect 38243 17493 38252 17527
rect 38200 17484 38252 17493
rect 38752 17484 38804 17536
rect 47676 17731 47728 17740
rect 47676 17697 47685 17731
rect 47685 17697 47719 17731
rect 47719 17697 47728 17731
rect 47676 17688 47728 17697
rect 48504 17688 48556 17740
rect 48688 17688 48740 17740
rect 49332 17731 49384 17740
rect 49332 17697 49341 17731
rect 49341 17697 49375 17731
rect 49375 17697 49384 17731
rect 49332 17688 49384 17697
rect 52460 17824 52512 17876
rect 57428 17867 57480 17876
rect 57428 17833 57437 17867
rect 57437 17833 57471 17867
rect 57471 17833 57480 17867
rect 57428 17824 57480 17833
rect 57888 17824 57940 17876
rect 48136 17663 48188 17672
rect 48136 17629 48145 17663
rect 48145 17629 48179 17663
rect 48179 17629 48188 17663
rect 48136 17620 48188 17629
rect 49056 17663 49108 17672
rect 49056 17629 49065 17663
rect 49065 17629 49099 17663
rect 49099 17629 49108 17663
rect 49056 17620 49108 17629
rect 40040 17484 40092 17536
rect 40684 17527 40736 17536
rect 40684 17493 40693 17527
rect 40693 17493 40727 17527
rect 40727 17493 40736 17527
rect 40684 17484 40736 17493
rect 41420 17527 41472 17536
rect 41420 17493 41429 17527
rect 41429 17493 41463 17527
rect 41463 17493 41472 17527
rect 41420 17484 41472 17493
rect 42156 17527 42208 17536
rect 42156 17493 42165 17527
rect 42165 17493 42199 17527
rect 42199 17493 42208 17527
rect 42156 17484 42208 17493
rect 43904 17527 43956 17536
rect 43904 17493 43913 17527
rect 43913 17493 43947 17527
rect 43947 17493 43956 17527
rect 43904 17484 43956 17493
rect 44640 17484 44692 17536
rect 44916 17484 44968 17536
rect 45468 17484 45520 17536
rect 46940 17527 46992 17536
rect 46940 17493 46949 17527
rect 46949 17493 46983 17527
rect 46983 17493 46992 17527
rect 46940 17484 46992 17493
rect 47308 17484 47360 17536
rect 47952 17484 48004 17536
rect 48044 17484 48096 17536
rect 57520 17688 57572 17740
rect 50068 17620 50120 17672
rect 51356 17620 51408 17672
rect 53472 17620 53524 17672
rect 56048 17663 56100 17672
rect 52736 17552 52788 17604
rect 50160 17527 50212 17536
rect 50160 17493 50169 17527
rect 50169 17493 50203 17527
rect 50203 17493 50212 17527
rect 50160 17484 50212 17493
rect 51908 17484 51960 17536
rect 53104 17527 53156 17536
rect 53104 17493 53113 17527
rect 53113 17493 53147 17527
rect 53147 17493 53156 17527
rect 53104 17484 53156 17493
rect 53564 17484 53616 17536
rect 56048 17629 56057 17663
rect 56057 17629 56091 17663
rect 56091 17629 56100 17663
rect 56048 17620 56100 17629
rect 55496 17595 55548 17604
rect 55496 17561 55505 17595
rect 55505 17561 55539 17595
rect 55539 17561 55548 17595
rect 56692 17620 56744 17672
rect 56876 17620 56928 17672
rect 58164 17620 58216 17672
rect 55496 17552 55548 17561
rect 57060 17552 57112 17604
rect 57796 17484 57848 17536
rect 58440 17484 58492 17536
rect 15394 17382 15446 17434
rect 15458 17382 15510 17434
rect 15522 17382 15574 17434
rect 15586 17382 15638 17434
rect 15650 17382 15702 17434
rect 29838 17382 29890 17434
rect 29902 17382 29954 17434
rect 29966 17382 30018 17434
rect 30030 17382 30082 17434
rect 30094 17382 30146 17434
rect 44282 17382 44334 17434
rect 44346 17382 44398 17434
rect 44410 17382 44462 17434
rect 44474 17382 44526 17434
rect 44538 17382 44590 17434
rect 58726 17382 58778 17434
rect 58790 17382 58842 17434
rect 58854 17382 58906 17434
rect 58918 17382 58970 17434
rect 58982 17382 59034 17434
rect 5632 17280 5684 17332
rect 5908 17280 5960 17332
rect 6644 17280 6696 17332
rect 6920 17280 6972 17332
rect 9220 17280 9272 17332
rect 2780 17212 2832 17264
rect 4804 17212 4856 17264
rect 4896 17212 4948 17264
rect 6828 17212 6880 17264
rect 8024 17255 8076 17264
rect 4160 17144 4212 17196
rect 6368 17144 6420 17196
rect 7104 17144 7156 17196
rect 8024 17221 8058 17255
rect 8058 17221 8076 17255
rect 8024 17212 8076 17221
rect 11336 17323 11388 17332
rect 11336 17289 11345 17323
rect 11345 17289 11379 17323
rect 11379 17289 11388 17323
rect 11336 17280 11388 17289
rect 11612 17280 11664 17332
rect 12900 17280 12952 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 15292 17280 15344 17332
rect 17592 17280 17644 17332
rect 2780 17076 2832 17128
rect 5264 17076 5316 17128
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 9220 17144 9272 17196
rect 9312 17076 9364 17128
rect 9588 17076 9640 17128
rect 10508 17187 10560 17196
rect 10508 17153 10542 17187
rect 10542 17153 10560 17187
rect 10508 17144 10560 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 4528 16940 4580 16992
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 5908 16940 5960 16992
rect 6828 16940 6880 16992
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 10876 17076 10928 17128
rect 11796 17076 11848 17128
rect 13728 17144 13780 17196
rect 13912 17212 13964 17264
rect 15936 17255 15988 17264
rect 15936 17221 15945 17255
rect 15945 17221 15979 17255
rect 15979 17221 15988 17255
rect 15936 17212 15988 17221
rect 16396 17212 16448 17264
rect 20260 17280 20312 17332
rect 19524 17255 19576 17264
rect 19524 17221 19533 17255
rect 19533 17221 19567 17255
rect 19567 17221 19576 17255
rect 19524 17212 19576 17221
rect 14832 17144 14884 17196
rect 19340 17144 19392 17196
rect 21456 17144 21508 17196
rect 22192 17280 22244 17332
rect 23848 17280 23900 17332
rect 24492 17280 24544 17332
rect 24768 17280 24820 17332
rect 24032 17255 24084 17264
rect 24032 17221 24041 17255
rect 24041 17221 24075 17255
rect 24075 17221 24084 17255
rect 24032 17212 24084 17221
rect 23756 17144 23808 17196
rect 23940 17144 23992 17196
rect 24400 17144 24452 17196
rect 25320 17212 25372 17264
rect 25596 17144 25648 17196
rect 9772 17008 9824 17060
rect 11428 16940 11480 16992
rect 12716 17076 12768 17128
rect 13360 17076 13412 17128
rect 12164 16940 12216 16992
rect 14004 17008 14056 17060
rect 14740 17076 14792 17128
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 24308 17119 24360 17128
rect 24308 17085 24317 17119
rect 24317 17085 24351 17119
rect 24351 17085 24360 17119
rect 24308 17076 24360 17085
rect 28632 17280 28684 17332
rect 29368 17280 29420 17332
rect 31852 17323 31904 17332
rect 26240 17076 26292 17128
rect 13820 16940 13872 16992
rect 14372 16940 14424 16992
rect 19800 16940 19852 16992
rect 23664 16983 23716 16992
rect 23664 16949 23673 16983
rect 23673 16949 23707 16983
rect 23707 16949 23716 16983
rect 23664 16940 23716 16949
rect 26608 16983 26660 16992
rect 26608 16949 26617 16983
rect 26617 16949 26651 16983
rect 26651 16949 26660 16983
rect 26608 16940 26660 16949
rect 27344 16940 27396 16992
rect 31852 17289 31861 17323
rect 31861 17289 31895 17323
rect 31895 17289 31904 17323
rect 31852 17280 31904 17289
rect 33140 17280 33192 17332
rect 33968 17280 34020 17332
rect 35348 17280 35400 17332
rect 40040 17280 40092 17332
rect 40684 17280 40736 17332
rect 40776 17280 40828 17332
rect 41512 17323 41564 17332
rect 41512 17289 41521 17323
rect 41521 17289 41555 17323
rect 41555 17289 41564 17323
rect 41512 17280 41564 17289
rect 44916 17323 44968 17332
rect 35256 17212 35308 17264
rect 32772 17144 32824 17196
rect 33324 17076 33376 17128
rect 34888 17076 34940 17128
rect 35440 17119 35492 17128
rect 35440 17085 35449 17119
rect 35449 17085 35483 17119
rect 35483 17085 35492 17119
rect 35440 17076 35492 17085
rect 35624 17119 35676 17128
rect 35624 17085 35633 17119
rect 35633 17085 35667 17119
rect 35667 17085 35676 17119
rect 35624 17076 35676 17085
rect 38108 17187 38160 17196
rect 38108 17153 38117 17187
rect 38117 17153 38151 17187
rect 38151 17153 38160 17187
rect 38108 17144 38160 17153
rect 44916 17289 44925 17323
rect 44925 17289 44959 17323
rect 44959 17289 44968 17323
rect 44916 17280 44968 17289
rect 47400 17323 47452 17332
rect 47400 17289 47409 17323
rect 47409 17289 47443 17323
rect 47443 17289 47452 17323
rect 47400 17280 47452 17289
rect 47492 17280 47544 17332
rect 48228 17280 48280 17332
rect 42708 17212 42760 17264
rect 48320 17212 48372 17264
rect 47124 17144 47176 17196
rect 47308 17144 47360 17196
rect 49516 17280 49568 17332
rect 49976 17280 50028 17332
rect 52828 17280 52880 17332
rect 53380 17280 53432 17332
rect 55404 17280 55456 17332
rect 56416 17280 56468 17332
rect 56692 17280 56744 17332
rect 58440 17280 58492 17332
rect 28080 16940 28132 16992
rect 28908 16940 28960 16992
rect 29552 16983 29604 16992
rect 29552 16949 29561 16983
rect 29561 16949 29595 16983
rect 29595 16949 29604 16983
rect 29552 16940 29604 16949
rect 33508 16983 33560 16992
rect 33508 16949 33517 16983
rect 33517 16949 33551 16983
rect 33551 16949 33560 16983
rect 33508 16940 33560 16949
rect 34336 16940 34388 16992
rect 35992 16940 36044 16992
rect 38660 17076 38712 17128
rect 39028 17076 39080 17128
rect 39488 17076 39540 17128
rect 41972 17119 42024 17128
rect 41972 17085 41981 17119
rect 41981 17085 42015 17119
rect 42015 17085 42024 17119
rect 41972 17076 42024 17085
rect 42064 17119 42116 17128
rect 42064 17085 42073 17119
rect 42073 17085 42107 17119
rect 42107 17085 42116 17119
rect 42064 17076 42116 17085
rect 42432 17119 42484 17128
rect 42432 17085 42441 17119
rect 42441 17085 42475 17119
rect 42475 17085 42484 17119
rect 42432 17076 42484 17085
rect 43444 17076 43496 17128
rect 45008 17119 45060 17128
rect 45008 17085 45017 17119
rect 45017 17085 45051 17119
rect 45051 17085 45060 17119
rect 45008 17076 45060 17085
rect 38660 16940 38712 16992
rect 39764 16983 39816 16992
rect 39764 16949 39773 16983
rect 39773 16949 39807 16983
rect 39807 16949 39816 16983
rect 39764 16940 39816 16949
rect 49148 17076 49200 17128
rect 42064 16940 42116 16992
rect 43444 16983 43496 16992
rect 43444 16949 43453 16983
rect 43453 16949 43487 16983
rect 43487 16949 43496 16983
rect 43444 16940 43496 16949
rect 50528 17119 50580 17128
rect 50528 17085 50537 17119
rect 50537 17085 50571 17119
rect 50571 17085 50580 17119
rect 50528 17076 50580 17085
rect 53012 17144 53064 17196
rect 53380 17076 53432 17128
rect 53564 17076 53616 17128
rect 49700 16940 49752 16992
rect 50436 16983 50488 16992
rect 50436 16949 50445 16983
rect 50445 16949 50479 16983
rect 50479 16949 50488 16983
rect 50436 16940 50488 16949
rect 55128 17119 55180 17128
rect 55128 17085 55137 17119
rect 55137 17085 55171 17119
rect 55171 17085 55180 17119
rect 55128 17076 55180 17085
rect 57428 17076 57480 17128
rect 53840 16940 53892 16992
rect 56324 16983 56376 16992
rect 56324 16949 56333 16983
rect 56333 16949 56367 16983
rect 56367 16949 56376 16983
rect 56324 16940 56376 16949
rect 56416 16983 56468 16992
rect 56416 16949 56425 16983
rect 56425 16949 56459 16983
rect 56459 16949 56468 16983
rect 56416 16940 56468 16949
rect 57428 16983 57480 16992
rect 57428 16949 57437 16983
rect 57437 16949 57471 16983
rect 57471 16949 57480 16983
rect 57428 16940 57480 16949
rect 8172 16838 8224 16890
rect 8236 16838 8288 16890
rect 8300 16838 8352 16890
rect 8364 16838 8416 16890
rect 8428 16838 8480 16890
rect 22616 16838 22668 16890
rect 22680 16838 22732 16890
rect 22744 16838 22796 16890
rect 22808 16838 22860 16890
rect 22872 16838 22924 16890
rect 37060 16838 37112 16890
rect 37124 16838 37176 16890
rect 37188 16838 37240 16890
rect 37252 16838 37304 16890
rect 37316 16838 37368 16890
rect 51504 16838 51556 16890
rect 51568 16838 51620 16890
rect 51632 16838 51684 16890
rect 51696 16838 51748 16890
rect 51760 16838 51812 16890
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 3332 16736 3384 16788
rect 4528 16736 4580 16788
rect 5908 16736 5960 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 8576 16668 8628 16720
rect 8760 16668 8812 16720
rect 10692 16736 10744 16788
rect 11428 16736 11480 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12164 16779 12216 16788
rect 12164 16745 12173 16779
rect 12173 16745 12207 16779
rect 12207 16745 12216 16779
rect 12164 16736 12216 16745
rect 9496 16668 9548 16720
rect 9772 16668 9824 16720
rect 3700 16600 3752 16652
rect 4896 16600 4948 16652
rect 4988 16600 5040 16652
rect 6368 16643 6420 16652
rect 6368 16609 6377 16643
rect 6377 16609 6411 16643
rect 6411 16609 6420 16643
rect 6368 16600 6420 16609
rect 8484 16600 8536 16652
rect 12072 16532 12124 16584
rect 14096 16736 14148 16788
rect 13912 16668 13964 16720
rect 14188 16600 14240 16652
rect 13452 16532 13504 16584
rect 14188 16396 14240 16448
rect 14372 16600 14424 16652
rect 16396 16668 16448 16720
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 18604 16736 18656 16788
rect 20168 16736 20220 16788
rect 20260 16736 20312 16788
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 19800 16600 19852 16652
rect 19892 16643 19944 16652
rect 19892 16609 19901 16643
rect 19901 16609 19935 16643
rect 19935 16609 19944 16643
rect 19892 16600 19944 16609
rect 20812 16600 20864 16652
rect 23296 16736 23348 16788
rect 23664 16736 23716 16788
rect 23756 16779 23808 16788
rect 23756 16745 23765 16779
rect 23765 16745 23799 16779
rect 23799 16745 23808 16779
rect 23756 16736 23808 16745
rect 24400 16736 24452 16788
rect 24860 16736 24912 16788
rect 25688 16736 25740 16788
rect 24032 16668 24084 16720
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 15108 16575 15160 16584
rect 15108 16541 15142 16575
rect 15142 16541 15160 16575
rect 15108 16532 15160 16541
rect 16120 16532 16172 16584
rect 18144 16532 18196 16584
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 15200 16396 15252 16448
rect 15292 16396 15344 16448
rect 19064 16439 19116 16448
rect 19064 16405 19073 16439
rect 19073 16405 19107 16439
rect 19107 16405 19116 16439
rect 19064 16396 19116 16405
rect 20168 16575 20220 16584
rect 20168 16541 20177 16575
rect 20177 16541 20211 16575
rect 20211 16541 20220 16575
rect 20168 16532 20220 16541
rect 20260 16575 20312 16584
rect 20260 16541 20294 16575
rect 20294 16541 20312 16575
rect 20260 16532 20312 16541
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 26608 16668 26660 16720
rect 28908 16736 28960 16788
rect 31668 16779 31720 16788
rect 29092 16668 29144 16720
rect 25688 16643 25740 16652
rect 25688 16609 25697 16643
rect 25697 16609 25731 16643
rect 25731 16609 25740 16643
rect 25688 16600 25740 16609
rect 26240 16600 26292 16652
rect 27344 16643 27396 16652
rect 27344 16609 27353 16643
rect 27353 16609 27387 16643
rect 27387 16609 27396 16643
rect 27344 16600 27396 16609
rect 28356 16600 28408 16652
rect 29368 16600 29420 16652
rect 31668 16745 31677 16779
rect 31677 16745 31711 16779
rect 31711 16745 31720 16779
rect 31668 16736 31720 16745
rect 31852 16736 31904 16788
rect 34520 16711 34572 16720
rect 34520 16677 34529 16711
rect 34529 16677 34563 16711
rect 34563 16677 34572 16711
rect 34520 16668 34572 16677
rect 34704 16643 34756 16652
rect 34704 16609 34713 16643
rect 34713 16609 34747 16643
rect 34747 16609 34756 16643
rect 34704 16600 34756 16609
rect 36636 16643 36688 16652
rect 36636 16609 36645 16643
rect 36645 16609 36679 16643
rect 36679 16609 36688 16643
rect 36636 16600 36688 16609
rect 26148 16532 26200 16584
rect 21088 16464 21140 16516
rect 26976 16464 27028 16516
rect 27896 16532 27948 16584
rect 30472 16532 30524 16584
rect 32128 16575 32180 16584
rect 32128 16541 32137 16575
rect 32137 16541 32171 16575
rect 32171 16541 32180 16575
rect 32128 16532 32180 16541
rect 34612 16532 34664 16584
rect 35992 16532 36044 16584
rect 38936 16779 38988 16788
rect 38936 16745 38945 16779
rect 38945 16745 38979 16779
rect 38979 16745 38988 16779
rect 38936 16736 38988 16745
rect 40132 16736 40184 16788
rect 38200 16600 38252 16652
rect 39488 16600 39540 16652
rect 42432 16736 42484 16788
rect 40040 16600 40092 16652
rect 40408 16643 40460 16652
rect 40408 16609 40417 16643
rect 40417 16609 40451 16643
rect 40451 16609 40460 16643
rect 40408 16600 40460 16609
rect 41788 16600 41840 16652
rect 42708 16643 42760 16652
rect 42708 16609 42717 16643
rect 42717 16609 42751 16643
rect 42751 16609 42760 16643
rect 42708 16600 42760 16609
rect 43260 16600 43312 16652
rect 44088 16736 44140 16788
rect 44640 16736 44692 16788
rect 45008 16779 45060 16788
rect 45008 16745 45017 16779
rect 45017 16745 45051 16779
rect 45051 16745 45060 16779
rect 45008 16736 45060 16745
rect 47492 16736 47544 16788
rect 48136 16736 48188 16788
rect 50528 16736 50580 16788
rect 20260 16396 20312 16448
rect 20904 16396 20956 16448
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25044 16396 25096 16405
rect 28080 16396 28132 16448
rect 33508 16464 33560 16516
rect 39028 16532 39080 16584
rect 42156 16532 42208 16584
rect 38200 16464 38252 16516
rect 28816 16396 28868 16448
rect 30380 16396 30432 16448
rect 31116 16396 31168 16448
rect 32680 16439 32732 16448
rect 32680 16405 32689 16439
rect 32689 16405 32723 16439
rect 32723 16405 32732 16439
rect 32680 16396 32732 16405
rect 34612 16396 34664 16448
rect 35624 16396 35676 16448
rect 38108 16439 38160 16448
rect 38108 16405 38117 16439
rect 38117 16405 38151 16439
rect 38151 16405 38160 16439
rect 38108 16396 38160 16405
rect 38476 16439 38528 16448
rect 38476 16405 38485 16439
rect 38485 16405 38519 16439
rect 38519 16405 38528 16439
rect 38476 16396 38528 16405
rect 38844 16396 38896 16448
rect 39304 16439 39356 16448
rect 39304 16405 39313 16439
rect 39313 16405 39347 16439
rect 39347 16405 39356 16439
rect 39304 16396 39356 16405
rect 39396 16439 39448 16448
rect 39396 16405 39405 16439
rect 39405 16405 39439 16439
rect 39439 16405 39448 16439
rect 39396 16396 39448 16405
rect 41420 16464 41472 16516
rect 40960 16396 41012 16448
rect 42524 16439 42576 16448
rect 42524 16405 42533 16439
rect 42533 16405 42567 16439
rect 42567 16405 42576 16439
rect 42524 16396 42576 16405
rect 43628 16575 43680 16584
rect 43628 16541 43637 16575
rect 43637 16541 43671 16575
rect 43671 16541 43680 16575
rect 43628 16532 43680 16541
rect 45468 16643 45520 16652
rect 45468 16609 45477 16643
rect 45477 16609 45511 16643
rect 45511 16609 45520 16643
rect 45468 16600 45520 16609
rect 46388 16600 46440 16652
rect 48320 16600 48372 16652
rect 51908 16736 51960 16788
rect 55128 16736 55180 16788
rect 56416 16736 56468 16788
rect 56692 16736 56744 16788
rect 57060 16779 57112 16788
rect 57060 16745 57069 16779
rect 57069 16745 57103 16779
rect 57103 16745 57112 16779
rect 57060 16736 57112 16745
rect 53840 16600 53892 16652
rect 54760 16643 54812 16652
rect 54760 16609 54769 16643
rect 54769 16609 54803 16643
rect 54803 16609 54812 16643
rect 54760 16600 54812 16609
rect 55404 16643 55456 16652
rect 55404 16609 55413 16643
rect 55413 16609 55447 16643
rect 55447 16609 55456 16643
rect 55404 16600 55456 16609
rect 46572 16532 46624 16584
rect 50436 16532 50488 16584
rect 53196 16575 53248 16584
rect 53196 16541 53205 16575
rect 53205 16541 53239 16575
rect 53239 16541 53248 16575
rect 53196 16532 53248 16541
rect 54852 16532 54904 16584
rect 44640 16464 44692 16516
rect 46940 16464 46992 16516
rect 49056 16464 49108 16516
rect 44916 16396 44968 16448
rect 48320 16396 48372 16448
rect 51908 16396 51960 16448
rect 15394 16294 15446 16346
rect 15458 16294 15510 16346
rect 15522 16294 15574 16346
rect 15586 16294 15638 16346
rect 15650 16294 15702 16346
rect 29838 16294 29890 16346
rect 29902 16294 29954 16346
rect 29966 16294 30018 16346
rect 30030 16294 30082 16346
rect 30094 16294 30146 16346
rect 44282 16294 44334 16346
rect 44346 16294 44398 16346
rect 44410 16294 44462 16346
rect 44474 16294 44526 16346
rect 44538 16294 44590 16346
rect 58726 16294 58778 16346
rect 58790 16294 58842 16346
rect 58854 16294 58906 16346
rect 58918 16294 58970 16346
rect 58982 16294 59034 16346
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 7932 16192 7984 16244
rect 11612 16192 11664 16244
rect 13728 16192 13780 16244
rect 14832 16192 14884 16244
rect 15936 16192 15988 16244
rect 18512 16192 18564 16244
rect 19064 16192 19116 16244
rect 20812 16192 20864 16244
rect 25596 16235 25648 16244
rect 25596 16201 25605 16235
rect 25605 16201 25639 16235
rect 25639 16201 25648 16235
rect 25596 16192 25648 16201
rect 26332 16192 26384 16244
rect 27436 16235 27488 16244
rect 27436 16201 27445 16235
rect 27445 16201 27479 16235
rect 27479 16201 27488 16235
rect 27436 16192 27488 16201
rect 27620 16235 27672 16244
rect 27620 16201 27629 16235
rect 27629 16201 27663 16235
rect 27663 16201 27672 16235
rect 27620 16192 27672 16201
rect 28080 16235 28132 16244
rect 28080 16201 28089 16235
rect 28089 16201 28123 16235
rect 28123 16201 28132 16235
rect 28080 16192 28132 16201
rect 13176 16124 13228 16176
rect 17960 16124 18012 16176
rect 19340 16124 19392 16176
rect 20260 16124 20312 16176
rect 13636 16056 13688 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 18512 16056 18564 16108
rect 21364 16056 21416 16108
rect 25044 16099 25096 16108
rect 25044 16065 25053 16099
rect 25053 16065 25087 16099
rect 25087 16065 25096 16099
rect 25044 16056 25096 16065
rect 27988 16099 28040 16108
rect 27988 16065 27997 16099
rect 27997 16065 28031 16099
rect 28031 16065 28040 16099
rect 27988 16056 28040 16065
rect 28356 16056 28408 16108
rect 28540 16056 28592 16108
rect 30380 16192 30432 16244
rect 30932 16192 30984 16244
rect 32128 16192 32180 16244
rect 32772 16192 32824 16244
rect 33324 16235 33376 16244
rect 33324 16201 33333 16235
rect 33333 16201 33367 16235
rect 33367 16201 33376 16235
rect 33324 16192 33376 16201
rect 28816 16056 28868 16108
rect 29644 16099 29696 16108
rect 29644 16065 29653 16099
rect 29653 16065 29687 16099
rect 29687 16065 29696 16099
rect 29644 16056 29696 16065
rect 33140 16056 33192 16108
rect 34520 16192 34572 16244
rect 36544 16192 36596 16244
rect 36636 16192 36688 16244
rect 34336 16099 34388 16108
rect 34336 16065 34345 16099
rect 34345 16065 34379 16099
rect 34379 16065 34388 16099
rect 34336 16056 34388 16065
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 14464 16031 14516 16040
rect 14464 15997 14473 16031
rect 14473 15997 14507 16031
rect 14507 15997 14516 16031
rect 14464 15988 14516 15997
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 9588 15852 9640 15904
rect 11060 15852 11112 15904
rect 11428 15852 11480 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 14280 15852 14332 15904
rect 15016 15920 15068 15972
rect 19524 16031 19576 16040
rect 19524 15997 19533 16031
rect 19533 15997 19567 16031
rect 19567 15997 19576 16031
rect 19524 15988 19576 15997
rect 20812 15988 20864 16040
rect 22468 15988 22520 16040
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 19156 15852 19208 15904
rect 26792 15963 26844 15972
rect 26792 15929 26801 15963
rect 26801 15929 26835 15963
rect 26835 15929 26844 15963
rect 26792 15920 26844 15929
rect 29000 15920 29052 15972
rect 21640 15895 21692 15904
rect 21640 15861 21649 15895
rect 21649 15861 21683 15895
rect 21683 15861 21692 15895
rect 21640 15852 21692 15861
rect 24308 15852 24360 15904
rect 26608 15852 26660 15904
rect 28080 15852 28132 15904
rect 33508 15988 33560 16040
rect 30196 15852 30248 15904
rect 30380 15895 30432 15904
rect 30380 15861 30389 15895
rect 30389 15861 30423 15895
rect 30423 15861 30432 15895
rect 30380 15852 30432 15861
rect 34428 16031 34480 16040
rect 34428 15997 34462 16031
rect 34462 15997 34480 16031
rect 34428 15988 34480 15997
rect 34980 15988 35032 16040
rect 36728 16056 36780 16108
rect 38660 16235 38712 16244
rect 38660 16201 38669 16235
rect 38669 16201 38703 16235
rect 38703 16201 38712 16235
rect 38660 16192 38712 16201
rect 39488 16192 39540 16244
rect 39764 16192 39816 16244
rect 40040 16192 40092 16244
rect 42800 16192 42852 16244
rect 43628 16192 43680 16244
rect 43996 16192 44048 16244
rect 44640 16192 44692 16244
rect 44916 16235 44968 16244
rect 44916 16201 44925 16235
rect 44925 16201 44959 16235
rect 44959 16201 44968 16235
rect 44916 16192 44968 16201
rect 45928 16235 45980 16244
rect 45928 16201 45937 16235
rect 45937 16201 45971 16235
rect 45971 16201 45980 16235
rect 45928 16192 45980 16201
rect 47952 16192 48004 16244
rect 51080 16235 51132 16244
rect 51080 16201 51089 16235
rect 51089 16201 51123 16235
rect 51123 16201 51132 16235
rect 51080 16192 51132 16201
rect 51172 16192 51224 16244
rect 52644 16192 52696 16244
rect 53196 16192 53248 16244
rect 54760 16192 54812 16244
rect 38752 16124 38804 16176
rect 40224 16124 40276 16176
rect 40316 16124 40368 16176
rect 56784 16124 56836 16176
rect 40960 16056 41012 16108
rect 48320 16056 48372 16108
rect 34060 15963 34112 15972
rect 34060 15929 34069 15963
rect 34069 15929 34103 15963
rect 34103 15929 34112 15963
rect 34060 15920 34112 15929
rect 34612 15852 34664 15904
rect 34796 15852 34848 15904
rect 36360 15852 36412 15904
rect 39488 15852 39540 15904
rect 42432 16031 42484 16040
rect 42432 15997 42441 16031
rect 42441 15997 42475 16031
rect 42475 15997 42484 16031
rect 42432 15988 42484 15997
rect 42524 15988 42576 16040
rect 45008 16031 45060 16040
rect 45008 15997 45017 16031
rect 45017 15997 45051 16031
rect 45051 15997 45060 16031
rect 45008 15988 45060 15997
rect 51908 15988 51960 16040
rect 53012 15988 53064 16040
rect 53196 16031 53248 16040
rect 53196 15997 53205 16031
rect 53205 15997 53239 16031
rect 53239 15997 53248 16031
rect 53196 15988 53248 15997
rect 53472 15988 53524 16040
rect 46572 15920 46624 15972
rect 47400 15920 47452 15972
rect 49792 15920 49844 15972
rect 50712 15920 50764 15972
rect 55680 16031 55732 16040
rect 55680 15997 55689 16031
rect 55689 15997 55723 16031
rect 55723 15997 55732 16031
rect 55680 15988 55732 15997
rect 57888 16031 57940 16040
rect 57888 15997 57897 16031
rect 57897 15997 57931 16031
rect 57931 15997 57940 16031
rect 57888 15988 57940 15997
rect 43352 15852 43404 15904
rect 43444 15895 43496 15904
rect 43444 15861 43453 15895
rect 43453 15861 43487 15895
rect 43487 15861 43496 15895
rect 43444 15852 43496 15861
rect 46388 15895 46440 15904
rect 46388 15861 46397 15895
rect 46397 15861 46431 15895
rect 46431 15861 46440 15895
rect 46388 15852 46440 15861
rect 49056 15852 49108 15904
rect 53472 15852 53524 15904
rect 55220 15895 55272 15904
rect 55220 15861 55229 15895
rect 55229 15861 55263 15895
rect 55263 15861 55272 15895
rect 55220 15852 55272 15861
rect 55864 15852 55916 15904
rect 57980 15852 58032 15904
rect 8172 15750 8224 15802
rect 8236 15750 8288 15802
rect 8300 15750 8352 15802
rect 8364 15750 8416 15802
rect 8428 15750 8480 15802
rect 22616 15750 22668 15802
rect 22680 15750 22732 15802
rect 22744 15750 22796 15802
rect 22808 15750 22860 15802
rect 22872 15750 22924 15802
rect 37060 15750 37112 15802
rect 37124 15750 37176 15802
rect 37188 15750 37240 15802
rect 37252 15750 37304 15802
rect 37316 15750 37368 15802
rect 51504 15750 51556 15802
rect 51568 15750 51620 15802
rect 51632 15750 51684 15802
rect 51696 15750 51748 15802
rect 51760 15750 51812 15802
rect 5448 15648 5500 15700
rect 9680 15648 9732 15700
rect 5816 15512 5868 15564
rect 6552 15512 6604 15564
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 9588 15512 9640 15564
rect 13544 15648 13596 15700
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 14004 15648 14056 15700
rect 14924 15648 14976 15700
rect 15752 15648 15804 15700
rect 18420 15648 18472 15700
rect 18512 15691 18564 15700
rect 18512 15657 18521 15691
rect 18521 15657 18555 15691
rect 18555 15657 18564 15691
rect 18512 15648 18564 15657
rect 19524 15691 19576 15700
rect 19524 15657 19533 15691
rect 19533 15657 19567 15691
rect 19567 15657 19576 15691
rect 19524 15648 19576 15657
rect 21364 15691 21416 15700
rect 21364 15657 21373 15691
rect 21373 15657 21407 15691
rect 21407 15657 21416 15691
rect 21364 15648 21416 15657
rect 21640 15648 21692 15700
rect 27436 15648 27488 15700
rect 14096 15512 14148 15564
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 8024 15444 8076 15496
rect 8576 15444 8628 15496
rect 8944 15487 8996 15496
rect 8944 15453 8953 15487
rect 8953 15453 8987 15487
rect 8987 15453 8996 15487
rect 8944 15444 8996 15453
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 20628 15512 20680 15564
rect 5816 15308 5868 15360
rect 9404 15376 9456 15428
rect 15200 15376 15252 15428
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 9588 15351 9640 15360
rect 9588 15317 9597 15351
rect 9597 15317 9631 15351
rect 9631 15317 9640 15351
rect 9588 15308 9640 15317
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 28080 15691 28132 15700
rect 28080 15657 28089 15691
rect 28089 15657 28123 15691
rect 28123 15657 28132 15691
rect 28080 15648 28132 15657
rect 32680 15648 32732 15700
rect 33140 15648 33192 15700
rect 34428 15648 34480 15700
rect 34704 15648 34756 15700
rect 38108 15648 38160 15700
rect 38200 15691 38252 15700
rect 38200 15657 38209 15691
rect 38209 15657 38243 15691
rect 38243 15657 38252 15691
rect 38200 15648 38252 15657
rect 38476 15648 38528 15700
rect 39028 15648 39080 15700
rect 39396 15648 39448 15700
rect 40316 15648 40368 15700
rect 41420 15691 41472 15700
rect 41420 15657 41429 15691
rect 41429 15657 41463 15691
rect 41463 15657 41472 15691
rect 41420 15648 41472 15657
rect 42432 15648 42484 15700
rect 45008 15648 45060 15700
rect 45928 15648 45980 15700
rect 29644 15580 29696 15632
rect 26240 15512 26292 15564
rect 26700 15555 26752 15564
rect 26700 15521 26709 15555
rect 26709 15521 26743 15555
rect 26743 15521 26752 15555
rect 26700 15512 26752 15521
rect 27988 15512 28040 15564
rect 23204 15444 23256 15496
rect 25688 15444 25740 15496
rect 27252 15444 27304 15496
rect 28264 15376 28316 15428
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 18512 15308 18564 15360
rect 19892 15308 19944 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 23388 15308 23440 15317
rect 26516 15308 26568 15360
rect 28172 15351 28224 15360
rect 28172 15317 28181 15351
rect 28181 15317 28215 15351
rect 28215 15317 28224 15351
rect 28172 15308 28224 15317
rect 28448 15444 28500 15496
rect 30196 15487 30248 15496
rect 29000 15376 29052 15428
rect 30196 15453 30205 15487
rect 30205 15453 30239 15487
rect 30239 15453 30248 15487
rect 30196 15444 30248 15453
rect 29276 15351 29328 15360
rect 29276 15317 29285 15351
rect 29285 15317 29319 15351
rect 29319 15317 29328 15351
rect 29276 15308 29328 15317
rect 31024 15308 31076 15360
rect 35440 15512 35492 15564
rect 36728 15512 36780 15564
rect 33324 15444 33376 15496
rect 37832 15444 37884 15496
rect 38660 15444 38712 15496
rect 47492 15648 47544 15700
rect 47860 15648 47912 15700
rect 47032 15580 47084 15632
rect 48412 15580 48464 15632
rect 49700 15648 49752 15700
rect 51172 15580 51224 15632
rect 42800 15512 42852 15564
rect 41144 15444 41196 15496
rect 44916 15512 44968 15564
rect 49792 15512 49844 15564
rect 50712 15487 50764 15496
rect 50712 15453 50721 15487
rect 50721 15453 50755 15487
rect 50755 15453 50764 15487
rect 50712 15444 50764 15453
rect 53104 15648 53156 15700
rect 56140 15648 56192 15700
rect 51448 15512 51500 15564
rect 51908 15512 51960 15564
rect 52552 15555 52604 15564
rect 52552 15521 52561 15555
rect 52561 15521 52595 15555
rect 52595 15521 52604 15555
rect 52552 15512 52604 15521
rect 53104 15512 53156 15564
rect 34060 15308 34112 15360
rect 35072 15308 35124 15360
rect 35256 15308 35308 15360
rect 36360 15308 36412 15360
rect 40408 15308 40460 15360
rect 52276 15487 52328 15496
rect 52276 15453 52285 15487
rect 52285 15453 52319 15487
rect 52319 15453 52328 15487
rect 52276 15444 52328 15453
rect 52368 15487 52420 15496
rect 52368 15453 52402 15487
rect 52402 15453 52420 15487
rect 52368 15444 52420 15453
rect 53288 15444 53340 15496
rect 55220 15444 55272 15496
rect 56048 15512 56100 15564
rect 42064 15376 42116 15428
rect 51356 15376 51408 15428
rect 58532 15376 58584 15428
rect 43996 15308 44048 15360
rect 47400 15351 47452 15360
rect 47400 15317 47409 15351
rect 47409 15317 47443 15351
rect 47443 15317 47452 15351
rect 47400 15308 47452 15317
rect 51264 15351 51316 15360
rect 51264 15317 51273 15351
rect 51273 15317 51307 15351
rect 51307 15317 51316 15351
rect 51264 15308 51316 15317
rect 52644 15308 52696 15360
rect 54576 15308 54628 15360
rect 55588 15308 55640 15360
rect 55772 15351 55824 15360
rect 55772 15317 55781 15351
rect 55781 15317 55815 15351
rect 55815 15317 55824 15351
rect 55772 15308 55824 15317
rect 57336 15308 57388 15360
rect 57888 15308 57940 15360
rect 15394 15206 15446 15258
rect 15458 15206 15510 15258
rect 15522 15206 15574 15258
rect 15586 15206 15638 15258
rect 15650 15206 15702 15258
rect 29838 15206 29890 15258
rect 29902 15206 29954 15258
rect 29966 15206 30018 15258
rect 30030 15206 30082 15258
rect 30094 15206 30146 15258
rect 44282 15206 44334 15258
rect 44346 15206 44398 15258
rect 44410 15206 44462 15258
rect 44474 15206 44526 15258
rect 44538 15206 44590 15258
rect 58726 15206 58778 15258
rect 58790 15206 58842 15258
rect 58854 15206 58906 15258
rect 58918 15206 58970 15258
rect 58982 15206 59034 15258
rect 5540 15104 5592 15156
rect 4712 14968 4764 15020
rect 6000 15036 6052 15088
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 6460 15036 6512 15088
rect 9864 15104 9916 15156
rect 9588 15036 9640 15088
rect 12624 15104 12676 15156
rect 12716 15104 12768 15156
rect 14188 15104 14240 15156
rect 15108 15147 15160 15156
rect 15108 15113 15117 15147
rect 15117 15113 15151 15147
rect 15151 15113 15160 15147
rect 15108 15104 15160 15113
rect 16856 15104 16908 15156
rect 18696 15104 18748 15156
rect 19156 15104 19208 15156
rect 19524 15104 19576 15156
rect 11244 15036 11296 15088
rect 7748 14943 7800 14952
rect 7748 14909 7782 14943
rect 7782 14909 7800 14943
rect 7748 14900 7800 14909
rect 8760 14968 8812 15020
rect 10876 14968 10928 15020
rect 11060 14968 11112 15020
rect 26700 15147 26752 15156
rect 26700 15113 26709 15147
rect 26709 15113 26743 15147
rect 26743 15113 26752 15147
rect 26700 15104 26752 15113
rect 28264 15147 28316 15156
rect 28264 15113 28273 15147
rect 28273 15113 28307 15147
rect 28307 15113 28316 15147
rect 28264 15104 28316 15113
rect 29000 15147 29052 15156
rect 29000 15113 29009 15147
rect 29009 15113 29043 15147
rect 29043 15113 29052 15147
rect 29000 15104 29052 15113
rect 33508 15104 33560 15156
rect 39580 15104 39632 15156
rect 41604 15104 41656 15156
rect 23388 15036 23440 15088
rect 23664 15036 23716 15088
rect 38200 15036 38252 15088
rect 38384 15036 38436 15088
rect 43352 15104 43404 15156
rect 45100 15104 45152 15156
rect 46296 15036 46348 15088
rect 46480 15036 46532 15088
rect 21732 14968 21784 15020
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 28172 14968 28224 15020
rect 8576 14900 8628 14952
rect 9956 14900 10008 14952
rect 14740 14900 14792 14952
rect 7472 14832 7524 14884
rect 15936 14900 15988 14952
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 8024 14764 8076 14816
rect 9312 14764 9364 14816
rect 13912 14764 13964 14816
rect 25872 14943 25924 14952
rect 25872 14909 25881 14943
rect 25881 14909 25915 14943
rect 25915 14909 25924 14943
rect 25872 14900 25924 14909
rect 28080 14900 28132 14952
rect 36544 14943 36596 14952
rect 36544 14909 36553 14943
rect 36553 14909 36587 14943
rect 36587 14909 36596 14943
rect 36544 14900 36596 14909
rect 18328 14764 18380 14816
rect 18972 14764 19024 14816
rect 20628 14764 20680 14816
rect 23756 14764 23808 14816
rect 24216 14764 24268 14816
rect 26792 14832 26844 14884
rect 41052 14832 41104 14884
rect 47400 14900 47452 14952
rect 50712 15147 50764 15156
rect 50712 15113 50721 15147
rect 50721 15113 50755 15147
rect 50755 15113 50764 15147
rect 50712 15104 50764 15113
rect 52460 15104 52512 15156
rect 53104 15147 53156 15156
rect 53104 15113 53113 15147
rect 53113 15113 53147 15147
rect 53147 15113 53156 15147
rect 53104 15104 53156 15113
rect 55496 15104 55548 15156
rect 52368 14968 52420 15020
rect 55404 14968 55456 15020
rect 57336 15104 57388 15156
rect 58532 15147 58584 15156
rect 58532 15113 58541 15147
rect 58541 15113 58575 15147
rect 58575 15113 58584 15147
rect 58532 15104 58584 15113
rect 56876 15011 56928 15020
rect 56876 14977 56885 15011
rect 56885 14977 56919 15011
rect 56919 14977 56928 15011
rect 56876 14968 56928 14977
rect 49240 14900 49292 14952
rect 51356 14943 51408 14952
rect 51356 14909 51365 14943
rect 51365 14909 51399 14943
rect 51399 14909 51408 14943
rect 51356 14900 51408 14909
rect 51908 14900 51960 14952
rect 53840 14900 53892 14952
rect 55956 14900 56008 14952
rect 56692 14943 56744 14952
rect 56692 14909 56726 14943
rect 56726 14909 56744 14943
rect 56692 14900 56744 14909
rect 57888 14943 57940 14952
rect 57888 14909 57897 14943
rect 57897 14909 57931 14943
rect 57931 14909 57940 14943
rect 57888 14900 57940 14909
rect 56140 14832 56192 14884
rect 56324 14875 56376 14884
rect 56324 14841 56333 14875
rect 56333 14841 56367 14875
rect 56367 14841 56376 14875
rect 56324 14832 56376 14841
rect 25688 14807 25740 14816
rect 25688 14773 25697 14807
rect 25697 14773 25731 14807
rect 25731 14773 25740 14807
rect 25688 14764 25740 14773
rect 26700 14764 26752 14816
rect 33324 14764 33376 14816
rect 34980 14764 35032 14816
rect 36268 14764 36320 14816
rect 37464 14807 37516 14816
rect 37464 14773 37473 14807
rect 37473 14773 37507 14807
rect 37507 14773 37516 14807
rect 37464 14764 37516 14773
rect 38660 14764 38712 14816
rect 39672 14807 39724 14816
rect 39672 14773 39681 14807
rect 39681 14773 39715 14807
rect 39715 14773 39724 14807
rect 39672 14764 39724 14773
rect 42064 14764 42116 14816
rect 44180 14807 44232 14816
rect 44180 14773 44189 14807
rect 44189 14773 44223 14807
rect 44223 14773 44232 14807
rect 44180 14764 44232 14773
rect 44916 14807 44968 14816
rect 44916 14773 44925 14807
rect 44925 14773 44959 14807
rect 44959 14773 44968 14807
rect 44916 14764 44968 14773
rect 46572 14807 46624 14816
rect 46572 14773 46581 14807
rect 46581 14773 46615 14807
rect 46615 14773 46624 14807
rect 46572 14764 46624 14773
rect 46756 14764 46808 14816
rect 49700 14807 49752 14816
rect 49700 14773 49709 14807
rect 49709 14773 49743 14807
rect 49743 14773 49752 14807
rect 49700 14764 49752 14773
rect 52000 14764 52052 14816
rect 55680 14764 55732 14816
rect 56692 14764 56744 14816
rect 57520 14807 57572 14816
rect 57520 14773 57529 14807
rect 57529 14773 57563 14807
rect 57563 14773 57572 14807
rect 57520 14764 57572 14773
rect 8172 14662 8224 14714
rect 8236 14662 8288 14714
rect 8300 14662 8352 14714
rect 8364 14662 8416 14714
rect 8428 14662 8480 14714
rect 22616 14662 22668 14714
rect 22680 14662 22732 14714
rect 22744 14662 22796 14714
rect 22808 14662 22860 14714
rect 22872 14662 22924 14714
rect 37060 14662 37112 14714
rect 37124 14662 37176 14714
rect 37188 14662 37240 14714
rect 37252 14662 37304 14714
rect 37316 14662 37368 14714
rect 51504 14662 51556 14714
rect 51568 14662 51620 14714
rect 51632 14662 51684 14714
rect 51696 14662 51748 14714
rect 51760 14662 51812 14714
rect 4712 14560 4764 14612
rect 6460 14560 6512 14612
rect 7748 14560 7800 14612
rect 8024 14560 8076 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 1952 14356 2004 14408
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 9404 14467 9456 14476
rect 9404 14433 9413 14467
rect 9413 14433 9447 14467
rect 9447 14433 9456 14467
rect 9404 14424 9456 14433
rect 11152 14560 11204 14612
rect 19156 14560 19208 14612
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 18328 14424 18380 14476
rect 19432 14424 19484 14476
rect 23204 14603 23256 14612
rect 23204 14569 23213 14603
rect 23213 14569 23247 14603
rect 23247 14569 23256 14603
rect 23204 14560 23256 14569
rect 25872 14560 25924 14612
rect 29276 14560 29328 14612
rect 31024 14603 31076 14612
rect 31024 14569 31033 14603
rect 31033 14569 31067 14603
rect 31067 14569 31076 14603
rect 31024 14560 31076 14569
rect 31668 14560 31720 14612
rect 34060 14560 34112 14612
rect 41696 14603 41748 14612
rect 41696 14569 41705 14603
rect 41705 14569 41739 14603
rect 41739 14569 41748 14603
rect 41696 14560 41748 14569
rect 44180 14560 44232 14612
rect 26424 14492 26476 14544
rect 21732 14467 21784 14476
rect 21732 14433 21741 14467
rect 21741 14433 21775 14467
rect 21775 14433 21784 14467
rect 21732 14424 21784 14433
rect 8576 14356 8628 14408
rect 12624 14356 12676 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 18052 14356 18104 14408
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 19984 14356 20036 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 22744 14424 22796 14476
rect 26516 14467 26568 14476
rect 26516 14433 26525 14467
rect 26525 14433 26559 14467
rect 26559 14433 26568 14467
rect 26516 14424 26568 14433
rect 31852 14535 31904 14544
rect 31852 14501 31861 14535
rect 31861 14501 31895 14535
rect 31895 14501 31904 14535
rect 31852 14492 31904 14501
rect 34796 14467 34848 14476
rect 34796 14433 34805 14467
rect 34805 14433 34839 14467
rect 34839 14433 34848 14467
rect 34796 14424 34848 14433
rect 35624 14424 35676 14476
rect 39672 14424 39724 14476
rect 24492 14356 24544 14408
rect 24676 14356 24728 14408
rect 5908 14288 5960 14340
rect 7840 14288 7892 14340
rect 22376 14288 22428 14340
rect 23664 14331 23716 14340
rect 23664 14297 23673 14331
rect 23673 14297 23707 14331
rect 23707 14297 23716 14331
rect 23664 14288 23716 14297
rect 23848 14288 23900 14340
rect 25688 14356 25740 14408
rect 25780 14288 25832 14340
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 2872 14220 2924 14229
rect 6184 14220 6236 14272
rect 7472 14220 7524 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 9128 14220 9180 14272
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 14924 14263 14976 14272
rect 14924 14229 14933 14263
rect 14933 14229 14967 14263
rect 14967 14229 14976 14263
rect 14924 14220 14976 14229
rect 16488 14220 16540 14272
rect 18144 14263 18196 14272
rect 18144 14229 18153 14263
rect 18153 14229 18187 14263
rect 18187 14229 18196 14263
rect 18144 14220 18196 14229
rect 18420 14220 18472 14272
rect 19616 14263 19668 14272
rect 19616 14229 19625 14263
rect 19625 14229 19659 14263
rect 19659 14229 19668 14263
rect 19616 14220 19668 14229
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 21456 14220 21508 14229
rect 23020 14220 23072 14272
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 23480 14220 23532 14272
rect 28080 14399 28132 14408
rect 28080 14365 28089 14399
rect 28089 14365 28123 14399
rect 28123 14365 28132 14399
rect 28080 14356 28132 14365
rect 28816 14399 28868 14408
rect 28816 14365 28825 14399
rect 28825 14365 28859 14399
rect 28859 14365 28868 14399
rect 28816 14356 28868 14365
rect 29736 14356 29788 14408
rect 35256 14356 35308 14408
rect 36636 14356 36688 14408
rect 38108 14288 38160 14340
rect 40684 14399 40736 14408
rect 40684 14365 40693 14399
rect 40693 14365 40727 14399
rect 40727 14365 40736 14399
rect 40684 14356 40736 14365
rect 43352 14467 43404 14476
rect 43352 14433 43361 14467
rect 43361 14433 43395 14467
rect 43395 14433 43404 14467
rect 43352 14424 43404 14433
rect 26148 14220 26200 14272
rect 27528 14263 27580 14272
rect 27528 14229 27537 14263
rect 27537 14229 27571 14263
rect 27571 14229 27580 14263
rect 27528 14220 27580 14229
rect 28632 14263 28684 14272
rect 28632 14229 28641 14263
rect 28641 14229 28675 14263
rect 28675 14229 28684 14263
rect 28632 14220 28684 14229
rect 29000 14220 29052 14272
rect 30564 14263 30616 14272
rect 30564 14229 30573 14263
rect 30573 14229 30607 14263
rect 30607 14229 30616 14263
rect 30564 14220 30616 14229
rect 30656 14220 30708 14272
rect 31392 14263 31444 14272
rect 31392 14229 31401 14263
rect 31401 14229 31435 14263
rect 31435 14229 31444 14263
rect 31392 14220 31444 14229
rect 35348 14263 35400 14272
rect 35348 14229 35357 14263
rect 35357 14229 35391 14263
rect 35391 14229 35400 14263
rect 35348 14220 35400 14229
rect 37556 14220 37608 14272
rect 38016 14263 38068 14272
rect 38016 14229 38025 14263
rect 38025 14229 38059 14263
rect 38059 14229 38068 14263
rect 38016 14220 38068 14229
rect 39672 14263 39724 14272
rect 39672 14229 39681 14263
rect 39681 14229 39715 14263
rect 39715 14229 39724 14263
rect 39672 14220 39724 14229
rect 40132 14220 40184 14272
rect 40592 14220 40644 14272
rect 42064 14288 42116 14340
rect 46572 14560 46624 14612
rect 49240 14603 49292 14612
rect 49240 14569 49249 14603
rect 49249 14569 49283 14603
rect 49283 14569 49292 14603
rect 49240 14560 49292 14569
rect 49700 14560 49752 14612
rect 51908 14560 51960 14612
rect 46756 14492 46808 14544
rect 47032 14424 47084 14476
rect 47860 14424 47912 14476
rect 48412 14424 48464 14476
rect 46480 14399 46532 14408
rect 46480 14365 46489 14399
rect 46489 14365 46523 14399
rect 46523 14365 46532 14399
rect 46480 14356 46532 14365
rect 41788 14220 41840 14272
rect 43076 14220 43128 14272
rect 44180 14263 44232 14272
rect 44180 14229 44189 14263
rect 44189 14229 44223 14263
rect 44223 14229 44232 14263
rect 44180 14220 44232 14229
rect 44732 14263 44784 14272
rect 44732 14229 44741 14263
rect 44741 14229 44775 14263
rect 44775 14229 44784 14263
rect 44732 14220 44784 14229
rect 47492 14399 47544 14408
rect 47492 14365 47526 14399
rect 47526 14365 47544 14399
rect 47492 14356 47544 14365
rect 49148 14356 49200 14408
rect 51356 14424 51408 14476
rect 52092 14424 52144 14476
rect 52184 14424 52236 14476
rect 54484 14560 54536 14612
rect 55956 14560 56008 14612
rect 56140 14560 56192 14612
rect 57888 14560 57940 14612
rect 50252 14356 50304 14408
rect 54760 14424 54812 14476
rect 55588 14424 55640 14476
rect 57704 14492 57756 14544
rect 57336 14424 57388 14476
rect 51264 14288 51316 14340
rect 51724 14288 51776 14340
rect 52276 14288 52328 14340
rect 53840 14356 53892 14408
rect 57980 14399 58032 14408
rect 57980 14365 57989 14399
rect 57989 14365 58023 14399
rect 58023 14365 58032 14399
rect 57980 14356 58032 14365
rect 54576 14288 54628 14340
rect 55864 14288 55916 14340
rect 57152 14288 57204 14340
rect 48228 14220 48280 14272
rect 48320 14263 48372 14272
rect 48320 14229 48329 14263
rect 48329 14229 48363 14263
rect 48363 14229 48372 14263
rect 48320 14220 48372 14229
rect 48412 14263 48464 14272
rect 48412 14229 48421 14263
rect 48421 14229 48455 14263
rect 48455 14229 48464 14263
rect 48412 14220 48464 14229
rect 48780 14263 48832 14272
rect 48780 14229 48789 14263
rect 48789 14229 48823 14263
rect 48823 14229 48832 14263
rect 48780 14220 48832 14229
rect 48964 14220 49016 14272
rect 51632 14263 51684 14272
rect 51632 14229 51641 14263
rect 51641 14229 51675 14263
rect 51675 14229 51684 14263
rect 51632 14220 51684 14229
rect 52000 14263 52052 14272
rect 52000 14229 52009 14263
rect 52009 14229 52043 14263
rect 52043 14229 52052 14263
rect 52000 14220 52052 14229
rect 55312 14263 55364 14272
rect 55312 14229 55321 14263
rect 55321 14229 55355 14263
rect 55355 14229 55364 14263
rect 55312 14220 55364 14229
rect 56876 14220 56928 14272
rect 15394 14118 15446 14170
rect 15458 14118 15510 14170
rect 15522 14118 15574 14170
rect 15586 14118 15638 14170
rect 15650 14118 15702 14170
rect 29838 14118 29890 14170
rect 29902 14118 29954 14170
rect 29966 14118 30018 14170
rect 30030 14118 30082 14170
rect 30094 14118 30146 14170
rect 44282 14118 44334 14170
rect 44346 14118 44398 14170
rect 44410 14118 44462 14170
rect 44474 14118 44526 14170
rect 44538 14118 44590 14170
rect 58726 14118 58778 14170
rect 58790 14118 58842 14170
rect 58854 14118 58906 14170
rect 58918 14118 58970 14170
rect 58982 14118 59034 14170
rect 2872 14016 2924 14068
rect 1952 13880 2004 13932
rect 5816 14016 5868 14068
rect 7840 14059 7892 14068
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 11152 14016 11204 14068
rect 12900 14016 12952 14068
rect 14924 14016 14976 14068
rect 18236 14016 18288 14068
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 7472 13880 7524 13932
rect 8024 13880 8076 13932
rect 11428 13880 11480 13932
rect 6460 13855 6512 13864
rect 6460 13821 6469 13855
rect 6469 13821 6503 13855
rect 6503 13821 6512 13855
rect 6460 13812 6512 13821
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 6092 13744 6144 13796
rect 13728 13812 13780 13864
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 16488 13812 16540 13864
rect 18144 13880 18196 13932
rect 18972 14016 19024 14068
rect 19064 14016 19116 14068
rect 19984 14059 20036 14068
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 20812 14016 20864 14068
rect 24584 14016 24636 14068
rect 24676 14016 24728 14068
rect 22744 13948 22796 14000
rect 23112 13948 23164 14000
rect 23480 13948 23532 14000
rect 27528 14016 27580 14068
rect 28080 14016 28132 14068
rect 29000 14016 29052 14068
rect 29276 14016 29328 14068
rect 30564 14016 30616 14068
rect 31024 14016 31076 14068
rect 34796 14016 34848 14068
rect 34980 14059 35032 14068
rect 34980 14025 34989 14059
rect 34989 14025 35023 14059
rect 35023 14025 35032 14059
rect 34980 14016 35032 14025
rect 36084 14016 36136 14068
rect 36544 14016 36596 14068
rect 38016 14016 38068 14068
rect 20168 13880 20220 13932
rect 23572 13880 23624 13932
rect 24584 13880 24636 13932
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 19616 13812 19668 13864
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 23020 13812 23072 13864
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 5448 13719 5500 13728
rect 5448 13685 5457 13719
rect 5457 13685 5491 13719
rect 5491 13685 5500 13719
rect 5448 13676 5500 13685
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 9864 13676 9916 13685
rect 13084 13676 13136 13728
rect 15752 13719 15804 13728
rect 15752 13685 15761 13719
rect 15761 13685 15795 13719
rect 15795 13685 15804 13719
rect 15752 13676 15804 13685
rect 18972 13676 19024 13728
rect 21548 13744 21600 13796
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 23388 13744 23440 13796
rect 23756 13812 23808 13864
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 25228 13812 25280 13864
rect 26148 13880 26200 13932
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 29184 13880 29236 13932
rect 30748 13880 30800 13932
rect 23848 13744 23900 13796
rect 24216 13744 24268 13796
rect 25964 13744 26016 13796
rect 28172 13744 28224 13796
rect 30932 13787 30984 13796
rect 30932 13753 30941 13787
rect 30941 13753 30975 13787
rect 30975 13753 30984 13787
rect 30932 13744 30984 13753
rect 25320 13719 25372 13728
rect 25320 13685 25329 13719
rect 25329 13685 25363 13719
rect 25363 13685 25372 13719
rect 25320 13676 25372 13685
rect 25412 13719 25464 13728
rect 25412 13685 25421 13719
rect 25421 13685 25455 13719
rect 25455 13685 25464 13719
rect 25412 13676 25464 13685
rect 28080 13719 28132 13728
rect 28080 13685 28089 13719
rect 28089 13685 28123 13719
rect 28123 13685 28132 13719
rect 28080 13676 28132 13685
rect 29368 13676 29420 13728
rect 30656 13676 30708 13728
rect 31668 13880 31720 13932
rect 37464 13948 37516 14000
rect 38292 13948 38344 14000
rect 36268 13880 36320 13932
rect 37648 13923 37700 13932
rect 37648 13889 37657 13923
rect 37657 13889 37691 13923
rect 37691 13889 37700 13923
rect 37648 13880 37700 13889
rect 34060 13855 34112 13864
rect 34060 13821 34069 13855
rect 34069 13821 34103 13855
rect 34103 13821 34112 13855
rect 34060 13812 34112 13821
rect 34612 13812 34664 13864
rect 35256 13855 35308 13864
rect 35256 13821 35265 13855
rect 35265 13821 35299 13855
rect 35299 13821 35308 13855
rect 35256 13812 35308 13821
rect 37832 13855 37884 13864
rect 37832 13821 37841 13855
rect 37841 13821 37875 13855
rect 37875 13821 37884 13855
rect 37832 13812 37884 13821
rect 38384 13812 38436 13864
rect 31576 13676 31628 13728
rect 33324 13676 33376 13728
rect 36176 13676 36228 13728
rect 36636 13719 36688 13728
rect 36636 13685 36645 13719
rect 36645 13685 36679 13719
rect 36679 13685 36688 13719
rect 36636 13676 36688 13685
rect 39948 13880 40000 13932
rect 40224 13812 40276 13864
rect 42064 14016 42116 14068
rect 42156 14016 42208 14068
rect 42800 14016 42852 14068
rect 44180 14016 44232 14068
rect 45652 14016 45704 14068
rect 46296 14059 46348 14068
rect 46296 14025 46305 14059
rect 46305 14025 46339 14059
rect 46339 14025 46348 14059
rect 46296 14016 46348 14025
rect 48228 14016 48280 14068
rect 48780 14016 48832 14068
rect 50252 14016 50304 14068
rect 51632 14016 51684 14068
rect 52000 14016 52052 14068
rect 53288 14016 53340 14068
rect 55312 14016 55364 14068
rect 55404 14059 55456 14068
rect 55404 14025 55413 14059
rect 55413 14025 55447 14059
rect 55447 14025 55456 14059
rect 55404 14016 55456 14025
rect 55772 14016 55824 14068
rect 56876 14059 56928 14068
rect 40592 13923 40644 13932
rect 40592 13889 40601 13923
rect 40601 13889 40635 13923
rect 40635 13889 40644 13923
rect 40592 13880 40644 13889
rect 41420 13855 41472 13864
rect 41420 13821 41454 13855
rect 41454 13821 41472 13855
rect 41420 13812 41472 13821
rect 41604 13855 41656 13864
rect 41604 13821 41613 13855
rect 41613 13821 41647 13855
rect 41647 13821 41656 13855
rect 41604 13812 41656 13821
rect 41052 13787 41104 13796
rect 41052 13753 41061 13787
rect 41061 13753 41095 13787
rect 41095 13753 41104 13787
rect 41052 13744 41104 13753
rect 45928 13880 45980 13932
rect 46296 13812 46348 13864
rect 40592 13676 40644 13728
rect 42432 13676 42484 13728
rect 43444 13676 43496 13728
rect 44088 13719 44140 13728
rect 44088 13685 44097 13719
rect 44097 13685 44131 13719
rect 44131 13685 44140 13719
rect 44088 13676 44140 13685
rect 45836 13719 45888 13728
rect 45836 13685 45845 13719
rect 45845 13685 45879 13719
rect 45879 13685 45888 13719
rect 45836 13676 45888 13685
rect 46848 13744 46900 13796
rect 47492 13880 47544 13932
rect 48780 13880 48832 13932
rect 47400 13812 47452 13864
rect 52092 13948 52144 14000
rect 54024 13880 54076 13932
rect 55956 13948 56008 14000
rect 56876 14025 56885 14059
rect 56885 14025 56919 14059
rect 56919 14025 56928 14059
rect 56876 14016 56928 14025
rect 53932 13812 53984 13864
rect 54760 13812 54812 13864
rect 55680 13812 55732 13864
rect 56692 13812 56744 13864
rect 51724 13744 51776 13796
rect 57336 13812 57388 13864
rect 57704 13812 57756 13864
rect 56324 13676 56376 13728
rect 56508 13719 56560 13728
rect 56508 13685 56517 13719
rect 56517 13685 56551 13719
rect 56551 13685 56560 13719
rect 56508 13676 56560 13685
rect 8172 13574 8224 13626
rect 8236 13574 8288 13626
rect 8300 13574 8352 13626
rect 8364 13574 8416 13626
rect 8428 13574 8480 13626
rect 22616 13574 22668 13626
rect 22680 13574 22732 13626
rect 22744 13574 22796 13626
rect 22808 13574 22860 13626
rect 22872 13574 22924 13626
rect 37060 13574 37112 13626
rect 37124 13574 37176 13626
rect 37188 13574 37240 13626
rect 37252 13574 37304 13626
rect 37316 13574 37368 13626
rect 51504 13574 51556 13626
rect 51568 13574 51620 13626
rect 51632 13574 51684 13626
rect 51696 13574 51748 13626
rect 51760 13574 51812 13626
rect 5908 13515 5960 13524
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 6092 13472 6144 13524
rect 7472 13472 7524 13524
rect 1952 13336 2004 13388
rect 5448 13336 5500 13388
rect 8576 13336 8628 13388
rect 11428 13472 11480 13524
rect 12624 13515 12676 13524
rect 12624 13481 12633 13515
rect 12633 13481 12667 13515
rect 12667 13481 12676 13515
rect 12624 13472 12676 13481
rect 13360 13472 13412 13524
rect 18052 13472 18104 13524
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 14096 13379 14148 13388
rect 14096 13345 14105 13379
rect 14105 13345 14139 13379
rect 14139 13345 14148 13379
rect 14096 13336 14148 13345
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 19064 13336 19116 13388
rect 19156 13336 19208 13388
rect 19984 13472 20036 13524
rect 22376 13472 22428 13524
rect 23388 13472 23440 13524
rect 23572 13472 23624 13524
rect 25780 13515 25832 13524
rect 25780 13481 25789 13515
rect 25789 13481 25823 13515
rect 25823 13481 25832 13515
rect 25780 13472 25832 13481
rect 25964 13472 26016 13524
rect 29368 13472 29420 13524
rect 3332 13200 3384 13252
rect 9864 13200 9916 13252
rect 11244 13268 11296 13320
rect 13912 13268 13964 13320
rect 14188 13268 14240 13320
rect 15752 13268 15804 13320
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 17776 13268 17828 13320
rect 4068 13132 4120 13184
rect 9588 13132 9640 13184
rect 12256 13200 12308 13252
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 12164 13132 12216 13184
rect 14464 13200 14516 13252
rect 17592 13200 17644 13252
rect 19892 13379 19944 13388
rect 19892 13345 19901 13379
rect 19901 13345 19935 13379
rect 19935 13345 19944 13379
rect 19892 13336 19944 13345
rect 20444 13379 20496 13388
rect 20444 13345 20453 13379
rect 20453 13345 20487 13379
rect 20487 13345 20496 13379
rect 20444 13336 20496 13345
rect 22468 13336 22520 13388
rect 23112 13379 23164 13388
rect 23112 13345 23121 13379
rect 23121 13345 23155 13379
rect 23155 13345 23164 13379
rect 23112 13336 23164 13345
rect 25412 13336 25464 13388
rect 30932 13472 30984 13524
rect 31852 13404 31904 13456
rect 31392 13336 31444 13388
rect 37556 13472 37608 13524
rect 38108 13515 38160 13524
rect 38108 13481 38117 13515
rect 38117 13481 38151 13515
rect 38151 13481 38160 13515
rect 38108 13472 38160 13481
rect 40684 13472 40736 13524
rect 41328 13472 41380 13524
rect 42064 13515 42116 13524
rect 42064 13481 42073 13515
rect 42073 13481 42107 13515
rect 42107 13481 42116 13515
rect 42064 13472 42116 13481
rect 45928 13515 45980 13524
rect 45928 13481 45937 13515
rect 45937 13481 45971 13515
rect 45971 13481 45980 13515
rect 45928 13472 45980 13481
rect 46296 13515 46348 13524
rect 46296 13481 46305 13515
rect 46305 13481 46339 13515
rect 46339 13481 46348 13515
rect 46296 13472 46348 13481
rect 48780 13515 48832 13524
rect 48780 13481 48789 13515
rect 48789 13481 48823 13515
rect 48823 13481 48832 13515
rect 48780 13472 48832 13481
rect 49148 13515 49200 13524
rect 49148 13481 49157 13515
rect 49157 13481 49191 13515
rect 49191 13481 49200 13515
rect 49148 13472 49200 13481
rect 35072 13336 35124 13388
rect 35624 13379 35676 13388
rect 35624 13345 35633 13379
rect 35633 13345 35667 13379
rect 35667 13345 35676 13379
rect 35624 13336 35676 13345
rect 35716 13336 35768 13388
rect 36084 13336 36136 13388
rect 36728 13336 36780 13388
rect 37648 13336 37700 13388
rect 38292 13379 38344 13388
rect 38292 13345 38301 13379
rect 38301 13345 38335 13379
rect 38335 13345 38344 13379
rect 38292 13336 38344 13345
rect 20168 13311 20220 13320
rect 20168 13277 20177 13311
rect 20177 13277 20211 13311
rect 20211 13277 20220 13311
rect 20168 13268 20220 13277
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 12532 13132 12584 13141
rect 13360 13132 13412 13184
rect 14096 13132 14148 13184
rect 14280 13132 14332 13184
rect 17868 13175 17920 13184
rect 17868 13141 17877 13175
rect 17877 13141 17911 13175
rect 17911 13141 17920 13175
rect 17868 13132 17920 13141
rect 18052 13132 18104 13184
rect 18972 13175 19024 13184
rect 18972 13141 18981 13175
rect 18981 13141 19015 13175
rect 19015 13141 19024 13175
rect 18972 13132 19024 13141
rect 19432 13132 19484 13184
rect 20720 13132 20772 13184
rect 22192 13132 22244 13184
rect 24124 13200 24176 13252
rect 24676 13200 24728 13252
rect 28632 13268 28684 13320
rect 24492 13132 24544 13184
rect 27252 13175 27304 13184
rect 27252 13141 27261 13175
rect 27261 13141 27295 13175
rect 27295 13141 27304 13175
rect 27252 13132 27304 13141
rect 28816 13175 28868 13184
rect 28816 13141 28825 13175
rect 28825 13141 28859 13175
rect 28859 13141 28868 13175
rect 28816 13132 28868 13141
rect 30472 13311 30524 13320
rect 30472 13277 30481 13311
rect 30481 13277 30515 13311
rect 30515 13277 30524 13311
rect 30472 13268 30524 13277
rect 30564 13311 30616 13320
rect 30564 13277 30598 13311
rect 30598 13277 30616 13311
rect 30564 13268 30616 13277
rect 30748 13311 30800 13320
rect 30748 13277 30757 13311
rect 30757 13277 30791 13311
rect 30791 13277 30800 13311
rect 30748 13268 30800 13277
rect 32312 13268 32364 13320
rect 34612 13268 34664 13320
rect 31668 13200 31720 13252
rect 30748 13132 30800 13184
rect 31484 13175 31536 13184
rect 31484 13141 31493 13175
rect 31493 13141 31527 13175
rect 31527 13141 31536 13175
rect 31484 13132 31536 13141
rect 31576 13132 31628 13184
rect 31852 13175 31904 13184
rect 31852 13141 31861 13175
rect 31861 13141 31895 13175
rect 31895 13141 31904 13175
rect 31852 13132 31904 13141
rect 33600 13200 33652 13252
rect 33876 13175 33928 13184
rect 33876 13141 33885 13175
rect 33885 13141 33919 13175
rect 33919 13141 33928 13175
rect 33876 13132 33928 13141
rect 36820 13268 36872 13320
rect 39672 13268 39724 13320
rect 40684 13379 40736 13388
rect 40684 13345 40693 13379
rect 40693 13345 40727 13379
rect 40727 13345 40736 13379
rect 40684 13336 40736 13345
rect 44916 13336 44968 13388
rect 45836 13336 45888 13388
rect 47216 13336 47268 13388
rect 47676 13404 47728 13456
rect 52184 13472 52236 13524
rect 57152 13515 57204 13524
rect 57152 13481 57161 13515
rect 57161 13481 57195 13515
rect 57195 13481 57204 13515
rect 57152 13472 57204 13481
rect 48412 13336 48464 13388
rect 56508 13379 56560 13388
rect 56508 13345 56517 13379
rect 56517 13345 56551 13379
rect 56551 13345 56560 13379
rect 56508 13336 56560 13345
rect 41880 13268 41932 13320
rect 41696 13200 41748 13252
rect 44088 13200 44140 13252
rect 36176 13132 36228 13184
rect 36544 13175 36596 13184
rect 36544 13141 36553 13175
rect 36553 13141 36587 13175
rect 36587 13141 36596 13175
rect 36544 13132 36596 13141
rect 37004 13175 37056 13184
rect 37004 13141 37013 13175
rect 37013 13141 37047 13175
rect 37047 13141 37056 13175
rect 37004 13132 37056 13141
rect 39120 13132 39172 13184
rect 39856 13175 39908 13184
rect 39856 13141 39865 13175
rect 39865 13141 39899 13175
rect 39899 13141 39908 13175
rect 39856 13132 39908 13141
rect 40132 13132 40184 13184
rect 40316 13175 40368 13184
rect 40316 13141 40325 13175
rect 40325 13141 40359 13175
rect 40359 13141 40368 13175
rect 40316 13132 40368 13141
rect 44732 13132 44784 13184
rect 47400 13175 47452 13184
rect 47400 13141 47409 13175
rect 47409 13141 47443 13175
rect 47443 13141 47452 13175
rect 47400 13132 47452 13141
rect 55680 13132 55732 13184
rect 56324 13175 56376 13184
rect 56324 13141 56333 13175
rect 56333 13141 56367 13175
rect 56367 13141 56376 13175
rect 56324 13132 56376 13141
rect 15394 13030 15446 13082
rect 15458 13030 15510 13082
rect 15522 13030 15574 13082
rect 15586 13030 15638 13082
rect 15650 13030 15702 13082
rect 29838 13030 29890 13082
rect 29902 13030 29954 13082
rect 29966 13030 30018 13082
rect 30030 13030 30082 13082
rect 30094 13030 30146 13082
rect 44282 13030 44334 13082
rect 44346 13030 44398 13082
rect 44410 13030 44462 13082
rect 44474 13030 44526 13082
rect 44538 13030 44590 13082
rect 58726 13030 58778 13082
rect 58790 13030 58842 13082
rect 58854 13030 58906 13082
rect 58918 13030 58970 13082
rect 58982 13030 59034 13082
rect 2228 12928 2280 12980
rect 3332 12971 3384 12980
rect 3332 12937 3341 12971
rect 3341 12937 3375 12971
rect 3375 12937 3384 12971
rect 3332 12928 3384 12937
rect 3976 12928 4028 12980
rect 6828 12928 6880 12980
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 9220 12971 9272 12980
rect 9220 12937 9229 12971
rect 9229 12937 9263 12971
rect 9263 12937 9272 12971
rect 9220 12928 9272 12937
rect 11060 12928 11112 12980
rect 11244 12928 11296 12980
rect 4068 12860 4120 12912
rect 7656 12860 7708 12912
rect 3056 12792 3108 12844
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 3424 12656 3476 12708
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 8668 12724 8720 12776
rect 9404 12724 9456 12776
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 12716 12928 12768 12980
rect 12440 12724 12492 12776
rect 14280 12928 14332 12980
rect 14464 12928 14516 12980
rect 17776 12928 17828 12980
rect 18604 12928 18656 12980
rect 19432 12928 19484 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 23940 12928 23992 12980
rect 24216 12928 24268 12980
rect 25320 12928 25372 12980
rect 28172 12928 28224 12980
rect 28816 12928 28868 12980
rect 30472 12928 30524 12980
rect 30564 12928 30616 12980
rect 31484 12928 31536 12980
rect 34060 12928 34112 12980
rect 35348 12928 35400 12980
rect 37004 12928 37056 12980
rect 21456 12860 21508 12912
rect 23112 12860 23164 12912
rect 23388 12860 23440 12912
rect 26332 12860 26384 12912
rect 28080 12860 28132 12912
rect 12532 12656 12584 12708
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 18880 12792 18932 12844
rect 20444 12792 20496 12844
rect 3148 12588 3200 12640
rect 7564 12631 7616 12640
rect 7564 12597 7573 12631
rect 7573 12597 7607 12631
rect 7607 12597 7616 12631
rect 7564 12588 7616 12597
rect 8576 12588 8628 12640
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 14188 12724 14240 12776
rect 14556 12724 14608 12776
rect 13544 12656 13596 12708
rect 15476 12656 15528 12708
rect 17408 12724 17460 12776
rect 17776 12724 17828 12776
rect 17868 12724 17920 12776
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 14740 12631 14792 12640
rect 14740 12597 14749 12631
rect 14749 12597 14783 12631
rect 14783 12597 14792 12631
rect 14740 12588 14792 12597
rect 17132 12631 17184 12640
rect 17132 12597 17141 12631
rect 17141 12597 17175 12631
rect 17175 12597 17184 12631
rect 17132 12588 17184 12597
rect 25136 12792 25188 12844
rect 29092 12835 29144 12844
rect 29092 12801 29101 12835
rect 29101 12801 29135 12835
rect 29135 12801 29144 12835
rect 29092 12792 29144 12801
rect 29184 12835 29236 12844
rect 29184 12801 29193 12835
rect 29193 12801 29227 12835
rect 29227 12801 29236 12835
rect 29184 12792 29236 12801
rect 22376 12767 22428 12776
rect 22376 12733 22385 12767
rect 22385 12733 22419 12767
rect 22419 12733 22428 12767
rect 22376 12724 22428 12733
rect 22192 12588 22244 12640
rect 22468 12588 22520 12640
rect 23480 12588 23532 12640
rect 25044 12724 25096 12776
rect 27252 12767 27304 12776
rect 23848 12656 23900 12708
rect 25504 12588 25556 12640
rect 26516 12588 26568 12640
rect 27252 12733 27261 12767
rect 27261 12733 27295 12767
rect 27295 12733 27304 12767
rect 27252 12724 27304 12733
rect 29276 12767 29328 12776
rect 29276 12733 29285 12767
rect 29285 12733 29319 12767
rect 29319 12733 29328 12767
rect 29276 12724 29328 12733
rect 30196 12835 30248 12844
rect 30196 12801 30205 12835
rect 30205 12801 30239 12835
rect 30239 12801 30248 12835
rect 30196 12792 30248 12801
rect 30288 12724 30340 12776
rect 28816 12656 28868 12708
rect 34336 12903 34388 12912
rect 34336 12869 34345 12903
rect 34345 12869 34379 12903
rect 34379 12869 34388 12903
rect 34336 12860 34388 12869
rect 35072 12903 35124 12912
rect 35072 12869 35081 12903
rect 35081 12869 35115 12903
rect 35115 12869 35124 12903
rect 35072 12860 35124 12869
rect 33968 12792 34020 12844
rect 34244 12792 34296 12844
rect 35716 12835 35768 12844
rect 35716 12801 35725 12835
rect 35725 12801 35759 12835
rect 35759 12801 35768 12835
rect 35716 12792 35768 12801
rect 37556 12792 37608 12844
rect 39856 12928 39908 12980
rect 39948 12971 40000 12980
rect 39948 12937 39957 12971
rect 39957 12937 39991 12971
rect 39991 12937 40000 12971
rect 39948 12928 40000 12937
rect 40316 12928 40368 12980
rect 40684 12928 40736 12980
rect 41696 12928 41748 12980
rect 42432 12928 42484 12980
rect 43076 12971 43128 12980
rect 43076 12937 43085 12971
rect 43085 12937 43119 12971
rect 43119 12937 43128 12971
rect 43076 12928 43128 12937
rect 47768 12928 47820 12980
rect 48044 12928 48096 12980
rect 53288 12971 53340 12980
rect 53288 12937 53297 12971
rect 53297 12937 53331 12971
rect 53331 12937 53340 12971
rect 53288 12928 53340 12937
rect 53380 12928 53432 12980
rect 56232 12928 56284 12980
rect 56692 12928 56744 12980
rect 40224 12835 40276 12844
rect 40224 12801 40233 12835
rect 40233 12801 40267 12835
rect 40267 12801 40276 12835
rect 40224 12792 40276 12801
rect 41788 12792 41840 12844
rect 42064 12792 42116 12844
rect 49608 12792 49660 12844
rect 53196 12835 53248 12844
rect 53196 12801 53205 12835
rect 53205 12801 53239 12835
rect 53239 12801 53248 12835
rect 53196 12792 53248 12801
rect 33508 12656 33560 12708
rect 47952 12724 48004 12776
rect 51172 12724 51224 12776
rect 51356 12724 51408 12776
rect 53012 12724 53064 12776
rect 35164 12656 35216 12708
rect 36728 12656 36780 12708
rect 57796 12724 57848 12776
rect 31484 12631 31536 12640
rect 31484 12597 31493 12631
rect 31493 12597 31527 12631
rect 31527 12597 31536 12631
rect 31484 12588 31536 12597
rect 32772 12631 32824 12640
rect 32772 12597 32781 12631
rect 32781 12597 32815 12631
rect 32815 12597 32824 12631
rect 32772 12588 32824 12597
rect 33140 12631 33192 12640
rect 33140 12597 33149 12631
rect 33149 12597 33183 12631
rect 33183 12597 33192 12631
rect 33140 12588 33192 12597
rect 34428 12588 34480 12640
rect 39120 12631 39172 12640
rect 39120 12597 39129 12631
rect 39129 12597 39163 12631
rect 39163 12597 39172 12631
rect 39120 12588 39172 12597
rect 48872 12631 48924 12640
rect 48872 12597 48881 12631
rect 48881 12597 48915 12631
rect 48915 12597 48924 12631
rect 48872 12588 48924 12597
rect 51080 12588 51132 12640
rect 52368 12631 52420 12640
rect 52368 12597 52377 12631
rect 52377 12597 52411 12631
rect 52411 12597 52420 12631
rect 52368 12588 52420 12597
rect 54116 12631 54168 12640
rect 54116 12597 54125 12631
rect 54125 12597 54159 12631
rect 54159 12597 54168 12631
rect 54116 12588 54168 12597
rect 56692 12588 56744 12640
rect 8172 12486 8224 12538
rect 8236 12486 8288 12538
rect 8300 12486 8352 12538
rect 8364 12486 8416 12538
rect 8428 12486 8480 12538
rect 22616 12486 22668 12538
rect 22680 12486 22732 12538
rect 22744 12486 22796 12538
rect 22808 12486 22860 12538
rect 22872 12486 22924 12538
rect 37060 12486 37112 12538
rect 37124 12486 37176 12538
rect 37188 12486 37240 12538
rect 37252 12486 37304 12538
rect 37316 12486 37368 12538
rect 51504 12486 51556 12538
rect 51568 12486 51620 12538
rect 51632 12486 51684 12538
rect 51696 12486 51748 12538
rect 51760 12486 51812 12538
rect 4160 12384 4212 12436
rect 7012 12427 7064 12436
rect 7012 12393 7021 12427
rect 7021 12393 7055 12427
rect 7055 12393 7064 12427
rect 7012 12384 7064 12393
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 12532 12384 12584 12436
rect 6184 12316 6236 12368
rect 6828 12316 6880 12368
rect 9128 12316 9180 12368
rect 9404 12316 9456 12368
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 17592 12427 17644 12436
rect 17592 12393 17601 12427
rect 17601 12393 17635 12427
rect 17635 12393 17644 12427
rect 17592 12384 17644 12393
rect 18512 12384 18564 12436
rect 19800 12384 19852 12436
rect 22192 12427 22244 12436
rect 22192 12393 22201 12427
rect 22201 12393 22235 12427
rect 22235 12393 22244 12427
rect 22192 12384 22244 12393
rect 22376 12427 22428 12436
rect 22376 12393 22385 12427
rect 22385 12393 22419 12427
rect 22419 12393 22428 12427
rect 22376 12384 22428 12393
rect 24492 12384 24544 12436
rect 26516 12384 26568 12436
rect 29092 12384 29144 12436
rect 17776 12316 17828 12368
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 3608 12180 3660 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 8760 12248 8812 12300
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 12256 12248 12308 12300
rect 12440 12248 12492 12300
rect 17132 12248 17184 12300
rect 21824 12248 21876 12300
rect 24768 12316 24820 12368
rect 23020 12248 23072 12300
rect 25228 12248 25280 12300
rect 25504 12291 25556 12300
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 25596 12291 25648 12300
rect 25596 12257 25605 12291
rect 25605 12257 25639 12291
rect 25639 12257 25648 12291
rect 25596 12248 25648 12257
rect 26332 12316 26384 12368
rect 29276 12316 29328 12368
rect 28816 12291 28868 12300
rect 28816 12257 28825 12291
rect 28825 12257 28859 12291
rect 28859 12257 28868 12291
rect 28816 12248 28868 12257
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 7932 12180 7984 12189
rect 8668 12180 8720 12232
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 3240 12155 3292 12164
rect 3240 12121 3249 12155
rect 3249 12121 3283 12155
rect 3283 12121 3292 12155
rect 3240 12112 3292 12121
rect 3884 12112 3936 12164
rect 4988 12112 5040 12164
rect 8024 12112 8076 12164
rect 8392 12112 8444 12164
rect 9588 12112 9640 12164
rect 15200 12112 15252 12164
rect 16488 12180 16540 12232
rect 17960 12180 18012 12232
rect 21088 12180 21140 12232
rect 23296 12223 23348 12232
rect 23296 12189 23305 12223
rect 23305 12189 23339 12223
rect 23339 12189 23348 12223
rect 23296 12180 23348 12189
rect 30656 12384 30708 12436
rect 30748 12384 30800 12436
rect 31852 12384 31904 12436
rect 33600 12427 33652 12436
rect 33600 12393 33609 12427
rect 33609 12393 33643 12427
rect 33643 12393 33652 12427
rect 33600 12384 33652 12393
rect 33968 12384 34020 12436
rect 40684 12384 40736 12436
rect 47860 12384 47912 12436
rect 49332 12384 49384 12436
rect 31116 12180 31168 12232
rect 20444 12112 20496 12164
rect 23480 12112 23532 12164
rect 24768 12112 24820 12164
rect 26700 12112 26752 12164
rect 32772 12316 32824 12368
rect 34336 12316 34388 12368
rect 36820 12316 36872 12368
rect 41696 12359 41748 12368
rect 41696 12325 41705 12359
rect 41705 12325 41739 12359
rect 41739 12325 41748 12359
rect 41696 12316 41748 12325
rect 42340 12316 42392 12368
rect 33140 12248 33192 12300
rect 33876 12291 33928 12300
rect 33876 12257 33885 12291
rect 33885 12257 33919 12291
rect 33919 12257 33928 12291
rect 33876 12248 33928 12257
rect 35808 12248 35860 12300
rect 41420 12248 41472 12300
rect 47768 12316 47820 12368
rect 34612 12180 34664 12232
rect 35992 12223 36044 12232
rect 35992 12189 36001 12223
rect 36001 12189 36035 12223
rect 36035 12189 36044 12223
rect 35992 12180 36044 12189
rect 36360 12180 36412 12232
rect 37464 12180 37516 12232
rect 42248 12180 42300 12232
rect 42984 12248 43036 12300
rect 45652 12248 45704 12300
rect 51448 12384 51500 12436
rect 52920 12384 52972 12436
rect 53748 12384 53800 12436
rect 57336 12384 57388 12436
rect 58440 12427 58492 12436
rect 58440 12393 58449 12427
rect 58449 12393 58483 12427
rect 58483 12393 58492 12427
rect 58440 12384 58492 12393
rect 45284 12223 45336 12232
rect 45284 12189 45293 12223
rect 45293 12189 45327 12223
rect 45327 12189 45336 12223
rect 45284 12180 45336 12189
rect 46020 12223 46072 12232
rect 46020 12189 46029 12223
rect 46029 12189 46063 12223
rect 46063 12189 46072 12223
rect 46020 12180 46072 12189
rect 45008 12112 45060 12164
rect 48320 12180 48372 12232
rect 48872 12180 48924 12232
rect 49608 12248 49660 12300
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 9220 12044 9272 12096
rect 9864 12044 9916 12096
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 13728 12044 13780 12096
rect 14188 12044 14240 12096
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 21824 12087 21876 12096
rect 21824 12053 21833 12087
rect 21833 12053 21867 12087
rect 21867 12053 21876 12087
rect 21824 12044 21876 12053
rect 24860 12087 24912 12096
rect 24860 12053 24869 12087
rect 24869 12053 24903 12087
rect 24903 12053 24912 12087
rect 24860 12044 24912 12053
rect 25228 12044 25280 12096
rect 26792 12087 26844 12096
rect 26792 12053 26801 12087
rect 26801 12053 26835 12087
rect 26835 12053 26844 12087
rect 26792 12044 26844 12053
rect 30380 12044 30432 12096
rect 31392 12044 31444 12096
rect 35348 12087 35400 12096
rect 35348 12053 35357 12087
rect 35357 12053 35391 12087
rect 35391 12053 35400 12087
rect 35348 12044 35400 12053
rect 36636 12087 36688 12096
rect 36636 12053 36645 12087
rect 36645 12053 36679 12087
rect 36679 12053 36688 12087
rect 36636 12044 36688 12053
rect 39028 12087 39080 12096
rect 39028 12053 39037 12087
rect 39037 12053 39071 12087
rect 39071 12053 39080 12087
rect 39028 12044 39080 12053
rect 42064 12087 42116 12096
rect 42064 12053 42073 12087
rect 42073 12053 42107 12087
rect 42107 12053 42116 12087
rect 42064 12044 42116 12053
rect 42156 12087 42208 12096
rect 42156 12053 42165 12087
rect 42165 12053 42199 12087
rect 42199 12053 42208 12087
rect 42156 12044 42208 12053
rect 43904 12044 43956 12096
rect 45560 12044 45612 12096
rect 46664 12087 46716 12096
rect 46664 12053 46673 12087
rect 46673 12053 46707 12087
rect 46707 12053 46716 12087
rect 46664 12044 46716 12053
rect 46848 12044 46900 12096
rect 47400 12087 47452 12096
rect 47400 12053 47409 12087
rect 47409 12053 47443 12087
rect 47443 12053 47452 12087
rect 47400 12044 47452 12053
rect 47768 12044 47820 12096
rect 48228 12044 48280 12096
rect 48964 12112 49016 12164
rect 53840 12316 53892 12368
rect 51080 12112 51132 12164
rect 54116 12248 54168 12300
rect 54576 12316 54628 12368
rect 55864 12316 55916 12368
rect 57888 12316 57940 12368
rect 49884 12087 49936 12096
rect 49884 12053 49893 12087
rect 49893 12053 49927 12087
rect 49927 12053 49936 12087
rect 49884 12044 49936 12053
rect 50160 12044 50212 12096
rect 52184 12044 52236 12096
rect 54484 12223 54536 12232
rect 54484 12189 54493 12223
rect 54493 12189 54527 12223
rect 54527 12189 54536 12223
rect 54484 12180 54536 12189
rect 55312 12223 55364 12232
rect 55312 12189 55321 12223
rect 55321 12189 55355 12223
rect 55355 12189 55364 12223
rect 55312 12180 55364 12189
rect 56692 12223 56744 12232
rect 56692 12189 56726 12223
rect 56726 12189 56744 12223
rect 56692 12180 56744 12189
rect 54392 12087 54444 12096
rect 54392 12053 54401 12087
rect 54401 12053 54435 12087
rect 54435 12053 54444 12087
rect 54392 12044 54444 12053
rect 55128 12087 55180 12096
rect 55128 12053 55137 12087
rect 55137 12053 55171 12087
rect 55171 12053 55180 12087
rect 55128 12044 55180 12053
rect 55956 12087 56008 12096
rect 55956 12053 55965 12087
rect 55965 12053 55999 12087
rect 55999 12053 56008 12087
rect 55956 12044 56008 12053
rect 56048 12044 56100 12096
rect 57336 12112 57388 12164
rect 58256 12112 58308 12164
rect 57152 12044 57204 12096
rect 57796 12087 57848 12096
rect 57796 12053 57805 12087
rect 57805 12053 57839 12087
rect 57839 12053 57848 12087
rect 57796 12044 57848 12053
rect 15394 11942 15446 11994
rect 15458 11942 15510 11994
rect 15522 11942 15574 11994
rect 15586 11942 15638 11994
rect 15650 11942 15702 11994
rect 29838 11942 29890 11994
rect 29902 11942 29954 11994
rect 29966 11942 30018 11994
rect 30030 11942 30082 11994
rect 30094 11942 30146 11994
rect 44282 11942 44334 11994
rect 44346 11942 44398 11994
rect 44410 11942 44462 11994
rect 44474 11942 44526 11994
rect 44538 11942 44590 11994
rect 58726 11942 58778 11994
rect 58790 11942 58842 11994
rect 58854 11942 58906 11994
rect 58918 11942 58970 11994
rect 58982 11942 59034 11994
rect 3056 11840 3108 11892
rect 3516 11840 3568 11892
rect 3608 11840 3660 11892
rect 3884 11840 3936 11892
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5172 11840 5224 11892
rect 5540 11840 5592 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3332 11704 3384 11756
rect 8576 11840 8628 11892
rect 10416 11883 10468 11892
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 12716 11840 12768 11892
rect 13544 11840 13596 11892
rect 15200 11883 15252 11892
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 16488 11840 16540 11892
rect 19340 11883 19392 11892
rect 19340 11849 19349 11883
rect 19349 11849 19383 11883
rect 19383 11849 19392 11883
rect 19340 11840 19392 11849
rect 7564 11772 7616 11824
rect 9864 11815 9916 11824
rect 9864 11781 9873 11815
rect 9873 11781 9907 11815
rect 9907 11781 9916 11815
rect 9864 11772 9916 11781
rect 12808 11772 12860 11824
rect 16304 11772 16356 11824
rect 17960 11772 18012 11824
rect 20720 11772 20772 11824
rect 7932 11704 7984 11756
rect 4252 11568 4304 11620
rect 8392 11704 8444 11756
rect 14740 11704 14792 11756
rect 23296 11840 23348 11892
rect 24216 11840 24268 11892
rect 24492 11840 24544 11892
rect 22468 11772 22520 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 21640 11704 21692 11756
rect 2872 11500 2924 11552
rect 3056 11500 3108 11552
rect 3608 11500 3660 11552
rect 4620 11500 4672 11552
rect 9128 11636 9180 11688
rect 9404 11636 9456 11688
rect 12440 11636 12492 11688
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 20444 11679 20496 11688
rect 20444 11645 20453 11679
rect 20453 11645 20487 11679
rect 20487 11645 20496 11679
rect 20444 11636 20496 11645
rect 8392 11568 8444 11620
rect 19800 11568 19852 11620
rect 20812 11568 20864 11620
rect 10324 11500 10376 11552
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 19524 11500 19576 11552
rect 23480 11679 23532 11688
rect 23480 11645 23489 11679
rect 23489 11645 23523 11679
rect 23523 11645 23532 11679
rect 23480 11636 23532 11645
rect 24216 11679 24268 11688
rect 24216 11645 24225 11679
rect 24225 11645 24259 11679
rect 24259 11645 24268 11679
rect 24216 11636 24268 11645
rect 24308 11679 24360 11688
rect 24308 11645 24342 11679
rect 24342 11645 24360 11679
rect 24308 11636 24360 11645
rect 24676 11636 24728 11688
rect 24860 11636 24912 11688
rect 25596 11840 25648 11892
rect 26792 11840 26844 11892
rect 29736 11840 29788 11892
rect 30380 11883 30432 11892
rect 30380 11849 30389 11883
rect 30389 11849 30423 11883
rect 30423 11849 30432 11883
rect 30380 11840 30432 11849
rect 31024 11840 31076 11892
rect 31116 11840 31168 11892
rect 32312 11840 32364 11892
rect 35348 11840 35400 11892
rect 35992 11883 36044 11892
rect 35992 11849 36001 11883
rect 36001 11849 36035 11883
rect 36035 11849 36044 11883
rect 35992 11840 36044 11849
rect 26424 11704 26476 11756
rect 28724 11636 28776 11688
rect 34336 11704 34388 11756
rect 42156 11840 42208 11892
rect 36820 11772 36872 11824
rect 38752 11772 38804 11824
rect 40224 11772 40276 11824
rect 36360 11747 36412 11756
rect 36360 11713 36369 11747
rect 36369 11713 36403 11747
rect 36403 11713 36412 11747
rect 36360 11704 36412 11713
rect 40500 11704 40552 11756
rect 42800 11883 42852 11892
rect 42800 11849 42809 11883
rect 42809 11849 42843 11883
rect 42843 11849 42852 11883
rect 42800 11840 42852 11849
rect 43904 11883 43956 11892
rect 43904 11849 43913 11883
rect 43913 11849 43947 11883
rect 43947 11849 43956 11883
rect 43904 11840 43956 11849
rect 45008 11883 45060 11892
rect 45008 11849 45017 11883
rect 45017 11849 45051 11883
rect 45051 11849 45060 11883
rect 45008 11840 45060 11849
rect 45284 11840 45336 11892
rect 45652 11883 45704 11892
rect 45652 11849 45661 11883
rect 45661 11849 45695 11883
rect 45695 11849 45704 11883
rect 46388 11883 46440 11892
rect 45652 11840 45704 11849
rect 46388 11849 46397 11883
rect 46397 11849 46431 11883
rect 46431 11849 46440 11883
rect 46388 11840 46440 11849
rect 47216 11840 47268 11892
rect 47400 11840 47452 11892
rect 49332 11883 49384 11892
rect 49332 11849 49341 11883
rect 49341 11849 49375 11883
rect 49375 11849 49384 11883
rect 49332 11840 49384 11849
rect 49884 11840 49936 11892
rect 43168 11772 43220 11824
rect 24032 11568 24084 11620
rect 34152 11636 34204 11688
rect 34428 11679 34480 11688
rect 34428 11645 34437 11679
rect 34437 11645 34471 11679
rect 34471 11645 34480 11679
rect 34428 11636 34480 11645
rect 25044 11500 25096 11552
rect 35072 11568 35124 11620
rect 36912 11636 36964 11688
rect 39028 11636 39080 11688
rect 40040 11679 40092 11688
rect 40040 11645 40049 11679
rect 40049 11645 40083 11679
rect 40083 11645 40092 11679
rect 40040 11636 40092 11645
rect 28908 11543 28960 11552
rect 28908 11509 28917 11543
rect 28917 11509 28951 11543
rect 28951 11509 28960 11543
rect 28908 11500 28960 11509
rect 29276 11543 29328 11552
rect 29276 11509 29285 11543
rect 29285 11509 29319 11543
rect 29319 11509 29328 11543
rect 29276 11500 29328 11509
rect 32956 11543 33008 11552
rect 32956 11509 32965 11543
rect 32965 11509 32999 11543
rect 32999 11509 33008 11543
rect 32956 11500 33008 11509
rect 33784 11500 33836 11552
rect 33876 11543 33928 11552
rect 33876 11509 33885 11543
rect 33885 11509 33919 11543
rect 33919 11509 33928 11543
rect 33876 11500 33928 11509
rect 34520 11500 34572 11552
rect 35440 11500 35492 11552
rect 36820 11500 36872 11552
rect 37004 11543 37056 11552
rect 37004 11509 37013 11543
rect 37013 11509 37047 11543
rect 37047 11509 37056 11543
rect 37004 11500 37056 11509
rect 39120 11543 39172 11552
rect 39120 11509 39129 11543
rect 39129 11509 39163 11543
rect 39163 11509 39172 11543
rect 39120 11500 39172 11509
rect 39672 11500 39724 11552
rect 40316 11568 40368 11620
rect 42800 11636 42852 11688
rect 42984 11679 43036 11688
rect 42984 11645 42993 11679
rect 42993 11645 43027 11679
rect 43027 11645 43036 11679
rect 42984 11636 43036 11645
rect 43812 11636 43864 11688
rect 47032 11704 47084 11756
rect 47308 11704 47360 11756
rect 50988 11840 51040 11892
rect 51172 11840 51224 11892
rect 52368 11840 52420 11892
rect 53012 11840 53064 11892
rect 54392 11840 54444 11892
rect 55128 11840 55180 11892
rect 51264 11704 51316 11756
rect 47216 11636 47268 11688
rect 47584 11679 47636 11688
rect 47584 11645 47593 11679
rect 47593 11645 47627 11679
rect 47627 11645 47636 11679
rect 47584 11636 47636 11645
rect 53472 11704 53524 11756
rect 53748 11747 53800 11756
rect 53748 11713 53757 11747
rect 53757 11713 53791 11747
rect 53791 11713 53800 11747
rect 53748 11704 53800 11713
rect 53840 11704 53892 11756
rect 52000 11679 52052 11688
rect 52000 11645 52009 11679
rect 52009 11645 52043 11679
rect 52043 11645 52052 11679
rect 52000 11636 52052 11645
rect 52092 11636 52144 11688
rect 53380 11679 53432 11688
rect 53380 11645 53389 11679
rect 53389 11645 53423 11679
rect 53423 11645 53432 11679
rect 53380 11636 53432 11645
rect 55312 11704 55364 11756
rect 57704 11840 57756 11892
rect 56692 11747 56744 11756
rect 56692 11713 56701 11747
rect 56701 11713 56735 11747
rect 56735 11713 56744 11747
rect 56692 11704 56744 11713
rect 56784 11747 56836 11756
rect 56784 11713 56818 11747
rect 56818 11713 56836 11747
rect 56784 11704 56836 11713
rect 55680 11636 55732 11688
rect 40684 11543 40736 11552
rect 40684 11509 40693 11543
rect 40693 11509 40727 11543
rect 40727 11509 40736 11543
rect 40684 11500 40736 11509
rect 41880 11500 41932 11552
rect 42248 11543 42300 11552
rect 42248 11509 42257 11543
rect 42257 11509 42291 11543
rect 42291 11509 42300 11543
rect 42248 11500 42300 11509
rect 42616 11500 42668 11552
rect 42892 11500 42944 11552
rect 43628 11500 43680 11552
rect 46020 11543 46072 11552
rect 46020 11509 46029 11543
rect 46029 11509 46063 11543
rect 46063 11509 46072 11543
rect 46020 11500 46072 11509
rect 46940 11500 46992 11552
rect 47952 11500 48004 11552
rect 49148 11500 49200 11552
rect 49608 11500 49660 11552
rect 51172 11500 51224 11552
rect 52276 11500 52328 11552
rect 52552 11543 52604 11552
rect 52552 11509 52561 11543
rect 52561 11509 52595 11543
rect 52595 11509 52604 11543
rect 52552 11500 52604 11509
rect 56140 11568 56192 11620
rect 55588 11543 55640 11552
rect 55588 11509 55597 11543
rect 55597 11509 55631 11543
rect 55631 11509 55640 11543
rect 55588 11500 55640 11509
rect 57336 11636 57388 11688
rect 57152 11500 57204 11552
rect 57612 11543 57664 11552
rect 57612 11509 57621 11543
rect 57621 11509 57655 11543
rect 57655 11509 57664 11543
rect 57612 11500 57664 11509
rect 8172 11398 8224 11450
rect 8236 11398 8288 11450
rect 8300 11398 8352 11450
rect 8364 11398 8416 11450
rect 8428 11398 8480 11450
rect 22616 11398 22668 11450
rect 22680 11398 22732 11450
rect 22744 11398 22796 11450
rect 22808 11398 22860 11450
rect 22872 11398 22924 11450
rect 37060 11398 37112 11450
rect 37124 11398 37176 11450
rect 37188 11398 37240 11450
rect 37252 11398 37304 11450
rect 37316 11398 37368 11450
rect 51504 11398 51556 11450
rect 51568 11398 51620 11450
rect 51632 11398 51684 11450
rect 51696 11398 51748 11450
rect 51760 11398 51812 11450
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 3240 11296 3292 11348
rect 3976 11339 4028 11348
rect 3976 11305 3985 11339
rect 3985 11305 4019 11339
rect 4019 11305 4028 11339
rect 3976 11296 4028 11305
rect 4160 11296 4212 11348
rect 4620 11296 4672 11348
rect 8024 11296 8076 11348
rect 9128 11296 9180 11348
rect 10324 11339 10376 11348
rect 10324 11305 10333 11339
rect 10333 11305 10367 11339
rect 10367 11305 10376 11339
rect 10324 11296 10376 11305
rect 10416 11296 10468 11348
rect 17316 11296 17368 11348
rect 19340 11296 19392 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 23388 11296 23440 11348
rect 24308 11296 24360 11348
rect 3148 11228 3200 11280
rect 3056 11160 3108 11212
rect 3516 11228 3568 11280
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 3608 11160 3660 11212
rect 3884 11160 3936 11212
rect 4252 11160 4304 11212
rect 3148 11024 3200 11076
rect 3516 11135 3568 11144
rect 3516 11101 3525 11135
rect 3525 11101 3559 11135
rect 3559 11101 3568 11135
rect 3516 11092 3568 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 8392 11203 8444 11212
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 8576 11160 8628 11212
rect 13820 11160 13872 11212
rect 6920 11092 6972 11144
rect 12256 11092 12308 11144
rect 3056 10956 3108 11008
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 7840 11024 7892 11076
rect 8576 11024 8628 11076
rect 10508 11024 10560 11076
rect 12440 11067 12492 11076
rect 12440 11033 12449 11067
rect 12449 11033 12483 11067
rect 12483 11033 12492 11067
rect 12440 11024 12492 11033
rect 13268 11024 13320 11076
rect 4988 10956 5040 11008
rect 7748 10999 7800 11008
rect 7748 10965 7757 10999
rect 7757 10965 7791 10999
rect 7791 10965 7800 10999
rect 7748 10956 7800 10965
rect 8668 10956 8720 11008
rect 9404 10956 9456 11008
rect 11060 10999 11112 11008
rect 11060 10965 11069 10999
rect 11069 10965 11103 10999
rect 11103 10965 11112 10999
rect 11060 10956 11112 10965
rect 12624 10956 12676 11008
rect 15108 11092 15160 11144
rect 15844 11092 15896 11144
rect 20444 11228 20496 11280
rect 23480 11228 23532 11280
rect 18788 11092 18840 11144
rect 23756 11203 23808 11212
rect 23756 11169 23765 11203
rect 23765 11169 23799 11203
rect 23799 11169 23808 11203
rect 23756 11160 23808 11169
rect 29000 11296 29052 11348
rect 29736 11339 29788 11348
rect 29736 11305 29745 11339
rect 29745 11305 29779 11339
rect 29779 11305 29788 11339
rect 29736 11296 29788 11305
rect 33784 11339 33836 11348
rect 33784 11305 33793 11339
rect 33793 11305 33827 11339
rect 33827 11305 33836 11339
rect 33784 11296 33836 11305
rect 33876 11296 33928 11348
rect 36268 11296 36320 11348
rect 37464 11296 37516 11348
rect 35072 11228 35124 11280
rect 34980 11160 35032 11212
rect 37556 11228 37608 11280
rect 35900 11203 35952 11212
rect 35900 11169 35909 11203
rect 35909 11169 35943 11203
rect 35943 11169 35952 11203
rect 35900 11160 35952 11169
rect 36084 11160 36136 11212
rect 36544 11160 36596 11212
rect 39672 11339 39724 11348
rect 39672 11305 39681 11339
rect 39681 11305 39715 11339
rect 39715 11305 39724 11339
rect 39672 11296 39724 11305
rect 40040 11296 40092 11348
rect 40316 11296 40368 11348
rect 40684 11296 40736 11348
rect 40960 11296 41012 11348
rect 38292 11203 38344 11212
rect 38292 11169 38301 11203
rect 38301 11169 38335 11203
rect 38335 11169 38344 11203
rect 38292 11160 38344 11169
rect 40408 11203 40460 11212
rect 40408 11169 40417 11203
rect 40417 11169 40451 11203
rect 40451 11169 40460 11203
rect 40408 11160 40460 11169
rect 24492 11092 24544 11144
rect 14280 10956 14332 11008
rect 14832 10999 14884 11008
rect 14832 10965 14841 10999
rect 14841 10965 14875 10999
rect 14875 10965 14884 10999
rect 14832 10956 14884 10965
rect 15200 10956 15252 11008
rect 21272 11024 21324 11076
rect 23296 11024 23348 11076
rect 25228 11092 25280 11144
rect 27804 11135 27856 11144
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 28632 11092 28684 11144
rect 32496 11092 32548 11144
rect 32956 11092 33008 11144
rect 35072 11092 35124 11144
rect 35624 11135 35676 11144
rect 35624 11101 35633 11135
rect 35633 11101 35667 11135
rect 35667 11101 35676 11135
rect 35624 11092 35676 11101
rect 37464 11135 37516 11144
rect 37464 11101 37473 11135
rect 37473 11101 37507 11135
rect 37507 11101 37516 11135
rect 37464 11092 37516 11101
rect 42800 11339 42852 11348
rect 42800 11305 42809 11339
rect 42809 11305 42843 11339
rect 42843 11305 42852 11339
rect 42800 11296 42852 11305
rect 43812 11296 43864 11348
rect 47584 11296 47636 11348
rect 50160 11296 50212 11348
rect 44088 11228 44140 11280
rect 46848 11228 46900 11280
rect 25688 11024 25740 11076
rect 29000 11024 29052 11076
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 23204 10999 23256 11008
rect 23204 10965 23213 10999
rect 23213 10965 23247 10999
rect 23247 10965 23256 10999
rect 23204 10956 23256 10965
rect 23572 10999 23624 11008
rect 23572 10965 23581 10999
rect 23581 10965 23615 10999
rect 23615 10965 23624 10999
rect 23572 10956 23624 10965
rect 26516 10999 26568 11008
rect 26516 10965 26525 10999
rect 26525 10965 26559 10999
rect 26559 10965 26568 10999
rect 26516 10956 26568 10965
rect 28356 10999 28408 11008
rect 28356 10965 28365 10999
rect 28365 10965 28399 10999
rect 28399 10965 28408 10999
rect 28356 10956 28408 10965
rect 30288 10956 30340 11008
rect 33600 11024 33652 11076
rect 34612 11024 34664 11076
rect 34428 10956 34480 11008
rect 35624 10956 35676 11008
rect 35716 10956 35768 11008
rect 38108 10999 38160 11008
rect 38108 10965 38117 10999
rect 38117 10965 38151 10999
rect 38151 10965 38160 10999
rect 38108 10956 38160 10965
rect 40224 11067 40276 11076
rect 40224 11033 40233 11067
rect 40233 11033 40267 11067
rect 40267 11033 40276 11067
rect 41880 11203 41932 11212
rect 41880 11169 41889 11203
rect 41889 11169 41923 11203
rect 41923 11169 41932 11203
rect 41880 11160 41932 11169
rect 42892 11203 42944 11212
rect 42892 11169 42901 11203
rect 42901 11169 42935 11203
rect 42935 11169 42944 11203
rect 42892 11160 42944 11169
rect 47124 11160 47176 11212
rect 47216 11203 47268 11212
rect 47216 11169 47225 11203
rect 47225 11169 47259 11203
rect 47259 11169 47268 11203
rect 47216 11160 47268 11169
rect 48228 11228 48280 11280
rect 47952 11160 48004 11212
rect 40224 11024 40276 11033
rect 38844 10956 38896 11008
rect 39856 10956 39908 11008
rect 40408 10956 40460 11008
rect 41328 11092 41380 11144
rect 41972 11135 42024 11144
rect 41972 11101 42006 11135
rect 42006 11101 42024 11135
rect 41972 11092 42024 11101
rect 42156 11135 42208 11144
rect 42156 11101 42165 11135
rect 42165 11101 42199 11135
rect 42199 11101 42208 11135
rect 42156 11092 42208 11101
rect 44180 11024 44232 11076
rect 45560 11092 45612 11144
rect 46940 11092 46992 11144
rect 47492 11135 47544 11144
rect 47492 11101 47501 11135
rect 47501 11101 47535 11135
rect 47535 11101 47544 11135
rect 47492 11092 47544 11101
rect 48964 11160 49016 11212
rect 49056 11203 49108 11212
rect 49056 11169 49065 11203
rect 49065 11169 49099 11203
rect 49099 11169 49108 11203
rect 49056 11160 49108 11169
rect 48872 11092 48924 11144
rect 52552 11296 52604 11348
rect 54484 11296 54536 11348
rect 51356 11160 51408 11212
rect 52184 11160 52236 11212
rect 52276 11203 52328 11212
rect 52276 11169 52285 11203
rect 52285 11169 52319 11203
rect 52319 11169 52328 11203
rect 52276 11160 52328 11169
rect 52552 11203 52604 11212
rect 52552 11169 52561 11203
rect 52561 11169 52595 11203
rect 52595 11169 52604 11203
rect 52552 11160 52604 11169
rect 52828 11203 52880 11212
rect 52828 11169 52837 11203
rect 52837 11169 52871 11203
rect 52871 11169 52880 11203
rect 52828 11160 52880 11169
rect 52644 11135 52696 11144
rect 52644 11101 52678 11135
rect 52678 11101 52696 11135
rect 52644 11092 52696 11101
rect 54024 11092 54076 11144
rect 55956 11296 56008 11348
rect 55496 11160 55548 11212
rect 55864 11203 55916 11212
rect 55864 11169 55873 11203
rect 55873 11169 55907 11203
rect 55907 11169 55916 11203
rect 55864 11160 55916 11169
rect 56876 11271 56928 11280
rect 56876 11237 56885 11271
rect 56885 11237 56919 11271
rect 56919 11237 56928 11271
rect 56876 11228 56928 11237
rect 57520 11092 57572 11144
rect 57612 11092 57664 11144
rect 44088 10956 44140 11008
rect 44732 10999 44784 11008
rect 44732 10965 44741 10999
rect 44741 10965 44775 10999
rect 44775 10965 44784 10999
rect 44732 10956 44784 10965
rect 49700 11024 49752 11076
rect 54668 11024 54720 11076
rect 55772 10999 55824 11008
rect 55772 10965 55781 10999
rect 55781 10965 55815 10999
rect 55815 10965 55824 10999
rect 55772 10956 55824 10965
rect 56784 10999 56836 11008
rect 56784 10965 56793 10999
rect 56793 10965 56827 10999
rect 56827 10965 56836 10999
rect 56784 10956 56836 10965
rect 56968 10956 57020 11008
rect 15394 10854 15446 10906
rect 15458 10854 15510 10906
rect 15522 10854 15574 10906
rect 15586 10854 15638 10906
rect 15650 10854 15702 10906
rect 29838 10854 29890 10906
rect 29902 10854 29954 10906
rect 29966 10854 30018 10906
rect 30030 10854 30082 10906
rect 30094 10854 30146 10906
rect 44282 10854 44334 10906
rect 44346 10854 44398 10906
rect 44410 10854 44462 10906
rect 44474 10854 44526 10906
rect 44538 10854 44590 10906
rect 58726 10854 58778 10906
rect 58790 10854 58842 10906
rect 58854 10854 58906 10906
rect 58918 10854 58970 10906
rect 58982 10854 59034 10906
rect 3148 10752 3200 10804
rect 3332 10752 3384 10804
rect 4528 10795 4580 10804
rect 4528 10761 4537 10795
rect 4537 10761 4571 10795
rect 4571 10761 4580 10795
rect 4528 10752 4580 10761
rect 6828 10752 6880 10804
rect 7196 10752 7248 10804
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 8392 10752 8444 10804
rect 8576 10795 8628 10804
rect 8576 10761 8585 10795
rect 8585 10761 8619 10795
rect 8619 10761 8628 10795
rect 8576 10752 8628 10761
rect 11060 10752 11112 10804
rect 11336 10752 11388 10804
rect 11704 10752 11756 10804
rect 12164 10752 12216 10804
rect 8852 10727 8904 10736
rect 2780 10616 2832 10668
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 3608 10616 3660 10668
rect 3332 10548 3384 10600
rect 4988 10616 5040 10668
rect 8852 10693 8861 10727
rect 8861 10693 8895 10727
rect 8895 10693 8904 10727
rect 8852 10684 8904 10693
rect 5448 10616 5500 10668
rect 5816 10659 5868 10668
rect 5816 10625 5829 10659
rect 5829 10625 5868 10659
rect 5816 10616 5868 10625
rect 5264 10480 5316 10532
rect 4068 10412 4120 10464
rect 4988 10412 5040 10464
rect 7748 10616 7800 10668
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 9956 10684 10008 10736
rect 10508 10727 10560 10736
rect 10508 10693 10517 10727
rect 10517 10693 10551 10727
rect 10551 10693 10560 10727
rect 10508 10684 10560 10693
rect 12072 10684 12124 10736
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 14832 10752 14884 10804
rect 12348 10591 12400 10600
rect 12348 10557 12357 10591
rect 12357 10557 12391 10591
rect 12391 10557 12400 10591
rect 12348 10548 12400 10557
rect 13820 10548 13872 10600
rect 15660 10616 15712 10668
rect 16672 10795 16724 10804
rect 16672 10761 16681 10795
rect 16681 10761 16715 10795
rect 16715 10761 16724 10795
rect 16672 10752 16724 10761
rect 18052 10752 18104 10804
rect 20352 10752 20404 10804
rect 21088 10795 21140 10804
rect 21088 10761 21097 10795
rect 21097 10761 21131 10795
rect 21131 10761 21140 10795
rect 21088 10752 21140 10761
rect 22192 10752 22244 10804
rect 29552 10752 29604 10804
rect 30656 10752 30708 10804
rect 31576 10795 31628 10804
rect 31576 10761 31585 10795
rect 31585 10761 31619 10795
rect 31619 10761 31628 10795
rect 31576 10752 31628 10761
rect 34612 10752 34664 10804
rect 34888 10752 34940 10804
rect 35072 10752 35124 10804
rect 36912 10752 36964 10804
rect 37464 10752 37516 10804
rect 38844 10795 38896 10804
rect 38844 10761 38853 10795
rect 38853 10761 38887 10795
rect 38887 10761 38896 10795
rect 38844 10752 38896 10761
rect 40960 10752 41012 10804
rect 41512 10795 41564 10804
rect 41512 10761 41521 10795
rect 41521 10761 41555 10795
rect 41555 10761 41564 10795
rect 41512 10752 41564 10761
rect 42156 10752 42208 10804
rect 43812 10795 43864 10804
rect 43812 10761 43821 10795
rect 43821 10761 43855 10795
rect 43855 10761 43864 10795
rect 43812 10752 43864 10761
rect 44180 10752 44232 10804
rect 47032 10795 47084 10804
rect 47032 10761 47041 10795
rect 47041 10761 47075 10795
rect 47075 10761 47084 10795
rect 47032 10752 47084 10761
rect 47124 10752 47176 10804
rect 16764 10616 16816 10668
rect 31484 10684 31536 10736
rect 17684 10616 17736 10668
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 12256 10480 12308 10532
rect 13544 10480 13596 10532
rect 18236 10616 18288 10668
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 23204 10616 23256 10668
rect 23296 10659 23348 10668
rect 23296 10625 23305 10659
rect 23305 10625 23339 10659
rect 23339 10625 23348 10659
rect 23296 10616 23348 10625
rect 23388 10659 23440 10668
rect 23388 10625 23397 10659
rect 23397 10625 23431 10659
rect 23431 10625 23440 10659
rect 23388 10616 23440 10625
rect 23572 10616 23624 10668
rect 24492 10616 24544 10668
rect 26516 10616 26568 10668
rect 27344 10616 27396 10668
rect 28356 10616 28408 10668
rect 29092 10659 29144 10668
rect 29092 10625 29101 10659
rect 29101 10625 29135 10659
rect 29135 10625 29144 10659
rect 29092 10616 29144 10625
rect 30288 10659 30340 10668
rect 30288 10625 30297 10659
rect 30297 10625 30331 10659
rect 30331 10625 30340 10659
rect 30288 10616 30340 10625
rect 30840 10616 30892 10668
rect 33600 10616 33652 10668
rect 35256 10616 35308 10668
rect 36636 10616 36688 10668
rect 37648 10659 37700 10668
rect 37648 10625 37657 10659
rect 37657 10625 37691 10659
rect 37691 10625 37700 10659
rect 37648 10616 37700 10625
rect 42524 10616 42576 10668
rect 43628 10616 43680 10668
rect 46664 10616 46716 10668
rect 48872 10616 48924 10668
rect 49700 10795 49752 10804
rect 49700 10761 49709 10795
rect 49709 10761 49743 10795
rect 49743 10761 49752 10795
rect 49700 10752 49752 10761
rect 51264 10752 51316 10804
rect 52000 10752 52052 10804
rect 52276 10752 52328 10804
rect 55220 10752 55272 10804
rect 56692 10752 56744 10804
rect 57704 10795 57756 10804
rect 57704 10761 57713 10795
rect 57713 10761 57747 10795
rect 57747 10761 57756 10795
rect 57704 10752 57756 10761
rect 51356 10684 51408 10736
rect 52092 10727 52144 10736
rect 52092 10693 52101 10727
rect 52101 10693 52135 10727
rect 52135 10693 52144 10727
rect 52092 10684 52144 10693
rect 51264 10616 51316 10668
rect 53840 10616 53892 10668
rect 17960 10548 18012 10600
rect 18604 10548 18656 10600
rect 19064 10591 19116 10600
rect 19064 10557 19073 10591
rect 19073 10557 19107 10591
rect 19107 10557 19116 10591
rect 19064 10548 19116 10557
rect 25044 10548 25096 10600
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 25320 10591 25372 10600
rect 25320 10557 25329 10591
rect 25329 10557 25363 10591
rect 25363 10557 25372 10591
rect 25320 10548 25372 10557
rect 8024 10412 8076 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 14096 10412 14148 10464
rect 15016 10412 15068 10464
rect 15844 10412 15896 10464
rect 16580 10412 16632 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18420 10480 18472 10532
rect 25688 10548 25740 10600
rect 20444 10412 20496 10464
rect 26700 10412 26752 10464
rect 28632 10523 28684 10532
rect 28632 10489 28641 10523
rect 28641 10489 28675 10523
rect 28675 10489 28684 10523
rect 29920 10548 29972 10600
rect 28632 10480 28684 10489
rect 28724 10455 28776 10464
rect 28724 10421 28733 10455
rect 28733 10421 28767 10455
rect 28767 10421 28776 10455
rect 28724 10412 28776 10421
rect 30288 10480 30340 10532
rect 30564 10412 30616 10464
rect 32496 10412 32548 10464
rect 34244 10455 34296 10464
rect 34244 10421 34253 10455
rect 34253 10421 34287 10455
rect 34287 10421 34296 10455
rect 34244 10412 34296 10421
rect 34336 10412 34388 10464
rect 36360 10412 36412 10464
rect 43904 10591 43956 10600
rect 43904 10557 43913 10591
rect 43913 10557 43947 10591
rect 43947 10557 43956 10591
rect 43904 10548 43956 10557
rect 42064 10480 42116 10532
rect 38200 10412 38252 10464
rect 40316 10455 40368 10464
rect 40316 10421 40325 10455
rect 40325 10421 40359 10455
rect 40359 10421 40368 10455
rect 40316 10412 40368 10421
rect 42708 10412 42760 10464
rect 44732 10412 44784 10464
rect 47492 10548 47544 10600
rect 52276 10591 52328 10600
rect 52276 10557 52285 10591
rect 52285 10557 52319 10591
rect 52319 10557 52328 10591
rect 52276 10548 52328 10557
rect 52552 10548 52604 10600
rect 56784 10684 56836 10736
rect 57888 10591 57940 10600
rect 57888 10557 57897 10591
rect 57897 10557 57931 10591
rect 57931 10557 57940 10591
rect 57888 10548 57940 10557
rect 52644 10480 52696 10532
rect 55312 10412 55364 10464
rect 55864 10412 55916 10464
rect 8172 10310 8224 10362
rect 8236 10310 8288 10362
rect 8300 10310 8352 10362
rect 8364 10310 8416 10362
rect 8428 10310 8480 10362
rect 22616 10310 22668 10362
rect 22680 10310 22732 10362
rect 22744 10310 22796 10362
rect 22808 10310 22860 10362
rect 22872 10310 22924 10362
rect 37060 10310 37112 10362
rect 37124 10310 37176 10362
rect 37188 10310 37240 10362
rect 37252 10310 37304 10362
rect 37316 10310 37368 10362
rect 51504 10310 51556 10362
rect 51568 10310 51620 10362
rect 51632 10310 51684 10362
rect 51696 10310 51748 10362
rect 51760 10310 51812 10362
rect 3424 10208 3476 10260
rect 4252 10208 4304 10260
rect 5816 10208 5868 10260
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 10784 10208 10836 10260
rect 12164 10208 12216 10260
rect 12348 10208 12400 10260
rect 2780 10072 2832 10124
rect 3332 10072 3384 10124
rect 12072 10140 12124 10192
rect 3148 9979 3200 9988
rect 3148 9945 3157 9979
rect 3157 9945 3191 9979
rect 3191 9945 3200 9979
rect 3148 9936 3200 9945
rect 3608 9936 3660 9988
rect 4068 10004 4120 10056
rect 7288 10004 7340 10056
rect 10416 10072 10468 10124
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 8668 10004 8720 10056
rect 9772 10004 9824 10056
rect 6828 9979 6880 9988
rect 6828 9945 6837 9979
rect 6837 9945 6871 9979
rect 6871 9945 6880 9979
rect 6828 9936 6880 9945
rect 11796 9936 11848 9988
rect 9680 9868 9732 9920
rect 10232 9868 10284 9920
rect 12624 10072 12676 10124
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 14280 10208 14332 10260
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 17316 10208 17368 10260
rect 18052 10208 18104 10260
rect 18236 10208 18288 10260
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 19984 10072 20036 10124
rect 20352 10115 20404 10124
rect 20352 10081 20361 10115
rect 20361 10081 20395 10115
rect 20395 10081 20404 10115
rect 20352 10072 20404 10081
rect 12440 10004 12492 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 14004 10004 14056 10056
rect 15108 10004 15160 10056
rect 13084 9868 13136 9920
rect 13268 9868 13320 9920
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 15200 9936 15252 9988
rect 14832 9868 14884 9920
rect 15844 9936 15896 9988
rect 18972 10004 19024 10056
rect 23756 10140 23808 10192
rect 30012 10140 30064 10192
rect 35900 10208 35952 10260
rect 36268 10208 36320 10260
rect 30288 10072 30340 10124
rect 30564 10115 30616 10124
rect 30564 10081 30598 10115
rect 30598 10081 30616 10115
rect 30564 10072 30616 10081
rect 30748 10115 30800 10124
rect 30748 10081 30757 10115
rect 30757 10081 30791 10115
rect 30791 10081 30800 10115
rect 30748 10072 30800 10081
rect 21548 10047 21600 10056
rect 21548 10013 21557 10047
rect 21557 10013 21591 10047
rect 21591 10013 21600 10047
rect 21548 10004 21600 10013
rect 18236 9936 18288 9988
rect 17592 9868 17644 9920
rect 18052 9868 18104 9920
rect 20352 9936 20404 9988
rect 25320 9936 25372 9988
rect 26424 9936 26476 9988
rect 28908 10004 28960 10056
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 29736 10004 29788 10013
rect 31576 10072 31628 10124
rect 37648 10208 37700 10260
rect 40500 10251 40552 10260
rect 40500 10217 40509 10251
rect 40509 10217 40543 10251
rect 40543 10217 40552 10251
rect 40500 10208 40552 10217
rect 41144 10208 41196 10260
rect 41788 10208 41840 10260
rect 38292 10115 38344 10124
rect 38292 10081 38301 10115
rect 38301 10081 38335 10115
rect 38335 10081 38344 10115
rect 38292 10072 38344 10081
rect 41972 10072 42024 10124
rect 43904 10208 43956 10260
rect 44732 10251 44784 10260
rect 42524 10140 42576 10192
rect 44732 10217 44741 10251
rect 44741 10217 44775 10251
rect 44775 10217 44784 10251
rect 44732 10208 44784 10217
rect 45836 10208 45888 10260
rect 47216 10208 47268 10260
rect 49516 10251 49568 10260
rect 49516 10217 49525 10251
rect 49525 10217 49559 10251
rect 49559 10217 49568 10251
rect 49516 10208 49568 10217
rect 50896 10140 50948 10192
rect 53932 10208 53984 10260
rect 55772 10208 55824 10260
rect 57888 10208 57940 10260
rect 44088 10072 44140 10124
rect 51356 10072 51408 10124
rect 52644 10072 52696 10124
rect 56692 10072 56744 10124
rect 31760 10004 31812 10056
rect 32680 10047 32732 10056
rect 32680 10013 32689 10047
rect 32689 10013 32723 10047
rect 32723 10013 32732 10047
rect 32680 10004 32732 10013
rect 33508 10004 33560 10056
rect 38108 10004 38160 10056
rect 39120 10004 39172 10056
rect 53564 10004 53616 10056
rect 57704 10115 57756 10124
rect 57704 10081 57713 10115
rect 57713 10081 57747 10115
rect 57747 10081 57756 10115
rect 57704 10072 57756 10081
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 22100 9868 22152 9920
rect 23756 9868 23808 9920
rect 26332 9868 26384 9920
rect 27344 9911 27396 9920
rect 27344 9877 27353 9911
rect 27353 9877 27387 9911
rect 27387 9877 27396 9911
rect 27344 9868 27396 9877
rect 29276 9868 29328 9920
rect 30288 9868 30340 9920
rect 31024 9868 31076 9920
rect 31668 9868 31720 9920
rect 33232 9911 33284 9920
rect 33232 9877 33241 9911
rect 33241 9877 33275 9911
rect 33275 9877 33284 9911
rect 33232 9868 33284 9877
rect 33968 9911 34020 9920
rect 33968 9877 33977 9911
rect 33977 9877 34011 9911
rect 34011 9877 34020 9911
rect 33968 9868 34020 9877
rect 34980 9868 35032 9920
rect 35532 9911 35584 9920
rect 35532 9877 35541 9911
rect 35541 9877 35575 9911
rect 35575 9877 35584 9911
rect 35532 9868 35584 9877
rect 37464 9868 37516 9920
rect 38200 9868 38252 9920
rect 41512 9868 41564 9920
rect 41880 9868 41932 9920
rect 48872 9868 48924 9920
rect 49056 9868 49108 9920
rect 50896 9911 50948 9920
rect 50896 9877 50905 9911
rect 50905 9877 50939 9911
rect 50939 9877 50948 9911
rect 50896 9868 50948 9877
rect 50988 9911 51040 9920
rect 50988 9877 50997 9911
rect 50997 9877 51031 9911
rect 51031 9877 51040 9911
rect 50988 9868 51040 9877
rect 52644 9868 52696 9920
rect 56876 9868 56928 9920
rect 56968 9868 57020 9920
rect 57704 9868 57756 9920
rect 15394 9766 15446 9818
rect 15458 9766 15510 9818
rect 15522 9766 15574 9818
rect 15586 9766 15638 9818
rect 15650 9766 15702 9818
rect 29838 9766 29890 9818
rect 29902 9766 29954 9818
rect 29966 9766 30018 9818
rect 30030 9766 30082 9818
rect 30094 9766 30146 9818
rect 44282 9766 44334 9818
rect 44346 9766 44398 9818
rect 44410 9766 44462 9818
rect 44474 9766 44526 9818
rect 44538 9766 44590 9818
rect 58726 9766 58778 9818
rect 58790 9766 58842 9818
rect 58854 9766 58906 9818
rect 58918 9766 58970 9818
rect 58982 9766 59034 9818
rect 3148 9664 3200 9716
rect 3332 9707 3384 9716
rect 3332 9673 3341 9707
rect 3341 9673 3375 9707
rect 3375 9673 3384 9707
rect 3332 9664 3384 9673
rect 8024 9664 8076 9716
rect 10416 9664 10468 9716
rect 6276 9596 6328 9648
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 2780 9460 2832 9512
rect 6368 9528 6420 9580
rect 6000 9435 6052 9444
rect 6000 9401 6009 9435
rect 6009 9401 6043 9435
rect 6043 9401 6052 9435
rect 6000 9392 6052 9401
rect 2964 9324 3016 9376
rect 3608 9324 3660 9376
rect 4712 9324 4764 9376
rect 6736 9392 6788 9444
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7472 9571 7524 9580
rect 7472 9537 7481 9571
rect 7481 9537 7515 9571
rect 7515 9537 7524 9571
rect 7472 9528 7524 9537
rect 9772 9639 9824 9648
rect 9772 9605 9781 9639
rect 9781 9605 9815 9639
rect 9815 9605 9824 9639
rect 9772 9596 9824 9605
rect 11336 9596 11388 9648
rect 13084 9664 13136 9716
rect 13912 9664 13964 9716
rect 17592 9664 17644 9716
rect 20168 9664 20220 9716
rect 29092 9664 29144 9716
rect 29552 9664 29604 9716
rect 30104 9664 30156 9716
rect 31484 9707 31536 9716
rect 31484 9673 31493 9707
rect 31493 9673 31527 9707
rect 31527 9673 31536 9707
rect 31484 9664 31536 9673
rect 32496 9664 32548 9716
rect 32680 9707 32732 9716
rect 32680 9673 32689 9707
rect 32689 9673 32723 9707
rect 32723 9673 32732 9707
rect 32680 9664 32732 9673
rect 33968 9664 34020 9716
rect 40500 9664 40552 9716
rect 40960 9664 41012 9716
rect 6920 9460 6972 9512
rect 8024 9460 8076 9512
rect 11704 9528 11756 9580
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 14004 9596 14056 9648
rect 16028 9596 16080 9648
rect 27068 9596 27120 9648
rect 27344 9596 27396 9648
rect 13728 9528 13780 9580
rect 14648 9528 14700 9580
rect 15752 9528 15804 9580
rect 16764 9528 16816 9580
rect 18052 9528 18104 9580
rect 20444 9528 20496 9580
rect 20720 9528 20772 9580
rect 21272 9528 21324 9580
rect 25780 9528 25832 9580
rect 26516 9528 26568 9580
rect 26700 9528 26752 9580
rect 27712 9528 27764 9580
rect 7196 9324 7248 9376
rect 11428 9460 11480 9512
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 12164 9392 12216 9444
rect 15936 9460 15988 9512
rect 17040 9460 17092 9512
rect 17868 9460 17920 9512
rect 18512 9460 18564 9512
rect 20536 9460 20588 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 20076 9392 20128 9444
rect 24216 9503 24268 9512
rect 24216 9469 24225 9503
rect 24225 9469 24259 9503
rect 24259 9469 24268 9503
rect 24216 9460 24268 9469
rect 24860 9460 24912 9512
rect 25504 9460 25556 9512
rect 26148 9460 26200 9512
rect 26240 9503 26292 9512
rect 26240 9469 26249 9503
rect 26249 9469 26283 9503
rect 26283 9469 26292 9503
rect 26240 9460 26292 9469
rect 26332 9460 26384 9512
rect 27160 9460 27212 9512
rect 28356 9503 28408 9512
rect 28356 9469 28365 9503
rect 28365 9469 28399 9503
rect 28399 9469 28408 9503
rect 28356 9460 28408 9469
rect 23112 9392 23164 9444
rect 28264 9392 28316 9444
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 20536 9324 20588 9376
rect 21640 9324 21692 9376
rect 22100 9324 22152 9376
rect 22468 9367 22520 9376
rect 22468 9333 22477 9367
rect 22477 9333 22511 9367
rect 22511 9333 22520 9367
rect 22468 9324 22520 9333
rect 23388 9367 23440 9376
rect 23388 9333 23397 9367
rect 23397 9333 23431 9367
rect 23431 9333 23440 9367
rect 23388 9324 23440 9333
rect 24032 9367 24084 9376
rect 24032 9333 24041 9367
rect 24041 9333 24075 9367
rect 24075 9333 24084 9367
rect 24032 9324 24084 9333
rect 24308 9324 24360 9376
rect 24768 9367 24820 9376
rect 24768 9333 24777 9367
rect 24777 9333 24811 9367
rect 24811 9333 24820 9367
rect 24768 9324 24820 9333
rect 25964 9324 26016 9376
rect 26516 9324 26568 9376
rect 27160 9367 27212 9376
rect 27160 9333 27169 9367
rect 27169 9333 27203 9367
rect 27203 9333 27212 9367
rect 27160 9324 27212 9333
rect 27804 9367 27856 9376
rect 27804 9333 27813 9367
rect 27813 9333 27847 9367
rect 27847 9333 27856 9367
rect 27804 9324 27856 9333
rect 29368 9528 29420 9580
rect 34152 9596 34204 9648
rect 34428 9596 34480 9648
rect 38752 9596 38804 9648
rect 39304 9596 39356 9648
rect 42524 9596 42576 9648
rect 43996 9596 44048 9648
rect 51264 9664 51316 9716
rect 44916 9639 44968 9648
rect 44916 9605 44925 9639
rect 44925 9605 44959 9639
rect 44959 9605 44968 9639
rect 44916 9596 44968 9605
rect 46388 9596 46440 9648
rect 52276 9664 52328 9716
rect 53840 9664 53892 9716
rect 52736 9639 52788 9648
rect 30656 9528 30708 9580
rect 29000 9324 29052 9376
rect 35440 9528 35492 9580
rect 34152 9460 34204 9512
rect 34336 9503 34388 9512
rect 34336 9469 34345 9503
rect 34345 9469 34379 9503
rect 34379 9469 34388 9503
rect 34336 9460 34388 9469
rect 35992 9503 36044 9512
rect 35992 9469 36001 9503
rect 36001 9469 36035 9503
rect 36035 9469 36044 9503
rect 35992 9460 36044 9469
rect 30288 9324 30340 9376
rect 30380 9324 30432 9376
rect 33324 9392 33376 9444
rect 35532 9392 35584 9444
rect 39764 9571 39816 9580
rect 39764 9537 39773 9571
rect 39773 9537 39807 9571
rect 39807 9537 39816 9571
rect 39764 9528 39816 9537
rect 44640 9528 44692 9580
rect 47676 9528 47728 9580
rect 50988 9528 51040 9580
rect 40408 9503 40460 9512
rect 40408 9469 40417 9503
rect 40417 9469 40451 9503
rect 40451 9469 40460 9503
rect 40408 9460 40460 9469
rect 41144 9503 41196 9512
rect 41144 9469 41153 9503
rect 41153 9469 41187 9503
rect 41187 9469 41196 9503
rect 41144 9460 41196 9469
rect 42432 9503 42484 9512
rect 42432 9469 42441 9503
rect 42441 9469 42475 9503
rect 42475 9469 42484 9503
rect 42432 9460 42484 9469
rect 44180 9460 44232 9512
rect 45468 9503 45520 9512
rect 45468 9469 45477 9503
rect 45477 9469 45511 9503
rect 45511 9469 45520 9503
rect 45468 9460 45520 9469
rect 48044 9503 48096 9512
rect 48044 9469 48053 9503
rect 48053 9469 48087 9503
rect 48087 9469 48096 9503
rect 48044 9460 48096 9469
rect 48780 9503 48832 9512
rect 48780 9469 48789 9503
rect 48789 9469 48823 9503
rect 48823 9469 48832 9503
rect 48780 9460 48832 9469
rect 49884 9460 49936 9512
rect 41328 9392 41380 9444
rect 42800 9392 42852 9444
rect 43260 9392 43312 9444
rect 52736 9605 52745 9639
rect 52745 9605 52779 9639
rect 52779 9605 52788 9639
rect 52736 9596 52788 9605
rect 57980 9596 58032 9648
rect 56140 9503 56192 9512
rect 56140 9469 56149 9503
rect 56149 9469 56183 9503
rect 56183 9469 56192 9503
rect 56140 9460 56192 9469
rect 55864 9392 55916 9444
rect 31760 9367 31812 9376
rect 31760 9333 31769 9367
rect 31769 9333 31803 9367
rect 31803 9333 31812 9367
rect 31760 9324 31812 9333
rect 36544 9367 36596 9376
rect 36544 9333 36553 9367
rect 36553 9333 36587 9367
rect 36587 9333 36596 9367
rect 36544 9324 36596 9333
rect 36820 9367 36872 9376
rect 36820 9333 36829 9367
rect 36829 9333 36863 9367
rect 36863 9333 36872 9367
rect 36820 9324 36872 9333
rect 37740 9367 37792 9376
rect 37740 9333 37749 9367
rect 37749 9333 37783 9367
rect 37783 9333 37792 9367
rect 37740 9324 37792 9333
rect 40132 9324 40184 9376
rect 41236 9324 41288 9376
rect 43076 9367 43128 9376
rect 43076 9333 43085 9367
rect 43085 9333 43119 9367
rect 43119 9333 43128 9367
rect 43076 9324 43128 9333
rect 43812 9324 43864 9376
rect 46296 9324 46348 9376
rect 46664 9324 46716 9376
rect 48136 9324 48188 9376
rect 49332 9367 49384 9376
rect 49332 9333 49341 9367
rect 49341 9333 49375 9367
rect 49375 9333 49384 9367
rect 49332 9324 49384 9333
rect 50068 9367 50120 9376
rect 50068 9333 50077 9367
rect 50077 9333 50111 9367
rect 50111 9333 50120 9367
rect 50068 9324 50120 9333
rect 54576 9324 54628 9376
rect 55220 9367 55272 9376
rect 55220 9333 55229 9367
rect 55229 9333 55263 9367
rect 55263 9333 55272 9367
rect 55220 9324 55272 9333
rect 56784 9367 56836 9376
rect 56784 9333 56793 9367
rect 56793 9333 56827 9367
rect 56827 9333 56836 9367
rect 56784 9324 56836 9333
rect 56876 9324 56928 9376
rect 57060 9367 57112 9376
rect 57060 9333 57069 9367
rect 57069 9333 57103 9367
rect 57103 9333 57112 9367
rect 57060 9324 57112 9333
rect 57428 9367 57480 9376
rect 57428 9333 57437 9367
rect 57437 9333 57471 9367
rect 57471 9333 57480 9367
rect 57428 9324 57480 9333
rect 58072 9367 58124 9376
rect 58072 9333 58081 9367
rect 58081 9333 58115 9367
rect 58115 9333 58124 9367
rect 58072 9324 58124 9333
rect 8172 9222 8224 9274
rect 8236 9222 8288 9274
rect 8300 9222 8352 9274
rect 8364 9222 8416 9274
rect 8428 9222 8480 9274
rect 22616 9222 22668 9274
rect 22680 9222 22732 9274
rect 22744 9222 22796 9274
rect 22808 9222 22860 9274
rect 22872 9222 22924 9274
rect 37060 9222 37112 9274
rect 37124 9222 37176 9274
rect 37188 9222 37240 9274
rect 37252 9222 37304 9274
rect 37316 9222 37368 9274
rect 51504 9222 51556 9274
rect 51568 9222 51620 9274
rect 51632 9222 51684 9274
rect 51696 9222 51748 9274
rect 51760 9222 51812 9274
rect 3516 9120 3568 9172
rect 3700 9120 3752 9172
rect 6368 9120 6420 9172
rect 3608 9052 3660 9104
rect 7104 9120 7156 9172
rect 7288 9120 7340 9172
rect 8484 9120 8536 9172
rect 9496 9120 9548 9172
rect 11152 9120 11204 9172
rect 11520 9120 11572 9172
rect 11796 9163 11848 9172
rect 11796 9129 11805 9163
rect 11805 9129 11839 9163
rect 11839 9129 11848 9163
rect 11796 9120 11848 9129
rect 11980 9120 12032 9172
rect 13728 9120 13780 9172
rect 17776 9120 17828 9172
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 20260 9120 20312 9172
rect 20720 9120 20772 9172
rect 2964 8984 3016 9036
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 4712 8916 4764 8968
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 5908 8984 5960 9036
rect 6736 8984 6788 9036
rect 3148 8780 3200 8832
rect 3884 8780 3936 8832
rect 6092 8848 6144 8900
rect 6184 8891 6236 8900
rect 6184 8857 6193 8891
rect 6193 8857 6227 8891
rect 6227 8857 6236 8891
rect 6184 8848 6236 8857
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9496 8916 9548 8968
rect 10140 8916 10192 8968
rect 11612 8984 11664 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 12348 8984 12400 9036
rect 19800 9095 19852 9104
rect 19800 9061 19809 9095
rect 19809 9061 19843 9095
rect 19843 9061 19852 9095
rect 19800 9052 19852 9061
rect 23388 9120 23440 9172
rect 11428 8916 11480 8968
rect 14648 8916 14700 8968
rect 19708 8916 19760 8968
rect 20720 8916 20772 8968
rect 22468 9052 22520 9104
rect 23112 9052 23164 9104
rect 24768 9052 24820 9104
rect 27344 9120 27396 9172
rect 29368 9163 29420 9172
rect 29368 9129 29377 9163
rect 29377 9129 29411 9163
rect 29411 9129 29420 9163
rect 29368 9120 29420 9129
rect 40408 9120 40460 9172
rect 8300 8848 8352 8900
rect 4712 8780 4764 8832
rect 4988 8780 5040 8832
rect 5632 8780 5684 8832
rect 6552 8780 6604 8832
rect 7840 8780 7892 8832
rect 8024 8780 8076 8832
rect 8576 8780 8628 8832
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 10324 8823 10376 8832
rect 10324 8789 10333 8823
rect 10333 8789 10367 8823
rect 10367 8789 10376 8823
rect 10324 8780 10376 8789
rect 11060 8848 11112 8900
rect 11704 8848 11756 8900
rect 15844 8848 15896 8900
rect 17316 8848 17368 8900
rect 13268 8780 13320 8832
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13820 8780 13872 8832
rect 17224 8780 17276 8832
rect 17868 8780 17920 8832
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 19616 8848 19668 8900
rect 20628 8848 20680 8900
rect 19800 8780 19852 8832
rect 19892 8780 19944 8832
rect 20352 8780 20404 8832
rect 21180 8848 21232 8900
rect 25780 8916 25832 8968
rect 23020 8823 23072 8832
rect 23020 8789 23029 8823
rect 23029 8789 23063 8823
rect 23063 8789 23072 8823
rect 23020 8780 23072 8789
rect 23480 8823 23532 8832
rect 23480 8789 23489 8823
rect 23489 8789 23523 8823
rect 23523 8789 23532 8823
rect 23480 8780 23532 8789
rect 24492 8780 24544 8832
rect 24768 8780 24820 8832
rect 28816 9052 28868 9104
rect 41236 9120 41288 9172
rect 41328 9120 41380 9172
rect 47400 9120 47452 9172
rect 48044 9163 48096 9172
rect 48044 9129 48053 9163
rect 48053 9129 48087 9163
rect 48087 9129 48096 9163
rect 48044 9120 48096 9129
rect 49332 9120 49384 9172
rect 56140 9120 56192 9172
rect 56876 9163 56928 9172
rect 56876 9129 56885 9163
rect 56885 9129 56919 9163
rect 56919 9129 56928 9163
rect 56876 9120 56928 9129
rect 26148 8848 26200 8900
rect 28816 8959 28868 8968
rect 28816 8925 28825 8959
rect 28825 8925 28859 8959
rect 28859 8925 28868 8959
rect 28816 8916 28868 8925
rect 28908 8916 28960 8968
rect 30380 8916 30432 8968
rect 30932 9027 30984 9036
rect 30932 8993 30941 9027
rect 30941 8993 30975 9027
rect 30975 8993 30984 9027
rect 30932 8984 30984 8993
rect 31484 8984 31536 9036
rect 32220 8916 32272 8968
rect 40316 8984 40368 9036
rect 29092 8848 29144 8900
rect 29736 8848 29788 8900
rect 27528 8823 27580 8832
rect 27528 8789 27537 8823
rect 27537 8789 27571 8823
rect 27571 8789 27580 8823
rect 27528 8780 27580 8789
rect 29644 8780 29696 8832
rect 30380 8823 30432 8832
rect 30380 8789 30389 8823
rect 30389 8789 30423 8823
rect 30423 8789 30432 8823
rect 30380 8780 30432 8789
rect 34244 8780 34296 8832
rect 34520 8780 34572 8832
rect 36084 8916 36136 8968
rect 36820 8916 36872 8968
rect 36912 8848 36964 8900
rect 37464 8848 37516 8900
rect 36728 8780 36780 8832
rect 38844 8959 38896 8968
rect 38844 8925 38853 8959
rect 38853 8925 38887 8959
rect 38887 8925 38896 8959
rect 38844 8916 38896 8925
rect 40776 9052 40828 9104
rect 40776 8848 40828 8900
rect 38292 8823 38344 8832
rect 38292 8789 38301 8823
rect 38301 8789 38335 8823
rect 38335 8789 38344 8823
rect 38292 8780 38344 8789
rect 38660 8780 38712 8832
rect 40224 8823 40276 8832
rect 40224 8789 40233 8823
rect 40233 8789 40267 8823
rect 40267 8789 40276 8823
rect 41788 9027 41840 9036
rect 41788 8993 41797 9027
rect 41797 8993 41831 9027
rect 41831 8993 41840 9027
rect 41788 8984 41840 8993
rect 43076 9052 43128 9104
rect 43812 9027 43864 9036
rect 43812 8993 43821 9027
rect 43821 8993 43855 9027
rect 43855 8993 43864 9027
rect 43812 8984 43864 8993
rect 43352 8916 43404 8968
rect 44916 8916 44968 8968
rect 45836 9027 45888 9036
rect 45836 8993 45845 9027
rect 45845 8993 45879 9027
rect 45879 8993 45888 9027
rect 45836 8984 45888 8993
rect 46296 8984 46348 9036
rect 46664 9027 46716 9036
rect 46664 8993 46673 9027
rect 46673 8993 46707 9027
rect 46707 8993 46716 9027
rect 46664 8984 46716 8993
rect 44732 8848 44784 8900
rect 40224 8780 40276 8789
rect 42340 8780 42392 8832
rect 42616 8823 42668 8832
rect 42616 8789 42625 8823
rect 42625 8789 42659 8823
rect 42659 8789 42668 8823
rect 42616 8780 42668 8789
rect 43904 8780 43956 8832
rect 46664 8848 46716 8900
rect 47952 8916 48004 8968
rect 46572 8780 46624 8832
rect 52276 8984 52328 9036
rect 53840 8984 53892 9036
rect 50160 8959 50212 8968
rect 50160 8925 50169 8959
rect 50169 8925 50203 8959
rect 50203 8925 50212 8959
rect 50160 8916 50212 8925
rect 52552 8916 52604 8968
rect 54024 8848 54076 8900
rect 57336 9052 57388 9104
rect 55496 8984 55548 9036
rect 56232 8984 56284 9036
rect 57060 8984 57112 9036
rect 54668 8959 54720 8968
rect 54668 8925 54677 8959
rect 54677 8925 54711 8959
rect 54711 8925 54720 8959
rect 54668 8916 54720 8925
rect 57612 8916 57664 8968
rect 48320 8780 48372 8832
rect 48412 8823 48464 8832
rect 48412 8789 48421 8823
rect 48421 8789 48455 8823
rect 48455 8789 48464 8823
rect 48412 8780 48464 8789
rect 48688 8780 48740 8832
rect 50804 8823 50856 8832
rect 50804 8789 50813 8823
rect 50813 8789 50847 8823
rect 50847 8789 50856 8823
rect 50804 8780 50856 8789
rect 54116 8780 54168 8832
rect 55772 8848 55824 8900
rect 54300 8823 54352 8832
rect 54300 8789 54309 8823
rect 54309 8789 54343 8823
rect 54343 8789 54352 8823
rect 54300 8780 54352 8789
rect 54576 8780 54628 8832
rect 55496 8823 55548 8832
rect 55496 8789 55505 8823
rect 55505 8789 55539 8823
rect 55539 8789 55548 8823
rect 55496 8780 55548 8789
rect 55588 8780 55640 8832
rect 15394 8678 15446 8730
rect 15458 8678 15510 8730
rect 15522 8678 15574 8730
rect 15586 8678 15638 8730
rect 15650 8678 15702 8730
rect 29838 8678 29890 8730
rect 29902 8678 29954 8730
rect 29966 8678 30018 8730
rect 30030 8678 30082 8730
rect 30094 8678 30146 8730
rect 44282 8678 44334 8730
rect 44346 8678 44398 8730
rect 44410 8678 44462 8730
rect 44474 8678 44526 8730
rect 44538 8678 44590 8730
rect 58726 8678 58778 8730
rect 58790 8678 58842 8730
rect 58854 8678 58906 8730
rect 58918 8678 58970 8730
rect 58982 8678 59034 8730
rect 2872 8576 2924 8628
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 4344 8576 4396 8628
rect 5172 8576 5224 8628
rect 6000 8576 6052 8628
rect 7472 8576 7524 8628
rect 7840 8576 7892 8628
rect 4712 8551 4764 8560
rect 4712 8517 4721 8551
rect 4721 8517 4755 8551
rect 4755 8517 4764 8551
rect 4712 8508 4764 8517
rect 5080 8508 5132 8560
rect 8300 8508 8352 8560
rect 8944 8576 8996 8628
rect 10324 8576 10376 8628
rect 11704 8576 11756 8628
rect 8668 8508 8720 8560
rect 4068 8372 4120 8424
rect 3608 8304 3660 8356
rect 4712 8304 4764 8356
rect 6184 8440 6236 8492
rect 6276 8440 6328 8492
rect 6368 8440 6420 8492
rect 6828 8440 6880 8492
rect 7012 8440 7064 8492
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 7196 8372 7248 8424
rect 8576 8440 8628 8492
rect 12992 8508 13044 8560
rect 13452 8576 13504 8628
rect 14556 8576 14608 8628
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 21180 8576 21232 8628
rect 21640 8576 21692 8628
rect 23296 8576 23348 8628
rect 23388 8576 23440 8628
rect 25780 8576 25832 8628
rect 26240 8576 26292 8628
rect 27528 8576 27580 8628
rect 29460 8576 29512 8628
rect 29736 8576 29788 8628
rect 30656 8576 30708 8628
rect 34888 8576 34940 8628
rect 36728 8619 36780 8628
rect 36728 8585 36737 8619
rect 36737 8585 36771 8619
rect 36771 8585 36780 8619
rect 36728 8576 36780 8585
rect 40040 8576 40092 8628
rect 40408 8576 40460 8628
rect 41144 8576 41196 8628
rect 8484 8372 8536 8424
rect 8668 8304 8720 8356
rect 9496 8372 9548 8424
rect 11796 8440 11848 8492
rect 23020 8440 23072 8492
rect 24216 8508 24268 8560
rect 24308 8508 24360 8560
rect 24676 8440 24728 8492
rect 24768 8483 24820 8492
rect 24768 8449 24777 8483
rect 24777 8449 24811 8483
rect 24811 8449 24820 8483
rect 24768 8440 24820 8449
rect 26608 8508 26660 8560
rect 13084 8372 13136 8424
rect 13268 8372 13320 8424
rect 12348 8304 12400 8356
rect 15844 8415 15896 8424
rect 15844 8381 15853 8415
rect 15853 8381 15887 8415
rect 15887 8381 15896 8415
rect 15844 8372 15896 8381
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 17960 8372 18012 8424
rect 18328 8415 18380 8424
rect 18328 8381 18337 8415
rect 18337 8381 18371 8415
rect 18371 8381 18380 8415
rect 18328 8372 18380 8381
rect 19800 8372 19852 8424
rect 19892 8372 19944 8424
rect 21272 8372 21324 8424
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 15936 8304 15988 8356
rect 16396 8304 16448 8356
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 25780 8483 25832 8492
rect 25780 8449 25814 8483
rect 25814 8449 25832 8483
rect 25780 8440 25832 8449
rect 25964 8483 26016 8492
rect 25964 8449 25973 8483
rect 25973 8449 26007 8483
rect 26007 8449 26016 8483
rect 25964 8440 26016 8449
rect 15476 8279 15528 8288
rect 15476 8245 15485 8279
rect 15485 8245 15519 8279
rect 15519 8245 15528 8279
rect 15476 8236 15528 8245
rect 16028 8236 16080 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 20444 8236 20496 8288
rect 21548 8236 21600 8288
rect 24768 8304 24820 8356
rect 25136 8304 25188 8356
rect 26332 8372 26384 8424
rect 33232 8508 33284 8560
rect 34244 8508 34296 8560
rect 29092 8483 29144 8492
rect 29092 8449 29101 8483
rect 29101 8449 29135 8483
rect 29135 8449 29144 8483
rect 29092 8440 29144 8449
rect 29552 8440 29604 8492
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 30288 8372 30340 8424
rect 30380 8415 30432 8424
rect 30380 8381 30389 8415
rect 30389 8381 30423 8415
rect 30423 8381 30432 8415
rect 30380 8372 30432 8381
rect 33416 8440 33468 8492
rect 32128 8415 32180 8424
rect 32128 8381 32137 8415
rect 32137 8381 32171 8415
rect 32171 8381 32180 8415
rect 32128 8372 32180 8381
rect 34428 8415 34480 8424
rect 34428 8381 34437 8415
rect 34437 8381 34471 8415
rect 34471 8381 34480 8415
rect 34428 8372 34480 8381
rect 26608 8347 26660 8356
rect 26608 8313 26617 8347
rect 26617 8313 26651 8347
rect 26651 8313 26660 8347
rect 26608 8304 26660 8313
rect 36544 8440 36596 8492
rect 37740 8440 37792 8492
rect 38660 8440 38712 8492
rect 39396 8508 39448 8560
rect 40132 8440 40184 8492
rect 41420 8508 41472 8560
rect 42616 8576 42668 8628
rect 43904 8576 43956 8628
rect 42156 8508 42208 8560
rect 42524 8440 42576 8492
rect 44824 8576 44876 8628
rect 46480 8576 46532 8628
rect 46572 8576 46624 8628
rect 47400 8576 47452 8628
rect 47216 8372 47268 8424
rect 47860 8576 47912 8628
rect 49884 8576 49936 8628
rect 50804 8576 50856 8628
rect 52276 8576 52328 8628
rect 53472 8619 53524 8628
rect 53472 8585 53481 8619
rect 53481 8585 53515 8619
rect 53515 8585 53524 8619
rect 53472 8576 53524 8585
rect 53840 8576 53892 8628
rect 47584 8483 47636 8492
rect 47584 8449 47593 8483
rect 47593 8449 47627 8483
rect 47627 8449 47636 8483
rect 47584 8440 47636 8449
rect 48688 8440 48740 8492
rect 54208 8508 54260 8560
rect 55772 8508 55824 8560
rect 56784 8576 56836 8628
rect 56876 8576 56928 8628
rect 57336 8619 57388 8628
rect 57336 8585 57345 8619
rect 57345 8585 57379 8619
rect 57379 8585 57388 8619
rect 57336 8576 57388 8585
rect 58072 8576 58124 8628
rect 49424 8440 49476 8492
rect 54392 8440 54444 8492
rect 55956 8483 56008 8492
rect 55956 8449 55965 8483
rect 55965 8449 55999 8483
rect 55999 8449 56008 8483
rect 55956 8440 56008 8449
rect 56048 8440 56100 8492
rect 33508 8279 33560 8288
rect 33508 8245 33517 8279
rect 33517 8245 33551 8279
rect 33551 8245 33560 8279
rect 33508 8236 33560 8245
rect 35348 8236 35400 8288
rect 36820 8236 36872 8288
rect 40776 8236 40828 8288
rect 42432 8304 42484 8356
rect 44180 8304 44232 8356
rect 44548 8304 44600 8356
rect 45468 8236 45520 8288
rect 51356 8372 51408 8424
rect 50252 8236 50304 8288
rect 50620 8236 50672 8288
rect 50712 8279 50764 8288
rect 50712 8245 50721 8279
rect 50721 8245 50755 8279
rect 50755 8245 50764 8279
rect 50712 8236 50764 8245
rect 52184 8279 52236 8288
rect 52184 8245 52193 8279
rect 52193 8245 52227 8279
rect 52227 8245 52236 8279
rect 52184 8236 52236 8245
rect 52276 8236 52328 8288
rect 53932 8372 53984 8424
rect 54116 8372 54168 8424
rect 54576 8372 54628 8424
rect 55036 8415 55088 8424
rect 55036 8381 55070 8415
rect 55070 8381 55088 8415
rect 55036 8372 55088 8381
rect 55404 8372 55456 8424
rect 53012 8279 53064 8288
rect 53012 8245 53021 8279
rect 53021 8245 53055 8279
rect 53055 8245 53064 8279
rect 53012 8236 53064 8245
rect 54668 8347 54720 8356
rect 54668 8313 54677 8347
rect 54677 8313 54711 8347
rect 54711 8313 54720 8347
rect 54668 8304 54720 8313
rect 57520 8304 57572 8356
rect 56324 8236 56376 8288
rect 8172 8134 8224 8186
rect 8236 8134 8288 8186
rect 8300 8134 8352 8186
rect 8364 8134 8416 8186
rect 8428 8134 8480 8186
rect 22616 8134 22668 8186
rect 22680 8134 22732 8186
rect 22744 8134 22796 8186
rect 22808 8134 22860 8186
rect 22872 8134 22924 8186
rect 37060 8134 37112 8186
rect 37124 8134 37176 8186
rect 37188 8134 37240 8186
rect 37252 8134 37304 8186
rect 37316 8134 37368 8186
rect 51504 8134 51556 8186
rect 51568 8134 51620 8186
rect 51632 8134 51684 8186
rect 51696 8134 51748 8186
rect 51760 8134 51812 8186
rect 3792 8032 3844 8084
rect 4068 8032 4120 8084
rect 5908 8032 5960 8084
rect 6092 8032 6144 8084
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 10140 8032 10192 8084
rect 10416 8032 10468 8084
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 15476 8032 15528 8084
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 3056 7871 3108 7880
rect 3056 7837 3066 7871
rect 3066 7837 3100 7871
rect 3100 7837 3108 7871
rect 3056 7828 3108 7837
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 17960 8032 18012 8084
rect 20720 8032 20772 8084
rect 24216 8075 24268 8084
rect 24216 8041 24225 8075
rect 24225 8041 24259 8075
rect 24259 8041 24268 8075
rect 24216 8032 24268 8041
rect 24952 8032 25004 8084
rect 29644 8032 29696 8084
rect 33508 8032 33560 8084
rect 35716 8032 35768 8084
rect 39396 8075 39448 8084
rect 39396 8041 39405 8075
rect 39405 8041 39439 8075
rect 39439 8041 39448 8075
rect 39396 8032 39448 8041
rect 17316 7896 17368 7948
rect 18236 7964 18288 8016
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 5632 7828 5684 7880
rect 5724 7803 5776 7812
rect 5724 7769 5733 7803
rect 5733 7769 5767 7803
rect 5767 7769 5776 7803
rect 5724 7760 5776 7769
rect 6920 7828 6972 7880
rect 7380 7828 7432 7880
rect 9680 7828 9732 7880
rect 10968 7828 11020 7880
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 12256 7828 12308 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 14464 7828 14516 7880
rect 14832 7828 14884 7880
rect 16212 7828 16264 7880
rect 17408 7828 17460 7880
rect 19064 7828 19116 7880
rect 19984 7896 20036 7948
rect 20628 7896 20680 7948
rect 20812 7896 20864 7948
rect 24492 7964 24544 8016
rect 24584 7896 24636 7948
rect 25872 7939 25924 7948
rect 25872 7905 25881 7939
rect 25881 7905 25915 7939
rect 25915 7905 25924 7939
rect 25872 7896 25924 7905
rect 33784 8007 33836 8016
rect 33784 7973 33793 8007
rect 33793 7973 33827 8007
rect 33827 7973 33836 8007
rect 33784 7964 33836 7973
rect 34888 7939 34940 7948
rect 34888 7905 34897 7939
rect 34897 7905 34931 7939
rect 34931 7905 34940 7939
rect 34888 7896 34940 7905
rect 34980 7896 35032 7948
rect 35716 7939 35768 7948
rect 35716 7905 35750 7939
rect 35750 7905 35768 7939
rect 35716 7896 35768 7905
rect 35900 7939 35952 7948
rect 35900 7905 35909 7939
rect 35909 7905 35943 7939
rect 35943 7905 35952 7939
rect 35900 7896 35952 7905
rect 36268 7896 36320 7948
rect 36820 7896 36872 7948
rect 36912 7896 36964 7948
rect 37740 7939 37792 7948
rect 37740 7905 37749 7939
rect 37749 7905 37783 7939
rect 37783 7905 37792 7939
rect 37740 7896 37792 7905
rect 40776 8032 40828 8084
rect 40960 8032 41012 8084
rect 42156 8032 42208 8084
rect 44088 8032 44140 8084
rect 40132 7964 40184 8016
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 22928 7828 22980 7880
rect 26240 7828 26292 7880
rect 28632 7871 28684 7880
rect 28632 7837 28641 7871
rect 28641 7837 28675 7871
rect 28675 7837 28684 7871
rect 28632 7828 28684 7837
rect 29736 7828 29788 7880
rect 32128 7828 32180 7880
rect 33048 7828 33100 7880
rect 33876 7871 33928 7880
rect 33876 7837 33885 7871
rect 33885 7837 33919 7871
rect 33919 7837 33928 7871
rect 33876 7828 33928 7837
rect 34704 7871 34756 7880
rect 34704 7837 34713 7871
rect 34713 7837 34747 7871
rect 34747 7837 34756 7871
rect 34704 7828 34756 7837
rect 40408 7896 40460 7948
rect 40500 7939 40552 7948
rect 40500 7905 40509 7939
rect 40509 7905 40543 7939
rect 40543 7905 40552 7939
rect 40500 7896 40552 7905
rect 41420 7896 41472 7948
rect 44732 7896 44784 7948
rect 44916 7896 44968 7948
rect 45468 7964 45520 8016
rect 45652 8007 45704 8016
rect 45652 7973 45661 8007
rect 45661 7973 45695 8007
rect 45695 7973 45704 8007
rect 45652 7964 45704 7973
rect 45560 7896 45612 7948
rect 47216 8075 47268 8084
rect 47216 8041 47225 8075
rect 47225 8041 47259 8075
rect 47259 8041 47268 8075
rect 47216 8032 47268 8041
rect 48780 8032 48832 8084
rect 50160 8032 50212 8084
rect 51356 8032 51408 8084
rect 54484 8032 54536 8084
rect 55036 8032 55088 8084
rect 55404 8032 55456 8084
rect 56048 8032 56100 8084
rect 56232 8032 56284 8084
rect 56324 8032 56376 8084
rect 46388 7896 46440 7948
rect 49148 7964 49200 8016
rect 49608 7964 49660 8016
rect 49424 7896 49476 7948
rect 40868 7871 40920 7880
rect 40868 7837 40902 7871
rect 40902 7837 40920 7871
rect 40868 7828 40920 7837
rect 41052 7871 41104 7880
rect 41052 7837 41061 7871
rect 41061 7837 41095 7871
rect 41095 7837 41104 7871
rect 41052 7828 41104 7837
rect 45928 7871 45980 7880
rect 45928 7837 45937 7871
rect 45937 7837 45971 7871
rect 45971 7837 45980 7871
rect 45928 7828 45980 7837
rect 47584 7828 47636 7880
rect 50804 7828 50856 7880
rect 52552 7828 52604 7880
rect 53472 7828 53524 7880
rect 55588 7964 55640 8016
rect 57612 8032 57664 8084
rect 54576 7939 54628 7948
rect 54576 7905 54585 7939
rect 54585 7905 54619 7939
rect 54619 7905 54628 7939
rect 54576 7896 54628 7905
rect 55312 7896 55364 7948
rect 55956 7896 56008 7948
rect 56416 7939 56468 7948
rect 56416 7905 56425 7939
rect 56425 7905 56459 7939
rect 56459 7905 56468 7939
rect 56416 7896 56468 7905
rect 55220 7828 55272 7880
rect 57520 7828 57572 7880
rect 9588 7760 9640 7812
rect 11520 7760 11572 7812
rect 6000 7692 6052 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 11244 7692 11296 7744
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 15292 7692 15344 7744
rect 17040 7692 17092 7744
rect 18144 7735 18196 7744
rect 18144 7701 18153 7735
rect 18153 7701 18187 7735
rect 18187 7701 18196 7735
rect 18144 7692 18196 7701
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 19708 7735 19760 7744
rect 19708 7701 19717 7735
rect 19717 7701 19751 7735
rect 19751 7701 19760 7735
rect 19708 7692 19760 7701
rect 19892 7760 19944 7812
rect 22284 7692 22336 7744
rect 23940 7760 23992 7812
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 24492 7692 24544 7744
rect 24860 7735 24912 7744
rect 24860 7701 24869 7735
rect 24869 7701 24903 7735
rect 24903 7701 24912 7735
rect 24860 7692 24912 7701
rect 25596 7692 25648 7744
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 26240 7692 26292 7744
rect 27620 7760 27672 7812
rect 29000 7760 29052 7812
rect 38936 7760 38988 7812
rect 43996 7760 44048 7812
rect 48136 7760 48188 7812
rect 49056 7760 49108 7812
rect 26884 7692 26936 7744
rect 29184 7735 29236 7744
rect 29184 7701 29193 7735
rect 29193 7701 29227 7735
rect 29227 7701 29236 7735
rect 29184 7692 29236 7701
rect 29368 7692 29420 7744
rect 30932 7692 30984 7744
rect 31300 7692 31352 7744
rect 33324 7692 33376 7744
rect 36452 7692 36504 7744
rect 36544 7735 36596 7744
rect 36544 7701 36553 7735
rect 36553 7701 36587 7735
rect 36587 7701 36596 7735
rect 36544 7692 36596 7701
rect 36636 7735 36688 7744
rect 36636 7701 36645 7735
rect 36645 7701 36679 7735
rect 36679 7701 36688 7735
rect 36636 7692 36688 7701
rect 37096 7735 37148 7744
rect 37096 7701 37105 7735
rect 37105 7701 37139 7735
rect 37139 7701 37148 7735
rect 37096 7692 37148 7701
rect 39120 7735 39172 7744
rect 39120 7701 39129 7735
rect 39129 7701 39163 7735
rect 39163 7701 39172 7735
rect 39120 7692 39172 7701
rect 40868 7692 40920 7744
rect 41696 7735 41748 7744
rect 41696 7701 41705 7735
rect 41705 7701 41739 7735
rect 41739 7701 41748 7735
rect 41696 7692 41748 7701
rect 43904 7735 43956 7744
rect 43904 7701 43913 7735
rect 43913 7701 43947 7735
rect 43947 7701 43956 7735
rect 43904 7692 43956 7701
rect 44180 7692 44232 7744
rect 44548 7692 44600 7744
rect 45928 7692 45980 7744
rect 46848 7735 46900 7744
rect 46848 7701 46857 7735
rect 46857 7701 46891 7735
rect 46891 7701 46900 7735
rect 46848 7692 46900 7701
rect 48412 7692 48464 7744
rect 49976 7692 50028 7744
rect 53564 7760 53616 7812
rect 51356 7692 51408 7744
rect 51448 7692 51500 7744
rect 53380 7692 53432 7744
rect 53932 7735 53984 7744
rect 53932 7701 53941 7735
rect 53941 7701 53975 7735
rect 53975 7701 53984 7735
rect 53932 7692 53984 7701
rect 54668 7692 54720 7744
rect 54944 7735 54996 7744
rect 54944 7701 54953 7735
rect 54953 7701 54987 7735
rect 54987 7701 54996 7735
rect 54944 7692 54996 7701
rect 55588 7692 55640 7744
rect 15394 7590 15446 7642
rect 15458 7590 15510 7642
rect 15522 7590 15574 7642
rect 15586 7590 15638 7642
rect 15650 7590 15702 7642
rect 29838 7590 29890 7642
rect 29902 7590 29954 7642
rect 29966 7590 30018 7642
rect 30030 7590 30082 7642
rect 30094 7590 30146 7642
rect 44282 7590 44334 7642
rect 44346 7590 44398 7642
rect 44410 7590 44462 7642
rect 44474 7590 44526 7642
rect 44538 7590 44590 7642
rect 58726 7590 58778 7642
rect 58790 7590 58842 7642
rect 58854 7590 58906 7642
rect 58918 7590 58970 7642
rect 58982 7590 59034 7642
rect 4068 7488 4120 7540
rect 6000 7488 6052 7540
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 7012 7420 7064 7472
rect 7104 7420 7156 7472
rect 8760 7420 8812 7472
rect 9312 7352 9364 7404
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 5724 7284 5776 7336
rect 7840 7284 7892 7336
rect 9496 7284 9548 7336
rect 11336 7352 11388 7404
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 13912 7488 13964 7540
rect 14832 7463 14884 7472
rect 14832 7429 14841 7463
rect 14841 7429 14875 7463
rect 14875 7429 14884 7463
rect 14832 7420 14884 7429
rect 3240 7191 3292 7200
rect 3240 7157 3249 7191
rect 3249 7157 3283 7191
rect 3283 7157 3292 7191
rect 3240 7148 3292 7157
rect 7380 7148 7432 7200
rect 9680 7216 9732 7268
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 9956 7148 10008 7200
rect 10968 7148 11020 7200
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 14832 7284 14884 7336
rect 15292 7395 15344 7404
rect 15292 7361 15326 7395
rect 15326 7361 15344 7395
rect 15292 7352 15344 7361
rect 15568 7352 15620 7404
rect 15844 7352 15896 7404
rect 18328 7420 18380 7472
rect 19708 7488 19760 7540
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 24400 7488 24452 7540
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 24860 7488 24912 7540
rect 25596 7488 25648 7540
rect 25688 7488 25740 7540
rect 27620 7531 27672 7540
rect 27620 7497 27629 7531
rect 27629 7497 27663 7531
rect 27663 7497 27672 7531
rect 27620 7488 27672 7497
rect 28632 7488 28684 7540
rect 29276 7488 29328 7540
rect 33876 7488 33928 7540
rect 34704 7488 34756 7540
rect 35992 7488 36044 7540
rect 36452 7488 36504 7540
rect 37096 7488 37148 7540
rect 37740 7488 37792 7540
rect 38292 7488 38344 7540
rect 38844 7488 38896 7540
rect 12256 7216 12308 7268
rect 14464 7259 14516 7268
rect 14464 7225 14473 7259
rect 14473 7225 14507 7259
rect 14507 7225 14516 7259
rect 18144 7352 18196 7404
rect 19432 7352 19484 7404
rect 23480 7352 23532 7404
rect 24768 7395 24820 7404
rect 24768 7361 24777 7395
rect 24777 7361 24811 7395
rect 24811 7361 24820 7395
rect 24768 7352 24820 7361
rect 25228 7420 25280 7472
rect 24952 7352 25004 7404
rect 25872 7420 25924 7472
rect 26148 7420 26200 7472
rect 26884 7420 26936 7472
rect 34520 7420 34572 7472
rect 33140 7352 33192 7404
rect 33324 7352 33376 7404
rect 14464 7216 14516 7225
rect 14556 7148 14608 7200
rect 17684 7216 17736 7268
rect 16028 7148 16080 7200
rect 16856 7148 16908 7200
rect 21180 7216 21232 7268
rect 29644 7327 29696 7336
rect 29644 7293 29653 7327
rect 29653 7293 29687 7327
rect 29687 7293 29696 7327
rect 29644 7284 29696 7293
rect 30288 7327 30340 7336
rect 30288 7293 30297 7327
rect 30297 7293 30331 7327
rect 30331 7293 30340 7327
rect 30288 7284 30340 7293
rect 32128 7327 32180 7336
rect 32128 7293 32137 7327
rect 32137 7293 32171 7327
rect 32171 7293 32180 7327
rect 32128 7284 32180 7293
rect 33600 7327 33652 7336
rect 33600 7293 33609 7327
rect 33609 7293 33643 7327
rect 33643 7293 33652 7327
rect 33600 7284 33652 7293
rect 34336 7352 34388 7404
rect 34704 7352 34756 7404
rect 35900 7352 35952 7404
rect 33048 7216 33100 7268
rect 40224 7488 40276 7540
rect 41420 7531 41472 7540
rect 41420 7497 41429 7531
rect 41429 7497 41463 7531
rect 41463 7497 41472 7531
rect 41420 7488 41472 7497
rect 42156 7531 42208 7540
rect 42156 7497 42165 7531
rect 42165 7497 42199 7531
rect 42199 7497 42208 7531
rect 42156 7488 42208 7497
rect 43260 7531 43312 7540
rect 43260 7497 43269 7531
rect 43269 7497 43303 7531
rect 43303 7497 43312 7531
rect 43260 7488 43312 7497
rect 40132 7420 40184 7472
rect 41052 7463 41104 7472
rect 41052 7429 41061 7463
rect 41061 7429 41095 7463
rect 41095 7429 41104 7463
rect 41052 7420 41104 7429
rect 38844 7395 38896 7404
rect 38844 7361 38853 7395
rect 38853 7361 38887 7395
rect 38887 7361 38896 7395
rect 38844 7352 38896 7361
rect 43904 7488 43956 7540
rect 43996 7531 44048 7540
rect 43996 7497 44005 7531
rect 44005 7497 44039 7531
rect 44039 7497 44048 7531
rect 43996 7488 44048 7497
rect 44088 7488 44140 7540
rect 44180 7488 44232 7540
rect 44456 7488 44508 7540
rect 44916 7488 44968 7540
rect 45560 7488 45612 7540
rect 46296 7488 46348 7540
rect 47952 7531 48004 7540
rect 47952 7497 47961 7531
rect 47961 7497 47995 7531
rect 47995 7497 48004 7531
rect 47952 7488 48004 7497
rect 48412 7531 48464 7540
rect 48412 7497 48421 7531
rect 48421 7497 48455 7531
rect 48455 7497 48464 7531
rect 48412 7488 48464 7497
rect 45652 7420 45704 7472
rect 45192 7352 45244 7404
rect 37188 7284 37240 7336
rect 39028 7327 39080 7336
rect 39028 7293 39037 7327
rect 39037 7293 39071 7327
rect 39071 7293 39080 7327
rect 39028 7284 39080 7293
rect 39856 7327 39908 7336
rect 39856 7293 39865 7327
rect 39865 7293 39899 7327
rect 39899 7293 39908 7327
rect 39856 7284 39908 7293
rect 40040 7284 40092 7336
rect 46572 7327 46624 7336
rect 46572 7293 46581 7327
rect 46581 7293 46615 7327
rect 46615 7293 46624 7327
rect 46572 7284 46624 7293
rect 20076 7148 20128 7200
rect 20996 7148 21048 7200
rect 21456 7148 21508 7200
rect 24400 7148 24452 7200
rect 24584 7148 24636 7200
rect 25228 7148 25280 7200
rect 29552 7148 29604 7200
rect 29736 7148 29788 7200
rect 32772 7191 32824 7200
rect 32772 7157 32781 7191
rect 32781 7157 32815 7191
rect 32815 7157 32824 7191
rect 32772 7148 32824 7157
rect 34612 7148 34664 7200
rect 35348 7148 35400 7200
rect 36728 7148 36780 7200
rect 38476 7191 38528 7200
rect 38476 7157 38485 7191
rect 38485 7157 38519 7191
rect 38519 7157 38528 7191
rect 38476 7148 38528 7157
rect 40040 7148 40092 7200
rect 41972 7148 42024 7200
rect 42432 7148 42484 7200
rect 42616 7191 42668 7200
rect 42616 7157 42625 7191
rect 42625 7157 42659 7191
rect 42659 7157 42668 7191
rect 42616 7148 42668 7157
rect 48780 7352 48832 7404
rect 50712 7488 50764 7540
rect 50804 7531 50856 7540
rect 50804 7497 50813 7531
rect 50813 7497 50847 7531
rect 50847 7497 50856 7531
rect 50804 7488 50856 7497
rect 52184 7488 52236 7540
rect 52736 7488 52788 7540
rect 53472 7488 53524 7540
rect 53564 7531 53616 7540
rect 53564 7497 53573 7531
rect 53573 7497 53607 7531
rect 53607 7497 53616 7531
rect 53564 7488 53616 7497
rect 53932 7488 53984 7540
rect 54024 7488 54076 7540
rect 54392 7488 54444 7540
rect 55312 7531 55364 7540
rect 55312 7497 55321 7531
rect 55321 7497 55355 7531
rect 55355 7497 55364 7531
rect 55312 7488 55364 7497
rect 55404 7488 55456 7540
rect 56232 7488 56284 7540
rect 56876 7531 56928 7540
rect 56876 7497 56885 7531
rect 56885 7497 56919 7531
rect 56919 7497 56928 7531
rect 56876 7488 56928 7497
rect 57428 7488 57480 7540
rect 57704 7488 57756 7540
rect 50620 7420 50672 7472
rect 49056 7395 49108 7404
rect 49056 7361 49065 7395
rect 49065 7361 49099 7395
rect 49099 7361 49108 7395
rect 49056 7352 49108 7361
rect 49884 7395 49936 7404
rect 49884 7361 49918 7395
rect 49918 7361 49936 7395
rect 49884 7352 49936 7361
rect 48504 7327 48556 7336
rect 48504 7293 48513 7327
rect 48513 7293 48547 7327
rect 48547 7293 48556 7327
rect 48504 7284 48556 7293
rect 50252 7284 50304 7336
rect 48596 7216 48648 7268
rect 49516 7259 49568 7268
rect 49516 7225 49525 7259
rect 49525 7225 49559 7259
rect 49559 7225 49568 7259
rect 49516 7216 49568 7225
rect 50068 7148 50120 7200
rect 50160 7148 50212 7200
rect 51356 7327 51408 7336
rect 51356 7293 51365 7327
rect 51365 7293 51399 7327
rect 51399 7293 51408 7327
rect 51356 7284 51408 7293
rect 53012 7395 53064 7404
rect 53012 7361 53021 7395
rect 53021 7361 53055 7395
rect 53055 7361 53064 7395
rect 53012 7352 53064 7361
rect 54484 7395 54536 7404
rect 54484 7361 54493 7395
rect 54493 7361 54527 7395
rect 54527 7361 54536 7395
rect 54484 7352 54536 7361
rect 55496 7420 55548 7472
rect 55864 7420 55916 7472
rect 58348 7395 58400 7404
rect 58348 7361 58357 7395
rect 58357 7361 58391 7395
rect 58391 7361 58400 7395
rect 58348 7352 58400 7361
rect 56692 7284 56744 7336
rect 50712 7191 50764 7200
rect 50712 7157 50721 7191
rect 50721 7157 50755 7191
rect 50755 7157 50764 7191
rect 50712 7148 50764 7157
rect 52184 7191 52236 7200
rect 52184 7157 52193 7191
rect 52193 7157 52227 7191
rect 52227 7157 52236 7191
rect 52184 7148 52236 7157
rect 55496 7148 55548 7200
rect 56784 7148 56836 7200
rect 57060 7148 57112 7200
rect 57704 7191 57756 7200
rect 57704 7157 57713 7191
rect 57713 7157 57747 7191
rect 57747 7157 57756 7191
rect 57704 7148 57756 7157
rect 58072 7191 58124 7200
rect 58072 7157 58081 7191
rect 58081 7157 58115 7191
rect 58115 7157 58124 7191
rect 58072 7148 58124 7157
rect 8172 7046 8224 7098
rect 8236 7046 8288 7098
rect 8300 7046 8352 7098
rect 8364 7046 8416 7098
rect 8428 7046 8480 7098
rect 22616 7046 22668 7098
rect 22680 7046 22732 7098
rect 22744 7046 22796 7098
rect 22808 7046 22860 7098
rect 22872 7046 22924 7098
rect 37060 7046 37112 7098
rect 37124 7046 37176 7098
rect 37188 7046 37240 7098
rect 37252 7046 37304 7098
rect 37316 7046 37368 7098
rect 51504 7046 51556 7098
rect 51568 7046 51620 7098
rect 51632 7046 51684 7098
rect 51696 7046 51748 7098
rect 51760 7046 51812 7098
rect 9496 6944 9548 6996
rect 1768 6740 1820 6792
rect 3332 6672 3384 6724
rect 5448 6740 5500 6792
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 9956 6876 10008 6928
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 10508 6944 10560 6996
rect 13268 6944 13320 6996
rect 14556 6944 14608 6996
rect 14096 6919 14148 6928
rect 14096 6885 14105 6919
rect 14105 6885 14139 6919
rect 14139 6885 14148 6919
rect 14096 6876 14148 6885
rect 15292 6876 15344 6928
rect 19432 6944 19484 6996
rect 13544 6808 13596 6860
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 15568 6808 15620 6860
rect 20076 6876 20128 6928
rect 22376 6876 22428 6928
rect 30288 6876 30340 6928
rect 32128 6944 32180 6996
rect 33140 6944 33192 6996
rect 33600 6944 33652 6996
rect 35348 6944 35400 6996
rect 35900 6944 35952 6996
rect 37740 6987 37792 6996
rect 37740 6953 37749 6987
rect 37749 6953 37783 6987
rect 37783 6953 37792 6987
rect 37740 6944 37792 6953
rect 38844 6944 38896 6996
rect 40500 6944 40552 6996
rect 40684 6944 40736 6996
rect 40960 6944 41012 6996
rect 44456 6944 44508 6996
rect 46572 6944 46624 6996
rect 48320 6944 48372 6996
rect 48596 6987 48648 6996
rect 48596 6953 48605 6987
rect 48605 6953 48639 6987
rect 48639 6953 48648 6987
rect 48596 6944 48648 6953
rect 49608 6944 49660 6996
rect 50252 6944 50304 6996
rect 16028 6851 16080 6860
rect 16028 6817 16062 6851
rect 16062 6817 16080 6851
rect 16028 6808 16080 6817
rect 16212 6851 16264 6860
rect 16212 6817 16221 6851
rect 16221 6817 16255 6851
rect 16255 6817 16264 6851
rect 16212 6808 16264 6817
rect 16856 6808 16908 6860
rect 18144 6808 18196 6860
rect 18972 6808 19024 6860
rect 19248 6851 19300 6860
rect 19248 6817 19257 6851
rect 19257 6817 19291 6851
rect 19291 6817 19300 6851
rect 19248 6808 19300 6817
rect 19984 6808 20036 6860
rect 21824 6808 21876 6860
rect 23388 6808 23440 6860
rect 25044 6851 25096 6860
rect 25044 6817 25053 6851
rect 25053 6817 25087 6851
rect 25087 6817 25096 6851
rect 25044 6808 25096 6817
rect 36084 6876 36136 6928
rect 36912 6876 36964 6928
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 4436 6647 4488 6656
rect 4436 6613 4445 6647
rect 4445 6613 4479 6647
rect 4479 6613 4488 6647
rect 4436 6604 4488 6613
rect 14924 6740 14976 6792
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 13084 6672 13136 6724
rect 14740 6672 14792 6724
rect 9312 6604 9364 6613
rect 11520 6604 11572 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 19800 6740 19852 6792
rect 16764 6604 16816 6656
rect 17408 6604 17460 6656
rect 17684 6604 17736 6656
rect 18880 6604 18932 6656
rect 20996 6672 21048 6724
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 21088 6604 21140 6656
rect 27528 6740 27580 6792
rect 27896 6740 27948 6792
rect 26516 6672 26568 6724
rect 31852 6808 31904 6860
rect 33784 6851 33836 6860
rect 33784 6817 33793 6851
rect 33793 6817 33827 6851
rect 33827 6817 33836 6851
rect 33784 6808 33836 6817
rect 36636 6808 36688 6860
rect 38476 6808 38528 6860
rect 38936 6851 38988 6860
rect 38936 6817 38945 6851
rect 38945 6817 38979 6851
rect 38979 6817 38988 6851
rect 38936 6808 38988 6817
rect 39120 6851 39172 6860
rect 39120 6817 39129 6851
rect 39129 6817 39163 6851
rect 39163 6817 39172 6851
rect 39120 6808 39172 6817
rect 39856 6808 39908 6860
rect 41512 6808 41564 6860
rect 41880 6851 41932 6860
rect 41880 6817 41889 6851
rect 41889 6817 41923 6851
rect 41923 6817 41932 6851
rect 41880 6808 41932 6817
rect 29184 6740 29236 6792
rect 30656 6740 30708 6792
rect 32772 6740 32824 6792
rect 32864 6783 32916 6792
rect 32864 6749 32873 6783
rect 32873 6749 32907 6783
rect 32907 6749 32916 6783
rect 32864 6740 32916 6749
rect 36360 6740 36412 6792
rect 37464 6783 37516 6792
rect 37464 6749 37473 6783
rect 37473 6749 37507 6783
rect 37507 6749 37516 6783
rect 37464 6740 37516 6749
rect 22836 6604 22888 6656
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 25136 6604 25188 6656
rect 27160 6604 27212 6656
rect 29644 6672 29696 6724
rect 35808 6715 35860 6724
rect 35808 6681 35817 6715
rect 35817 6681 35851 6715
rect 35851 6681 35860 6715
rect 35808 6672 35860 6681
rect 30288 6604 30340 6656
rect 30472 6647 30524 6656
rect 30472 6613 30481 6647
rect 30481 6613 30515 6647
rect 30515 6613 30524 6647
rect 30472 6604 30524 6613
rect 30840 6604 30892 6656
rect 31208 6604 31260 6656
rect 31944 6647 31996 6656
rect 31944 6613 31953 6647
rect 31953 6613 31987 6647
rect 31987 6613 31996 6647
rect 31944 6604 31996 6613
rect 32404 6647 32456 6656
rect 32404 6613 32413 6647
rect 32413 6613 32447 6647
rect 32447 6613 32456 6647
rect 32404 6604 32456 6613
rect 34704 6604 34756 6656
rect 40500 6740 40552 6792
rect 41604 6740 41656 6792
rect 43352 6808 43404 6860
rect 44824 6808 44876 6860
rect 46112 6851 46164 6860
rect 42432 6740 42484 6792
rect 46112 6817 46121 6851
rect 46121 6817 46155 6851
rect 46155 6817 46164 6851
rect 46112 6808 46164 6817
rect 49148 6876 49200 6928
rect 49884 6876 49936 6928
rect 51356 6944 51408 6996
rect 51632 6987 51684 6996
rect 51632 6953 51641 6987
rect 51641 6953 51675 6987
rect 51675 6953 51684 6987
rect 51632 6944 51684 6953
rect 53104 6944 53156 6996
rect 54576 6944 54628 6996
rect 54944 6944 54996 6996
rect 55404 6944 55456 6996
rect 50896 6876 50948 6928
rect 52828 6876 52880 6928
rect 56232 6919 56284 6928
rect 56232 6885 56241 6919
rect 56241 6885 56275 6919
rect 56275 6885 56284 6919
rect 56232 6876 56284 6885
rect 48504 6808 48556 6860
rect 54208 6851 54260 6860
rect 54208 6817 54217 6851
rect 54217 6817 54251 6851
rect 54251 6817 54260 6851
rect 54208 6808 54260 6817
rect 54944 6808 54996 6860
rect 46296 6783 46348 6792
rect 46296 6749 46305 6783
rect 46305 6749 46339 6783
rect 46339 6749 46348 6783
rect 46296 6740 46348 6749
rect 38752 6672 38804 6724
rect 39396 6672 39448 6724
rect 38200 6647 38252 6656
rect 38200 6613 38209 6647
rect 38209 6613 38243 6647
rect 38243 6613 38252 6647
rect 38200 6604 38252 6613
rect 39028 6604 39080 6656
rect 40040 6604 40092 6656
rect 41144 6647 41196 6656
rect 41144 6613 41153 6647
rect 41153 6613 41187 6647
rect 41187 6613 41196 6647
rect 41144 6604 41196 6613
rect 42248 6672 42300 6724
rect 42524 6647 42576 6656
rect 42524 6613 42533 6647
rect 42533 6613 42567 6647
rect 42567 6613 42576 6647
rect 42524 6604 42576 6613
rect 42708 6672 42760 6724
rect 45192 6672 45244 6724
rect 44456 6604 44508 6656
rect 44732 6604 44784 6656
rect 45468 6604 45520 6656
rect 46940 6604 46992 6656
rect 48228 6647 48280 6656
rect 48228 6613 48237 6647
rect 48237 6613 48271 6647
rect 48271 6613 48280 6647
rect 48228 6604 48280 6613
rect 53288 6783 53340 6792
rect 53288 6749 53297 6783
rect 53297 6749 53331 6783
rect 53331 6749 53340 6783
rect 53288 6740 53340 6749
rect 56416 6808 56468 6860
rect 56692 6740 56744 6792
rect 57336 6740 57388 6792
rect 58072 6740 58124 6792
rect 58440 6783 58492 6792
rect 58440 6749 58449 6783
rect 58449 6749 58483 6783
rect 58483 6749 58492 6783
rect 58440 6740 58492 6749
rect 53932 6604 53984 6656
rect 54116 6647 54168 6656
rect 54116 6613 54125 6647
rect 54125 6613 54159 6647
rect 54159 6613 54168 6647
rect 54116 6604 54168 6613
rect 54208 6604 54260 6656
rect 55772 6604 55824 6656
rect 58532 6672 58584 6724
rect 58256 6647 58308 6656
rect 58256 6613 58265 6647
rect 58265 6613 58299 6647
rect 58299 6613 58308 6647
rect 58256 6604 58308 6613
rect 15394 6502 15446 6554
rect 15458 6502 15510 6554
rect 15522 6502 15574 6554
rect 15586 6502 15638 6554
rect 15650 6502 15702 6554
rect 29838 6502 29890 6554
rect 29902 6502 29954 6554
rect 29966 6502 30018 6554
rect 30030 6502 30082 6554
rect 30094 6502 30146 6554
rect 44282 6502 44334 6554
rect 44346 6502 44398 6554
rect 44410 6502 44462 6554
rect 44474 6502 44526 6554
rect 44538 6502 44590 6554
rect 58726 6502 58778 6554
rect 58790 6502 58842 6554
rect 58854 6502 58906 6554
rect 58918 6502 58970 6554
rect 58982 6502 59034 6554
rect 2596 6400 2648 6452
rect 3332 6443 3384 6452
rect 3332 6409 3341 6443
rect 3341 6409 3375 6443
rect 3375 6409 3384 6443
rect 3332 6400 3384 6409
rect 4436 6400 4488 6452
rect 6736 6400 6788 6452
rect 9864 6400 9916 6452
rect 11428 6400 11480 6452
rect 5448 6375 5500 6384
rect 5448 6341 5457 6375
rect 5457 6341 5491 6375
rect 5491 6341 5500 6375
rect 5448 6332 5500 6341
rect 5632 6332 5684 6384
rect 8760 6332 8812 6384
rect 9404 6332 9456 6384
rect 11796 6332 11848 6384
rect 13084 6443 13136 6452
rect 13084 6409 13093 6443
rect 13093 6409 13127 6443
rect 13127 6409 13136 6443
rect 13084 6400 13136 6409
rect 14556 6400 14608 6452
rect 15936 6400 15988 6452
rect 18052 6400 18104 6452
rect 20720 6400 20772 6452
rect 21548 6443 21600 6452
rect 21548 6409 21557 6443
rect 21557 6409 21591 6443
rect 21591 6409 21600 6443
rect 21548 6400 21600 6409
rect 22192 6443 22244 6452
rect 22192 6409 22201 6443
rect 22201 6409 22235 6443
rect 22235 6409 22244 6443
rect 22192 6400 22244 6409
rect 24400 6400 24452 6452
rect 25596 6400 25648 6452
rect 25964 6400 26016 6452
rect 26424 6443 26476 6452
rect 26424 6409 26433 6443
rect 26433 6409 26467 6443
rect 26467 6409 26476 6443
rect 26424 6400 26476 6409
rect 29368 6400 29420 6452
rect 29552 6443 29604 6452
rect 29552 6409 29561 6443
rect 29561 6409 29595 6443
rect 29595 6409 29604 6443
rect 29552 6400 29604 6409
rect 30288 6400 30340 6452
rect 31668 6400 31720 6452
rect 34428 6400 34480 6452
rect 37740 6400 37792 6452
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 3240 6264 3292 6316
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 9588 6264 9640 6316
rect 7748 6196 7800 6248
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 14832 6332 14884 6384
rect 14740 6264 14792 6316
rect 2228 6060 2280 6112
rect 7564 6128 7616 6180
rect 8024 6128 8076 6180
rect 10508 6196 10560 6248
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 18880 6375 18932 6384
rect 18880 6341 18889 6375
rect 18889 6341 18923 6375
rect 18923 6341 18932 6375
rect 18880 6332 18932 6341
rect 18512 6264 18564 6316
rect 16672 6196 16724 6248
rect 19432 6196 19484 6248
rect 22836 6332 22888 6384
rect 32404 6332 32456 6384
rect 33324 6332 33376 6384
rect 34060 6332 34112 6384
rect 35072 6332 35124 6384
rect 39856 6400 39908 6452
rect 40224 6400 40276 6452
rect 41236 6400 41288 6452
rect 41512 6400 41564 6452
rect 40500 6332 40552 6384
rect 41604 6332 41656 6384
rect 20720 6307 20772 6316
rect 20720 6273 20729 6307
rect 20729 6273 20763 6307
rect 20763 6273 20772 6307
rect 20720 6264 20772 6273
rect 19708 6196 19760 6248
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 5172 6060 5224 6112
rect 14648 6060 14700 6112
rect 17776 6171 17828 6180
rect 17776 6137 17785 6171
rect 17785 6137 17819 6171
rect 17819 6137 17828 6171
rect 17776 6128 17828 6137
rect 20076 6128 20128 6180
rect 23112 6264 23164 6316
rect 27896 6264 27948 6316
rect 28908 6264 28960 6316
rect 29736 6264 29788 6316
rect 24400 6196 24452 6248
rect 25136 6196 25188 6248
rect 15660 6060 15712 6112
rect 16764 6060 16816 6112
rect 16948 6060 17000 6112
rect 19340 6060 19392 6112
rect 19800 6060 19852 6112
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 29644 6128 29696 6180
rect 30840 6307 30892 6316
rect 30840 6273 30849 6307
rect 30849 6273 30883 6307
rect 30883 6273 30892 6307
rect 30840 6264 30892 6273
rect 33508 6264 33560 6316
rect 34888 6307 34940 6316
rect 34888 6273 34897 6307
rect 34897 6273 34931 6307
rect 34931 6273 34940 6307
rect 34888 6264 34940 6273
rect 22376 6060 22428 6112
rect 23388 6103 23440 6112
rect 23388 6069 23397 6103
rect 23397 6069 23431 6103
rect 23431 6069 23440 6103
rect 23388 6060 23440 6069
rect 24124 6060 24176 6112
rect 25044 6060 25096 6112
rect 26148 6060 26200 6112
rect 30012 6060 30064 6112
rect 31484 6196 31536 6248
rect 30564 6171 30616 6180
rect 30564 6137 30573 6171
rect 30573 6137 30607 6171
rect 30607 6137 30616 6171
rect 30564 6128 30616 6137
rect 31944 6196 31996 6248
rect 31760 6103 31812 6112
rect 31760 6069 31769 6103
rect 31769 6069 31803 6103
rect 31803 6069 31812 6103
rect 31760 6060 31812 6069
rect 32956 6060 33008 6112
rect 34980 6196 35032 6248
rect 35624 6196 35676 6248
rect 40684 6264 40736 6316
rect 41512 6264 41564 6316
rect 42708 6400 42760 6452
rect 45468 6400 45520 6452
rect 48596 6400 48648 6452
rect 49148 6400 49200 6452
rect 52184 6400 52236 6452
rect 53748 6400 53800 6452
rect 56876 6400 56928 6452
rect 46112 6332 46164 6384
rect 49884 6332 49936 6384
rect 51632 6332 51684 6384
rect 52828 6332 52880 6384
rect 38568 6239 38620 6248
rect 38568 6205 38577 6239
rect 38577 6205 38611 6239
rect 38611 6205 38620 6239
rect 38568 6196 38620 6205
rect 40132 6196 40184 6248
rect 45560 6264 45612 6316
rect 48228 6264 48280 6316
rect 43904 6196 43956 6248
rect 44916 6239 44968 6248
rect 44916 6205 44925 6239
rect 44925 6205 44959 6239
rect 44959 6205 44968 6239
rect 44916 6196 44968 6205
rect 47124 6239 47176 6248
rect 47124 6205 47133 6239
rect 47133 6205 47167 6239
rect 47167 6205 47176 6239
rect 47124 6196 47176 6205
rect 49608 6239 49660 6248
rect 49608 6205 49617 6239
rect 49617 6205 49651 6239
rect 49651 6205 49660 6239
rect 49608 6196 49660 6205
rect 50068 6307 50120 6316
rect 50068 6273 50077 6307
rect 50077 6273 50111 6307
rect 50111 6273 50120 6307
rect 50068 6264 50120 6273
rect 52276 6196 52328 6248
rect 38200 6171 38252 6180
rect 34704 6060 34756 6112
rect 35164 6060 35216 6112
rect 35532 6060 35584 6112
rect 38200 6137 38209 6171
rect 38209 6137 38243 6171
rect 38243 6137 38252 6171
rect 38200 6128 38252 6137
rect 41236 6128 41288 6180
rect 42340 6128 42392 6180
rect 46940 6128 46992 6180
rect 36728 6060 36780 6112
rect 38384 6060 38436 6112
rect 39120 6103 39172 6112
rect 39120 6069 39129 6103
rect 39129 6069 39163 6103
rect 39163 6069 39172 6103
rect 39120 6060 39172 6069
rect 39948 6060 40000 6112
rect 41328 6060 41380 6112
rect 42616 6060 42668 6112
rect 45468 6103 45520 6112
rect 45468 6069 45477 6103
rect 45477 6069 45511 6103
rect 45511 6069 45520 6103
rect 45468 6060 45520 6069
rect 45652 6060 45704 6112
rect 48872 6060 48924 6112
rect 50344 6103 50396 6112
rect 50344 6069 50353 6103
rect 50353 6069 50387 6103
rect 50387 6069 50396 6103
rect 50344 6060 50396 6069
rect 50528 6060 50580 6112
rect 52552 6264 52604 6316
rect 54944 6307 54996 6316
rect 54944 6273 54953 6307
rect 54953 6273 54987 6307
rect 54987 6273 54996 6307
rect 54944 6264 54996 6273
rect 55772 6307 55824 6316
rect 55772 6273 55806 6307
rect 55806 6273 55824 6307
rect 55772 6264 55824 6273
rect 56784 6264 56836 6316
rect 57796 6264 57848 6316
rect 52736 6128 52788 6180
rect 55036 6196 55088 6248
rect 56140 6196 56192 6248
rect 55312 6128 55364 6180
rect 55404 6171 55456 6180
rect 55404 6137 55413 6171
rect 55413 6137 55447 6171
rect 55447 6137 55456 6171
rect 55404 6128 55456 6137
rect 54024 6060 54076 6112
rect 55772 6060 55824 6112
rect 55864 6060 55916 6112
rect 56600 6196 56652 6248
rect 57152 6239 57204 6248
rect 57152 6205 57161 6239
rect 57161 6205 57195 6239
rect 57195 6205 57204 6239
rect 57152 6196 57204 6205
rect 57244 6239 57296 6248
rect 57244 6205 57253 6239
rect 57253 6205 57287 6239
rect 57287 6205 57296 6239
rect 57244 6196 57296 6205
rect 56600 6103 56652 6112
rect 56600 6069 56609 6103
rect 56609 6069 56643 6103
rect 56643 6069 56652 6103
rect 56600 6060 56652 6069
rect 57520 6103 57572 6112
rect 57520 6069 57529 6103
rect 57529 6069 57563 6103
rect 57563 6069 57572 6103
rect 57520 6060 57572 6069
rect 8172 5958 8224 6010
rect 8236 5958 8288 6010
rect 8300 5958 8352 6010
rect 8364 5958 8416 6010
rect 8428 5958 8480 6010
rect 22616 5958 22668 6010
rect 22680 5958 22732 6010
rect 22744 5958 22796 6010
rect 22808 5958 22860 6010
rect 22872 5958 22924 6010
rect 37060 5958 37112 6010
rect 37124 5958 37176 6010
rect 37188 5958 37240 6010
rect 37252 5958 37304 6010
rect 37316 5958 37368 6010
rect 51504 5958 51556 6010
rect 51568 5958 51620 6010
rect 51632 5958 51684 6010
rect 51696 5958 51748 6010
rect 51760 5958 51812 6010
rect 2504 5856 2556 5908
rect 3976 5856 4028 5908
rect 5172 5856 5224 5908
rect 8024 5856 8076 5908
rect 9588 5899 9640 5908
rect 9588 5865 9597 5899
rect 9597 5865 9631 5899
rect 9631 5865 9640 5899
rect 9588 5856 9640 5865
rect 9680 5856 9732 5908
rect 10784 5856 10836 5908
rect 11888 5856 11940 5908
rect 12808 5856 12860 5908
rect 13544 5856 13596 5908
rect 14096 5856 14148 5908
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 14924 5856 14976 5908
rect 15108 5856 15160 5908
rect 17684 5856 17736 5908
rect 17776 5899 17828 5908
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 22376 5856 22428 5908
rect 22652 5856 22704 5908
rect 26148 5856 26200 5908
rect 28264 5899 28316 5908
rect 28264 5865 28273 5899
rect 28273 5865 28307 5899
rect 28307 5865 28316 5899
rect 28264 5856 28316 5865
rect 29552 5856 29604 5908
rect 8576 5788 8628 5840
rect 5172 5720 5224 5772
rect 12164 5788 12216 5840
rect 3884 5652 3936 5704
rect 5632 5695 5684 5704
rect 2596 5584 2648 5636
rect 3332 5584 3384 5636
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 4620 5516 4672 5568
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 5540 5584 5592 5636
rect 10692 5652 10744 5704
rect 15844 5720 15896 5772
rect 16948 5720 17000 5772
rect 19432 5720 19484 5772
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 16396 5652 16448 5704
rect 17776 5652 17828 5704
rect 18144 5652 18196 5704
rect 8852 5584 8904 5636
rect 9312 5584 9364 5636
rect 6184 5516 6236 5568
rect 7840 5516 7892 5568
rect 9772 5584 9824 5636
rect 10140 5584 10192 5636
rect 15292 5584 15344 5636
rect 12348 5516 12400 5568
rect 12532 5516 12584 5568
rect 14188 5516 14240 5568
rect 15660 5516 15712 5568
rect 15936 5584 15988 5636
rect 16672 5584 16724 5636
rect 16120 5516 16172 5568
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 17132 5516 17184 5525
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 19064 5559 19116 5568
rect 19064 5525 19073 5559
rect 19073 5525 19107 5559
rect 19107 5525 19116 5559
rect 19064 5516 19116 5525
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 26240 5720 26292 5772
rect 26424 5763 26476 5772
rect 26424 5729 26433 5763
rect 26433 5729 26467 5763
rect 26467 5729 26476 5763
rect 26424 5720 26476 5729
rect 27712 5720 27764 5772
rect 21732 5652 21784 5704
rect 22192 5652 22244 5704
rect 23020 5652 23072 5704
rect 23388 5695 23440 5704
rect 23388 5661 23397 5695
rect 23397 5661 23431 5695
rect 23431 5661 23440 5695
rect 23388 5652 23440 5661
rect 23664 5695 23716 5704
rect 23664 5661 23673 5695
rect 23673 5661 23707 5695
rect 23707 5661 23716 5695
rect 23664 5652 23716 5661
rect 25320 5584 25372 5636
rect 19800 5516 19852 5568
rect 20720 5516 20772 5568
rect 21916 5516 21968 5568
rect 22008 5516 22060 5568
rect 22376 5516 22428 5568
rect 23940 5516 23992 5568
rect 24400 5516 24452 5568
rect 25872 5559 25924 5568
rect 25872 5525 25881 5559
rect 25881 5525 25915 5559
rect 25915 5525 25924 5559
rect 25872 5516 25924 5525
rect 26332 5652 26384 5704
rect 29276 5652 29328 5704
rect 30656 5720 30708 5772
rect 32864 5856 32916 5908
rect 32956 5856 33008 5908
rect 34612 5856 34664 5908
rect 35808 5856 35860 5908
rect 38568 5856 38620 5908
rect 32220 5720 32272 5772
rect 29552 5584 29604 5636
rect 28448 5559 28500 5568
rect 28448 5525 28457 5559
rect 28457 5525 28491 5559
rect 28491 5525 28500 5559
rect 28448 5516 28500 5525
rect 40224 5856 40276 5908
rect 44916 5856 44968 5908
rect 45652 5856 45704 5908
rect 46940 5856 46992 5908
rect 49608 5899 49660 5908
rect 49608 5865 49617 5899
rect 49617 5865 49651 5899
rect 49651 5865 49660 5899
rect 49608 5856 49660 5865
rect 54208 5856 54260 5908
rect 55036 5856 55088 5908
rect 55312 5856 55364 5908
rect 57060 5856 57112 5908
rect 57428 5899 57480 5908
rect 57428 5865 57437 5899
rect 57437 5865 57471 5899
rect 57471 5865 57480 5899
rect 57428 5856 57480 5865
rect 58348 5856 58400 5908
rect 39396 5763 39448 5772
rect 39396 5729 39405 5763
rect 39405 5729 39439 5763
rect 39439 5729 39448 5763
rect 39396 5720 39448 5729
rect 31852 5695 31904 5704
rect 31852 5661 31861 5695
rect 31861 5661 31895 5695
rect 31895 5661 31904 5695
rect 31852 5652 31904 5661
rect 33600 5695 33652 5704
rect 33600 5661 33609 5695
rect 33609 5661 33643 5695
rect 33643 5661 33652 5695
rect 33600 5652 33652 5661
rect 34704 5695 34756 5704
rect 34704 5661 34713 5695
rect 34713 5661 34747 5695
rect 34747 5661 34756 5695
rect 34704 5652 34756 5661
rect 36912 5652 36964 5704
rect 37464 5652 37516 5704
rect 40592 5720 40644 5772
rect 41880 5720 41932 5772
rect 50344 5720 50396 5772
rect 52552 5720 52604 5772
rect 39856 5695 39908 5704
rect 39856 5661 39865 5695
rect 39865 5661 39899 5695
rect 39899 5661 39908 5695
rect 39856 5652 39908 5661
rect 39948 5652 40000 5704
rect 30564 5627 30616 5636
rect 30564 5593 30573 5627
rect 30573 5593 30607 5627
rect 30607 5593 30616 5627
rect 30564 5584 30616 5593
rect 30748 5584 30800 5636
rect 31300 5627 31352 5636
rect 31300 5593 31309 5627
rect 31309 5593 31343 5627
rect 31343 5593 31352 5627
rect 31300 5584 31352 5593
rect 31484 5584 31536 5636
rect 34612 5584 34664 5636
rect 35532 5627 35584 5636
rect 35532 5593 35541 5627
rect 35541 5593 35575 5627
rect 35575 5593 35584 5627
rect 35532 5584 35584 5593
rect 40684 5652 40736 5704
rect 43352 5652 43404 5704
rect 43996 5695 44048 5704
rect 43996 5661 44005 5695
rect 44005 5661 44039 5695
rect 44039 5661 44048 5695
rect 43996 5652 44048 5661
rect 44180 5652 44232 5704
rect 45376 5695 45428 5704
rect 45376 5661 45385 5695
rect 45385 5661 45419 5695
rect 45419 5661 45428 5695
rect 45376 5652 45428 5661
rect 45836 5695 45888 5704
rect 45836 5661 45845 5695
rect 45845 5661 45879 5695
rect 45879 5661 45888 5695
rect 45836 5652 45888 5661
rect 48688 5695 48740 5704
rect 48688 5661 48697 5695
rect 48697 5661 48731 5695
rect 48731 5661 48740 5695
rect 48688 5652 48740 5661
rect 50160 5652 50212 5704
rect 50988 5695 51040 5704
rect 50988 5661 50997 5695
rect 50997 5661 51031 5695
rect 51031 5661 51040 5695
rect 50988 5652 51040 5661
rect 53932 5652 53984 5704
rect 55128 5695 55180 5704
rect 55128 5661 55137 5695
rect 55137 5661 55171 5695
rect 55171 5661 55180 5695
rect 55128 5652 55180 5661
rect 55496 5695 55548 5704
rect 55496 5661 55505 5695
rect 55505 5661 55539 5695
rect 55539 5661 55548 5695
rect 55496 5652 55548 5661
rect 55864 5652 55916 5704
rect 57520 5720 57572 5772
rect 57980 5763 58032 5772
rect 57980 5729 57989 5763
rect 57989 5729 58023 5763
rect 58023 5729 58032 5763
rect 57980 5720 58032 5729
rect 41420 5584 41472 5636
rect 43076 5584 43128 5636
rect 31116 5516 31168 5568
rect 31208 5559 31260 5568
rect 31208 5525 31217 5559
rect 31217 5525 31251 5559
rect 31251 5525 31260 5559
rect 31208 5516 31260 5525
rect 34152 5559 34204 5568
rect 34152 5525 34161 5559
rect 34161 5525 34195 5559
rect 34195 5525 34204 5559
rect 34152 5516 34204 5525
rect 36268 5516 36320 5568
rect 40132 5516 40184 5568
rect 40776 5559 40828 5568
rect 40776 5525 40785 5559
rect 40785 5525 40819 5559
rect 40819 5525 40828 5559
rect 40776 5516 40828 5525
rect 41972 5516 42024 5568
rect 43812 5559 43864 5568
rect 43812 5525 43821 5559
rect 43821 5525 43855 5559
rect 43855 5525 43864 5559
rect 43812 5516 43864 5525
rect 43904 5516 43956 5568
rect 44088 5516 44140 5568
rect 55036 5584 55088 5636
rect 57704 5652 57756 5704
rect 57888 5652 57940 5704
rect 48504 5516 48556 5568
rect 49424 5516 49476 5568
rect 52368 5559 52420 5568
rect 52368 5525 52377 5559
rect 52377 5525 52411 5559
rect 52411 5525 52420 5559
rect 52368 5516 52420 5525
rect 54944 5559 54996 5568
rect 54944 5525 54953 5559
rect 54953 5525 54987 5559
rect 54987 5525 54996 5559
rect 54944 5516 54996 5525
rect 56508 5516 56560 5568
rect 56784 5516 56836 5568
rect 15394 5414 15446 5466
rect 15458 5414 15510 5466
rect 15522 5414 15574 5466
rect 15586 5414 15638 5466
rect 15650 5414 15702 5466
rect 29838 5414 29890 5466
rect 29902 5414 29954 5466
rect 29966 5414 30018 5466
rect 30030 5414 30082 5466
rect 30094 5414 30146 5466
rect 44282 5414 44334 5466
rect 44346 5414 44398 5466
rect 44410 5414 44462 5466
rect 44474 5414 44526 5466
rect 44538 5414 44590 5466
rect 58726 5414 58778 5466
rect 58790 5414 58842 5466
rect 58854 5414 58906 5466
rect 58918 5414 58970 5466
rect 58982 5414 59034 5466
rect 3332 5312 3384 5364
rect 3608 5244 3660 5296
rect 5448 5244 5500 5296
rect 5632 5244 5684 5296
rect 5172 5176 5224 5228
rect 5724 5176 5776 5228
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 10508 5312 10560 5364
rect 11704 5312 11756 5364
rect 12348 5312 12400 5364
rect 13084 5312 13136 5364
rect 13820 5312 13872 5364
rect 12072 5244 12124 5296
rect 1768 5108 1820 5160
rect 2872 5108 2924 5160
rect 5080 5108 5132 5160
rect 5448 5108 5500 5160
rect 7840 5176 7892 5228
rect 3884 5040 3936 5092
rect 5632 5040 5684 5092
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 9036 5108 9088 5160
rect 11704 5176 11756 5228
rect 15752 5312 15804 5364
rect 17684 5244 17736 5296
rect 13728 5176 13780 5228
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 15752 5219 15804 5228
rect 15752 5185 15761 5219
rect 15761 5185 15795 5219
rect 15795 5185 15804 5219
rect 15752 5176 15804 5185
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 19524 5312 19576 5364
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 18420 5244 18472 5296
rect 19064 5244 19116 5296
rect 21456 5312 21508 5364
rect 22284 5355 22336 5364
rect 22284 5321 22293 5355
rect 22293 5321 22327 5355
rect 22327 5321 22336 5355
rect 22284 5312 22336 5321
rect 23664 5312 23716 5364
rect 21916 5244 21968 5296
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 10968 5108 11020 5160
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 17776 5108 17828 5160
rect 11152 5040 11204 5092
rect 5448 4972 5500 5024
rect 6000 4972 6052 5024
rect 7564 4972 7616 5024
rect 7932 4972 7984 5024
rect 8668 4972 8720 5024
rect 11796 5040 11848 5092
rect 14740 5040 14792 5092
rect 18052 5040 18104 5092
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 22928 5244 22980 5296
rect 23572 5176 23624 5228
rect 26608 5312 26660 5364
rect 28908 5355 28960 5364
rect 28908 5321 28917 5355
rect 28917 5321 28951 5355
rect 28951 5321 28960 5355
rect 28908 5312 28960 5321
rect 29092 5312 29144 5364
rect 29552 5312 29604 5364
rect 30656 5312 30708 5364
rect 31116 5312 31168 5364
rect 27068 5244 27120 5296
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 11888 4972 11940 5024
rect 14464 4972 14516 5024
rect 15108 4972 15160 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 17040 4972 17092 5024
rect 20260 5040 20312 5092
rect 19340 4972 19392 5024
rect 19708 4972 19760 5024
rect 20812 5151 20864 5160
rect 20812 5117 20846 5151
rect 20846 5117 20864 5151
rect 20812 5108 20864 5117
rect 21548 5108 21600 5160
rect 24400 5151 24452 5160
rect 24400 5117 24409 5151
rect 24409 5117 24443 5151
rect 24443 5117 24452 5151
rect 24400 5108 24452 5117
rect 25596 5219 25648 5228
rect 25596 5185 25605 5219
rect 25605 5185 25639 5219
rect 25639 5185 25648 5219
rect 25596 5176 25648 5185
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 25412 5151 25464 5160
rect 32036 5244 32088 5296
rect 34152 5244 34204 5296
rect 28448 5176 28500 5228
rect 29276 5176 29328 5228
rect 29644 5219 29696 5228
rect 29644 5185 29653 5219
rect 29653 5185 29687 5219
rect 29687 5185 29696 5219
rect 29644 5176 29696 5185
rect 31024 5176 31076 5228
rect 31576 5176 31628 5228
rect 33048 5219 33100 5228
rect 33048 5185 33057 5219
rect 33057 5185 33091 5219
rect 33091 5185 33100 5219
rect 33048 5176 33100 5185
rect 34796 5219 34848 5228
rect 34796 5185 34805 5219
rect 34805 5185 34839 5219
rect 34839 5185 34848 5219
rect 34796 5176 34848 5185
rect 37464 5312 37516 5364
rect 37556 5312 37608 5364
rect 39856 5312 39908 5364
rect 40408 5312 40460 5364
rect 41696 5312 41748 5364
rect 44916 5312 44968 5364
rect 45560 5312 45612 5364
rect 45652 5355 45704 5364
rect 45652 5321 45661 5355
rect 45661 5321 45695 5355
rect 45695 5321 45704 5355
rect 45652 5312 45704 5321
rect 45836 5312 45888 5364
rect 46848 5312 46900 5364
rect 48412 5312 48464 5364
rect 35440 5176 35492 5228
rect 35992 5219 36044 5228
rect 35992 5185 36001 5219
rect 36001 5185 36035 5219
rect 36035 5185 36044 5219
rect 35992 5176 36044 5185
rect 36268 5219 36320 5228
rect 36268 5185 36277 5219
rect 36277 5185 36311 5219
rect 36311 5185 36320 5219
rect 36268 5176 36320 5185
rect 39120 5244 39172 5296
rect 42524 5244 42576 5296
rect 40316 5219 40368 5228
rect 40316 5185 40325 5219
rect 40325 5185 40359 5219
rect 40359 5185 40368 5219
rect 40316 5176 40368 5185
rect 40408 5219 40460 5228
rect 40408 5185 40442 5219
rect 40442 5185 40460 5219
rect 40408 5176 40460 5185
rect 25412 5117 25446 5151
rect 25446 5117 25464 5151
rect 25412 5108 25464 5117
rect 29736 5108 29788 5160
rect 24768 5040 24820 5092
rect 26148 5040 26200 5092
rect 34704 5108 34756 5160
rect 36452 5108 36504 5160
rect 37556 5108 37608 5160
rect 39396 5151 39448 5160
rect 39396 5117 39405 5151
rect 39405 5117 39439 5151
rect 39439 5117 39448 5151
rect 39396 5108 39448 5117
rect 39580 5151 39632 5160
rect 39580 5117 39589 5151
rect 39589 5117 39623 5151
rect 39623 5117 39632 5151
rect 39580 5108 39632 5117
rect 40132 5108 40184 5160
rect 41420 5108 41472 5160
rect 42708 5219 42760 5228
rect 42708 5185 42717 5219
rect 42717 5185 42751 5219
rect 42751 5185 42760 5219
rect 42708 5176 42760 5185
rect 43812 5244 43864 5296
rect 45468 5244 45520 5296
rect 26332 4972 26384 5024
rect 28172 5015 28224 5024
rect 28172 4981 28181 5015
rect 28181 4981 28215 5015
rect 28215 4981 28224 5015
rect 28172 4972 28224 4981
rect 29644 4972 29696 5024
rect 30288 4972 30340 5024
rect 30656 5015 30708 5024
rect 30656 4981 30665 5015
rect 30665 4981 30699 5015
rect 30699 4981 30708 5015
rect 30656 4972 30708 4981
rect 32680 5015 32732 5024
rect 32680 4981 32689 5015
rect 32689 4981 32723 5015
rect 32723 4981 32732 5015
rect 32680 4972 32732 4981
rect 34152 4972 34204 5024
rect 34336 4972 34388 5024
rect 35624 5040 35676 5092
rect 36728 5040 36780 5092
rect 37648 5040 37700 5092
rect 36912 5015 36964 5024
rect 36912 4981 36921 5015
rect 36921 4981 36955 5015
rect 36955 4981 36964 5015
rect 36912 4972 36964 4981
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 40684 4972 40736 5024
rect 41420 4972 41472 5024
rect 43996 4972 44048 5024
rect 46204 5151 46256 5160
rect 46204 5117 46213 5151
rect 46213 5117 46247 5151
rect 46247 5117 46256 5151
rect 46204 5108 46256 5117
rect 47124 5040 47176 5092
rect 48228 5151 48280 5160
rect 48228 5117 48237 5151
rect 48237 5117 48271 5151
rect 48271 5117 48280 5151
rect 48228 5108 48280 5117
rect 50988 5312 51040 5364
rect 53748 5355 53800 5364
rect 53748 5321 53757 5355
rect 53757 5321 53791 5355
rect 53791 5321 53800 5355
rect 53748 5312 53800 5321
rect 54116 5312 54168 5364
rect 57152 5312 57204 5364
rect 57888 5312 57940 5364
rect 58532 5355 58584 5364
rect 58532 5321 58541 5355
rect 58541 5321 58575 5355
rect 58575 5321 58584 5355
rect 58532 5312 58584 5321
rect 52092 5244 52144 5296
rect 49424 5219 49476 5228
rect 49424 5185 49433 5219
rect 49433 5185 49467 5219
rect 49467 5185 49476 5219
rect 49424 5176 49476 5185
rect 49700 5219 49752 5228
rect 49700 5185 49709 5219
rect 49709 5185 49743 5219
rect 49743 5185 49752 5219
rect 49700 5176 49752 5185
rect 50528 5176 50580 5228
rect 52368 5176 52420 5228
rect 54484 5176 54536 5228
rect 56692 5176 56744 5228
rect 48596 5040 48648 5092
rect 48780 5108 48832 5160
rect 52276 5108 52328 5160
rect 53656 5108 53708 5160
rect 54208 5151 54260 5160
rect 54208 5117 54217 5151
rect 54217 5117 54251 5151
rect 54251 5117 54260 5151
rect 54208 5108 54260 5117
rect 45192 4972 45244 5024
rect 47032 4972 47084 5024
rect 47216 4972 47268 5024
rect 49148 5083 49200 5092
rect 49148 5049 49157 5083
rect 49157 5049 49191 5083
rect 49191 5049 49200 5083
rect 49148 5040 49200 5049
rect 55680 5151 55732 5160
rect 55680 5117 55689 5151
rect 55689 5117 55723 5151
rect 55723 5117 55732 5151
rect 55680 5108 55732 5117
rect 56324 5151 56376 5160
rect 56324 5117 56333 5151
rect 56333 5117 56367 5151
rect 56367 5117 56376 5151
rect 56324 5108 56376 5117
rect 49792 4972 49844 5024
rect 50344 5015 50396 5024
rect 50344 4981 50353 5015
rect 50353 4981 50387 5015
rect 50387 4981 50396 5015
rect 50344 4972 50396 4981
rect 51080 4972 51132 5024
rect 52092 5015 52144 5024
rect 52092 4981 52101 5015
rect 52101 4981 52135 5015
rect 52135 4981 52144 5015
rect 52092 4972 52144 4981
rect 52920 5015 52972 5024
rect 52920 4981 52929 5015
rect 52929 4981 52963 5015
rect 52963 4981 52972 5015
rect 52920 4972 52972 4981
rect 53840 5015 53892 5024
rect 53840 4981 53849 5015
rect 53849 4981 53883 5015
rect 53883 4981 53892 5015
rect 53840 4972 53892 4981
rect 56692 5040 56744 5092
rect 57060 5219 57112 5228
rect 57060 5185 57069 5219
rect 57069 5185 57103 5219
rect 57103 5185 57112 5219
rect 57060 5176 57112 5185
rect 57428 5176 57480 5228
rect 57060 5040 57112 5092
rect 55588 4972 55640 5024
rect 56232 5015 56284 5024
rect 56232 4981 56241 5015
rect 56241 4981 56275 5015
rect 56275 4981 56284 5015
rect 56232 4972 56284 4981
rect 56968 5015 57020 5024
rect 56968 4981 56977 5015
rect 56977 4981 57011 5015
rect 57011 4981 57020 5015
rect 56968 4972 57020 4981
rect 8172 4870 8224 4922
rect 8236 4870 8288 4922
rect 8300 4870 8352 4922
rect 8364 4870 8416 4922
rect 8428 4870 8480 4922
rect 22616 4870 22668 4922
rect 22680 4870 22732 4922
rect 22744 4870 22796 4922
rect 22808 4870 22860 4922
rect 22872 4870 22924 4922
rect 37060 4870 37112 4922
rect 37124 4870 37176 4922
rect 37188 4870 37240 4922
rect 37252 4870 37304 4922
rect 37316 4870 37368 4922
rect 51504 4870 51556 4922
rect 51568 4870 51620 4922
rect 51632 4870 51684 4922
rect 51696 4870 51748 4922
rect 51760 4870 51812 4922
rect 2228 4768 2280 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3424 4768 3476 4820
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 7656 4768 7708 4820
rect 2596 4700 2648 4752
rect 4528 4700 4580 4752
rect 5448 4700 5500 4752
rect 3332 4632 3384 4684
rect 5080 4632 5132 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2596 4564 2648 4616
rect 2872 4564 2924 4616
rect 3056 4496 3108 4548
rect 3976 4539 4028 4548
rect 3976 4505 4001 4539
rect 4001 4505 4028 4539
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 6276 4700 6328 4752
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 10232 4743 10284 4752
rect 10232 4709 10241 4743
rect 10241 4709 10275 4743
rect 10275 4709 10284 4743
rect 10232 4700 10284 4709
rect 10876 4632 10928 4684
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 9128 4607 9180 4616
rect 7564 4564 7616 4573
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 10692 4564 10744 4616
rect 11152 4564 11204 4616
rect 11796 4564 11848 4616
rect 3976 4496 4028 4505
rect 7748 4496 7800 4548
rect 8024 4496 8076 4548
rect 11612 4496 11664 4548
rect 14832 4632 14884 4684
rect 17500 4768 17552 4820
rect 18420 4768 18472 4820
rect 19984 4768 20036 4820
rect 21916 4768 21968 4820
rect 26332 4768 26384 4820
rect 14096 4564 14148 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 17132 4564 17184 4616
rect 16028 4496 16080 4548
rect 17224 4496 17276 4548
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4804 4428 4856 4480
rect 5908 4428 5960 4480
rect 11244 4428 11296 4480
rect 11796 4428 11848 4480
rect 13912 4471 13964 4480
rect 13912 4437 13921 4471
rect 13921 4437 13955 4471
rect 13955 4437 13964 4471
rect 13912 4428 13964 4437
rect 14832 4471 14884 4480
rect 14832 4437 14841 4471
rect 14841 4437 14875 4471
rect 14875 4437 14884 4471
rect 14832 4428 14884 4437
rect 15200 4428 15252 4480
rect 15844 4428 15896 4480
rect 17684 4564 17736 4616
rect 18052 4564 18104 4616
rect 23020 4632 23072 4684
rect 23940 4675 23992 4684
rect 23940 4641 23949 4675
rect 23949 4641 23983 4675
rect 23983 4641 23992 4675
rect 23940 4632 23992 4641
rect 24124 4675 24176 4684
rect 24124 4641 24133 4675
rect 24133 4641 24167 4675
rect 24167 4641 24176 4675
rect 24124 4632 24176 4641
rect 24400 4632 24452 4684
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 20720 4564 20772 4616
rect 22008 4564 22060 4616
rect 17776 4428 17828 4480
rect 19064 4471 19116 4480
rect 19064 4437 19073 4471
rect 19073 4437 19107 4471
rect 19107 4437 19116 4471
rect 19064 4428 19116 4437
rect 19984 4496 20036 4548
rect 24768 4496 24820 4548
rect 26240 4564 26292 4616
rect 20812 4428 20864 4480
rect 23480 4471 23532 4480
rect 23480 4437 23489 4471
rect 23489 4437 23523 4471
rect 23523 4437 23532 4471
rect 23480 4428 23532 4437
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 25504 4496 25556 4548
rect 26424 4496 26476 4548
rect 26332 4428 26384 4480
rect 26608 4428 26660 4480
rect 29736 4768 29788 4820
rect 27620 4700 27672 4752
rect 31208 4743 31260 4752
rect 31208 4709 31217 4743
rect 31217 4709 31251 4743
rect 31251 4709 31260 4743
rect 31208 4700 31260 4709
rect 27712 4632 27764 4684
rect 33232 4768 33284 4820
rect 33600 4811 33652 4820
rect 33600 4777 33609 4811
rect 33609 4777 33643 4811
rect 33643 4777 33652 4811
rect 33600 4768 33652 4777
rect 34704 4768 34756 4820
rect 32036 4700 32088 4752
rect 27988 4564 28040 4616
rect 29184 4564 29236 4616
rect 29552 4564 29604 4616
rect 30564 4607 30616 4616
rect 30564 4573 30573 4607
rect 30573 4573 30607 4607
rect 30607 4573 30616 4607
rect 30564 4564 30616 4573
rect 31392 4564 31444 4616
rect 31484 4496 31536 4548
rect 31760 4496 31812 4548
rect 34060 4675 34112 4684
rect 34060 4641 34069 4675
rect 34069 4641 34103 4675
rect 34103 4641 34112 4675
rect 34060 4632 34112 4641
rect 34612 4700 34664 4752
rect 35992 4768 36044 4820
rect 36452 4700 36504 4752
rect 34428 4632 34480 4684
rect 36912 4768 36964 4820
rect 36820 4700 36872 4752
rect 38292 4700 38344 4752
rect 32680 4564 32732 4616
rect 33324 4539 33376 4548
rect 33324 4505 33333 4539
rect 33333 4505 33367 4539
rect 33367 4505 33376 4539
rect 33324 4496 33376 4505
rect 35808 4564 35860 4616
rect 36544 4607 36596 4616
rect 36544 4573 36553 4607
rect 36553 4573 36587 4607
rect 36587 4573 36596 4607
rect 36544 4564 36596 4573
rect 29368 4471 29420 4480
rect 29368 4437 29377 4471
rect 29377 4437 29411 4471
rect 29411 4437 29420 4471
rect 29368 4428 29420 4437
rect 30288 4428 30340 4480
rect 31116 4471 31168 4480
rect 31116 4437 31125 4471
rect 31125 4437 31159 4471
rect 31159 4437 31168 4471
rect 31116 4428 31168 4437
rect 31944 4428 31996 4480
rect 33416 4471 33468 4480
rect 33416 4437 33425 4471
rect 33425 4437 33459 4471
rect 33459 4437 33468 4471
rect 33416 4428 33468 4437
rect 33968 4471 34020 4480
rect 33968 4437 33977 4471
rect 33977 4437 34011 4471
rect 34011 4437 34020 4471
rect 33968 4428 34020 4437
rect 35900 4496 35952 4548
rect 37280 4632 37332 4684
rect 39580 4768 39632 4820
rect 40040 4768 40092 4820
rect 40316 4768 40368 4820
rect 39948 4632 40000 4684
rect 40500 4675 40552 4684
rect 40500 4641 40509 4675
rect 40509 4641 40543 4675
rect 40543 4641 40552 4675
rect 40500 4632 40552 4641
rect 36820 4564 36872 4616
rect 38016 4607 38068 4616
rect 38016 4573 38025 4607
rect 38025 4573 38059 4607
rect 38059 4573 38068 4607
rect 38016 4564 38068 4573
rect 40776 4632 40828 4684
rect 43076 4811 43128 4820
rect 43076 4777 43085 4811
rect 43085 4777 43119 4811
rect 43119 4777 43128 4811
rect 43076 4768 43128 4777
rect 43352 4811 43404 4820
rect 43352 4777 43361 4811
rect 43361 4777 43395 4811
rect 43395 4777 43404 4811
rect 43352 4768 43404 4777
rect 43996 4768 44048 4820
rect 37556 4496 37608 4548
rect 40868 4607 40920 4616
rect 40868 4573 40877 4607
rect 40877 4573 40911 4607
rect 40911 4573 40920 4607
rect 40868 4564 40920 4573
rect 43904 4675 43956 4684
rect 43904 4641 43913 4675
rect 43913 4641 43947 4675
rect 43947 4641 43956 4675
rect 43904 4632 43956 4641
rect 44088 4632 44140 4684
rect 44916 4700 44968 4752
rect 44640 4632 44692 4684
rect 45468 4700 45520 4752
rect 45560 4632 45612 4684
rect 45652 4675 45704 4684
rect 45652 4641 45661 4675
rect 45661 4641 45695 4675
rect 45695 4641 45704 4675
rect 45652 4632 45704 4641
rect 46204 4768 46256 4820
rect 48228 4700 48280 4752
rect 48688 4768 48740 4820
rect 48780 4768 48832 4820
rect 46388 4632 46440 4684
rect 46940 4675 46992 4684
rect 46940 4641 46949 4675
rect 46949 4641 46983 4675
rect 46983 4641 46992 4675
rect 46940 4632 46992 4641
rect 48504 4632 48556 4684
rect 50068 4768 50120 4820
rect 50344 4768 50396 4820
rect 52276 4768 52328 4820
rect 54024 4768 54076 4820
rect 56324 4811 56376 4820
rect 56324 4777 56333 4811
rect 56333 4777 56367 4811
rect 56367 4777 56376 4811
rect 56324 4768 56376 4777
rect 56508 4768 56560 4820
rect 49424 4632 49476 4684
rect 42708 4564 42760 4616
rect 44180 4564 44232 4616
rect 39212 4496 39264 4548
rect 40224 4539 40276 4548
rect 40224 4505 40233 4539
rect 40233 4505 40267 4539
rect 40267 4505 40276 4539
rect 40224 4496 40276 4505
rect 41972 4496 42024 4548
rect 42064 4496 42116 4548
rect 36084 4428 36136 4480
rect 36268 4428 36320 4480
rect 37464 4471 37516 4480
rect 37464 4437 37473 4471
rect 37473 4437 37507 4471
rect 37507 4437 37516 4471
rect 37464 4428 37516 4437
rect 38200 4471 38252 4480
rect 38200 4437 38209 4471
rect 38209 4437 38243 4471
rect 38243 4437 38252 4471
rect 38200 4428 38252 4437
rect 39856 4471 39908 4480
rect 39856 4437 39865 4471
rect 39865 4437 39899 4471
rect 39899 4437 39908 4471
rect 39856 4428 39908 4437
rect 40316 4471 40368 4480
rect 40316 4437 40325 4471
rect 40325 4437 40359 4471
rect 40359 4437 40368 4471
rect 40316 4428 40368 4437
rect 41880 4428 41932 4480
rect 45376 4564 45428 4616
rect 46020 4607 46072 4616
rect 46020 4573 46054 4607
rect 46054 4573 46072 4607
rect 47216 4607 47268 4616
rect 46020 4564 46072 4573
rect 47216 4573 47250 4607
rect 47250 4573 47268 4607
rect 47216 4564 47268 4573
rect 48412 4564 48464 4616
rect 49240 4564 49292 4616
rect 52920 4632 52972 4684
rect 53104 4675 53156 4684
rect 53104 4641 53113 4675
rect 53113 4641 53147 4675
rect 53147 4641 53156 4675
rect 53104 4632 53156 4641
rect 43628 4428 43680 4480
rect 47124 4496 47176 4548
rect 51448 4607 51500 4616
rect 51448 4573 51457 4607
rect 51457 4573 51491 4607
rect 51491 4573 51500 4607
rect 51448 4564 51500 4573
rect 50712 4496 50764 4548
rect 53288 4564 53340 4616
rect 54024 4607 54076 4616
rect 54024 4573 54033 4607
rect 54033 4573 54067 4607
rect 54067 4573 54076 4607
rect 54024 4564 54076 4573
rect 54116 4607 54168 4616
rect 54116 4573 54125 4607
rect 54125 4573 54159 4607
rect 54159 4573 54168 4607
rect 54116 4564 54168 4573
rect 56784 4675 56836 4684
rect 56784 4641 56793 4675
rect 56793 4641 56827 4675
rect 56827 4641 56836 4675
rect 56784 4632 56836 4641
rect 57060 4632 57112 4684
rect 56048 4564 56100 4616
rect 56232 4564 56284 4616
rect 45652 4428 45704 4480
rect 50160 4471 50212 4480
rect 50160 4437 50169 4471
rect 50169 4437 50203 4471
rect 50203 4437 50212 4471
rect 50160 4428 50212 4437
rect 51264 4471 51316 4480
rect 51264 4437 51273 4471
rect 51273 4437 51307 4471
rect 51307 4437 51316 4471
rect 51264 4428 51316 4437
rect 52092 4471 52144 4480
rect 52092 4437 52101 4471
rect 52101 4437 52135 4471
rect 52135 4437 52144 4471
rect 52092 4428 52144 4437
rect 55312 4471 55364 4480
rect 55312 4437 55321 4471
rect 55321 4437 55355 4471
rect 55355 4437 55364 4471
rect 55312 4428 55364 4437
rect 55772 4471 55824 4480
rect 55772 4437 55781 4471
rect 55781 4437 55815 4471
rect 55815 4437 55824 4471
rect 55772 4428 55824 4437
rect 59084 4496 59136 4548
rect 58532 4428 58584 4480
rect 15394 4326 15446 4378
rect 15458 4326 15510 4378
rect 15522 4326 15574 4378
rect 15586 4326 15638 4378
rect 15650 4326 15702 4378
rect 29838 4326 29890 4378
rect 29902 4326 29954 4378
rect 29966 4326 30018 4378
rect 30030 4326 30082 4378
rect 30094 4326 30146 4378
rect 44282 4326 44334 4378
rect 44346 4326 44398 4378
rect 44410 4326 44462 4378
rect 44474 4326 44526 4378
rect 44538 4326 44590 4378
rect 58726 4326 58778 4378
rect 58790 4326 58842 4378
rect 58854 4326 58906 4378
rect 58918 4326 58970 4378
rect 58982 4326 59034 4378
rect 3976 4224 4028 4276
rect 7840 4224 7892 4276
rect 8852 4224 8904 4276
rect 2688 4156 2740 4208
rect 3884 4199 3936 4208
rect 3884 4165 3893 4199
rect 3893 4165 3927 4199
rect 3927 4165 3936 4199
rect 3884 4156 3936 4165
rect 2964 4088 3016 4140
rect 3148 4088 3200 4140
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 6368 4156 6420 4165
rect 7932 4156 7984 4208
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 7012 4088 7064 4140
rect 9680 4224 9732 4276
rect 14280 4224 14332 4276
rect 15200 4267 15252 4276
rect 15200 4233 15209 4267
rect 15209 4233 15243 4267
rect 15243 4233 15252 4267
rect 15200 4224 15252 4233
rect 15752 4224 15804 4276
rect 10784 4156 10836 4208
rect 6276 4020 6328 4072
rect 6828 4020 6880 4072
rect 7380 4020 7432 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 11428 4088 11480 4140
rect 14832 4156 14884 4208
rect 11796 4131 11848 4140
rect 11796 4097 11830 4131
rect 11830 4097 11848 4131
rect 11796 4088 11848 4097
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 13268 4131 13320 4140
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 10140 4020 10192 4072
rect 10416 4020 10468 4072
rect 11060 4020 11112 4072
rect 14464 4020 14516 4072
rect 14556 4020 14608 4072
rect 17408 4156 17460 4208
rect 19064 4224 19116 4276
rect 21548 4224 21600 4276
rect 21824 4224 21876 4276
rect 2872 3884 2924 3936
rect 4160 3884 4212 3936
rect 4712 3884 4764 3936
rect 5908 3884 5960 3936
rect 6000 3884 6052 3936
rect 6184 3884 6236 3936
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 9588 3952 9640 4004
rect 9772 3952 9824 4004
rect 10232 3884 10284 3936
rect 10876 3927 10928 3936
rect 10876 3893 10885 3927
rect 10885 3893 10919 3927
rect 10919 3893 10928 3927
rect 10876 3884 10928 3893
rect 11704 3884 11756 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 15016 3952 15068 4004
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 17776 4088 17828 4140
rect 18144 4088 18196 4140
rect 19800 4088 19852 4140
rect 15384 4020 15436 4072
rect 16304 4020 16356 4072
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 17316 4020 17368 4072
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 19432 4020 19484 4072
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 20996 4063 21048 4072
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 21088 4063 21140 4072
rect 21088 4029 21097 4063
rect 21097 4029 21131 4063
rect 21131 4029 21140 4063
rect 21088 4020 21140 4029
rect 22100 4088 22152 4140
rect 22376 4088 22428 4140
rect 23112 4224 23164 4276
rect 23572 4224 23624 4276
rect 26424 4267 26476 4276
rect 26424 4233 26433 4267
rect 26433 4233 26467 4267
rect 26467 4233 26476 4267
rect 26424 4224 26476 4233
rect 29552 4224 29604 4276
rect 29736 4224 29788 4276
rect 21732 4020 21784 4072
rect 21916 4063 21968 4072
rect 21916 4029 21925 4063
rect 21925 4029 21959 4063
rect 21959 4029 21968 4063
rect 21916 4020 21968 4029
rect 23480 4088 23532 4140
rect 25688 4156 25740 4208
rect 26608 4156 26660 4208
rect 27344 4199 27396 4208
rect 27344 4165 27353 4199
rect 27353 4165 27387 4199
rect 27387 4165 27396 4199
rect 27344 4156 27396 4165
rect 29368 4156 29420 4208
rect 23572 4020 23624 4072
rect 24584 4088 24636 4140
rect 25320 4131 25372 4140
rect 25320 4097 25329 4131
rect 25329 4097 25363 4131
rect 25363 4097 25372 4131
rect 25320 4088 25372 4097
rect 25596 4131 25648 4140
rect 25596 4097 25605 4131
rect 25605 4097 25639 4131
rect 25639 4097 25648 4131
rect 25596 4088 25648 4097
rect 25872 4131 25924 4140
rect 25872 4097 25881 4131
rect 25881 4097 25915 4131
rect 25915 4097 25924 4131
rect 25872 4088 25924 4097
rect 26148 4020 26200 4072
rect 18328 3952 18380 4004
rect 22192 3952 22244 4004
rect 23388 3952 23440 4004
rect 26332 4020 26384 4072
rect 27252 4088 27304 4140
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 30564 4224 30616 4276
rect 31944 4267 31996 4276
rect 31944 4233 31953 4267
rect 31953 4233 31987 4267
rect 31987 4233 31996 4267
rect 31944 4224 31996 4233
rect 34060 4224 34112 4276
rect 35900 4224 35952 4276
rect 36820 4224 36872 4276
rect 37464 4224 37516 4276
rect 39212 4224 39264 4276
rect 40316 4224 40368 4276
rect 29736 4131 29788 4140
rect 29736 4097 29745 4131
rect 29745 4097 29779 4131
rect 29779 4097 29788 4131
rect 29736 4088 29788 4097
rect 36268 4156 36320 4208
rect 42064 4224 42116 4276
rect 43628 4267 43680 4276
rect 43628 4233 43637 4267
rect 43637 4233 43671 4267
rect 43671 4233 43680 4267
rect 43628 4224 43680 4233
rect 45192 4267 45244 4276
rect 45192 4233 45201 4267
rect 45201 4233 45235 4267
rect 45235 4233 45244 4267
rect 45192 4224 45244 4233
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 32220 4131 32272 4140
rect 32220 4097 32229 4131
rect 32229 4097 32263 4131
rect 32263 4097 32272 4131
rect 32220 4088 32272 4097
rect 33232 4131 33284 4140
rect 33232 4097 33241 4131
rect 33241 4097 33275 4131
rect 33275 4097 33284 4131
rect 33232 4088 33284 4097
rect 26516 3952 26568 4004
rect 27068 3952 27120 4004
rect 27896 3952 27948 4004
rect 15568 3884 15620 3936
rect 16396 3884 16448 3936
rect 17684 3884 17736 3936
rect 19156 3927 19208 3936
rect 19156 3893 19165 3927
rect 19165 3893 19199 3927
rect 19199 3893 19208 3927
rect 19156 3884 19208 3893
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 21640 3884 21692 3936
rect 23756 3884 23808 3936
rect 25136 3884 25188 3936
rect 25780 3884 25832 3936
rect 26976 3927 27028 3936
rect 26976 3893 26985 3927
rect 26985 3893 27019 3927
rect 27019 3893 27028 3927
rect 26976 3884 27028 3893
rect 27344 3927 27396 3936
rect 27344 3893 27353 3927
rect 27353 3893 27387 3927
rect 27387 3893 27396 3927
rect 27344 3884 27396 3893
rect 27804 3927 27856 3936
rect 27804 3893 27813 3927
rect 27813 3893 27847 3927
rect 27847 3893 27856 3927
rect 27804 3884 27856 3893
rect 29552 3884 29604 3936
rect 31208 4020 31260 4072
rect 31484 4020 31536 4072
rect 31852 4020 31904 4072
rect 32956 4063 33008 4072
rect 32956 4029 32965 4063
rect 32965 4029 32999 4063
rect 32999 4029 33008 4063
rect 32956 4020 33008 4029
rect 34428 4020 34480 4072
rect 35072 4063 35124 4072
rect 35072 4029 35081 4063
rect 35081 4029 35115 4063
rect 35115 4029 35124 4063
rect 35072 4020 35124 4029
rect 30748 3995 30800 4004
rect 30748 3961 30757 3995
rect 30757 3961 30791 3995
rect 30791 3961 30800 3995
rect 30748 3952 30800 3961
rect 35532 4020 35584 4072
rect 35992 4088 36044 4140
rect 38660 4088 38712 4140
rect 39028 4131 39080 4140
rect 39028 4097 39037 4131
rect 39037 4097 39071 4131
rect 39071 4097 39080 4131
rect 39028 4088 39080 4097
rect 39856 4088 39908 4140
rect 40040 4131 40092 4140
rect 40040 4097 40049 4131
rect 40049 4097 40083 4131
rect 40083 4097 40092 4131
rect 40040 4088 40092 4097
rect 37372 4063 37424 4072
rect 37372 4029 37381 4063
rect 37381 4029 37415 4063
rect 37415 4029 37424 4063
rect 37372 4020 37424 4029
rect 39764 4020 39816 4072
rect 39488 3952 39540 4004
rect 41880 4156 41932 4208
rect 41420 4131 41472 4140
rect 41420 4097 41429 4131
rect 41429 4097 41463 4131
rect 41463 4097 41472 4131
rect 41420 4088 41472 4097
rect 42340 4156 42392 4208
rect 43260 4156 43312 4208
rect 48596 4224 48648 4276
rect 49240 4224 49292 4276
rect 49424 4267 49476 4276
rect 49424 4233 49433 4267
rect 49433 4233 49467 4267
rect 49467 4233 49476 4267
rect 49424 4224 49476 4233
rect 53748 4224 53800 4276
rect 45836 4156 45888 4208
rect 54024 4156 54076 4208
rect 43168 4088 43220 4140
rect 43536 4131 43588 4140
rect 43536 4097 43545 4131
rect 43545 4097 43579 4131
rect 43579 4097 43588 4131
rect 43536 4088 43588 4097
rect 41328 4020 41380 4072
rect 33140 3884 33192 3936
rect 33600 3884 33652 3936
rect 35256 3884 35308 3936
rect 37740 3884 37792 3936
rect 40040 3884 40092 3936
rect 41604 3927 41656 3936
rect 41604 3893 41613 3927
rect 41613 3893 41647 3927
rect 41647 3893 41656 3927
rect 41604 3884 41656 3893
rect 41972 3884 42024 3936
rect 42800 4063 42852 4072
rect 42800 4029 42809 4063
rect 42809 4029 42843 4063
rect 42843 4029 42852 4063
rect 42800 4020 42852 4029
rect 42892 4063 42944 4072
rect 42892 4029 42901 4063
rect 42901 4029 42935 4063
rect 42935 4029 42944 4063
rect 42892 4020 42944 4029
rect 42984 4020 43036 4072
rect 45560 4088 45612 4140
rect 46480 4088 46532 4140
rect 47860 4131 47912 4140
rect 47860 4097 47869 4131
rect 47869 4097 47903 4131
rect 47903 4097 47912 4131
rect 47860 4088 47912 4097
rect 48228 4131 48280 4140
rect 48228 4097 48237 4131
rect 48237 4097 48271 4131
rect 48271 4097 48280 4131
rect 48228 4088 48280 4097
rect 52736 4131 52788 4140
rect 52736 4097 52745 4131
rect 52745 4097 52779 4131
rect 52779 4097 52788 4131
rect 52736 4088 52788 4097
rect 55680 4224 55732 4276
rect 44088 4020 44140 4072
rect 46020 4020 46072 4072
rect 44824 3952 44876 4004
rect 45284 3952 45336 4004
rect 42432 3927 42484 3936
rect 42432 3893 42441 3927
rect 42441 3893 42475 3927
rect 42475 3893 42484 3927
rect 42432 3884 42484 3893
rect 43076 3884 43128 3936
rect 43260 3927 43312 3936
rect 43260 3893 43269 3927
rect 43269 3893 43303 3927
rect 43303 3893 43312 3927
rect 43260 3884 43312 3893
rect 43352 3927 43404 3936
rect 43352 3893 43361 3927
rect 43361 3893 43395 3927
rect 43395 3893 43404 3927
rect 43352 3884 43404 3893
rect 43720 3884 43772 3936
rect 49332 4020 49384 4072
rect 49884 4020 49936 4072
rect 52000 4063 52052 4072
rect 52000 4029 52009 4063
rect 52009 4029 52043 4063
rect 52043 4029 52052 4063
rect 52000 4020 52052 4029
rect 47676 3927 47728 3936
rect 47676 3893 47685 3927
rect 47685 3893 47719 3927
rect 47719 3893 47728 3927
rect 47676 3884 47728 3893
rect 49516 3884 49568 3936
rect 52552 3927 52604 3936
rect 52552 3893 52561 3927
rect 52561 3893 52595 3927
rect 52595 3893 52604 3927
rect 52552 3884 52604 3893
rect 53104 3884 53156 3936
rect 54576 4020 54628 4072
rect 54116 3995 54168 4004
rect 54116 3961 54125 3995
rect 54125 3961 54159 3995
rect 54159 3961 54168 3995
rect 55496 4063 55548 4072
rect 55496 4029 55530 4063
rect 55530 4029 55548 4063
rect 55496 4020 55548 4029
rect 54116 3952 54168 3961
rect 54852 3952 54904 4004
rect 56140 3952 56192 4004
rect 56600 4224 56652 4276
rect 56416 4088 56468 4140
rect 57888 4131 57940 4140
rect 57888 4097 57897 4131
rect 57897 4097 57931 4131
rect 57931 4097 57940 4131
rect 57888 4088 57940 4097
rect 57152 4020 57204 4072
rect 57244 4063 57296 4072
rect 57244 4029 57253 4063
rect 57253 4029 57287 4063
rect 57287 4029 57296 4063
rect 57244 4020 57296 4029
rect 54208 3927 54260 3936
rect 54208 3893 54217 3927
rect 54217 3893 54251 3927
rect 54251 3893 54260 3927
rect 54208 3884 54260 3893
rect 54300 3884 54352 3936
rect 55496 3884 55548 3936
rect 55588 3884 55640 3936
rect 56324 3884 56376 3936
rect 56416 3927 56468 3936
rect 56416 3893 56425 3927
rect 56425 3893 56459 3927
rect 56459 3893 56468 3927
rect 56416 3884 56468 3893
rect 56600 3884 56652 3936
rect 57244 3884 57296 3936
rect 57612 3927 57664 3936
rect 57612 3893 57621 3927
rect 57621 3893 57655 3927
rect 57655 3893 57664 3927
rect 57612 3884 57664 3893
rect 58256 3884 58308 3936
rect 8172 3782 8224 3834
rect 8236 3782 8288 3834
rect 8300 3782 8352 3834
rect 8364 3782 8416 3834
rect 8428 3782 8480 3834
rect 22616 3782 22668 3834
rect 22680 3782 22732 3834
rect 22744 3782 22796 3834
rect 22808 3782 22860 3834
rect 22872 3782 22924 3834
rect 37060 3782 37112 3834
rect 37124 3782 37176 3834
rect 37188 3782 37240 3834
rect 37252 3782 37304 3834
rect 37316 3782 37368 3834
rect 51504 3782 51556 3834
rect 51568 3782 51620 3834
rect 51632 3782 51684 3834
rect 51696 3782 51748 3834
rect 51760 3782 51812 3834
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 5448 3680 5500 3732
rect 6644 3680 6696 3732
rect 6828 3680 6880 3732
rect 8944 3680 8996 3732
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 10140 3680 10192 3732
rect 10784 3680 10836 3732
rect 12992 3680 13044 3732
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 3976 3612 4028 3664
rect 4804 3612 4856 3664
rect 8760 3612 8812 3664
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 4252 3476 4304 3528
rect 2780 3408 2832 3460
rect 3056 3408 3108 3460
rect 3332 3408 3384 3460
rect 4712 3476 4764 3528
rect 6184 3544 6236 3596
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6460 3476 6512 3528
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 4896 3408 4948 3460
rect 5908 3408 5960 3460
rect 7380 3476 7432 3528
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9036 3476 9088 3528
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 4804 3340 4856 3392
rect 4988 3383 5040 3392
rect 4988 3349 4997 3383
rect 4997 3349 5031 3383
rect 5031 3349 5040 3383
rect 4988 3340 5040 3349
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 7748 3408 7800 3460
rect 9312 3408 9364 3460
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 11336 3408 11388 3460
rect 12532 3408 12584 3460
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 15752 3544 15804 3596
rect 15476 3519 15528 3528
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 15568 3476 15620 3528
rect 16120 3655 16172 3664
rect 16120 3621 16129 3655
rect 16129 3621 16163 3655
rect 16163 3621 16172 3655
rect 16120 3612 16172 3621
rect 17316 3723 17368 3732
rect 17316 3689 17325 3723
rect 17325 3689 17359 3723
rect 17359 3689 17368 3723
rect 17316 3680 17368 3689
rect 18328 3680 18380 3732
rect 19156 3680 19208 3732
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 20996 3680 21048 3732
rect 22284 3723 22336 3732
rect 22284 3689 22293 3723
rect 22293 3689 22327 3723
rect 22327 3689 22336 3723
rect 22284 3680 22336 3689
rect 16212 3544 16264 3596
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 21456 3655 21508 3664
rect 21456 3621 21465 3655
rect 21465 3621 21499 3655
rect 21499 3621 21508 3655
rect 21456 3612 21508 3621
rect 24308 3680 24360 3732
rect 24400 3680 24452 3732
rect 26608 3680 26660 3732
rect 26700 3723 26752 3732
rect 26700 3689 26709 3723
rect 26709 3689 26743 3723
rect 26743 3689 26752 3723
rect 26700 3680 26752 3689
rect 22744 3655 22796 3664
rect 22744 3621 22753 3655
rect 22753 3621 22787 3655
rect 22787 3621 22796 3655
rect 22744 3612 22796 3621
rect 27252 3680 27304 3732
rect 29184 3680 29236 3732
rect 22836 3587 22888 3596
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 24768 3544 24820 3596
rect 25044 3587 25096 3596
rect 25044 3553 25053 3587
rect 25053 3553 25087 3587
rect 25087 3553 25096 3587
rect 25044 3544 25096 3553
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 17500 3476 17552 3528
rect 19616 3476 19668 3528
rect 20720 3476 20772 3528
rect 17776 3408 17828 3460
rect 9864 3340 9916 3392
rect 14648 3340 14700 3392
rect 16304 3340 16356 3392
rect 16672 3340 16724 3392
rect 21364 3408 21416 3460
rect 21548 3340 21600 3392
rect 22744 3476 22796 3528
rect 25780 3544 25832 3596
rect 26240 3544 26292 3596
rect 27068 3587 27120 3596
rect 27068 3553 27077 3587
rect 27077 3553 27111 3587
rect 27111 3553 27120 3587
rect 27068 3544 27120 3553
rect 28172 3544 28224 3596
rect 26424 3476 26476 3528
rect 26884 3519 26936 3528
rect 26884 3485 26893 3519
rect 26893 3485 26927 3519
rect 26927 3485 26936 3519
rect 26884 3476 26936 3485
rect 30288 3544 30340 3596
rect 31668 3680 31720 3732
rect 31392 3612 31444 3664
rect 33600 3723 33652 3732
rect 33600 3689 33609 3723
rect 33609 3689 33643 3723
rect 33643 3689 33652 3723
rect 33600 3680 33652 3689
rect 33968 3680 34020 3732
rect 35164 3723 35216 3732
rect 35164 3689 35173 3723
rect 35173 3689 35207 3723
rect 35207 3689 35216 3723
rect 35164 3680 35216 3689
rect 35900 3680 35952 3732
rect 37556 3680 37608 3732
rect 39028 3680 39080 3732
rect 24124 3408 24176 3460
rect 26608 3451 26660 3460
rect 26608 3417 26617 3451
rect 26617 3417 26651 3451
rect 26651 3417 26660 3451
rect 26608 3408 26660 3417
rect 28356 3408 28408 3460
rect 31208 3408 31260 3460
rect 31300 3408 31352 3460
rect 24032 3340 24084 3392
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 25044 3340 25096 3392
rect 28172 3340 28224 3392
rect 28448 3383 28500 3392
rect 28448 3349 28457 3383
rect 28457 3349 28491 3383
rect 28491 3349 28500 3383
rect 28448 3340 28500 3349
rect 28540 3383 28592 3392
rect 28540 3349 28549 3383
rect 28549 3349 28583 3383
rect 28583 3349 28592 3383
rect 28540 3340 28592 3349
rect 28908 3383 28960 3392
rect 28908 3349 28917 3383
rect 28917 3349 28951 3383
rect 28951 3349 28960 3383
rect 28908 3340 28960 3349
rect 29092 3340 29144 3392
rect 30748 3340 30800 3392
rect 30840 3340 30892 3392
rect 32036 3519 32088 3528
rect 32036 3485 32045 3519
rect 32045 3485 32079 3519
rect 32079 3485 32088 3519
rect 32036 3476 32088 3485
rect 34336 3544 34388 3596
rect 39396 3612 39448 3664
rect 34796 3476 34848 3528
rect 34888 3519 34940 3528
rect 34888 3485 34897 3519
rect 34897 3485 34931 3519
rect 34931 3485 34940 3519
rect 34888 3476 34940 3485
rect 34980 3519 35032 3528
rect 34980 3485 34989 3519
rect 34989 3485 35023 3519
rect 35023 3485 35032 3519
rect 34980 3476 35032 3485
rect 35992 3476 36044 3528
rect 34244 3408 34296 3460
rect 37372 3519 37424 3528
rect 37372 3485 37381 3519
rect 37381 3485 37415 3519
rect 37415 3485 37424 3519
rect 37372 3476 37424 3485
rect 40960 3544 41012 3596
rect 42248 3544 42300 3596
rect 42708 3680 42760 3732
rect 43076 3680 43128 3732
rect 44088 3612 44140 3664
rect 44180 3544 44232 3596
rect 44456 3587 44508 3596
rect 44456 3553 44465 3587
rect 44465 3553 44499 3587
rect 44499 3553 44508 3587
rect 44456 3544 44508 3553
rect 38936 3476 38988 3528
rect 39212 3408 39264 3460
rect 33508 3340 33560 3392
rect 35624 3383 35676 3392
rect 35624 3349 35633 3383
rect 35633 3349 35667 3383
rect 35667 3349 35676 3383
rect 35624 3340 35676 3349
rect 35716 3340 35768 3392
rect 38384 3340 38436 3392
rect 43352 3476 43404 3528
rect 40224 3451 40276 3460
rect 40224 3417 40233 3451
rect 40233 3417 40267 3451
rect 40267 3417 40276 3451
rect 40224 3408 40276 3417
rect 43904 3408 43956 3460
rect 39856 3383 39908 3392
rect 39856 3349 39865 3383
rect 39865 3349 39899 3383
rect 39899 3349 39908 3383
rect 39856 3340 39908 3349
rect 41880 3340 41932 3392
rect 43720 3340 43772 3392
rect 43812 3383 43864 3392
rect 43812 3349 43821 3383
rect 43821 3349 43855 3383
rect 43855 3349 43864 3383
rect 43812 3340 43864 3349
rect 44180 3383 44232 3392
rect 44180 3349 44189 3383
rect 44189 3349 44223 3383
rect 44223 3349 44232 3383
rect 44180 3340 44232 3349
rect 44824 3680 44876 3732
rect 45836 3680 45888 3732
rect 46480 3723 46532 3732
rect 46480 3689 46489 3723
rect 46489 3689 46523 3723
rect 46523 3689 46532 3723
rect 46480 3680 46532 3689
rect 47400 3723 47452 3732
rect 47400 3689 47409 3723
rect 47409 3689 47443 3723
rect 47443 3689 47452 3723
rect 47400 3680 47452 3689
rect 47768 3680 47820 3732
rect 49424 3680 49476 3732
rect 49792 3723 49844 3732
rect 49792 3689 49801 3723
rect 49801 3689 49835 3723
rect 49835 3689 49844 3723
rect 49792 3680 49844 3689
rect 50712 3723 50764 3732
rect 50712 3689 50721 3723
rect 50721 3689 50755 3723
rect 50755 3689 50764 3723
rect 50712 3680 50764 3689
rect 47676 3612 47728 3664
rect 47584 3587 47636 3596
rect 47584 3553 47593 3587
rect 47593 3553 47627 3587
rect 47627 3553 47636 3587
rect 47584 3544 47636 3553
rect 44824 3519 44876 3528
rect 44824 3485 44833 3519
rect 44833 3485 44867 3519
rect 44867 3485 44876 3519
rect 44824 3476 44876 3485
rect 45192 3476 45244 3528
rect 48044 3519 48096 3528
rect 48044 3485 48053 3519
rect 48053 3485 48087 3519
rect 48087 3485 48096 3519
rect 48044 3476 48096 3485
rect 50528 3544 50580 3596
rect 50988 3519 51040 3528
rect 50988 3485 50997 3519
rect 50997 3485 51031 3519
rect 51031 3485 51040 3519
rect 50988 3476 51040 3485
rect 52736 3544 52788 3596
rect 54208 3680 54260 3732
rect 53840 3544 53892 3596
rect 54116 3544 54168 3596
rect 58256 3655 58308 3664
rect 58256 3621 58265 3655
rect 58265 3621 58299 3655
rect 58299 3621 58308 3655
rect 58256 3612 58308 3621
rect 56876 3587 56928 3596
rect 56876 3553 56885 3587
rect 56885 3553 56919 3587
rect 56919 3553 56928 3587
rect 56876 3544 56928 3553
rect 48320 3383 48372 3392
rect 48320 3349 48329 3383
rect 48329 3349 48363 3383
rect 48363 3349 48372 3383
rect 48320 3340 48372 3349
rect 49516 3408 49568 3460
rect 50252 3451 50304 3460
rect 50252 3417 50261 3451
rect 50261 3417 50295 3451
rect 50295 3417 50304 3451
rect 50252 3408 50304 3417
rect 50436 3408 50488 3460
rect 52552 3408 52604 3460
rect 49700 3340 49752 3392
rect 51264 3383 51316 3392
rect 51264 3349 51273 3383
rect 51273 3349 51307 3383
rect 51307 3349 51316 3383
rect 51264 3340 51316 3349
rect 55036 3476 55088 3528
rect 55312 3519 55364 3528
rect 55312 3485 55321 3519
rect 55321 3485 55355 3519
rect 55355 3485 55364 3519
rect 55312 3476 55364 3485
rect 56968 3476 57020 3528
rect 57428 3476 57480 3528
rect 52828 3383 52880 3392
rect 52828 3349 52837 3383
rect 52837 3349 52871 3383
rect 52871 3349 52880 3383
rect 52828 3340 52880 3349
rect 53288 3383 53340 3392
rect 53288 3349 53297 3383
rect 53297 3349 53331 3383
rect 53331 3349 53340 3383
rect 53288 3340 53340 3349
rect 54576 3340 54628 3392
rect 55128 3383 55180 3392
rect 55128 3349 55137 3383
rect 55137 3349 55171 3383
rect 55171 3349 55180 3383
rect 55128 3340 55180 3349
rect 15394 3238 15446 3290
rect 15458 3238 15510 3290
rect 15522 3238 15574 3290
rect 15586 3238 15638 3290
rect 15650 3238 15702 3290
rect 29838 3238 29890 3290
rect 29902 3238 29954 3290
rect 29966 3238 30018 3290
rect 30030 3238 30082 3290
rect 30094 3238 30146 3290
rect 44282 3238 44334 3290
rect 44346 3238 44398 3290
rect 44410 3238 44462 3290
rect 44474 3238 44526 3290
rect 44538 3238 44590 3290
rect 58726 3238 58778 3290
rect 58790 3238 58842 3290
rect 58854 3238 58906 3290
rect 58918 3238 58970 3290
rect 58982 3238 59034 3290
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 2780 3136 2832 3145
rect 2596 3068 2648 3120
rect 4620 3136 4672 3188
rect 4712 3136 4764 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7748 3179 7800 3188
rect 7748 3145 7757 3179
rect 7757 3145 7791 3179
rect 7791 3145 7800 3179
rect 7748 3136 7800 3145
rect 8024 3136 8076 3188
rect 9220 3136 9272 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10876 3136 10928 3188
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 11520 3136 11572 3188
rect 11612 3136 11664 3188
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 14648 3179 14700 3188
rect 14648 3145 14657 3179
rect 14657 3145 14691 3179
rect 14691 3145 14700 3179
rect 14648 3136 14700 3145
rect 16120 3136 16172 3188
rect 16856 3136 16908 3188
rect 17684 3136 17736 3188
rect 17776 3136 17828 3188
rect 20536 3136 20588 3188
rect 21364 3179 21416 3188
rect 21364 3145 21373 3179
rect 21373 3145 21407 3179
rect 21407 3145 21416 3179
rect 21364 3136 21416 3145
rect 21548 3136 21600 3188
rect 21640 3136 21692 3188
rect 21732 3136 21784 3188
rect 23112 3136 23164 3188
rect 23388 3179 23440 3188
rect 23388 3145 23397 3179
rect 23397 3145 23431 3179
rect 23431 3145 23440 3179
rect 23388 3136 23440 3145
rect 24124 3179 24176 3188
rect 24124 3145 24133 3179
rect 24133 3145 24167 3179
rect 24167 3145 24176 3179
rect 24124 3136 24176 3145
rect 24400 3136 24452 3188
rect 26884 3136 26936 3188
rect 28356 3179 28408 3188
rect 28356 3145 28365 3179
rect 28365 3145 28399 3179
rect 28399 3145 28408 3179
rect 28356 3136 28408 3145
rect 28540 3136 28592 3188
rect 28908 3136 28960 3188
rect 29552 3136 29604 3188
rect 30840 3136 30892 3188
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 3976 3000 4028 3052
rect 5356 3000 5408 3052
rect 5908 3000 5960 3052
rect 4804 2975 4856 2984
rect 4804 2941 4813 2975
rect 4813 2941 4847 2975
rect 4847 2941 4856 2975
rect 4804 2932 4856 2941
rect 4344 2864 4396 2916
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 13912 3068 13964 3120
rect 13268 3043 13320 3052
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 14740 3043 14792 3052
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 16396 3043 16448 3052
rect 16396 3009 16405 3043
rect 16405 3009 16439 3043
rect 16439 3009 16448 3043
rect 16396 3000 16448 3009
rect 16672 3000 16724 3052
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 17040 3000 17092 3052
rect 20168 3068 20220 3120
rect 18144 3000 18196 3052
rect 7012 2932 7064 2984
rect 3608 2796 3660 2848
rect 3700 2796 3752 2848
rect 8760 2975 8812 2984
rect 8760 2941 8769 2975
rect 8769 2941 8803 2975
rect 8803 2941 8812 2975
rect 8760 2932 8812 2941
rect 9312 2864 9364 2916
rect 4712 2796 4764 2848
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 6828 2796 6880 2848
rect 10508 2975 10560 2984
rect 10508 2941 10517 2975
rect 10517 2941 10551 2975
rect 10551 2941 10560 2975
rect 10508 2932 10560 2941
rect 12532 2932 12584 2984
rect 14280 2932 14332 2984
rect 13268 2864 13320 2916
rect 14924 2864 14976 2916
rect 16764 2932 16816 2984
rect 20904 3000 20956 3052
rect 21364 3000 21416 3052
rect 27712 3068 27764 3120
rect 23756 3000 23808 3052
rect 25688 3043 25740 3052
rect 25688 3009 25697 3043
rect 25697 3009 25731 3043
rect 25731 3009 25740 3043
rect 25688 3000 25740 3009
rect 25872 3043 25924 3052
rect 25872 3009 25881 3043
rect 25881 3009 25915 3043
rect 25915 3009 25924 3043
rect 25872 3000 25924 3009
rect 31116 3136 31168 3188
rect 31484 3136 31536 3188
rect 31852 3136 31904 3188
rect 32312 3179 32364 3188
rect 32312 3145 32321 3179
rect 32321 3145 32355 3179
rect 32355 3145 32364 3179
rect 32312 3136 32364 3145
rect 18512 2864 18564 2916
rect 18972 2907 19024 2916
rect 18972 2873 18981 2907
rect 18981 2873 19015 2907
rect 19015 2873 19024 2907
rect 18972 2864 19024 2873
rect 19156 2864 19208 2916
rect 24124 2932 24176 2984
rect 26884 2932 26936 2984
rect 28356 2932 28408 2984
rect 28448 2975 28500 2984
rect 28448 2941 28457 2975
rect 28457 2941 28491 2975
rect 28491 2941 28500 2975
rect 28448 2932 28500 2941
rect 29092 2932 29144 2984
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 29276 2864 29328 2916
rect 30932 3000 30984 3052
rect 31484 2975 31536 2984
rect 31484 2941 31493 2975
rect 31493 2941 31527 2975
rect 31527 2941 31536 2975
rect 31484 2932 31536 2941
rect 31668 3000 31720 3052
rect 34244 3136 34296 3188
rect 37372 3136 37424 3188
rect 37464 3136 37516 3188
rect 36268 3068 36320 3120
rect 37740 3068 37792 3120
rect 34060 3000 34112 3052
rect 34612 3043 34664 3052
rect 34612 3009 34621 3043
rect 34621 3009 34655 3043
rect 34655 3009 34664 3043
rect 34612 3000 34664 3009
rect 32864 2975 32916 2984
rect 32864 2941 32873 2975
rect 32873 2941 32907 2975
rect 32907 2941 32916 2975
rect 32864 2932 32916 2941
rect 32956 2864 33008 2916
rect 33140 2975 33192 2984
rect 33140 2941 33149 2975
rect 33149 2941 33183 2975
rect 33183 2941 33192 2975
rect 33140 2932 33192 2941
rect 35348 2975 35400 2984
rect 35348 2941 35357 2975
rect 35357 2941 35391 2975
rect 35391 2941 35400 2975
rect 35348 2932 35400 2941
rect 23480 2796 23532 2848
rect 31760 2839 31812 2848
rect 31760 2805 31769 2839
rect 31769 2805 31803 2839
rect 31803 2805 31812 2839
rect 31760 2796 31812 2805
rect 33508 2864 33560 2916
rect 36176 3000 36228 3052
rect 37832 3000 37884 3052
rect 38936 3179 38988 3188
rect 38936 3145 38945 3179
rect 38945 3145 38979 3179
rect 38979 3145 38988 3179
rect 38936 3136 38988 3145
rect 39212 3136 39264 3188
rect 39856 3136 39908 3188
rect 40592 3179 40644 3188
rect 40592 3145 40601 3179
rect 40601 3145 40635 3179
rect 40635 3145 40644 3179
rect 40592 3136 40644 3145
rect 34428 2796 34480 2848
rect 36636 2864 36688 2916
rect 37648 2932 37700 2984
rect 39948 3068 40000 3120
rect 36820 2864 36872 2916
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 35992 2796 36044 2805
rect 36268 2796 36320 2848
rect 37464 2796 37516 2848
rect 41604 3136 41656 3188
rect 43536 3136 43588 3188
rect 43812 3136 43864 3188
rect 43904 3179 43956 3188
rect 43904 3145 43913 3179
rect 43913 3145 43947 3179
rect 43947 3145 43956 3179
rect 43904 3136 43956 3145
rect 45560 3136 45612 3188
rect 47032 3136 47084 3188
rect 47860 3136 47912 3188
rect 45100 3068 45152 3120
rect 45284 3068 45336 3120
rect 40684 2932 40736 2984
rect 41788 2932 41840 2984
rect 43996 2932 44048 2984
rect 44824 3000 44876 3052
rect 46388 3043 46440 3052
rect 46388 3009 46397 3043
rect 46397 3009 46431 3043
rect 46431 3009 46440 3043
rect 46388 3000 46440 3009
rect 46480 3043 46532 3052
rect 46480 3009 46489 3043
rect 46489 3009 46523 3043
rect 46523 3009 46532 3043
rect 46480 3000 46532 3009
rect 46756 3043 46808 3052
rect 46756 3009 46765 3043
rect 46765 3009 46799 3043
rect 46799 3009 46808 3043
rect 46756 3000 46808 3009
rect 48044 3068 48096 3120
rect 51080 3136 51132 3188
rect 52552 3136 52604 3188
rect 52828 3136 52880 3188
rect 54392 3136 54444 3188
rect 54576 3136 54628 3188
rect 55772 3136 55824 3188
rect 56324 3136 56376 3188
rect 57428 3136 57480 3188
rect 57612 3136 57664 3188
rect 57980 3136 58032 3188
rect 47124 3043 47176 3052
rect 47124 3009 47133 3043
rect 47133 3009 47167 3043
rect 47167 3009 47176 3043
rect 47124 3000 47176 3009
rect 50160 3068 50212 3120
rect 45100 2932 45152 2984
rect 46848 2932 46900 2984
rect 44732 2864 44784 2916
rect 47860 2932 47912 2984
rect 49240 2932 49292 2984
rect 50068 2932 50120 2984
rect 52460 3000 52512 3052
rect 41144 2796 41196 2848
rect 41880 2796 41932 2848
rect 41972 2796 42024 2848
rect 47676 2796 47728 2848
rect 51908 2975 51960 2984
rect 51908 2941 51917 2975
rect 51917 2941 51951 2975
rect 51951 2941 51960 2975
rect 51908 2932 51960 2941
rect 53656 3043 53708 3052
rect 53656 3009 53665 3043
rect 53665 3009 53699 3043
rect 53699 3009 53708 3043
rect 53656 3000 53708 3009
rect 54208 2932 54260 2984
rect 57244 2975 57296 2984
rect 57244 2941 57253 2975
rect 57253 2941 57287 2975
rect 57287 2941 57296 2975
rect 57244 2932 57296 2941
rect 55036 2864 55088 2916
rect 51172 2839 51224 2848
rect 51172 2805 51181 2839
rect 51181 2805 51215 2839
rect 51215 2805 51224 2839
rect 51172 2796 51224 2805
rect 52460 2796 52512 2848
rect 55404 2796 55456 2848
rect 8172 2694 8224 2746
rect 8236 2694 8288 2746
rect 8300 2694 8352 2746
rect 8364 2694 8416 2746
rect 8428 2694 8480 2746
rect 22616 2694 22668 2746
rect 22680 2694 22732 2746
rect 22744 2694 22796 2746
rect 22808 2694 22860 2746
rect 22872 2694 22924 2746
rect 37060 2694 37112 2746
rect 37124 2694 37176 2746
rect 37188 2694 37240 2746
rect 37252 2694 37304 2746
rect 37316 2694 37368 2746
rect 51504 2694 51556 2746
rect 51568 2694 51620 2746
rect 51632 2694 51684 2746
rect 51696 2694 51748 2746
rect 51760 2694 51812 2746
rect 3608 2592 3660 2644
rect 2688 2524 2740 2576
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 4988 2592 5040 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 9036 2592 9088 2644
rect 11152 2592 11204 2644
rect 14740 2592 14792 2644
rect 16396 2592 16448 2644
rect 16856 2592 16908 2644
rect 20168 2635 20220 2644
rect 20168 2601 20177 2635
rect 20177 2601 20211 2635
rect 20211 2601 20220 2635
rect 20168 2592 20220 2601
rect 22100 2592 22152 2644
rect 24032 2635 24084 2644
rect 24032 2601 24041 2635
rect 24041 2601 24075 2635
rect 24075 2601 24084 2635
rect 24032 2592 24084 2601
rect 24400 2635 24452 2644
rect 24400 2601 24409 2635
rect 24409 2601 24443 2635
rect 24443 2601 24452 2635
rect 24400 2592 24452 2601
rect 25596 2592 25648 2644
rect 27068 2635 27120 2644
rect 27068 2601 27077 2635
rect 27077 2601 27111 2635
rect 27111 2601 27120 2635
rect 27068 2592 27120 2601
rect 27436 2635 27488 2644
rect 27436 2601 27445 2635
rect 27445 2601 27479 2635
rect 27479 2601 27488 2635
rect 27436 2592 27488 2601
rect 29000 2592 29052 2644
rect 31576 2592 31628 2644
rect 34796 2592 34848 2644
rect 34980 2592 35032 2644
rect 38660 2592 38712 2644
rect 39488 2635 39540 2644
rect 39488 2601 39497 2635
rect 39497 2601 39531 2635
rect 39531 2601 39540 2635
rect 39488 2592 39540 2601
rect 41512 2592 41564 2644
rect 44180 2592 44232 2644
rect 45560 2592 45612 2644
rect 47400 2592 47452 2644
rect 49700 2592 49752 2644
rect 50252 2635 50304 2644
rect 50252 2601 50261 2635
rect 50261 2601 50295 2635
rect 50295 2601 50304 2635
rect 50252 2592 50304 2601
rect 52736 2592 52788 2644
rect 53288 2592 53340 2644
rect 55312 2592 55364 2644
rect 56416 2592 56468 2644
rect 58532 2635 58584 2644
rect 58532 2601 58541 2635
rect 58541 2601 58575 2635
rect 58575 2601 58584 2635
rect 58532 2592 58584 2601
rect 4528 2524 4580 2576
rect 2044 2456 2096 2508
rect 15752 2524 15804 2576
rect 22284 2524 22336 2576
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5908 2388 5960 2440
rect 1676 2363 1728 2372
rect 1676 2329 1685 2363
rect 1685 2329 1719 2363
rect 1719 2329 1728 2363
rect 1676 2320 1728 2329
rect 4160 2363 4212 2372
rect 4160 2329 4169 2363
rect 4169 2329 4203 2363
rect 4203 2329 4212 2363
rect 4160 2320 4212 2329
rect 5264 2320 5316 2372
rect 7196 2388 7248 2440
rect 7564 2456 7616 2508
rect 9956 2456 10008 2508
rect 11612 2499 11664 2508
rect 11612 2465 11621 2499
rect 11621 2465 11655 2499
rect 11655 2465 11664 2499
rect 11612 2456 11664 2465
rect 8760 2388 8812 2440
rect 8392 2320 8444 2372
rect 9772 2388 9824 2440
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 12348 2456 12400 2508
rect 15844 2499 15896 2508
rect 15844 2465 15853 2499
rect 15853 2465 15887 2499
rect 15887 2465 15896 2499
rect 15844 2456 15896 2465
rect 17868 2456 17920 2508
rect 14004 2388 14056 2440
rect 11152 2320 11204 2372
rect 14740 2320 14792 2372
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16580 2320 16632 2372
rect 18236 2388 18288 2440
rect 19340 2388 19392 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20076 2388 20128 2440
rect 20812 2499 20864 2508
rect 20812 2465 20821 2499
rect 20821 2465 20855 2499
rect 20855 2465 20864 2499
rect 20812 2456 20864 2465
rect 22468 2456 22520 2508
rect 25872 2499 25924 2508
rect 25872 2465 25881 2499
rect 25881 2465 25915 2499
rect 25915 2465 25924 2499
rect 25872 2456 25924 2465
rect 27436 2456 27488 2508
rect 21916 2431 21968 2440
rect 21916 2397 21925 2431
rect 21925 2397 21959 2431
rect 21959 2397 21968 2431
rect 21916 2388 21968 2397
rect 22192 2388 22244 2440
rect 23388 2388 23440 2440
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25228 2388 25280 2440
rect 25320 2388 25372 2440
rect 27528 2388 27580 2440
rect 27712 2431 27764 2440
rect 27712 2397 27721 2431
rect 27721 2397 27755 2431
rect 27755 2397 27764 2431
rect 27712 2388 27764 2397
rect 30748 2456 30800 2508
rect 31760 2456 31812 2508
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 30196 2388 30248 2440
rect 30656 2431 30708 2440
rect 30656 2397 30665 2431
rect 30665 2397 30699 2431
rect 30699 2397 30708 2431
rect 30656 2388 30708 2397
rect 35992 2524 36044 2576
rect 32680 2456 32732 2508
rect 18604 2320 18656 2372
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 35624 2456 35676 2508
rect 35716 2456 35768 2508
rect 38752 2499 38804 2508
rect 38752 2465 38761 2499
rect 38761 2465 38795 2499
rect 38795 2465 38804 2499
rect 38752 2456 38804 2465
rect 39028 2456 39080 2508
rect 42616 2456 42668 2508
rect 44088 2499 44140 2508
rect 44088 2465 44097 2499
rect 44097 2465 44131 2499
rect 44131 2465 44140 2499
rect 44088 2456 44140 2465
rect 45652 2456 45704 2508
rect 47492 2456 47544 2508
rect 50620 2456 50672 2508
rect 52368 2456 52420 2508
rect 55588 2456 55640 2508
rect 36176 2431 36228 2440
rect 36176 2397 36185 2431
rect 36185 2397 36219 2431
rect 36219 2397 36228 2431
rect 36176 2388 36228 2397
rect 34428 2320 34480 2372
rect 37556 2388 37608 2440
rect 34060 2252 34112 2304
rect 34796 2252 34848 2304
rect 38016 2320 38068 2372
rect 40040 2388 40092 2440
rect 40132 2388 40184 2440
rect 43260 2388 43312 2440
rect 43904 2320 43956 2372
rect 47124 2388 47176 2440
rect 46204 2320 46256 2372
rect 48320 2388 48372 2440
rect 48412 2388 48464 2440
rect 49700 2388 49752 2440
rect 51080 2388 51132 2440
rect 51172 2388 51224 2440
rect 52460 2388 52512 2440
rect 54944 2388 54996 2440
rect 55404 2431 55456 2440
rect 55404 2397 55413 2431
rect 55413 2397 55447 2431
rect 55447 2397 55456 2431
rect 55404 2388 55456 2397
rect 57152 2431 57204 2440
rect 57152 2397 57161 2431
rect 57161 2397 57195 2431
rect 57195 2397 57204 2431
rect 57152 2388 57204 2397
rect 57888 2499 57940 2508
rect 57888 2465 57897 2499
rect 57897 2465 57931 2499
rect 57931 2465 57940 2499
rect 57888 2456 57940 2465
rect 35808 2252 35860 2304
rect 53196 2252 53248 2304
rect 15394 2150 15446 2202
rect 15458 2150 15510 2202
rect 15522 2150 15574 2202
rect 15586 2150 15638 2202
rect 15650 2150 15702 2202
rect 29838 2150 29890 2202
rect 29902 2150 29954 2202
rect 29966 2150 30018 2202
rect 30030 2150 30082 2202
rect 30094 2150 30146 2202
rect 44282 2150 44334 2202
rect 44346 2150 44398 2202
rect 44410 2150 44462 2202
rect 44474 2150 44526 2202
rect 44538 2150 44590 2202
rect 58726 2150 58778 2202
rect 58790 2150 58842 2202
rect 58854 2150 58906 2202
rect 58918 2150 58970 2202
rect 58982 2150 59034 2202
rect 32036 2048 32088 2100
rect 34060 2048 34112 2100
rect 38200 2048 38252 2100
rect 35808 1980 35860 2032
rect 31852 1504 31904 1556
rect 35348 1504 35400 1556
<< metal2 >>
rect 8172 27772 8480 27781
rect 8172 27770 8178 27772
rect 8234 27770 8258 27772
rect 8314 27770 8338 27772
rect 8394 27770 8418 27772
rect 8474 27770 8480 27772
rect 8234 27718 8236 27770
rect 8416 27718 8418 27770
rect 8172 27716 8178 27718
rect 8234 27716 8258 27718
rect 8314 27716 8338 27718
rect 8394 27716 8418 27718
rect 8474 27716 8480 27718
rect 8172 27707 8480 27716
rect 22616 27772 22924 27781
rect 22616 27770 22622 27772
rect 22678 27770 22702 27772
rect 22758 27770 22782 27772
rect 22838 27770 22862 27772
rect 22918 27770 22924 27772
rect 22678 27718 22680 27770
rect 22860 27718 22862 27770
rect 22616 27716 22622 27718
rect 22678 27716 22702 27718
rect 22758 27716 22782 27718
rect 22838 27716 22862 27718
rect 22918 27716 22924 27718
rect 22616 27707 22924 27716
rect 37060 27772 37368 27781
rect 37060 27770 37066 27772
rect 37122 27770 37146 27772
rect 37202 27770 37226 27772
rect 37282 27770 37306 27772
rect 37362 27770 37368 27772
rect 37122 27718 37124 27770
rect 37304 27718 37306 27770
rect 37060 27716 37066 27718
rect 37122 27716 37146 27718
rect 37202 27716 37226 27718
rect 37282 27716 37306 27718
rect 37362 27716 37368 27718
rect 37060 27707 37368 27716
rect 51504 27772 51812 27781
rect 51504 27770 51510 27772
rect 51566 27770 51590 27772
rect 51646 27770 51670 27772
rect 51726 27770 51750 27772
rect 51806 27770 51812 27772
rect 51566 27718 51568 27770
rect 51748 27718 51750 27770
rect 51504 27716 51510 27718
rect 51566 27716 51590 27718
rect 51646 27716 51670 27718
rect 51726 27716 51750 27718
rect 51806 27716 51812 27718
rect 51504 27707 51812 27716
rect 15394 27228 15702 27237
rect 15394 27226 15400 27228
rect 15456 27226 15480 27228
rect 15536 27226 15560 27228
rect 15616 27226 15640 27228
rect 15696 27226 15702 27228
rect 15456 27174 15458 27226
rect 15638 27174 15640 27226
rect 15394 27172 15400 27174
rect 15456 27172 15480 27174
rect 15536 27172 15560 27174
rect 15616 27172 15640 27174
rect 15696 27172 15702 27174
rect 15394 27163 15702 27172
rect 29838 27228 30146 27237
rect 29838 27226 29844 27228
rect 29900 27226 29924 27228
rect 29980 27226 30004 27228
rect 30060 27226 30084 27228
rect 30140 27226 30146 27228
rect 29900 27174 29902 27226
rect 30082 27174 30084 27226
rect 29838 27172 29844 27174
rect 29900 27172 29924 27174
rect 29980 27172 30004 27174
rect 30060 27172 30084 27174
rect 30140 27172 30146 27174
rect 29838 27163 30146 27172
rect 44282 27228 44590 27237
rect 44282 27226 44288 27228
rect 44344 27226 44368 27228
rect 44424 27226 44448 27228
rect 44504 27226 44528 27228
rect 44584 27226 44590 27228
rect 44344 27174 44346 27226
rect 44526 27174 44528 27226
rect 44282 27172 44288 27174
rect 44344 27172 44368 27174
rect 44424 27172 44448 27174
rect 44504 27172 44528 27174
rect 44584 27172 44590 27174
rect 44282 27163 44590 27172
rect 58726 27228 59034 27237
rect 58726 27226 58732 27228
rect 58788 27226 58812 27228
rect 58868 27226 58892 27228
rect 58948 27226 58972 27228
rect 59028 27226 59034 27228
rect 58788 27174 58790 27226
rect 58970 27174 58972 27226
rect 58726 27172 58732 27174
rect 58788 27172 58812 27174
rect 58868 27172 58892 27174
rect 58948 27172 58972 27174
rect 59028 27172 59034 27174
rect 58726 27163 59034 27172
rect 8172 26684 8480 26693
rect 8172 26682 8178 26684
rect 8234 26682 8258 26684
rect 8314 26682 8338 26684
rect 8394 26682 8418 26684
rect 8474 26682 8480 26684
rect 8234 26630 8236 26682
rect 8416 26630 8418 26682
rect 8172 26628 8178 26630
rect 8234 26628 8258 26630
rect 8314 26628 8338 26630
rect 8394 26628 8418 26630
rect 8474 26628 8480 26630
rect 8172 26619 8480 26628
rect 22616 26684 22924 26693
rect 22616 26682 22622 26684
rect 22678 26682 22702 26684
rect 22758 26682 22782 26684
rect 22838 26682 22862 26684
rect 22918 26682 22924 26684
rect 22678 26630 22680 26682
rect 22860 26630 22862 26682
rect 22616 26628 22622 26630
rect 22678 26628 22702 26630
rect 22758 26628 22782 26630
rect 22838 26628 22862 26630
rect 22918 26628 22924 26630
rect 22616 26619 22924 26628
rect 37060 26684 37368 26693
rect 37060 26682 37066 26684
rect 37122 26682 37146 26684
rect 37202 26682 37226 26684
rect 37282 26682 37306 26684
rect 37362 26682 37368 26684
rect 37122 26630 37124 26682
rect 37304 26630 37306 26682
rect 37060 26628 37066 26630
rect 37122 26628 37146 26630
rect 37202 26628 37226 26630
rect 37282 26628 37306 26630
rect 37362 26628 37368 26630
rect 37060 26619 37368 26628
rect 51504 26684 51812 26693
rect 51504 26682 51510 26684
rect 51566 26682 51590 26684
rect 51646 26682 51670 26684
rect 51726 26682 51750 26684
rect 51806 26682 51812 26684
rect 51566 26630 51568 26682
rect 51748 26630 51750 26682
rect 51504 26628 51510 26630
rect 51566 26628 51590 26630
rect 51646 26628 51670 26630
rect 51726 26628 51750 26630
rect 51806 26628 51812 26630
rect 51504 26619 51812 26628
rect 15394 26140 15702 26149
rect 15394 26138 15400 26140
rect 15456 26138 15480 26140
rect 15536 26138 15560 26140
rect 15616 26138 15640 26140
rect 15696 26138 15702 26140
rect 15456 26086 15458 26138
rect 15638 26086 15640 26138
rect 15394 26084 15400 26086
rect 15456 26084 15480 26086
rect 15536 26084 15560 26086
rect 15616 26084 15640 26086
rect 15696 26084 15702 26086
rect 15394 26075 15702 26084
rect 29838 26140 30146 26149
rect 29838 26138 29844 26140
rect 29900 26138 29924 26140
rect 29980 26138 30004 26140
rect 30060 26138 30084 26140
rect 30140 26138 30146 26140
rect 29900 26086 29902 26138
rect 30082 26086 30084 26138
rect 29838 26084 29844 26086
rect 29900 26084 29924 26086
rect 29980 26084 30004 26086
rect 30060 26084 30084 26086
rect 30140 26084 30146 26086
rect 29838 26075 30146 26084
rect 44282 26140 44590 26149
rect 44282 26138 44288 26140
rect 44344 26138 44368 26140
rect 44424 26138 44448 26140
rect 44504 26138 44528 26140
rect 44584 26138 44590 26140
rect 44344 26086 44346 26138
rect 44526 26086 44528 26138
rect 44282 26084 44288 26086
rect 44344 26084 44368 26086
rect 44424 26084 44448 26086
rect 44504 26084 44528 26086
rect 44584 26084 44590 26086
rect 44282 26075 44590 26084
rect 58726 26140 59034 26149
rect 58726 26138 58732 26140
rect 58788 26138 58812 26140
rect 58868 26138 58892 26140
rect 58948 26138 58972 26140
rect 59028 26138 59034 26140
rect 58788 26086 58790 26138
rect 58970 26086 58972 26138
rect 58726 26084 58732 26086
rect 58788 26084 58812 26086
rect 58868 26084 58892 26086
rect 58948 26084 58972 26086
rect 59028 26084 59034 26086
rect 58726 26075 59034 26084
rect 8172 25596 8480 25605
rect 8172 25594 8178 25596
rect 8234 25594 8258 25596
rect 8314 25594 8338 25596
rect 8394 25594 8418 25596
rect 8474 25594 8480 25596
rect 8234 25542 8236 25594
rect 8416 25542 8418 25594
rect 8172 25540 8178 25542
rect 8234 25540 8258 25542
rect 8314 25540 8338 25542
rect 8394 25540 8418 25542
rect 8474 25540 8480 25542
rect 8172 25531 8480 25540
rect 22616 25596 22924 25605
rect 22616 25594 22622 25596
rect 22678 25594 22702 25596
rect 22758 25594 22782 25596
rect 22838 25594 22862 25596
rect 22918 25594 22924 25596
rect 22678 25542 22680 25594
rect 22860 25542 22862 25594
rect 22616 25540 22622 25542
rect 22678 25540 22702 25542
rect 22758 25540 22782 25542
rect 22838 25540 22862 25542
rect 22918 25540 22924 25542
rect 22616 25531 22924 25540
rect 37060 25596 37368 25605
rect 37060 25594 37066 25596
rect 37122 25594 37146 25596
rect 37202 25594 37226 25596
rect 37282 25594 37306 25596
rect 37362 25594 37368 25596
rect 37122 25542 37124 25594
rect 37304 25542 37306 25594
rect 37060 25540 37066 25542
rect 37122 25540 37146 25542
rect 37202 25540 37226 25542
rect 37282 25540 37306 25542
rect 37362 25540 37368 25542
rect 37060 25531 37368 25540
rect 51504 25596 51812 25605
rect 51504 25594 51510 25596
rect 51566 25594 51590 25596
rect 51646 25594 51670 25596
rect 51726 25594 51750 25596
rect 51806 25594 51812 25596
rect 51566 25542 51568 25594
rect 51748 25542 51750 25594
rect 51504 25540 51510 25542
rect 51566 25540 51590 25542
rect 51646 25540 51670 25542
rect 51726 25540 51750 25542
rect 51806 25540 51812 25542
rect 51504 25531 51812 25540
rect 15394 25052 15702 25061
rect 15394 25050 15400 25052
rect 15456 25050 15480 25052
rect 15536 25050 15560 25052
rect 15616 25050 15640 25052
rect 15696 25050 15702 25052
rect 15456 24998 15458 25050
rect 15638 24998 15640 25050
rect 15394 24996 15400 24998
rect 15456 24996 15480 24998
rect 15536 24996 15560 24998
rect 15616 24996 15640 24998
rect 15696 24996 15702 24998
rect 15394 24987 15702 24996
rect 29838 25052 30146 25061
rect 29838 25050 29844 25052
rect 29900 25050 29924 25052
rect 29980 25050 30004 25052
rect 30060 25050 30084 25052
rect 30140 25050 30146 25052
rect 29900 24998 29902 25050
rect 30082 24998 30084 25050
rect 29838 24996 29844 24998
rect 29900 24996 29924 24998
rect 29980 24996 30004 24998
rect 30060 24996 30084 24998
rect 30140 24996 30146 24998
rect 29838 24987 30146 24996
rect 44282 25052 44590 25061
rect 44282 25050 44288 25052
rect 44344 25050 44368 25052
rect 44424 25050 44448 25052
rect 44504 25050 44528 25052
rect 44584 25050 44590 25052
rect 44344 24998 44346 25050
rect 44526 24998 44528 25050
rect 44282 24996 44288 24998
rect 44344 24996 44368 24998
rect 44424 24996 44448 24998
rect 44504 24996 44528 24998
rect 44584 24996 44590 24998
rect 44282 24987 44590 24996
rect 58726 25052 59034 25061
rect 58726 25050 58732 25052
rect 58788 25050 58812 25052
rect 58868 25050 58892 25052
rect 58948 25050 58972 25052
rect 59028 25050 59034 25052
rect 58788 24998 58790 25050
rect 58970 24998 58972 25050
rect 58726 24996 58732 24998
rect 58788 24996 58812 24998
rect 58868 24996 58892 24998
rect 58948 24996 58972 24998
rect 59028 24996 59034 24998
rect 58726 24987 59034 24996
rect 8172 24508 8480 24517
rect 8172 24506 8178 24508
rect 8234 24506 8258 24508
rect 8314 24506 8338 24508
rect 8394 24506 8418 24508
rect 8474 24506 8480 24508
rect 8234 24454 8236 24506
rect 8416 24454 8418 24506
rect 8172 24452 8178 24454
rect 8234 24452 8258 24454
rect 8314 24452 8338 24454
rect 8394 24452 8418 24454
rect 8474 24452 8480 24454
rect 8172 24443 8480 24452
rect 22616 24508 22924 24517
rect 22616 24506 22622 24508
rect 22678 24506 22702 24508
rect 22758 24506 22782 24508
rect 22838 24506 22862 24508
rect 22918 24506 22924 24508
rect 22678 24454 22680 24506
rect 22860 24454 22862 24506
rect 22616 24452 22622 24454
rect 22678 24452 22702 24454
rect 22758 24452 22782 24454
rect 22838 24452 22862 24454
rect 22918 24452 22924 24454
rect 22616 24443 22924 24452
rect 37060 24508 37368 24517
rect 37060 24506 37066 24508
rect 37122 24506 37146 24508
rect 37202 24506 37226 24508
rect 37282 24506 37306 24508
rect 37362 24506 37368 24508
rect 37122 24454 37124 24506
rect 37304 24454 37306 24506
rect 37060 24452 37066 24454
rect 37122 24452 37146 24454
rect 37202 24452 37226 24454
rect 37282 24452 37306 24454
rect 37362 24452 37368 24454
rect 37060 24443 37368 24452
rect 51504 24508 51812 24517
rect 51504 24506 51510 24508
rect 51566 24506 51590 24508
rect 51646 24506 51670 24508
rect 51726 24506 51750 24508
rect 51806 24506 51812 24508
rect 51566 24454 51568 24506
rect 51748 24454 51750 24506
rect 51504 24452 51510 24454
rect 51566 24452 51590 24454
rect 51646 24452 51670 24454
rect 51726 24452 51750 24454
rect 51806 24452 51812 24454
rect 51504 24443 51812 24452
rect 15394 23964 15702 23973
rect 15394 23962 15400 23964
rect 15456 23962 15480 23964
rect 15536 23962 15560 23964
rect 15616 23962 15640 23964
rect 15696 23962 15702 23964
rect 15456 23910 15458 23962
rect 15638 23910 15640 23962
rect 15394 23908 15400 23910
rect 15456 23908 15480 23910
rect 15536 23908 15560 23910
rect 15616 23908 15640 23910
rect 15696 23908 15702 23910
rect 15394 23899 15702 23908
rect 29838 23964 30146 23973
rect 29838 23962 29844 23964
rect 29900 23962 29924 23964
rect 29980 23962 30004 23964
rect 30060 23962 30084 23964
rect 30140 23962 30146 23964
rect 29900 23910 29902 23962
rect 30082 23910 30084 23962
rect 29838 23908 29844 23910
rect 29900 23908 29924 23910
rect 29980 23908 30004 23910
rect 30060 23908 30084 23910
rect 30140 23908 30146 23910
rect 29838 23899 30146 23908
rect 44282 23964 44590 23973
rect 44282 23962 44288 23964
rect 44344 23962 44368 23964
rect 44424 23962 44448 23964
rect 44504 23962 44528 23964
rect 44584 23962 44590 23964
rect 44344 23910 44346 23962
rect 44526 23910 44528 23962
rect 44282 23908 44288 23910
rect 44344 23908 44368 23910
rect 44424 23908 44448 23910
rect 44504 23908 44528 23910
rect 44584 23908 44590 23910
rect 44282 23899 44590 23908
rect 58726 23964 59034 23973
rect 58726 23962 58732 23964
rect 58788 23962 58812 23964
rect 58868 23962 58892 23964
rect 58948 23962 58972 23964
rect 59028 23962 59034 23964
rect 58788 23910 58790 23962
rect 58970 23910 58972 23962
rect 58726 23908 58732 23910
rect 58788 23908 58812 23910
rect 58868 23908 58892 23910
rect 58948 23908 58972 23910
rect 59028 23908 59034 23910
rect 58726 23899 59034 23908
rect 8172 23420 8480 23429
rect 8172 23418 8178 23420
rect 8234 23418 8258 23420
rect 8314 23418 8338 23420
rect 8394 23418 8418 23420
rect 8474 23418 8480 23420
rect 8234 23366 8236 23418
rect 8416 23366 8418 23418
rect 8172 23364 8178 23366
rect 8234 23364 8258 23366
rect 8314 23364 8338 23366
rect 8394 23364 8418 23366
rect 8474 23364 8480 23366
rect 8172 23355 8480 23364
rect 22616 23420 22924 23429
rect 22616 23418 22622 23420
rect 22678 23418 22702 23420
rect 22758 23418 22782 23420
rect 22838 23418 22862 23420
rect 22918 23418 22924 23420
rect 22678 23366 22680 23418
rect 22860 23366 22862 23418
rect 22616 23364 22622 23366
rect 22678 23364 22702 23366
rect 22758 23364 22782 23366
rect 22838 23364 22862 23366
rect 22918 23364 22924 23366
rect 22616 23355 22924 23364
rect 37060 23420 37368 23429
rect 37060 23418 37066 23420
rect 37122 23418 37146 23420
rect 37202 23418 37226 23420
rect 37282 23418 37306 23420
rect 37362 23418 37368 23420
rect 37122 23366 37124 23418
rect 37304 23366 37306 23418
rect 37060 23364 37066 23366
rect 37122 23364 37146 23366
rect 37202 23364 37226 23366
rect 37282 23364 37306 23366
rect 37362 23364 37368 23366
rect 37060 23355 37368 23364
rect 51504 23420 51812 23429
rect 51504 23418 51510 23420
rect 51566 23418 51590 23420
rect 51646 23418 51670 23420
rect 51726 23418 51750 23420
rect 51806 23418 51812 23420
rect 51566 23366 51568 23418
rect 51748 23366 51750 23418
rect 51504 23364 51510 23366
rect 51566 23364 51590 23366
rect 51646 23364 51670 23366
rect 51726 23364 51750 23366
rect 51806 23364 51812 23366
rect 51504 23355 51812 23364
rect 38844 23112 38896 23118
rect 38844 23054 38896 23060
rect 47860 23112 47912 23118
rect 47860 23054 47912 23060
rect 15394 22876 15702 22885
rect 15394 22874 15400 22876
rect 15456 22874 15480 22876
rect 15536 22874 15560 22876
rect 15616 22874 15640 22876
rect 15696 22874 15702 22876
rect 15456 22822 15458 22874
rect 15638 22822 15640 22874
rect 15394 22820 15400 22822
rect 15456 22820 15480 22822
rect 15536 22820 15560 22822
rect 15616 22820 15640 22822
rect 15696 22820 15702 22822
rect 15394 22811 15702 22820
rect 29838 22876 30146 22885
rect 29838 22874 29844 22876
rect 29900 22874 29924 22876
rect 29980 22874 30004 22876
rect 30060 22874 30084 22876
rect 30140 22874 30146 22876
rect 29900 22822 29902 22874
rect 30082 22822 30084 22874
rect 29838 22820 29844 22822
rect 29900 22820 29924 22822
rect 29980 22820 30004 22822
rect 30060 22820 30084 22822
rect 30140 22820 30146 22822
rect 29838 22811 30146 22820
rect 38292 22636 38344 22642
rect 38292 22578 38344 22584
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 8172 22332 8480 22341
rect 8172 22330 8178 22332
rect 8234 22330 8258 22332
rect 8314 22330 8338 22332
rect 8394 22330 8418 22332
rect 8474 22330 8480 22332
rect 8234 22278 8236 22330
rect 8416 22278 8418 22330
rect 8172 22276 8178 22278
rect 8234 22276 8258 22278
rect 8314 22276 8338 22278
rect 8394 22276 8418 22278
rect 8474 22276 8480 22278
rect 8172 22267 8480 22276
rect 22616 22332 22924 22341
rect 22616 22330 22622 22332
rect 22678 22330 22702 22332
rect 22758 22330 22782 22332
rect 22838 22330 22862 22332
rect 22918 22330 22924 22332
rect 22678 22278 22680 22330
rect 22860 22278 22862 22330
rect 22616 22276 22622 22278
rect 22678 22276 22702 22278
rect 22758 22276 22782 22278
rect 22838 22276 22862 22278
rect 22918 22276 22924 22278
rect 22616 22267 22924 22276
rect 24320 22098 24348 22374
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2792 19854 2820 20470
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2884 19786 2912 20742
rect 3160 20058 3188 21422
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3148 20052 3200 20058
rect 3148 19994 3200 20000
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2516 17610 2544 18022
rect 3068 17882 3096 18702
rect 3252 18306 3280 20742
rect 3344 19514 3372 20742
rect 3712 20466 3740 21286
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20466 4016 20878
rect 4080 20602 4108 21422
rect 4448 21146 4476 21626
rect 5368 21486 5396 21830
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 5368 20942 5396 21422
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 4172 20398 4200 20742
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4448 20482 4476 20538
rect 4356 20454 4476 20482
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 3516 19984 3568 19990
rect 3516 19926 3568 19932
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3528 19378 3556 19926
rect 4356 19718 4384 20454
rect 4436 20324 4488 20330
rect 4436 20266 4488 20272
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3620 18426 3648 18566
rect 4264 18426 4292 18702
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 3252 18290 3372 18306
rect 3252 18284 3384 18290
rect 3252 18278 3332 18284
rect 3332 18226 3384 18232
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2792 17270 2820 17546
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2792 16794 2820 17070
rect 3344 16794 3372 18226
rect 4356 18154 4384 19654
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 4448 18086 4476 20266
rect 4540 19854 4568 20742
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 5000 20058 5028 20402
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4724 19514 4752 19722
rect 5276 19718 5304 20334
rect 5368 19854 5396 20878
rect 5460 20806 5488 21422
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4448 17746 4476 18022
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4724 17678 4752 17818
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4172 17202 4200 17614
rect 4816 17270 4844 18566
rect 5000 17678 5028 19654
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 18222 5120 18566
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5276 17762 5304 18158
rect 5184 17746 5304 17762
rect 5172 17740 5304 17746
rect 5224 17734 5304 17740
rect 5172 17682 5224 17688
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4908 17270 4936 17614
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4540 16794 4568 16934
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3712 16250 3740 16594
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 1964 13938 1992 14350
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1964 13394 1992 13874
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2240 12986 2268 14350
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 14074 2912 14214
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3344 12986 3372 13194
rect 3988 12986 4016 13670
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3068 11898 3096 12786
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3068 11558 3096 11698
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2884 11354 2912 11494
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3068 11218 3096 11494
rect 3160 11286 3188 12582
rect 3436 12238 3464 12650
rect 3620 12434 3648 12786
rect 3528 12406 3648 12434
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 3252 11354 3280 12106
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2792 10674 2820 11086
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3068 10674 3096 10950
rect 3160 10810 3188 11018
rect 3344 10810 3372 11698
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2792 10130 2820 10610
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10130 3372 10542
rect 3436 10266 3464 12174
rect 3528 11898 3556 12406
rect 3804 12322 3832 12786
rect 3620 12294 3832 12322
rect 3620 12238 3648 12294
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11898 3648 12038
rect 3896 11898 3924 12106
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3528 11150 3556 11222
rect 3620 11218 3648 11494
rect 3896 11218 3924 11834
rect 3988 11354 4016 12922
rect 4080 12918 4108 13126
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4080 11234 4108 12854
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4172 11354 4200 12378
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3988 11206 4108 11234
rect 4264 11218 4292 11562
rect 4252 11212 4304 11218
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 2792 9518 2820 10066
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3160 9722 3188 9930
rect 3344 9722 3372 10066
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2884 8634 2912 9522
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9042 3004 9318
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3068 7886 3096 8910
rect 3160 8838 3188 9658
rect 3528 9178 3556 11086
rect 3620 10674 3648 11154
rect 3988 11150 4016 11206
rect 4252 11154 4304 11160
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 9994 3648 10610
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10062 4108 10406
rect 4264 10266 4292 11154
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3608 9988 3660 9994
rect 3608 9930 3660 9936
rect 3620 9466 3648 9930
rect 3620 9438 3740 9466
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3620 9110 3648 9318
rect 3712 9178 3740 9438
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3620 8634 3648 9046
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1780 5166 1808 6734
rect 2608 6458 2636 7278
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 3602 1808 5102
rect 2240 4826 2268 6054
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2332 4622 2360 6258
rect 2516 5914 2544 6258
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 3068 5658 3096 7822
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6322 3280 7142
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 6458 3372 6666
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 2596 5636 2648 5642
rect 3068 5630 3188 5658
rect 2596 5578 2648 5584
rect 2608 4758 2636 5578
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2884 4826 2912 5102
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2596 4616 2648 4622
rect 2872 4616 2924 4622
rect 2648 4564 2728 4570
rect 2596 4558 2728 4564
rect 2872 4558 2924 4564
rect 2608 4542 2728 4558
rect 2700 4214 2728 4542
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 952 800 980 3431
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 1688 1170 1716 2314
rect 1504 1142 1716 1170
rect 1504 800 1532 1142
rect 2056 800 2084 2450
rect 2608 800 2636 3062
rect 2700 2582 2728 4150
rect 2884 3942 2912 4558
rect 3068 4554 3096 5510
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2976 4146 3004 4422
rect 3160 4146 3188 5630
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3344 5370 3372 5578
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3344 4690 3372 5306
rect 3620 5302 3648 8298
rect 3804 8090 3832 8910
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3896 5710 3924 8774
rect 4356 8634 4384 10950
rect 4540 10810 4568 16730
rect 4908 16658 4936 17206
rect 5000 16658 5028 17614
rect 5276 17134 5304 17734
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4724 14618 4752 14962
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 5000 11898 5028 12106
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11898 5212 12038
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4632 11354 4660 11494
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 5000 10674 5028 10950
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5000 10470 5028 10610
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8974 4752 9318
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 4724 8838 4752 8910
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4724 8566 4752 8774
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 8090 4108 8366
rect 4724 8362 4752 8502
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4080 7546 4108 8026
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4448 6458 4476 6598
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5914 4016 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3896 5098 3924 5646
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3436 4570 3464 4762
rect 3344 4542 3464 4570
rect 3344 4486 3372 4542
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2792 3194 2820 3402
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2884 3058 2912 3878
rect 3160 3738 3188 4082
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3344 3466 3372 4422
rect 3896 4214 3924 5034
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3988 4282 4016 4490
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3988 3670 4016 4218
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3068 3058 3096 3402
rect 3988 3058 4016 3606
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3620 2938 3648 2994
rect 3160 2910 3648 2938
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 3160 800 3188 2910
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3620 2650 3648 2790
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3712 800 3740 2790
rect 4172 2378 4200 3878
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4264 800 4292 3470
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4356 2650 4384 2858
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4540 2582 4568 4694
rect 4632 4146 4660 5510
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4724 3534 4752 3878
rect 4816 3670 4844 4422
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3194 4660 3334
rect 4724 3194 4752 3470
rect 4816 3398 4844 3606
rect 4908 3466 4936 8230
rect 5000 7954 5028 8774
rect 5092 8566 5120 8910
rect 5184 8634 5212 8910
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5914 5212 6054
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5184 5778 5212 5850
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5184 5234 5212 5714
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5092 4690 5120 5102
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4724 2446 4752 2790
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4816 800 4844 2926
rect 5000 2650 5028 3334
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5276 2378 5304 10474
rect 5368 3058 5396 16934
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5460 15706 5488 15982
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5552 15162 5580 17478
rect 5644 17338 5672 17478
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5828 15570 5856 21626
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 21146 6224 21286
rect 6288 21146 6316 21422
rect 7576 21418 7604 21830
rect 10520 21690 10548 21966
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7116 21146 7144 21286
rect 7576 21146 7604 21354
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 20602 6684 20742
rect 7576 20602 7604 21082
rect 7852 20874 7880 21422
rect 8172 21244 8480 21253
rect 8172 21242 8178 21244
rect 8234 21242 8258 21244
rect 8314 21242 8338 21244
rect 8394 21242 8418 21244
rect 8474 21242 8480 21244
rect 8234 21190 8236 21242
rect 8416 21190 8418 21242
rect 8172 21188 8178 21190
rect 8234 21188 8258 21190
rect 8314 21188 8338 21190
rect 8394 21188 8418 21190
rect 8474 21188 8480 21190
rect 8172 21179 8480 21188
rect 8680 20874 8708 21422
rect 8772 21146 8800 21490
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8956 21146 8984 21286
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 5920 17338 5948 20198
rect 6380 20058 6408 20198
rect 6656 20058 6684 20266
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5920 16998 5948 17070
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5920 16794 5948 16934
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5828 14074 5856 15302
rect 6012 15094 6040 15846
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5460 13394 5488 13670
rect 5920 13530 5948 14282
rect 6104 13802 6132 19790
rect 6656 19378 6684 19994
rect 6748 19514 6776 20402
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7300 19514 7328 20334
rect 7576 20058 7604 20538
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6196 18630 6224 19110
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6196 18086 6224 18566
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 14278 6224 18022
rect 6656 17338 6684 18158
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6840 17270 6868 17614
rect 7300 17610 7328 18022
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6380 16658 6408 17138
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 15094 6500 15438
rect 6564 15162 6592 15506
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 15088 6512 15094
rect 6460 15030 6512 15036
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6472 13870 6500 14554
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6104 13530 6132 13738
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11898 5580 12174
rect 6196 11898 6224 12310
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5460 6798 5488 10610
rect 5828 10266 5856 10610
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 7886 5672 8774
rect 5920 8090 5948 8978
rect 6012 8634 6040 9386
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7342 5764 7754
rect 6012 7750 6040 8366
rect 6104 8090 6132 8842
rect 6196 8498 6224 8842
rect 6288 8498 6316 9590
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6380 9178 6408 9522
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6380 8498 6408 9114
rect 6564 8838 6592 15098
rect 6840 12986 6868 16934
rect 6932 16794 6960 17274
rect 7116 17202 7144 17478
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 13938 7328 15302
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7484 14278 7512 14826
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13938 7512 14214
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 12442 7052 12718
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6840 10810 6868 12310
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6826 10024 6882 10033
rect 6826 9959 6828 9968
rect 6880 9959 6882 9968
rect 6828 9930 6880 9936
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 9042 6776 9386
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6840 8498 6868 9930
rect 6932 9518 6960 11086
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7208 9586 7236 10746
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6920 9512 6972 9518
rect 7208 9466 7236 9522
rect 6920 9454 6972 9460
rect 6932 8974 6960 9454
rect 7116 9438 7236 9466
rect 7116 9178 7144 9438
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7546 6040 7686
rect 6196 7546 6224 8434
rect 6932 7886 6960 8910
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 7024 7478 7052 8434
rect 7116 7478 7144 9114
rect 7208 8430 7236 9318
rect 7300 9178 7328 9998
rect 7484 9738 7512 13466
rect 7668 12918 7696 18294
rect 7852 17490 7880 20810
rect 9416 20806 9444 21422
rect 9876 21350 9904 21626
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9692 20942 9720 21286
rect 9784 21146 9812 21286
rect 9876 21146 9904 21286
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8172 20156 8480 20165
rect 8172 20154 8178 20156
rect 8234 20154 8258 20156
rect 8314 20154 8338 20156
rect 8394 20154 8418 20156
rect 8474 20154 8480 20156
rect 8234 20102 8236 20154
rect 8416 20102 8418 20154
rect 8172 20100 8178 20102
rect 8234 20100 8258 20102
rect 8314 20100 8338 20102
rect 8394 20100 8418 20102
rect 8474 20100 8480 20102
rect 8172 20091 8480 20100
rect 8772 20058 8800 20402
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 9048 20058 9076 20198
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9416 19718 9444 20742
rect 9876 20466 9904 20742
rect 10428 20466 10456 21490
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10980 20806 11008 21422
rect 11072 20874 11100 21830
rect 11348 21622 11376 21830
rect 11336 21616 11388 21622
rect 11336 21558 11388 21564
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13740 20534 13768 20742
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 9680 20392 9732 20398
rect 11520 20392 11572 20398
rect 9680 20334 9732 20340
rect 11518 20360 11520 20369
rect 11572 20360 11574 20369
rect 9692 20058 9720 20334
rect 9864 20324 9916 20330
rect 11518 20295 11574 20304
rect 9864 20266 9916 20272
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 8172 19068 8480 19077
rect 8172 19066 8178 19068
rect 8234 19066 8258 19068
rect 8314 19066 8338 19068
rect 8394 19066 8418 19068
rect 8474 19066 8480 19068
rect 8234 19014 8236 19066
rect 8416 19014 8418 19066
rect 8172 19012 8178 19014
rect 8234 19012 8258 19014
rect 8314 19012 8338 19014
rect 8394 19012 8418 19014
rect 8474 19012 8480 19014
rect 8172 19003 8480 19012
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7944 17610 7972 18022
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7852 17462 7972 17490
rect 7944 16250 7972 17462
rect 8036 17270 8064 18566
rect 8772 18290 8800 19654
rect 9692 19174 9720 19858
rect 9876 19242 9904 20266
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11348 19514 11376 19722
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8956 18426 8984 18702
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8172 17980 8480 17989
rect 8172 17978 8178 17980
rect 8234 17978 8258 17980
rect 8314 17978 8338 17980
rect 8394 17978 8418 17980
rect 8474 17978 8480 17980
rect 8234 17926 8236 17978
rect 8416 17926 8418 17978
rect 8172 17924 8178 17926
rect 8234 17924 8258 17926
rect 8314 17924 8338 17926
rect 8394 17924 8418 17926
rect 8474 17924 8480 17926
rect 8172 17915 8480 17924
rect 8588 17882 8616 18158
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8172 16892 8480 16901
rect 8172 16890 8178 16892
rect 8234 16890 8258 16892
rect 8314 16890 8338 16892
rect 8394 16890 8418 16892
rect 8474 16890 8480 16892
rect 8234 16838 8236 16890
rect 8416 16838 8418 16890
rect 8172 16836 8178 16838
rect 8234 16836 8258 16838
rect 8314 16836 8338 16838
rect 8394 16836 8418 16838
rect 8474 16836 8480 16838
rect 8172 16827 8480 16836
rect 8588 16726 8616 17682
rect 8772 17542 8800 18226
rect 9048 18222 9076 18634
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 9232 17338 9260 18158
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9232 17202 9260 17274
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9324 17134 9352 17818
rect 9416 17746 9444 18022
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9508 16726 9536 19110
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9588 17128 9640 17134
rect 9640 17088 9720 17116
rect 9588 17070 9640 17076
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16538 8524 16594
rect 8772 16538 8800 16662
rect 8496 16510 8800 16538
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7944 15570 7972 16186
rect 8172 15804 8480 15813
rect 8172 15802 8178 15804
rect 8234 15802 8258 15804
rect 8314 15802 8338 15804
rect 8394 15802 8418 15804
rect 8474 15802 8480 15804
rect 8234 15750 8236 15802
rect 8416 15750 8418 15802
rect 8172 15748 8178 15750
rect 8234 15748 8258 15750
rect 8314 15748 8338 15750
rect 8394 15748 8418 15750
rect 8474 15748 8480 15750
rect 8172 15739 8480 15748
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14618 7788 14894
rect 8036 14822 8064 15438
rect 8588 14958 8616 15438
rect 8772 15026 8800 16510
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14618 8064 14758
rect 8172 14716 8480 14725
rect 8172 14714 8178 14716
rect 8234 14714 8258 14716
rect 8314 14714 8338 14716
rect 8394 14714 8418 14716
rect 8474 14714 8480 14716
rect 8234 14662 8236 14714
rect 8416 14662 8418 14714
rect 8172 14660 8178 14662
rect 8234 14660 8258 14662
rect 8314 14660 8338 14662
rect 8394 14660 8418 14662
rect 8474 14660 8480 14662
rect 8172 14651 8480 14660
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8588 14414 8616 14894
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7852 14074 7880 14282
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 11830 7604 12582
rect 7668 12306 7696 12854
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7484 9710 7604 9738
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7484 8634 7512 9522
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 7392 7206 7420 7822
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 6798 7420 7142
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 5460 6390 5488 6734
rect 6748 6458 6776 6734
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5460 5624 5488 6326
rect 5644 5710 5672 6326
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5540 5636 5592 5642
rect 5460 5596 5540 5624
rect 5460 5302 5488 5596
rect 5540 5578 5592 5584
rect 5644 5302 5672 5646
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5460 5166 5488 5238
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 4758 5488 4966
rect 5644 4758 5672 5034
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5736 4690 5764 5170
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4826 6040 4966
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5446 4176 5502 4185
rect 5446 4111 5448 4120
rect 5500 4111 5502 4120
rect 5448 4082 5500 4088
rect 5460 3738 5488 4082
rect 5920 3942 5948 4422
rect 6196 4146 6224 5510
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6288 4078 6316 4694
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5920 3466 5948 3878
rect 6012 3641 6040 3878
rect 5998 3632 6054 3641
rect 6196 3602 6224 3878
rect 5998 3567 6054 3576
rect 6184 3596 6236 3602
rect 6012 3534 6040 3567
rect 6184 3538 6236 3544
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 3058 5948 3402
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5552 1442 5580 2450
rect 5920 2446 5948 2790
rect 6380 2650 6408 4150
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3738 6684 3878
rect 6840 3738 6868 4014
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 5368 1414 5580 1442
rect 5368 800 5396 1414
rect 6472 800 6500 3470
rect 6840 2854 6868 3470
rect 7024 3194 7052 4082
rect 7392 4078 7420 6734
rect 7576 6186 7604 9710
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7576 4622 7604 4966
rect 7668 4826 7696 12242
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7944 11762 7972 12174
rect 8036 12170 8064 13874
rect 8172 13628 8480 13637
rect 8172 13626 8178 13628
rect 8234 13626 8258 13628
rect 8314 13626 8338 13628
rect 8394 13626 8418 13628
rect 8474 13626 8480 13628
rect 8234 13574 8236 13626
rect 8416 13574 8418 13626
rect 8172 13572 8178 13574
rect 8234 13572 8258 13574
rect 8314 13572 8338 13574
rect 8394 13572 8418 13574
rect 8474 13572 8480 13574
rect 8172 13563 8480 13572
rect 8588 13394 8616 14350
rect 8772 14278 8800 14962
rect 8956 14618 8984 15438
rect 9404 15428 9456 15434
rect 9404 15370 9456 15376
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8172 12540 8480 12549
rect 8172 12538 8178 12540
rect 8234 12538 8258 12540
rect 8314 12538 8338 12540
rect 8394 12538 8418 12540
rect 8474 12538 8480 12540
rect 8234 12486 8236 12538
rect 8416 12486 8418 12538
rect 8172 12484 8178 12486
rect 8234 12484 8258 12486
rect 8314 12484 8338 12486
rect 8394 12484 8418 12486
rect 8474 12484 8480 12486
rect 8172 12475 8480 12484
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8036 11642 8064 12106
rect 8404 11762 8432 12106
rect 8588 11898 8616 12582
rect 8680 12238 8708 12718
rect 8772 12306 8800 12922
rect 9140 12374 9168 14214
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9232 12986 9260 13806
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8390 11656 8446 11665
rect 8036 11614 8390 11642
rect 8390 11591 8392 11600
rect 8444 11591 8446 11600
rect 8392 11562 8444 11568
rect 8172 11452 8480 11461
rect 8172 11450 8178 11452
rect 8234 11450 8258 11452
rect 8314 11450 8338 11452
rect 8394 11450 8418 11452
rect 8474 11450 8480 11452
rect 8234 11398 8236 11450
rect 8416 11398 8418 11450
rect 8172 11396 8178 11398
rect 8234 11396 8258 11398
rect 8314 11396 8338 11398
rect 8394 11396 8418 11398
rect 8474 11396 8480 11398
rect 8172 11387 8480 11396
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10674 7788 10950
rect 7852 10810 7880 11018
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 8036 10674 8064 11290
rect 8588 11218 8616 11834
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8404 10810 8432 11154
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8588 10810 8616 11018
rect 8680 11014 8708 12174
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 10062 8064 10406
rect 8172 10364 8480 10373
rect 8172 10362 8178 10364
rect 8234 10362 8258 10364
rect 8314 10362 8338 10364
rect 8394 10362 8418 10364
rect 8474 10362 8480 10364
rect 8234 10310 8236 10362
rect 8416 10310 8418 10362
rect 8172 10308 8178 10310
rect 8234 10308 8258 10310
rect 8314 10308 8338 10310
rect 8394 10308 8418 10310
rect 8474 10308 8480 10310
rect 8172 10299 8480 10308
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8668 10056 8720 10062
rect 8772 10044 8800 12242
rect 9324 12238 9352 14758
rect 9416 14482 9444 15370
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9416 12782 9444 14418
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11354 9168 11630
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8720 10016 8800 10044
rect 8668 9998 8720 10004
rect 8036 9722 8064 9998
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8036 9602 8064 9658
rect 7944 9574 8064 9602
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8634 7880 8774
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7944 8498 7972 9574
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 8922 8064 9454
rect 8172 9276 8480 9285
rect 8172 9274 8178 9276
rect 8234 9274 8258 9276
rect 8314 9274 8338 9276
rect 8394 9274 8418 9276
rect 8474 9274 8480 9276
rect 8234 9222 8236 9274
rect 8416 9222 8418 9274
rect 8172 9220 8178 9222
rect 8234 9220 8258 9222
rect 8314 9220 8338 9222
rect 8394 9220 8418 9222
rect 8474 9220 8480 9222
rect 8172 9211 8480 9220
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8036 8894 8248 8922
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8498 8064 8774
rect 8220 8498 8248 8894
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8312 8566 8340 8842
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7944 8090 7972 8434
rect 8496 8430 8524 9114
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8498 8616 8774
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8172 8188 8480 8197
rect 8172 8186 8178 8188
rect 8234 8186 8258 8188
rect 8314 8186 8338 8188
rect 8394 8186 8418 8188
rect 8474 8186 8480 8188
rect 8234 8134 8236 8186
rect 8416 8134 8418 8186
rect 8172 8132 8178 8134
rect 8234 8132 8258 8134
rect 8314 8132 8338 8134
rect 8394 8132 8418 8134
rect 8474 8132 8480 8134
rect 8172 8123 8480 8132
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7760 4554 7788 6190
rect 7852 5574 7880 7278
rect 8172 7100 8480 7109
rect 8172 7098 8178 7100
rect 8234 7098 8258 7100
rect 8314 7098 8338 7100
rect 8394 7098 8418 7100
rect 8474 7098 8480 7100
rect 8234 7046 8236 7098
rect 8416 7046 8418 7098
rect 8172 7044 8178 7046
rect 8234 7044 8258 7046
rect 8314 7044 8338 7046
rect 8394 7044 8418 7046
rect 8474 7044 8480 7046
rect 8172 7035 8480 7044
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5914 8064 6122
rect 8172 6012 8480 6021
rect 8172 6010 8178 6012
rect 8234 6010 8258 6012
rect 8314 6010 8338 6012
rect 8394 6010 8418 6012
rect 8474 6010 8480 6012
rect 8234 5958 8236 6010
rect 8416 5958 8418 6010
rect 8172 5956 8178 5958
rect 8234 5956 8258 5958
rect 8314 5956 8338 5958
rect 8394 5956 8418 5958
rect 8474 5956 8480 5958
rect 8172 5947 8480 5956
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8588 5846 8616 8434
rect 8680 8362 8708 8502
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8680 8090 8708 8298
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8772 6390 8800 7414
rect 8760 6384 8812 6390
rect 8666 6352 8722 6361
rect 8760 6326 8812 6332
rect 8666 6287 8668 6296
rect 8720 6287 8722 6296
rect 8668 6258 8720 6264
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8864 5642 8892 10678
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8634 8984 8910
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 5370 7880 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7852 4282 7880 5170
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7944 4214 7972 4966
rect 8036 4826 8064 5102
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8172 4924 8480 4933
rect 8172 4922 8178 4924
rect 8234 4922 8258 4924
rect 8314 4922 8338 4924
rect 8394 4922 8418 4924
rect 8474 4922 8480 4924
rect 8234 4870 8236 4922
rect 8416 4870 8418 4922
rect 8172 4868 8178 4870
rect 8234 4868 8258 4870
rect 8314 4868 8338 4870
rect 8394 4868 8418 4870
rect 8474 4868 8480 4870
rect 8172 4859 8480 4868
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8680 4706 8708 4966
rect 8496 4690 8708 4706
rect 8484 4684 8708 4690
rect 8536 4678 8708 4684
rect 8484 4626 8536 4632
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7392 3534 7420 4014
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 7024 800 7052 2926
rect 7208 2446 7236 3334
rect 7760 3194 7788 3402
rect 8036 3194 8064 4490
rect 8864 4282 8892 5102
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8172 3836 8480 3845
rect 8172 3834 8178 3836
rect 8234 3834 8258 3836
rect 8314 3834 8338 3836
rect 8394 3834 8418 3836
rect 8474 3834 8480 3836
rect 8234 3782 8236 3834
rect 8416 3782 8418 3834
rect 8172 3780 8178 3782
rect 8234 3780 8258 3782
rect 8314 3780 8338 3782
rect 8394 3780 8418 3782
rect 8474 3780 8480 3782
rect 8172 3771 8480 3780
rect 8956 3738 8984 5743
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9048 4078 9076 5102
rect 9126 4720 9182 4729
rect 9126 4655 9182 4664
rect 9140 4622 9168 4655
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8772 2990 8800 3606
rect 8956 3534 8984 3674
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8172 2748 8480 2757
rect 8172 2746 8178 2748
rect 8234 2746 8258 2748
rect 8314 2746 8338 2748
rect 8394 2746 8418 2748
rect 8474 2746 8480 2748
rect 8234 2694 8236 2746
rect 8416 2694 8418 2746
rect 8172 2692 8178 2694
rect 8234 2692 8258 2694
rect 8314 2692 8338 2694
rect 8394 2692 8418 2694
rect 8474 2692 8480 2694
rect 8172 2683 8480 2692
rect 9048 2650 9076 3470
rect 9232 3194 9260 12038
rect 9416 11694 9444 12310
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10674 9444 10950
rect 9508 10713 9536 16662
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9600 15570 9628 15846
rect 9692 15706 9720 17088
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9784 16726 9812 17002
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9600 15094 9628 15302
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9876 14482 9904 15098
rect 9968 14958 9996 18090
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17678 10824 18022
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10520 17202 10548 17546
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10888 17134 10916 17478
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10704 16794 10732 17070
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10888 15026 10916 17070
rect 11072 15910 11100 17614
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13258 9904 13670
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12170 9628 13126
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9876 11830 9904 12038
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 9586 11656 9642 11665
rect 9642 11614 9720 11642
rect 9586 11591 9642 11600
rect 9494 10704 9550 10713
rect 9404 10668 9456 10674
rect 9494 10639 9550 10648
rect 9404 10610 9456 10616
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 6662 9352 7346
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9416 6390 9444 10610
rect 9508 9178 9536 10639
rect 9692 9926 9720 11614
rect 9968 10742 9996 14894
rect 11072 13274 11100 14962
rect 11164 14618 11192 19246
rect 11532 17678 11560 20198
rect 12084 19922 12112 20198
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11348 17338 11376 17546
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11440 16998 11468 17478
rect 11624 17338 11652 18158
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11808 17134 11836 19314
rect 12084 18970 12112 19858
rect 12360 19310 12388 19994
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12176 18902 12204 19246
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12912 18970 12940 19178
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12164 18896 12216 18902
rect 12164 18838 12216 18844
rect 13096 18834 13124 19110
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 16794 11468 16934
rect 11900 16794 11928 17138
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 15094 11284 15438
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11164 14074 11192 14554
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11164 13954 11192 14010
rect 11164 13926 11376 13954
rect 11440 13938 11468 15846
rect 11244 13320 11296 13326
rect 11072 13246 11192 13274
rect 11244 13262 11296 13268
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12986 11100 13126
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11354 10364 11494
rect 10428 11354 10456 11834
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9968 10266 9996 10678
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10428 10130 10456 11290
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10520 10742 10548 11018
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10810 11100 10950
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9784 9654 9812 9998
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 9772 9648 9824 9654
rect 9770 9616 9772 9625
rect 9824 9616 9826 9625
rect 9770 9551 9826 9560
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9508 8430 9536 8910
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9600 7818 9628 8774
rect 10152 8090 10180 8910
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 7002 9536 7278
rect 9692 7274 9720 7822
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 5914 9628 6258
rect 9692 5914 9720 6734
rect 9876 6458 9904 7142
rect 9968 6934 9996 7142
rect 9956 6928 10008 6934
rect 10244 6882 10272 9862
rect 10428 9722 10456 10066
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 8634 10364 8774
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 9956 6870 10008 6876
rect 10152 6866 10272 6882
rect 10140 6860 10272 6866
rect 10192 6854 10272 6860
rect 10140 6802 10192 6808
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9324 3466 9352 5578
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9692 4026 9720 4218
rect 9600 4010 9720 4026
rect 9784 4010 9812 5578
rect 9588 4004 9720 4010
rect 9640 3998 9720 4004
rect 9772 4004 9824 4010
rect 9588 3946 9640 3952
rect 9772 3946 9824 3952
rect 10060 3738 10088 6258
rect 10152 5642 10180 6802
rect 10428 6798 10456 8026
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10520 6254 10548 6938
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5930 10548 6190
rect 10428 5902 10548 5930
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10152 3738 10180 4014
rect 10244 3942 10272 4694
rect 10428 4078 10456 5902
rect 10704 5710 10732 7686
rect 10796 5914 10824 10202
rect 11164 9178 11192 13246
rect 11256 12986 11284 13262
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11348 10810 11376 13926
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11440 13530 11468 13874
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 9654 11376 10406
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11440 8974 11468 9454
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 9178 11560 9318
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11624 9042 11652 16186
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 12306 11744 12582
rect 11992 12434 12020 17478
rect 12728 17134 12756 18566
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12912 17814 12940 18022
rect 12900 17808 12952 17814
rect 12898 17776 12900 17785
rect 12952 17776 12954 17785
rect 12898 17711 12954 17720
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12912 17338 12940 17614
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16794 12204 16934
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12084 16046 12112 16526
rect 13188 16182 13216 20402
rect 13832 20398 13860 20742
rect 13924 20602 13952 21422
rect 14740 21412 14792 21418
rect 14740 21354 14792 21360
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14476 21146 14504 21286
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 14660 20466 14688 21286
rect 14752 21010 14780 21354
rect 14844 21146 14872 21898
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 15394 21788 15702 21797
rect 15394 21786 15400 21788
rect 15456 21786 15480 21788
rect 15536 21786 15560 21788
rect 15616 21786 15640 21788
rect 15696 21786 15702 21788
rect 15456 21734 15458 21786
rect 15638 21734 15640 21786
rect 15394 21732 15400 21734
rect 15456 21732 15480 21734
rect 15536 21732 15560 21734
rect 15616 21732 15640 21734
rect 15696 21732 15702 21734
rect 15394 21723 15702 21732
rect 23032 21622 23060 21830
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 18696 21480 18748 21486
rect 18696 21422 18748 21428
rect 15212 21146 15240 21422
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13832 20058 13860 20334
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13648 18970 13676 19722
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13176 16176 13228 16182
rect 13176 16118 13228 16124
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 15162 12664 15302
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 13530 12664 14350
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12782 12204 13126
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11900 12406 12020 12434
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11716 9586 11744 10746
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11716 8906 11744 9522
rect 11808 9178 11836 9930
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7206 11008 7822
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9324 2922 9352 3402
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 3194 9904 3334
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9494 3088 9550 3097
rect 9494 3023 9496 3032
rect 9548 3023 9550 3032
rect 9496 2994 9548 3000
rect 10520 2990 10548 5306
rect 10796 5250 10824 5850
rect 10796 5222 10916 5250
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7576 800 7604 2450
rect 9784 2446 9812 2790
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 8392 2372 8444 2378
rect 8444 2332 8708 2360
rect 8392 2314 8444 2320
rect 8680 800 8708 2332
rect 8772 898 8800 2382
rect 9968 1170 9996 2450
rect 10704 2360 10732 4558
rect 10796 4214 10824 5102
rect 10888 4690 10916 5222
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10980 4690 11008 5102
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10796 3738 10824 4150
rect 11072 4078 11100 8842
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7750 11284 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11150 5128 11206 5137
rect 11150 5063 11152 5072
rect 11204 5063 11206 5072
rect 11152 5034 11204 5040
rect 11164 4622 11192 5034
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11256 4486 11284 7686
rect 11348 7410 11376 8230
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11532 7410 11560 7754
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 6458 11468 6734
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11440 4146 11468 6394
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10888 3194 10916 3878
rect 11348 3618 11376 4082
rect 11164 3590 11376 3618
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11164 2650 11192 3590
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 11348 3194 11376 3402
rect 11532 3194 11560 6598
rect 11716 5370 11744 8570
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 6390 11836 8434
rect 11900 6440 11928 12406
rect 12176 10810 12204 12718
rect 12268 12442 12296 13194
rect 12532 13184 12584 13190
rect 12452 13144 12532 13172
rect 12452 12782 12480 13144
rect 12532 13126 12584 13132
rect 12728 12986 12756 15098
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 14074 12940 14214
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13096 13394 13124 13670
rect 13372 13530 13400 17070
rect 13464 16590 13492 17478
rect 13740 17202 13768 19382
rect 13832 18086 13860 19654
rect 14108 19310 14136 19926
rect 14292 19922 14320 20198
rect 14936 20058 14964 20742
rect 15394 20700 15702 20709
rect 15394 20698 15400 20700
rect 15456 20698 15480 20700
rect 15536 20698 15560 20700
rect 15616 20698 15640 20700
rect 15696 20698 15702 20700
rect 15456 20646 15458 20698
rect 15638 20646 15640 20698
rect 15394 20644 15400 20646
rect 15456 20644 15480 20646
rect 15536 20644 15560 20646
rect 15616 20644 15640 20646
rect 15696 20644 15702 20646
rect 15394 20635 15702 20644
rect 15856 20534 15884 21286
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14936 19446 14964 19994
rect 15028 19446 15056 20334
rect 15120 19938 15148 20402
rect 15120 19910 15240 19938
rect 15212 19854 15240 19910
rect 15200 19848 15252 19854
rect 15476 19848 15528 19854
rect 15200 19790 15252 19796
rect 15304 19796 15476 19802
rect 15304 19790 15528 19796
rect 15304 19774 15516 19790
rect 16500 19786 16528 20878
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 19854 16620 20742
rect 16684 20262 16712 20878
rect 18142 20360 18198 20369
rect 18142 20295 18144 20304
rect 18196 20295 18198 20304
rect 18144 20266 18196 20272
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 16868 19922 16896 20198
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16488 19780 16540 19786
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 15028 18970 15056 19382
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15304 18834 15332 19774
rect 16488 19722 16540 19728
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 15394 19612 15702 19621
rect 15394 19610 15400 19612
rect 15456 19610 15480 19612
rect 15536 19610 15560 19612
rect 15616 19610 15640 19612
rect 15696 19610 15702 19612
rect 15456 19558 15458 19610
rect 15638 19558 15640 19610
rect 15394 19556 15400 19558
rect 15456 19556 15480 19558
rect 15536 19556 15560 19558
rect 15616 19556 15640 19558
rect 15696 19556 15702 19558
rect 15394 19547 15702 19556
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 14188 18216 14240 18222
rect 15304 18170 15332 18770
rect 15394 18524 15702 18533
rect 15394 18522 15400 18524
rect 15456 18522 15480 18524
rect 15536 18522 15560 18524
rect 15616 18522 15640 18524
rect 15696 18522 15702 18524
rect 15456 18470 15458 18522
rect 15638 18470 15640 18522
rect 15394 18468 15400 18470
rect 15456 18468 15480 18470
rect 15536 18468 15560 18470
rect 15616 18468 15640 18470
rect 15696 18468 15702 18470
rect 15394 18459 15702 18468
rect 14188 18158 14240 18164
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17542 13860 18022
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13740 16250 13768 17138
rect 13832 16998 13860 17478
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15706 13584 15846
rect 13648 15706 13676 16050
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13372 13190 13400 13466
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12452 12306 12480 12718
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12544 12442 12572 12650
rect 12532 12436 12584 12442
rect 12728 12434 12756 12922
rect 13740 12850 13768 13806
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13832 12730 13860 16934
rect 13924 16726 13952 17206
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14016 15858 14044 17002
rect 14108 16794 14136 17614
rect 14200 17542 14228 18158
rect 15212 18142 15332 18170
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 13924 15830 14044 15858
rect 13924 14822 13952 15830
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 13326 13952 14758
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 14016 12850 14044 15642
rect 14108 15570 14136 16730
rect 14200 16658 14228 17478
rect 14752 17338 14780 17614
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16658 14412 16934
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 16046 14228 16390
rect 14188 16040 14240 16046
rect 14464 16040 14516 16046
rect 14188 15982 14240 15988
rect 14292 16000 14464 16028
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 13394 14136 15506
rect 14200 15162 14228 15982
rect 14292 15910 14320 16000
rect 14464 15982 14516 15988
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14752 14958 14780 17070
rect 14844 16250 14872 17138
rect 15212 16674 15240 18142
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 17338 15332 18022
rect 15934 17776 15990 17785
rect 15934 17711 15990 17720
rect 15394 17436 15702 17445
rect 15394 17434 15400 17436
rect 15456 17434 15480 17436
rect 15536 17434 15560 17436
rect 15616 17434 15640 17436
rect 15696 17434 15702 17436
rect 15456 17382 15458 17434
rect 15638 17382 15640 17434
rect 15394 17380 15400 17382
rect 15456 17380 15480 17382
rect 15536 17380 15560 17382
rect 15616 17380 15640 17382
rect 15696 17380 15702 17382
rect 15394 17371 15702 17380
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15948 17270 15976 17711
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 14936 16646 15240 16674
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14936 15706 14964 16646
rect 15212 16640 15240 16646
rect 15292 16652 15344 16658
rect 15212 16612 15292 16640
rect 15292 16594 15344 16600
rect 16132 16590 16160 19654
rect 16224 18834 16252 19654
rect 16500 19514 16528 19722
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16868 18970 16896 19858
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17328 19378 17356 19790
rect 17972 19786 18000 20198
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 18248 19514 18276 20878
rect 18708 20058 18736 21422
rect 18984 20806 19012 21558
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 16960 18970 16988 19314
rect 18616 19242 18644 19926
rect 18800 19446 18828 20742
rect 18984 20398 19012 20742
rect 19352 20602 19380 21286
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16408 16726 16436 17206
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15120 16130 15148 16526
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15028 16102 15148 16130
rect 15028 15978 15056 16102
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15120 15162 15148 15982
rect 15212 15434 15240 16390
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13556 12714 13860 12730
rect 13544 12708 13860 12714
rect 13596 12702 13860 12708
rect 13544 12650 13596 12656
rect 12728 12406 12848 12434
rect 12532 12378 12584 12384
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12268 11150 12296 12242
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12084 10418 12112 10678
rect 12268 10538 12296 11086
rect 12452 11082 12480 11630
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12084 10390 12296 10418
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11992 9178 12020 9522
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 12084 9042 12112 10134
rect 12176 9450 12204 10202
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12268 8514 12296 10390
rect 12360 10266 12388 10542
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12636 10130 12664 10950
rect 12728 10130 12756 11834
rect 12820 11830 12848 12406
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 13280 11082 13308 12038
rect 13556 11898 13584 12650
rect 14016 12628 14044 12786
rect 13832 12600 14044 12628
rect 13832 12434 13860 12600
rect 13740 12406 13860 12434
rect 13740 12102 13768 12406
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12440 10056 12492 10062
rect 12728 10010 12756 10066
rect 13280 10062 13308 11018
rect 13832 10810 13860 11154
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 12492 10004 12756 10010
rect 12440 9998 12756 10004
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12452 9982 12756 9998
rect 13280 9926 13308 9998
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13096 9722 13124 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12176 8486 12296 8514
rect 12176 7342 12204 8486
rect 12360 8362 12388 8978
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12360 7970 12388 8298
rect 13004 8090 13032 8502
rect 13096 8430 13124 9658
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13280 8430 13308 8774
rect 13464 8634 13492 8774
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12268 7942 12388 7970
rect 12268 7886 12296 7942
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 11900 6412 12020 6440
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 3194 11652 4490
rect 11716 3942 11744 5170
rect 11808 5098 11836 6326
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11900 5914 11928 6258
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11808 4622 11836 5034
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11808 4146 11836 4422
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11900 3194 11928 4966
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11610 3088 11666 3097
rect 11610 3023 11666 3032
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11624 2514 11652 3023
rect 11992 2774 12020 6412
rect 12176 6254 12204 7278
rect 12268 7274 12296 7822
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 13280 7002 13308 7822
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13556 6866 13584 10474
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13740 9178 13768 9522
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13832 8838 13860 10542
rect 14108 10470 14136 13126
rect 14200 12782 14228 13262
rect 14292 13190 14320 14350
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 13258 14504 13874
rect 14752 13870 14780 14894
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 14074 14964 14214
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12986 14320 13126
rect 14476 12986 14504 13194
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12434 14596 12718
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14200 12406 14596 12434
rect 14200 12102 14228 12406
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9722 13952 9862
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14016 9654 14044 9998
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13912 9376 13964 9382
rect 13964 9336 14044 9364
rect 13912 9318 13964 9324
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12176 5846 12204 6190
rect 12820 5914 12848 6598
rect 13096 6458 13124 6666
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13556 5914 13584 6802
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12360 5370 12388 5510
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12084 3534 12112 5238
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12360 3097 12388 5306
rect 12544 3466 12572 5510
rect 13832 5370 13860 8774
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13924 7546 13952 7686
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13096 5166 13124 5306
rect 13726 5264 13782 5273
rect 13726 5199 13728 5208
rect 13780 5199 13782 5208
rect 13728 5170 13780 5176
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3738 13032 3878
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12346 3088 12402 3097
rect 12346 3023 12402 3032
rect 12544 2990 12572 3402
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 11808 2746 12020 2774
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11808 2446 11836 2746
rect 12268 2514 12388 2530
rect 12268 2508 12400 2514
rect 12268 2502 12348 2508
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11152 2372 11204 2378
rect 10704 2332 10916 2360
rect 9784 1142 9996 1170
rect 8772 870 8892 898
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 8864 762 8892 870
rect 9140 870 9260 898
rect 9140 762 9168 870
rect 9232 800 9260 870
rect 9784 800 9812 1142
rect 10888 800 10916 2332
rect 11152 2314 11204 2320
rect 8864 734 9168 762
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11164 762 11192 2314
rect 11348 870 11468 898
rect 11348 762 11376 870
rect 11440 800 11468 870
rect 11992 870 12112 898
rect 11992 800 12020 870
rect 11164 734 11376 762
rect 11426 0 11482 800
rect 11978 0 12034 800
rect 12084 762 12112 870
rect 12268 762 12296 2502
rect 12348 2450 12400 2456
rect 13188 2122 13216 4082
rect 13280 3058 13308 4082
rect 13924 3126 13952 4422
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 13096 2094 13216 2122
rect 13096 800 13124 2094
rect 12084 734 12296 762
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13280 762 13308 2858
rect 14016 2446 14044 9336
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14108 5914 14136 6870
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5574 14228 12038
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10266 14320 10950
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14660 9586 14688 12582
rect 14752 11762 14780 12582
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15212 11898 15240 12106
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 10810 14872 10950
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14832 9920 14884 9926
rect 15028 9908 15056 10406
rect 15120 10062 15148 11086
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15212 9994 15240 10950
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15028 9880 15148 9908
rect 14832 9862 14884 9868
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14568 8634 14596 9454
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14476 7274 14504 7822
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 7002 14596 7142
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14660 6866 14688 8910
rect 14844 7886 14872 9862
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14476 5930 14504 6598
rect 14568 6458 14596 6598
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 6118 14688 6802
rect 14752 6730 14780 7686
rect 14844 7478 14872 7822
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14844 6390 14872 7278
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14476 5902 14596 5930
rect 14752 5914 14780 6258
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14108 3670 14136 4558
rect 14292 4282 14320 4558
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14476 4078 14504 4966
rect 14568 4078 14596 5902
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14568 3602 14596 4014
rect 14752 3602 14780 5034
rect 14844 4690 14872 6326
rect 14936 5914 14964 6734
rect 15120 5914 15148 9880
rect 15304 8786 15332 16390
rect 15394 16348 15702 16357
rect 15394 16346 15400 16348
rect 15456 16346 15480 16348
rect 15536 16346 15560 16348
rect 15616 16346 15640 16348
rect 15696 16346 15702 16348
rect 15456 16294 15458 16346
rect 15638 16294 15640 16346
rect 15394 16292 15400 16294
rect 15456 16292 15480 16294
rect 15536 16292 15560 16294
rect 15616 16292 15640 16294
rect 15696 16292 15702 16294
rect 15394 16283 15702 16292
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15706 15792 15846
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15394 15260 15702 15269
rect 15394 15258 15400 15260
rect 15456 15258 15480 15260
rect 15536 15258 15560 15260
rect 15616 15258 15640 15260
rect 15696 15258 15702 15260
rect 15456 15206 15458 15258
rect 15638 15206 15640 15258
rect 15394 15204 15400 15206
rect 15456 15204 15480 15206
rect 15536 15204 15560 15206
rect 15616 15204 15640 15206
rect 15696 15204 15702 15206
rect 15394 15195 15702 15204
rect 15948 14958 15976 16186
rect 16960 16114 16988 16594
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 15162 16896 15302
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15394 14172 15702 14181
rect 15394 14170 15400 14172
rect 15456 14170 15480 14172
rect 15536 14170 15560 14172
rect 15616 14170 15640 14172
rect 15696 14170 15702 14172
rect 15456 14118 15458 14170
rect 15638 14118 15640 14170
rect 15394 14116 15400 14118
rect 15456 14116 15480 14118
rect 15536 14116 15560 14118
rect 15616 14116 15640 14118
rect 15696 14116 15702 14118
rect 15394 14107 15702 14116
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15764 13326 15792 13670
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15394 13084 15702 13093
rect 15394 13082 15400 13084
rect 15456 13082 15480 13084
rect 15536 13082 15560 13084
rect 15616 13082 15640 13084
rect 15696 13082 15702 13084
rect 15456 13030 15458 13082
rect 15638 13030 15640 13082
rect 15394 13028 15400 13030
rect 15456 13028 15480 13030
rect 15536 13028 15560 13030
rect 15616 13028 15640 13030
rect 15696 13028 15702 13030
rect 15394 13019 15702 13028
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 12442 15516 12650
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15394 11996 15702 12005
rect 15394 11994 15400 11996
rect 15456 11994 15480 11996
rect 15536 11994 15560 11996
rect 15616 11994 15640 11996
rect 15696 11994 15702 11996
rect 15456 11942 15458 11994
rect 15638 11942 15640 11994
rect 15394 11940 15400 11942
rect 15456 11940 15480 11942
rect 15536 11940 15560 11942
rect 15616 11940 15640 11942
rect 15696 11940 15702 11942
rect 15394 11931 15702 11940
rect 15856 11150 15884 12038
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15394 10908 15702 10917
rect 15394 10906 15400 10908
rect 15456 10906 15480 10908
rect 15536 10906 15560 10908
rect 15616 10906 15640 10908
rect 15696 10906 15702 10908
rect 15456 10854 15458 10906
rect 15638 10854 15640 10906
rect 15394 10852 15400 10854
rect 15456 10852 15480 10854
rect 15536 10852 15560 10854
rect 15616 10852 15640 10854
rect 15696 10852 15702 10854
rect 15394 10843 15702 10852
rect 15672 10674 15792 10690
rect 15660 10668 15792 10674
rect 15712 10662 15792 10668
rect 15660 10610 15712 10616
rect 15764 9874 15792 10662
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 9994 15884 10406
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15764 9846 15884 9874
rect 15394 9820 15702 9829
rect 15394 9818 15400 9820
rect 15456 9818 15480 9820
rect 15536 9818 15560 9820
rect 15616 9818 15640 9820
rect 15696 9818 15702 9820
rect 15456 9766 15458 9818
rect 15638 9766 15640 9818
rect 15394 9764 15400 9766
rect 15456 9764 15480 9766
rect 15536 9764 15560 9766
rect 15616 9764 15640 9766
rect 15696 9764 15702 9766
rect 15394 9755 15702 9764
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15212 8758 15332 8786
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4214 14872 4422
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14660 3194 14688 3334
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14292 1578 14320 2926
rect 14752 2650 14780 2994
rect 14936 2922 14964 5170
rect 15120 5030 15148 5850
rect 15212 5234 15240 8758
rect 15394 8732 15702 8741
rect 15394 8730 15400 8732
rect 15456 8730 15480 8732
rect 15536 8730 15560 8732
rect 15616 8730 15640 8732
rect 15696 8730 15702 8732
rect 15456 8678 15458 8730
rect 15638 8678 15640 8730
rect 15394 8676 15400 8678
rect 15456 8676 15480 8678
rect 15536 8676 15560 8678
rect 15616 8676 15640 8678
rect 15696 8676 15702 8678
rect 15394 8667 15702 8676
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 8090 15516 8230
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7410 15332 7686
rect 15394 7644 15702 7653
rect 15394 7642 15400 7644
rect 15456 7642 15480 7644
rect 15536 7642 15560 7644
rect 15616 7642 15640 7644
rect 15696 7642 15702 7644
rect 15456 7590 15458 7642
rect 15638 7590 15640 7642
rect 15394 7588 15400 7590
rect 15456 7588 15480 7590
rect 15536 7588 15560 7590
rect 15616 7588 15640 7590
rect 15696 7588 15702 7590
rect 15394 7579 15702 7588
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15304 5642 15332 6870
rect 15580 6866 15608 7346
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15394 6556 15702 6565
rect 15394 6554 15400 6556
rect 15456 6554 15480 6556
rect 15536 6554 15560 6556
rect 15616 6554 15640 6556
rect 15696 6554 15702 6556
rect 15456 6502 15458 6554
rect 15638 6502 15640 6554
rect 15394 6500 15400 6502
rect 15456 6500 15480 6502
rect 15536 6500 15560 6502
rect 15616 6500 15640 6502
rect 15696 6500 15702 6502
rect 15394 6491 15702 6500
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15672 5574 15700 6054
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15394 5468 15702 5477
rect 15394 5466 15400 5468
rect 15456 5466 15480 5468
rect 15536 5466 15560 5468
rect 15616 5466 15640 5468
rect 15696 5466 15702 5468
rect 15456 5414 15458 5466
rect 15638 5414 15640 5466
rect 15394 5412 15400 5414
rect 15456 5412 15480 5414
rect 15536 5412 15560 5414
rect 15616 5412 15640 5414
rect 15696 5412 15702 5414
rect 15394 5403 15702 5412
rect 15764 5370 15792 9522
rect 15856 8906 15884 9846
rect 15948 9518 15976 14894
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13870 16528 14214
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16500 13326 16528 13806
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16500 12238 16528 13262
rect 17420 12782 17448 19110
rect 18616 18766 18644 19178
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18708 18970 18736 19110
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 17338 17632 17614
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 18156 16590 18184 17478
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16794 18644 17070
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 16250 18552 16526
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 18984 16130 19012 20334
rect 19168 19378 19196 20402
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19352 19854 19380 20198
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19076 18970 19104 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19352 17202 19380 19246
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19076 16250 19104 16390
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19352 16182 19380 17138
rect 19340 16176 19392 16182
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17144 12306 17172 12582
rect 17604 12442 17632 13194
rect 17788 12986 17816 13262
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17788 12866 17816 12922
rect 17696 12838 17816 12866
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11898 16528 12174
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16316 10606 16344 11766
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 10810 16712 11630
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11354 17356 11494
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 17696 10674 17724 12838
rect 17880 12782 17908 13126
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17788 12374 17816 12718
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17972 12238 18000 16118
rect 18512 16108 18564 16114
rect 18984 16102 19104 16130
rect 19340 16118 19392 16124
rect 18512 16050 18564 16056
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15706 18460 15846
rect 18524 15706 18552 16050
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14482 18368 14758
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18064 13530 18092 14350
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 13938 18184 14214
rect 18248 14074 18276 14350
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18064 12434 18092 13126
rect 18064 12406 18184 12434
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17972 11830 18000 12174
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10810 18092 10950
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16028 9648 16080 9654
rect 16026 9616 16028 9625
rect 16080 9616 16082 9625
rect 16592 9602 16620 10406
rect 16026 9551 16082 9560
rect 16408 9574 16620 9602
rect 16776 9586 16804 10610
rect 17960 10600 18012 10606
rect 17682 10568 17738 10577
rect 17960 10542 18012 10548
rect 17682 10503 17738 10512
rect 17696 10470 17724 10503
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17038 10296 17094 10305
rect 17038 10231 17040 10240
rect 17092 10231 17094 10240
rect 17316 10260 17368 10266
rect 17040 10202 17092 10208
rect 17316 10202 17368 10208
rect 16764 9580 16816 9586
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15856 7410 15884 8366
rect 16408 8362 16436 9574
rect 16764 9522 16816 9528
rect 17052 9518 17080 10202
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17328 8906 17356 10202
rect 17592 9920 17644 9926
rect 17972 9908 18000 10542
rect 18052 10260 18104 10266
rect 18156 10248 18184 12406
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18248 10266 18276 10610
rect 18104 10220 18184 10248
rect 18236 10260 18288 10266
rect 18052 10202 18104 10208
rect 18236 10202 18288 10208
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18052 9920 18104 9926
rect 17972 9880 18052 9908
rect 17592 9862 17644 9868
rect 18052 9862 18104 9868
rect 17604 9722 17632 9862
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 18064 9586 18092 9862
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9178 17816 9318
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15948 6882 15976 8298
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 7954 16068 8230
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15856 6854 15976 6882
rect 16040 6866 16068 7142
rect 16224 6866 16252 7822
rect 16776 7188 16804 8366
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16856 7200 16908 7206
rect 16776 7160 16856 7188
rect 16028 6860 16080 6866
rect 15856 5778 15884 6854
rect 16028 6802 16080 6808
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15948 6458 15976 6734
rect 16776 6662 16804 7160
rect 16856 7142 16908 7148
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16868 6474 16896 6802
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16776 6446 16896 6474
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15856 5624 15884 5714
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 15936 5636 15988 5642
rect 15856 5596 15936 5624
rect 15936 5578 15988 5584
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15108 5024 15160 5030
rect 15384 5024 15436 5030
rect 15108 4966 15160 4972
rect 15304 4984 15384 5012
rect 15016 4616 15068 4622
rect 15304 4570 15332 4984
rect 15384 4966 15436 4972
rect 15016 4558 15068 4564
rect 15028 4010 15056 4558
rect 15120 4542 15332 4570
rect 15120 4162 15148 4542
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4282 15240 4422
rect 15394 4380 15702 4389
rect 15394 4378 15400 4380
rect 15456 4378 15480 4380
rect 15536 4378 15560 4380
rect 15616 4378 15640 4380
rect 15696 4378 15702 4380
rect 15456 4326 15458 4378
rect 15638 4326 15640 4378
rect 15394 4324 15400 4326
rect 15456 4324 15480 4326
rect 15536 4324 15560 4326
rect 15616 4324 15640 4326
rect 15696 4324 15702 4326
rect 15394 4315 15702 4324
rect 15764 4282 15792 5170
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16040 4554 16068 4966
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15856 4162 15884 4422
rect 15120 4134 15240 4162
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15120 2961 15148 3470
rect 15106 2952 15162 2961
rect 14924 2916 14976 2922
rect 15106 2887 15162 2896
rect 14924 2858 14976 2864
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 15212 2446 15240 4134
rect 15304 4134 15424 4162
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 14200 1550 14320 1578
rect 13556 870 13676 898
rect 13556 762 13584 870
rect 13648 800 13676 870
rect 14200 800 14228 1550
rect 14752 800 14780 2314
rect 15304 800 15332 4134
rect 15396 4078 15424 4134
rect 15488 4134 15884 4162
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15488 3534 15516 4134
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3534 15608 3878
rect 16132 3670 16160 5510
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15394 3292 15702 3301
rect 15394 3290 15400 3292
rect 15456 3290 15480 3292
rect 15536 3290 15560 3292
rect 15616 3290 15640 3292
rect 15696 3290 15702 3292
rect 15456 3238 15458 3290
rect 15638 3238 15640 3290
rect 15394 3236 15400 3238
rect 15456 3236 15480 3238
rect 15536 3236 15560 3238
rect 15616 3236 15640 3238
rect 15696 3236 15702 3238
rect 15394 3227 15702 3236
rect 15764 2582 15792 3538
rect 16120 3188 16172 3194
rect 16224 3176 16252 3538
rect 16316 3516 16344 4014
rect 16408 3942 16436 5646
rect 16684 5642 16712 6190
rect 16776 6118 16804 6446
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16396 3528 16448 3534
rect 16316 3488 16396 3516
rect 16396 3470 16448 3476
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16172 3148 16252 3176
rect 16120 3130 16172 3136
rect 16316 3097 16344 3334
rect 16302 3088 16358 3097
rect 16302 3023 16358 3032
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16408 2650 16436 2994
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15394 2204 15702 2213
rect 15394 2202 15400 2204
rect 15456 2202 15480 2204
rect 15536 2202 15560 2204
rect 15616 2202 15640 2204
rect 15696 2202 15702 2204
rect 15456 2150 15458 2202
rect 15638 2150 15640 2202
rect 15394 2148 15400 2150
rect 15456 2148 15480 2150
rect 15536 2148 15560 2150
rect 15616 2148 15640 2150
rect 15696 2148 15702 2150
rect 15394 2139 15702 2148
rect 15856 800 15884 2450
rect 16500 2122 16528 4082
rect 16684 3602 16712 5578
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3058 16712 3334
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16776 2990 16804 6054
rect 16960 5778 16988 6054
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16868 3194 16896 5170
rect 17052 5030 17080 7686
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17052 4146 17080 4966
rect 17144 4622 17172 5510
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 17236 4554 17264 8774
rect 17328 7954 17356 8842
rect 17880 8838 17908 9454
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17328 7732 17356 7890
rect 17420 7886 17448 8230
rect 17972 8090 18000 8366
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17328 7704 17724 7732
rect 17696 7274 17724 7704
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17052 3058 17080 4082
rect 17236 4078 17264 4490
rect 17420 4214 17448 6598
rect 17696 5914 17724 6598
rect 18064 6458 18092 9522
rect 18248 9178 18276 9930
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18340 8514 18368 14418
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13394 18460 14214
rect 18524 13870 18552 15302
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18524 12442 18552 13806
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18616 12986 18644 13330
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12436 18564 12442
rect 18432 12406 18512 12434
rect 18432 11014 18460 12406
rect 18512 12378 18564 12384
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10713 18460 10950
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18432 10538 18460 10639
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18616 10305 18644 10542
rect 18602 10296 18658 10305
rect 18512 10260 18564 10266
rect 18602 10231 18658 10240
rect 18512 10202 18564 10208
rect 18524 9518 18552 10202
rect 18708 10146 18736 15098
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18984 14074 19012 14758
rect 19076 14074 19104 16102
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19168 15162 19196 15846
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19168 14618 19196 14894
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19444 14482 19472 18566
rect 19536 17814 19564 20538
rect 19628 20534 19656 21286
rect 22616 21244 22924 21253
rect 22616 21242 22622 21244
rect 22678 21242 22702 21244
rect 22758 21242 22782 21244
rect 22838 21242 22862 21244
rect 22918 21242 22924 21244
rect 22678 21190 22680 21242
rect 22860 21190 22862 21242
rect 22616 21188 22622 21190
rect 22678 21188 22702 21190
rect 22758 21188 22782 21190
rect 22838 21188 22862 21190
rect 22918 21188 22924 21190
rect 22616 21179 22924 21188
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19628 19854 19656 20470
rect 19812 19922 19840 20742
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19628 19378 19656 19790
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19628 18426 19656 19314
rect 19812 18850 19840 19858
rect 19904 18970 19932 20878
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20456 20602 20484 20742
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20180 19854 20208 19994
rect 20456 19922 20484 20538
rect 20548 20466 20576 20742
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20640 20262 20668 20878
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 21192 19854 21220 20198
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19812 18822 19932 18850
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19536 17270 19564 17750
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19812 16998 19840 18158
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19812 16658 19840 16934
rect 19904 16658 19932 18822
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 17542 20392 18566
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19536 15706 19564 15982
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19536 15162 19564 15642
rect 19904 15366 19932 16594
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13190 19012 13670
rect 19076 13394 19104 14010
rect 19628 13870 19656 14214
rect 19996 14074 20024 14350
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 19156 13388 19208 13394
rect 19628 13376 19656 13806
rect 19996 13530 20024 14010
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20088 13410 20116 17478
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20272 16794 20300 17274
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20180 16590 20208 16730
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20272 16454 20300 16526
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20364 16266 20392 17478
rect 20456 16590 20484 17818
rect 20534 17776 20590 17785
rect 20534 17711 20536 17720
rect 20588 17711 20590 17720
rect 20536 17682 20588 17688
rect 20732 17678 20760 18022
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20272 16238 20392 16266
rect 20272 16182 20300 16238
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20272 15366 20300 16118
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 19892 13388 19944 13394
rect 19208 13348 19656 13376
rect 19812 13348 19892 13376
rect 19156 13330 19208 13336
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12986 19472 13126
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18892 12434 18920 12786
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 12434 19656 12718
rect 19812 12442 19840 13348
rect 19892 13330 19944 13336
rect 19996 13382 20116 13410
rect 18892 12406 19104 12434
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18800 10674 18828 11086
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 19076 10606 19104 12406
rect 19352 12406 19656 12434
rect 19800 12436 19852 12442
rect 19352 11898 19380 12406
rect 19800 12378 19852 12384
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19352 11354 19380 11834
rect 19812 11626 19840 12378
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19064 10600 19116 10606
rect 19062 10568 19064 10577
rect 19116 10568 19118 10577
rect 19062 10503 19118 10512
rect 18708 10118 19012 10146
rect 18984 10062 19012 10118
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18248 8486 18368 8514
rect 18248 8022 18276 8486
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7410 18184 7686
rect 18340 7478 18368 8366
rect 18984 7954 19012 9998
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18984 6866 19012 7890
rect 19076 7886 19104 8774
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 6866 19288 7686
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19444 7002 19472 7346
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5914 17816 6122
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17788 5710 17816 5850
rect 18156 5794 18184 6802
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6390 18920 6598
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18064 5766 18184 5794
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3738 17356 4014
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17512 3534 17540 4762
rect 17696 4622 17724 5238
rect 17788 5166 17816 5646
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 18064 5098 18092 5766
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4146 17816 4422
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 18064 4078 18092 4558
rect 18156 4146 18184 5646
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17696 3194 17724 3878
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17788 3194 17816 3402
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16868 2650 16896 2994
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17788 2514 17908 2530
rect 17788 2508 17920 2514
rect 17788 2502 17868 2508
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16408 2094 16528 2122
rect 16408 800 16436 2094
rect 13280 734 13584 762
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16592 762 16620 2314
rect 16868 870 16988 898
rect 16868 762 16896 870
rect 16960 800 16988 870
rect 17512 870 17632 898
rect 17512 800 17540 870
rect 16592 734 16896 762
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 17604 762 17632 870
rect 17788 762 17816 2502
rect 17868 2450 17920 2456
rect 18156 1578 18184 2994
rect 18248 2446 18276 5510
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18432 4826 18460 5238
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 18340 3738 18368 3946
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18524 2922 18552 6258
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19076 5302 19104 5510
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 19352 5114 19380 6054
rect 19444 5778 19472 6190
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19536 5370 19564 11494
rect 19996 10130 20024 13382
rect 20180 13326 20208 13874
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9722 20208 9862
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19352 5086 19472 5114
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19076 4282 19104 4422
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19168 3738 19196 3878
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18970 2952 19026 2961
rect 18512 2916 18564 2922
rect 18970 2887 18972 2896
rect 18512 2858 18564 2864
rect 19024 2887 19026 2896
rect 19156 2916 19208 2922
rect 18972 2858 19024 2864
rect 19156 2858 19208 2864
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18064 1550 18184 1578
rect 18064 800 18092 1550
rect 18616 800 18644 2314
rect 19168 800 19196 2858
rect 19352 2446 19380 4966
rect 19444 4078 19472 5086
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19628 3534 19656 8842
rect 19720 8634 19748 8910
rect 19812 8838 19840 9046
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19904 8650 19932 8774
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19812 8622 19932 8650
rect 20088 8634 20116 9386
rect 20272 9178 20300 15302
rect 20456 13394 20484 16526
rect 20824 16250 20852 16594
rect 21100 16522 21128 19654
rect 21192 19514 21220 19790
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21284 18834 21312 20742
rect 22204 20602 22232 20946
rect 23032 20942 23060 21286
rect 23676 21078 23704 21966
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24228 21690 24256 21830
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23952 20942 23980 21422
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23952 20602 23980 20878
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 21652 20058 21680 20198
rect 22616 20156 22924 20165
rect 22616 20154 22622 20156
rect 22678 20154 22702 20156
rect 22758 20154 22782 20156
rect 22838 20154 22862 20156
rect 22918 20154 22924 20156
rect 22678 20102 22680 20154
rect 22860 20102 22862 20154
rect 22616 20100 22622 20102
rect 22678 20100 22702 20102
rect 22758 20100 22782 20102
rect 22838 20100 22862 20102
rect 22918 20100 22924 20102
rect 22616 20091 22924 20100
rect 23768 20058 23796 20198
rect 23860 20058 23888 20402
rect 24044 20398 24072 21286
rect 24320 21146 24348 22034
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24308 21140 24360 21146
rect 24308 21082 24360 21088
rect 24412 21010 24440 21830
rect 24688 21434 24716 22374
rect 24780 21690 24808 22510
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 37924 22432 37976 22438
rect 37924 22374 37976 22380
rect 25424 22030 25452 22374
rect 37060 22332 37368 22341
rect 37060 22330 37066 22332
rect 37122 22330 37146 22332
rect 37202 22330 37226 22332
rect 37282 22330 37306 22332
rect 37362 22330 37368 22332
rect 37122 22278 37124 22330
rect 37304 22278 37306 22330
rect 37060 22276 37066 22278
rect 37122 22276 37146 22278
rect 37202 22276 37226 22278
rect 37282 22276 37306 22278
rect 37362 22276 37368 22278
rect 37060 22267 37368 22276
rect 37936 22094 37964 22374
rect 37844 22066 37964 22094
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26528 21690 26556 21830
rect 29838 21788 30146 21797
rect 29838 21786 29844 21788
rect 29900 21786 29924 21788
rect 29980 21786 30004 21788
rect 30060 21786 30084 21788
rect 30140 21786 30146 21788
rect 29900 21734 29902 21786
rect 30082 21734 30084 21786
rect 29838 21732 29844 21734
rect 29900 21732 29924 21734
rect 29980 21732 30004 21734
rect 30060 21732 30084 21734
rect 30140 21732 30146 21734
rect 29838 21723 30146 21732
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 26516 21684 26568 21690
rect 26516 21626 26568 21632
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 24860 21480 24912 21486
rect 24688 21428 24860 21434
rect 24688 21422 24912 21428
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 24688 21406 24900 21422
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 24306 20904 24362 20913
rect 24306 20839 24308 20848
rect 24360 20839 24362 20848
rect 24308 20810 24360 20816
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 21640 19916 21692 19922
rect 21560 19876 21640 19904
rect 21560 19174 21588 19876
rect 21640 19858 21692 19864
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17202 21496 17478
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21088 16516 21140 16522
rect 21088 16458 21140 16464
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20824 16046 20852 16186
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 14822 20668 15506
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20456 12850 20484 13330
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11694 20484 12106
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20364 10810 20392 11630
rect 20456 11370 20484 11630
rect 20456 11342 20576 11370
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20456 10470 20484 11222
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20364 9994 20392 10066
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20364 8838 20392 9930
rect 20456 9586 20484 10406
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20548 9518 20576 11342
rect 20640 9674 20668 14758
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14074 20852 14350
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 11830 20760 13126
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20640 9646 20760 9674
rect 20732 9586 20760 9646
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20536 9512 20588 9518
rect 20456 9460 20536 9466
rect 20456 9454 20588 9460
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20456 9438 20576 9454
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20076 8628 20128 8634
rect 19812 8430 19840 8622
rect 20076 8570 20128 8576
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 20456 8378 20484 9438
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 8634 20576 9318
rect 20640 8906 20668 9454
rect 20732 9178 20760 9522
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 7546 19748 7686
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19812 6798 19840 8366
rect 19904 7818 19932 8366
rect 20456 8350 20576 8378
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19720 5370 19748 6190
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19812 5778 19840 6054
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19800 5568 19852 5574
rect 19904 5556 19932 7754
rect 19996 6866 20024 7890
rect 20456 7886 20484 8230
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 6934 20116 7142
rect 20076 6928 20128 6934
rect 20548 6914 20576 8350
rect 20640 7954 20668 8842
rect 20732 8090 20760 8910
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20824 7954 20852 11562
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20548 6886 20760 6914
rect 20076 6870 20128 6876
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 19852 5528 19932 5556
rect 19800 5510 19852 5516
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19720 5030 19748 5306
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19812 4146 19840 5510
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19996 4826 20024 5102
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19996 3738 20024 4490
rect 20088 4078 20116 6122
rect 20272 5681 20300 6598
rect 20732 6458 20760 6886
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20720 6316 20772 6322
rect 20916 6304 20944 16390
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21376 15706 21404 16050
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21008 12986 21036 13806
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21468 12918 21496 14214
rect 21560 13802 21588 19110
rect 21652 18630 21680 19654
rect 22664 19514 22692 19654
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 22616 19068 22924 19077
rect 22616 19066 22622 19068
rect 22678 19066 22702 19068
rect 22758 19066 22782 19068
rect 22838 19066 22862 19068
rect 22918 19066 22924 19068
rect 22678 19014 22680 19066
rect 22860 19014 22862 19066
rect 22616 19012 22622 19014
rect 22678 19012 22702 19014
rect 22758 19012 22782 19014
rect 22838 19012 22862 19014
rect 22918 19012 22924 19014
rect 22616 19003 22924 19012
rect 23492 18970 23520 19246
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 22756 18426 22784 18702
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22204 17338 22232 17478
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22480 16046 22508 18022
rect 22616 17980 22924 17989
rect 22616 17978 22622 17980
rect 22678 17978 22702 17980
rect 22758 17978 22782 17980
rect 22838 17978 22862 17980
rect 22918 17978 22924 17980
rect 22678 17926 22680 17978
rect 22860 17926 22862 17978
rect 22616 17924 22622 17926
rect 22678 17924 22702 17926
rect 22758 17924 22782 17926
rect 22838 17924 22862 17926
rect 22918 17924 22924 17926
rect 22616 17915 22924 17924
rect 23308 17678 23336 18566
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 22616 16892 22924 16901
rect 22616 16890 22622 16892
rect 22678 16890 22702 16892
rect 22758 16890 22782 16892
rect 22838 16890 22862 16892
rect 22918 16890 22924 16892
rect 22678 16838 22680 16890
rect 22860 16838 22862 16890
rect 22616 16836 22622 16838
rect 22678 16836 22702 16838
rect 22758 16836 22782 16838
rect 22838 16836 22862 16838
rect 22918 16836 22924 16838
rect 22616 16827 22924 16836
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21652 15706 21680 15846
rect 22616 15804 22924 15813
rect 22616 15802 22622 15804
rect 22678 15802 22702 15804
rect 22758 15802 22782 15804
rect 22838 15802 22862 15804
rect 22918 15802 22924 15804
rect 22678 15750 22680 15802
rect 22860 15750 22862 15802
rect 22616 15748 22622 15750
rect 22678 15748 22702 15750
rect 22758 15748 22782 15750
rect 22838 15748 22862 15750
rect 22918 15748 22924 15750
rect 22616 15739 22924 15748
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21744 14482 21772 14962
rect 22616 14716 22924 14725
rect 22616 14714 22622 14716
rect 22678 14714 22702 14716
rect 22758 14714 22782 14716
rect 22838 14714 22862 14716
rect 22918 14714 22924 14716
rect 22678 14662 22680 14714
rect 22860 14662 22862 14714
rect 22616 14660 22622 14662
rect 22678 14660 22702 14662
rect 22758 14660 22782 14662
rect 22838 14660 22862 14662
rect 22918 14660 22924 14662
rect 22616 14651 22924 14660
rect 23216 14618 23244 15438
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 22388 13530 22416 14282
rect 22756 14006 22784 14418
rect 23020 14272 23072 14278
rect 23020 14214 23072 14220
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 23032 13870 23060 14214
rect 23124 14006 23152 14214
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22480 13394 22508 13670
rect 22616 13628 22924 13637
rect 22616 13626 22622 13628
rect 22678 13626 22702 13628
rect 22758 13626 22782 13628
rect 22838 13626 22862 13628
rect 22918 13626 22924 13628
rect 22678 13574 22680 13626
rect 22860 13574 22862 13626
rect 22616 13572 22622 13574
rect 22678 13572 22702 13574
rect 22758 13572 22782 13574
rect 22838 13572 22862 13574
rect 22918 13572 22924 13574
rect 22616 13563 22924 13572
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 22204 12646 22232 13126
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22204 12442 22232 12582
rect 22388 12442 22416 12718
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21100 10810 21128 12174
rect 21836 12102 21864 12242
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21652 11354 21680 11698
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21284 10266 21312 11018
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8634 21220 8842
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21284 8430 21312 9522
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21560 8294 21588 9998
rect 21836 9674 21864 12038
rect 22480 11830 22508 12582
rect 22616 12540 22924 12549
rect 22616 12538 22622 12540
rect 22678 12538 22702 12540
rect 22758 12538 22782 12540
rect 22838 12538 22862 12540
rect 22918 12538 22924 12540
rect 22678 12486 22680 12538
rect 22860 12486 22862 12538
rect 22616 12484 22622 12486
rect 22678 12484 22702 12486
rect 22758 12484 22782 12486
rect 22838 12484 22862 12486
rect 22918 12484 22924 12486
rect 22616 12475 22924 12484
rect 23032 12306 23060 13806
rect 23124 13394 23152 13942
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23112 12912 23164 12918
rect 23112 12854 23164 12860
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22616 11452 22924 11461
rect 22616 11450 22622 11452
rect 22678 11450 22702 11452
rect 22758 11450 22782 11452
rect 22838 11450 22862 11452
rect 22918 11450 22924 11452
rect 22678 11398 22680 11450
rect 22860 11398 22862 11450
rect 22616 11396 22622 11398
rect 22678 11396 22702 11398
rect 22758 11396 22782 11398
rect 22838 11396 22862 11398
rect 22918 11396 22924 11398
rect 22616 11387 22924 11396
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21744 9646 21864 9674
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21652 8634 21680 9318
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21192 7274 21220 7822
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21468 7206 21496 7822
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21008 6730 21036 7142
rect 21744 6848 21772 9646
rect 22112 9382 22140 9862
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 21824 6860 21876 6866
rect 21744 6820 21824 6848
rect 21824 6802 21876 6808
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20772 6276 20944 6304
rect 20720 6258 20772 6264
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20258 5672 20314 5681
rect 20258 5607 20314 5616
rect 20272 5098 20300 5607
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20732 4622 20760 5510
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 20548 3194 20576 3878
rect 20732 3534 20760 4558
rect 20824 4486 20852 5102
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 20180 2650 20208 3062
rect 20916 3058 20944 6054
rect 21008 5234 21036 6666
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21100 4078 21128 6598
rect 22204 6458 22232 10746
rect 22616 10364 22924 10373
rect 22616 10362 22622 10364
rect 22678 10362 22702 10364
rect 22758 10362 22782 10364
rect 22838 10362 22862 10364
rect 22918 10362 22924 10364
rect 22678 10310 22680 10362
rect 22860 10310 22862 10362
rect 22616 10308 22622 10310
rect 22678 10308 22702 10310
rect 22758 10308 22782 10310
rect 22838 10308 22862 10310
rect 22918 10308 22924 10310
rect 22616 10299 22924 10308
rect 23124 9450 23152 12854
rect 23308 12730 23336 16730
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 15094 23428 15302
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23492 14362 23520 18906
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23584 17814 23612 18702
rect 24044 18222 24072 20334
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 24228 19718 24256 20198
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24228 18970 24256 19654
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 24136 18426 24164 18566
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 23860 17338 23888 18158
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23952 17202 23980 17478
rect 24044 17270 24072 18158
rect 24320 17542 24348 20810
rect 24596 20602 24624 21286
rect 24584 20596 24636 20602
rect 24584 20538 24636 20544
rect 24780 18902 24808 21406
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25792 21146 25820 21286
rect 26068 21146 26096 21422
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25780 21140 25832 21146
rect 25780 21082 25832 21088
rect 26056 21140 26108 21146
rect 26056 21082 26108 21088
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24858 20360 24914 20369
rect 24964 20346 24992 20946
rect 25332 20942 25360 21082
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25412 20936 25464 20942
rect 25596 20936 25648 20942
rect 25412 20878 25464 20884
rect 25502 20904 25558 20913
rect 25424 20806 25452 20878
rect 25558 20884 25596 20890
rect 25558 20878 25648 20884
rect 25558 20862 25636 20878
rect 25502 20839 25558 20848
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 24914 20318 24992 20346
rect 24858 20295 24860 20304
rect 24912 20295 24914 20304
rect 24860 20266 24912 20272
rect 24768 18896 24820 18902
rect 24768 18838 24820 18844
rect 24872 18426 24900 20266
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23676 16794 23704 16934
rect 23768 16794 23796 17138
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 24044 16726 24072 17206
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23400 14334 23520 14362
rect 23676 14346 23704 15030
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23664 14340 23716 14346
rect 23400 13802 23428 14334
rect 23664 14282 23716 14288
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23492 14006 23520 14214
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23400 13530 23428 13738
rect 23584 13530 23612 13874
rect 23768 13870 23796 14758
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23860 13802 23888 14282
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23400 12918 23428 13466
rect 24136 13258 24164 17478
rect 24504 17338 24532 18022
rect 24964 17746 24992 18022
rect 25056 17746 25084 18362
rect 25332 18290 25360 20198
rect 25792 19854 25820 21082
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 26160 18766 26188 20742
rect 26620 20466 26648 21286
rect 26804 21010 26832 21490
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26712 20602 26740 20946
rect 27908 20602 27936 21558
rect 30196 21480 30248 21486
rect 30196 21422 30248 21428
rect 30012 21412 30064 21418
rect 30012 21354 30064 21360
rect 30024 21146 30052 21354
rect 30208 21146 30236 21422
rect 35348 21412 35400 21418
rect 35348 21354 35400 21360
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30012 21140 30064 21146
rect 30012 21082 30064 21088
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28000 20602 28028 20878
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 27988 20596 28040 20602
rect 27988 20538 28040 20544
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27356 19854 27384 20198
rect 28552 19854 28580 20742
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 27356 19514 27384 19790
rect 28644 19514 28672 20198
rect 28828 20058 28856 20878
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 30564 20800 30616 20806
rect 30564 20742 30616 20748
rect 28920 20602 28948 20742
rect 29838 20700 30146 20709
rect 29838 20698 29844 20700
rect 29900 20698 29924 20700
rect 29980 20698 30004 20700
rect 30060 20698 30084 20700
rect 30140 20698 30146 20700
rect 29900 20646 29902 20698
rect 30082 20646 30084 20698
rect 29838 20644 29844 20646
rect 29900 20644 29924 20646
rect 29980 20644 30004 20646
rect 30060 20644 30084 20646
rect 30140 20644 30146 20646
rect 29838 20635 30146 20644
rect 30576 20602 30604 20742
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 30564 20596 30616 20602
rect 30564 20538 30616 20544
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 29460 20528 29512 20534
rect 29460 20470 29512 20476
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 29012 19514 29040 19654
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 28724 19168 28776 19174
rect 28724 19110 28776 19116
rect 28736 18834 28764 19110
rect 28828 18970 28856 19314
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 25148 17746 25176 18090
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24780 17338 24808 17614
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24320 15910 24348 17070
rect 24412 16794 24440 17138
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24412 15722 24440 16730
rect 24872 16658 24900 16730
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24320 15694 24440 15722
rect 24320 15026 24348 15694
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24228 13802 24256 14758
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24216 13796 24268 13802
rect 24216 13738 24268 13744
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 24228 12986 24256 13738
rect 24504 13190 24532 14350
rect 24688 14074 24716 14350
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24596 13938 24624 14010
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 13258 24716 13806
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23308 12702 23520 12730
rect 23492 12646 23520 12702
rect 23848 12708 23900 12714
rect 23848 12650 23900 12656
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23308 11898 23336 12174
rect 23492 12170 23520 12582
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23204 11008 23256 11014
rect 23204 10950 23256 10956
rect 23216 10674 23244 10950
rect 23308 10674 23336 11018
rect 23400 10674 23428 11290
rect 23492 11286 23520 11630
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 23584 10674 23612 10950
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23768 10198 23796 11154
rect 23756 10192 23808 10198
rect 23756 10134 23808 10140
rect 23768 9926 23796 10134
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23112 9444 23164 9450
rect 23112 9386 23164 9392
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22480 9110 22508 9318
rect 22616 9276 22924 9285
rect 22616 9274 22622 9276
rect 22678 9274 22702 9276
rect 22758 9274 22782 9276
rect 22838 9274 22862 9276
rect 22918 9274 22924 9276
rect 22678 9222 22680 9274
rect 22860 9222 22862 9274
rect 22616 9220 22622 9222
rect 22678 9220 22702 9222
rect 22758 9220 22782 9222
rect 22838 9220 22862 9222
rect 22918 9220 22924 9222
rect 22616 9211 22924 9220
rect 23124 9110 23152 9386
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23400 9178 23428 9318
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 23294 8800 23350 8809
rect 23032 8498 23060 8774
rect 23294 8735 23350 8744
rect 23308 8634 23336 8735
rect 23400 8634 23428 9114
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 22616 8188 22924 8197
rect 22616 8186 22622 8188
rect 22678 8186 22702 8188
rect 22758 8186 22782 8188
rect 22838 8186 22862 8188
rect 22918 8186 22924 8188
rect 22678 8134 22680 8186
rect 22860 8134 22862 8186
rect 22616 8132 22622 8134
rect 22678 8132 22702 8134
rect 22758 8132 22782 8134
rect 22838 8132 22862 8134
rect 22918 8132 22924 8134
rect 22616 8123 22924 8132
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22940 7698 22968 7822
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 20996 4072 21048 4078
rect 20996 4014 21048 4020
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 21008 3738 21036 4014
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 21468 3670 21496 5306
rect 21560 5166 21588 6394
rect 22204 5710 22232 6394
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21560 4282 21588 5102
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21744 4078 21772 5646
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 21928 5302 21956 5510
rect 21916 5296 21968 5302
rect 21916 5238 21968 5244
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21836 4282 21864 4966
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 21928 4078 21956 4762
rect 22020 4622 22048 5510
rect 22296 5370 22324 7686
rect 22940 7670 23060 7698
rect 22616 7100 22924 7109
rect 22616 7098 22622 7100
rect 22678 7098 22702 7100
rect 22758 7098 22782 7100
rect 22838 7098 22862 7100
rect 22918 7098 22924 7100
rect 22678 7046 22680 7098
rect 22860 7046 22862 7098
rect 22616 7044 22622 7046
rect 22678 7044 22702 7046
rect 22758 7044 22782 7046
rect 22838 7044 22862 7046
rect 22918 7044 22924 7046
rect 22616 7035 22924 7044
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22388 6118 22416 6870
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 6390 22876 6598
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22388 5914 22416 6054
rect 22616 6012 22924 6021
rect 22616 6010 22622 6012
rect 22678 6010 22702 6012
rect 22758 6010 22782 6012
rect 22838 6010 22862 6012
rect 22918 6010 22924 6012
rect 22678 5958 22680 6010
rect 22860 5958 22862 6010
rect 22616 5956 22622 5958
rect 22678 5956 22702 5958
rect 22758 5956 22782 5958
rect 22838 5956 22862 5958
rect 22918 5956 22924 5958
rect 22616 5947 22924 5956
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22652 5908 22704 5914
rect 22652 5850 22704 5856
rect 22664 5778 22692 5850
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 23032 5710 23060 7670
rect 23492 7410 23520 8774
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22388 4146 22416 5510
rect 22928 5296 22980 5302
rect 23032 5284 23060 5646
rect 22980 5256 23060 5284
rect 22928 5238 22980 5244
rect 22616 4924 22924 4933
rect 22616 4922 22622 4924
rect 22678 4922 22702 4924
rect 22758 4922 22782 4924
rect 22838 4922 22862 4924
rect 22918 4922 22924 4924
rect 22678 4870 22680 4922
rect 22860 4870 22862 4922
rect 22616 4868 22622 4870
rect 22678 4868 22702 4870
rect 22758 4868 22782 4870
rect 22838 4868 22862 4870
rect 22918 4868 22924 4870
rect 22616 4859 22924 4868
rect 23032 4690 23060 5256
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21376 3194 21404 3402
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 3194 21588 3334
rect 21652 3194 21680 3878
rect 21744 3194 21772 4014
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 17604 734 17816 762
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19444 762 19472 2382
rect 20088 1306 20116 2382
rect 20088 1278 20300 1306
rect 19628 870 19748 898
rect 19628 762 19656 870
rect 19720 800 19748 870
rect 20272 800 20300 1278
rect 20824 800 20852 2450
rect 21376 800 21404 2994
rect 22112 2650 22140 4082
rect 22192 4004 22244 4010
rect 22192 3946 22244 3952
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22204 2446 22232 3946
rect 22616 3836 22924 3845
rect 22616 3834 22622 3836
rect 22678 3834 22702 3836
rect 22758 3834 22782 3836
rect 22838 3834 22862 3836
rect 22918 3834 22924 3836
rect 22678 3782 22680 3834
rect 22860 3782 22862 3834
rect 22616 3780 22622 3782
rect 22678 3780 22702 3782
rect 22758 3780 22782 3782
rect 22838 3780 22862 3782
rect 22918 3780 22924 3782
rect 22616 3771 22924 3780
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22296 2582 22324 3674
rect 22744 3664 22796 3670
rect 22744 3606 22796 3612
rect 22756 3534 22784 3606
rect 22836 3596 22888 3602
rect 23032 3584 23060 4626
rect 23124 4282 23152 6258
rect 23400 6118 23428 6802
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23388 5704 23440 5710
rect 23386 5672 23388 5681
rect 23664 5704 23716 5710
rect 23440 5672 23442 5681
rect 23664 5646 23716 5652
rect 23386 5607 23442 5616
rect 23676 5370 23704 5646
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 22888 3556 23060 3584
rect 22836 3538 22888 3544
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 23124 3194 23152 4218
rect 23492 4146 23520 4422
rect 23584 4282 23612 5170
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23572 4072 23624 4078
rect 23860 4060 23888 12650
rect 23952 12434 23980 12922
rect 24504 12442 24532 13126
rect 24492 12436 24544 12442
rect 23952 12406 24072 12434
rect 24044 11626 24072 12406
rect 24492 12378 24544 12384
rect 24504 11898 24532 12378
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24228 11694 24256 11834
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 24044 9382 24072 11562
rect 24320 11354 24348 11630
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24504 11150 24532 11834
rect 24688 11694 24716 13194
rect 24768 12368 24820 12374
rect 24768 12310 24820 12316
rect 24780 12170 24808 12310
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24872 12102 24900 16594
rect 25056 16574 25084 17682
rect 25332 17270 25360 18226
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25424 17746 25452 17818
rect 25412 17740 25464 17746
rect 25412 17682 25464 17688
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25608 17542 25636 17614
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 24964 16546 25084 16574
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24872 11694 24900 12038
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24504 10674 24532 11086
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24872 9518 24900 11630
rect 24964 10690 24992 16546
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 25056 16114 25084 16390
rect 25608 16250 25636 17138
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 25700 16658 25728 16730
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25688 15496 25740 15502
rect 25688 15438 25740 15444
rect 25700 14822 25728 15438
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25700 14414 25728 14758
rect 25884 14618 25912 14894
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25780 14340 25832 14346
rect 25780 14282 25832 14288
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25056 11558 25084 12718
rect 25148 11830 25176 12786
rect 25240 12306 25268 13806
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 25332 12986 25360 13670
rect 25424 13394 25452 13670
rect 25792 13530 25820 14282
rect 25964 13796 26016 13802
rect 25964 13738 26016 13744
rect 25976 13530 26004 13738
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 25412 13388 25464 13394
rect 25412 13330 25464 13336
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25516 12306 25544 12582
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25596 12300 25648 12306
rect 25596 12242 25648 12248
rect 25240 12102 25268 12242
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 25240 11150 25268 12038
rect 25608 11898 25636 12242
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25228 11144 25280 11150
rect 25228 11086 25280 11092
rect 24964 10662 25176 10690
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24228 8566 24256 9454
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24320 8566 24348 9318
rect 24780 9110 24808 9318
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24308 8560 24360 8566
rect 24308 8502 24360 8508
rect 24228 8090 24256 8502
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 24504 8022 24532 8774
rect 24780 8498 24808 8774
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 23952 7546 23980 7754
rect 24504 7750 24532 7958
rect 24584 7948 24636 7954
rect 24584 7890 24636 7896
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24412 7546 24440 7686
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24596 7206 24624 7890
rect 24688 7546 24716 8434
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24780 7410 24808 8298
rect 24964 8090 24992 8366
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24872 7546 24900 7686
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 24964 7410 24992 8026
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24412 6458 24440 7142
rect 24596 6662 24624 7142
rect 25056 6866 25084 10542
rect 25148 8514 25176 10662
rect 25240 10606 25268 11086
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25700 10606 25728 11018
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25332 9994 25360 10542
rect 25320 9988 25372 9994
rect 25320 9930 25372 9936
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25148 8486 25268 8514
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 25148 6746 25176 8298
rect 25240 7478 25268 8486
rect 25228 7472 25280 7478
rect 25228 7414 25280 7420
rect 25240 7206 25268 7414
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 24964 6718 25176 6746
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 23952 4690 23980 5510
rect 24136 4690 24164 6054
rect 24412 5574 24440 6190
rect 24766 5672 24822 5681
rect 24964 5658 24992 6718
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6254 25176 6598
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 24822 5630 24992 5658
rect 24766 5607 24822 5616
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24412 5166 24440 5510
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 24780 5098 24808 5607
rect 24768 5092 24820 5098
rect 24768 5034 24820 5040
rect 25056 4690 25084 6054
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 23624 4032 23888 4060
rect 23572 4014 23624 4020
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23400 3194 23428 3946
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23768 3058 23796 3878
rect 24412 3738 24440 4626
rect 25148 4570 25176 6190
rect 25320 5636 25372 5642
rect 25320 5578 25372 5584
rect 24768 4548 24820 4554
rect 24768 4490 24820 4496
rect 25056 4542 25176 4570
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24596 4146 24624 4422
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 22616 2748 22924 2757
rect 22616 2746 22622 2748
rect 22678 2746 22702 2748
rect 22758 2746 22782 2748
rect 22838 2746 22862 2748
rect 22918 2746 22924 2748
rect 22678 2694 22680 2746
rect 22860 2694 22862 2746
rect 22616 2692 22622 2694
rect 22678 2692 22702 2694
rect 22758 2692 22782 2694
rect 22838 2692 22862 2694
rect 22918 2692 22924 2694
rect 22616 2683 22924 2692
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 21928 800 21956 2382
rect 22480 800 22508 2450
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23032 870 23152 898
rect 23032 800 23060 870
rect 19444 734 19656 762
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23124 762 23152 870
rect 23400 762 23428 2382
rect 23492 1578 23520 2790
rect 24044 2650 24072 3334
rect 24136 3194 24164 3402
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 23492 1550 23612 1578
rect 23584 800 23612 1550
rect 24136 800 24164 2926
rect 24320 2774 24348 3674
rect 24780 3602 24808 4490
rect 25056 3602 25084 4542
rect 25332 4146 25360 5578
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25424 4026 25452 5102
rect 25516 4554 25544 9454
rect 25792 8974 25820 9522
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25792 8498 25820 8570
rect 25976 8498 26004 9318
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25872 7948 25924 7954
rect 25872 7890 25924 7896
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25608 7546 25636 7686
rect 25700 7546 25728 7686
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25884 7478 25912 7890
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 25976 6458 26004 8434
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25608 5234 25636 6394
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25332 3998 25452 4026
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25056 3398 25084 3538
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 24412 3194 24440 3334
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 25148 2774 25176 3878
rect 25332 3602 25360 3998
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 24320 2746 24440 2774
rect 25148 2746 25360 2774
rect 24412 2650 24440 2746
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 25332 2446 25360 2746
rect 25608 2650 25636 4082
rect 25700 3058 25728 4150
rect 25884 4146 25912 5510
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 26068 4026 26096 18566
rect 26252 17882 26280 18566
rect 26620 17882 26648 18702
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 26148 17808 26200 17814
rect 26148 17750 26200 17756
rect 26974 17776 27030 17785
rect 26160 16590 26188 17750
rect 26332 17740 26384 17746
rect 26974 17711 26976 17720
rect 26332 17682 26384 17688
rect 27028 17711 27030 17720
rect 26976 17682 27028 17688
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26252 16658 26280 17070
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26252 15570 26280 16594
rect 26344 16250 26372 17682
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26620 16726 26648 16934
rect 26608 16720 26660 16726
rect 26608 16662 26660 16668
rect 26988 16522 27016 17682
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 13938 26188 14214
rect 26436 13938 26464 14486
rect 26528 14482 26556 15302
rect 26620 15042 26648 15846
rect 26700 15564 26752 15570
rect 26700 15506 26752 15512
rect 26712 15162 26740 15506
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26620 15014 26740 15042
rect 26712 14822 26740 15014
rect 26804 14890 26832 15914
rect 27080 15450 27108 18770
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 27264 18426 27292 18566
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 17814 27660 18022
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27356 16998 27384 17478
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 27356 16658 27384 16934
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27632 16250 27660 17614
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27896 17536 27948 17542
rect 27896 17478 27948 17484
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27448 15706 27476 16186
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27252 15496 27304 15502
rect 27080 15444 27252 15450
rect 27080 15438 27304 15444
rect 27080 15422 27292 15438
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26332 12912 26384 12918
rect 26332 12854 26384 12860
rect 26344 12374 26372 12854
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26436 11762 26464 13874
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26528 12442 26556 12582
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26712 12170 26740 14758
rect 26700 12164 26752 12170
rect 26700 12106 26752 12112
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26436 10146 26464 11698
rect 26516 11008 26568 11014
rect 26516 10950 26568 10956
rect 26528 10674 26556 10950
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26712 10470 26740 12106
rect 26792 12096 26844 12102
rect 26792 12038 26844 12044
rect 26804 11898 26832 12038
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26436 10118 26648 10146
rect 26424 9988 26476 9994
rect 26424 9930 26476 9936
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26344 9518 26372 9862
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26160 8906 26188 9454
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 26252 8634 26280 9454
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26332 8424 26384 8430
rect 26252 8384 26332 8412
rect 26252 7886 26280 8384
rect 26332 8366 26384 8372
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26252 7750 26280 7822
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 26148 7472 26200 7478
rect 26148 7414 26200 7420
rect 26160 6118 26188 7414
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26160 5914 26188 6054
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 26252 5778 26280 7686
rect 26436 6458 26464 9930
rect 26516 9580 26568 9586
rect 26516 9522 26568 9528
rect 26528 9382 26556 9522
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26620 8566 26648 10118
rect 27080 9654 27108 15422
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27540 14074 27568 14214
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27264 12782 27292 13126
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27356 9926 27384 10610
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 27356 9654 27384 9862
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26608 8356 26660 8362
rect 26608 8298 26660 8304
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 26424 6452 26476 6458
rect 26424 6394 26476 6400
rect 26436 5778 26464 6394
rect 26240 5772 26292 5778
rect 26240 5714 26292 5720
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26148 5092 26200 5098
rect 26148 5034 26200 5040
rect 26160 4078 26188 5034
rect 26252 4706 26280 5714
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26344 5030 26372 5646
rect 26332 5024 26384 5030
rect 26332 4966 26384 4972
rect 26344 4826 26372 4966
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26252 4678 26372 4706
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 25884 3998 26096 4026
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 25792 3602 25820 3878
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 25884 3058 25912 3998
rect 26252 3602 26280 4558
rect 26344 4486 26372 4678
rect 26424 4548 26476 4554
rect 26424 4490 26476 4496
rect 26332 4480 26384 4486
rect 26332 4422 26384 4428
rect 26344 4162 26372 4422
rect 26436 4282 26464 4490
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 26344 4134 26464 4162
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25872 2508 25924 2514
rect 25872 2450 25924 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25320 2440 25372 2446
rect 25320 2382 25372 2388
rect 24596 1306 24624 2382
rect 24596 1278 24716 1306
rect 24688 800 24716 1278
rect 25240 800 25268 2382
rect 25884 1306 25912 2450
rect 25792 1278 25912 1306
rect 25792 800 25820 1278
rect 26344 800 26372 4014
rect 26436 3534 26464 4134
rect 26528 4010 26556 6666
rect 26620 5370 26648 8298
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 26620 4214 26648 4422
rect 26608 4208 26660 4214
rect 26608 4150 26660 4156
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26712 3738 26740 9522
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26896 7478 26924 7686
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 27080 5302 27108 9590
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 27172 9382 27200 9454
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 27172 6662 27200 9318
rect 27356 9178 27384 9590
rect 27724 9586 27752 17478
rect 27908 16590 27936 17478
rect 28092 16998 28120 18566
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28644 17338 28672 18158
rect 28632 17332 28684 17338
rect 28632 17274 28684 17280
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 28092 16250 28120 16390
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 28368 16114 28396 16594
rect 28644 16574 28672 17274
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28920 16794 28948 16934
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28552 16546 28672 16574
rect 28552 16114 28580 16546
rect 28816 16448 28868 16454
rect 28816 16390 28868 16396
rect 28828 16114 28856 16390
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28540 16108 28592 16114
rect 28540 16050 28592 16056
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28000 15570 28028 16050
rect 29012 15978 29040 19450
rect 29472 19310 29500 20470
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29564 19514 29592 20198
rect 29748 19990 29776 20334
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29736 19984 29788 19990
rect 29736 19926 29788 19932
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29748 19378 29776 19926
rect 30116 19922 30144 20198
rect 30576 19922 30604 20402
rect 30760 19922 30788 20538
rect 30852 20534 30880 21286
rect 31668 21072 31720 21078
rect 31668 21014 31720 21020
rect 31024 20936 31076 20942
rect 31024 20878 31076 20884
rect 30840 20528 30892 20534
rect 30840 20470 30892 20476
rect 31036 20262 31064 20878
rect 31680 20602 31708 21014
rect 35360 20942 35388 21354
rect 37060 21244 37368 21253
rect 37060 21242 37066 21244
rect 37122 21242 37146 21244
rect 37202 21242 37226 21244
rect 37282 21242 37306 21244
rect 37362 21242 37368 21244
rect 37122 21190 37124 21242
rect 37304 21190 37306 21242
rect 37060 21188 37066 21190
rect 37122 21188 37146 21190
rect 37202 21188 37226 21190
rect 37282 21188 37306 21190
rect 37362 21188 37368 21190
rect 37060 21179 37368 21188
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 35348 20936 35400 20942
rect 35348 20878 35400 20884
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 32876 20602 32904 20878
rect 33416 20800 33468 20806
rect 33416 20742 33468 20748
rect 31668 20596 31720 20602
rect 31588 20556 31668 20584
rect 31024 20256 31076 20262
rect 31024 20198 31076 20204
rect 30104 19916 30156 19922
rect 30104 19858 30156 19864
rect 30196 19916 30248 19922
rect 30196 19858 30248 19864
rect 30564 19916 30616 19922
rect 30564 19858 30616 19864
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30932 19916 30984 19922
rect 30932 19858 30984 19864
rect 29838 19612 30146 19621
rect 29838 19610 29844 19612
rect 29900 19610 29924 19612
rect 29980 19610 30004 19612
rect 30060 19610 30084 19612
rect 30140 19610 30146 19612
rect 29900 19558 29902 19610
rect 30082 19558 30084 19610
rect 29838 19556 29844 19558
rect 29900 19556 29924 19558
rect 29980 19556 30004 19558
rect 30060 19556 30084 19558
rect 30140 19556 30146 19558
rect 29838 19547 30146 19556
rect 30208 19446 30236 19858
rect 30196 19440 30248 19446
rect 30196 19382 30248 19388
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29460 19304 29512 19310
rect 29460 19246 29512 19252
rect 29288 18970 29316 19246
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29092 18624 29144 18630
rect 29092 18566 29144 18572
rect 29104 18222 29132 18566
rect 29472 18290 29500 19246
rect 30852 18970 30880 19314
rect 30840 18964 30892 18970
rect 30840 18906 30892 18912
rect 30656 18828 30708 18834
rect 30656 18770 30708 18776
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 29838 18524 30146 18533
rect 29838 18522 29844 18524
rect 29900 18522 29924 18524
rect 29980 18522 30004 18524
rect 30060 18522 30084 18524
rect 30140 18522 30146 18524
rect 29900 18470 29902 18522
rect 30082 18470 30084 18522
rect 29838 18468 29844 18470
rect 29900 18468 29924 18470
rect 29980 18468 30004 18470
rect 30060 18468 30084 18470
rect 30140 18468 30146 18470
rect 29838 18459 30146 18468
rect 30392 18290 30420 18566
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 29104 16726 29132 18158
rect 29276 18080 29328 18086
rect 29276 18022 29328 18028
rect 29288 17746 29316 18022
rect 29276 17740 29328 17746
rect 29276 17682 29328 17688
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 29380 17338 29408 17478
rect 29368 17332 29420 17338
rect 29368 17274 29420 17280
rect 29092 16720 29144 16726
rect 29472 16674 29500 18226
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30208 17882 30236 18158
rect 30196 17876 30248 17882
rect 30196 17818 30248 17824
rect 30392 17678 30420 18226
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 29838 17436 30146 17445
rect 29838 17434 29844 17436
rect 29900 17434 29924 17436
rect 29980 17434 30004 17436
rect 30060 17434 30084 17436
rect 30140 17434 30146 17436
rect 29900 17382 29902 17434
rect 30082 17382 30084 17434
rect 29838 17380 29844 17382
rect 29900 17380 29924 17382
rect 29980 17380 30004 17382
rect 30060 17380 30084 17382
rect 30140 17380 30146 17382
rect 29838 17371 30146 17380
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 29092 16662 29144 16668
rect 29380 16658 29500 16674
rect 29368 16652 29500 16658
rect 29420 16646 29500 16652
rect 29368 16594 29420 16600
rect 29000 15972 29052 15978
rect 29052 15932 29132 15960
rect 29000 15914 29052 15920
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 28092 15706 28120 15846
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 27988 15564 28040 15570
rect 27988 15506 28040 15512
rect 28092 14958 28120 15642
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28184 15026 28212 15302
rect 28276 15162 28304 15370
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 28080 14952 28132 14958
rect 28080 14894 28132 14900
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28092 14074 28120 14350
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 28092 12918 28120 13670
rect 28184 12986 28212 13738
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 28080 12912 28132 12918
rect 28080 12854 28132 12860
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27816 9382 27844 11086
rect 28356 11008 28408 11014
rect 28356 10950 28408 10956
rect 28368 10674 28396 10950
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28460 9602 28488 15438
rect 29000 15428 29052 15434
rect 29000 15370 29052 15376
rect 29012 15162 29040 15370
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28644 13326 28672 14214
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28828 13190 28856 14350
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 29012 14074 29040 14214
rect 29000 14068 29052 14074
rect 29000 14010 29052 14016
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28828 12986 28856 13126
rect 28816 12980 28868 12986
rect 29104 12968 29132 15932
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29288 14618 29316 15302
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29288 14074 29316 14554
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 28816 12922 28868 12928
rect 29012 12940 29132 12968
rect 28816 12708 28868 12714
rect 28816 12650 28868 12656
rect 28828 12306 28856 12650
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28644 10538 28672 11086
rect 28632 10532 28684 10538
rect 28632 10474 28684 10480
rect 28736 10470 28764 11630
rect 28908 11552 28960 11558
rect 28908 11494 28960 11500
rect 28724 10464 28776 10470
rect 28724 10406 28776 10412
rect 28920 10062 28948 11494
rect 29012 11354 29040 12940
rect 29196 12850 29224 13874
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29380 13530 29408 13670
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29104 12442 29132 12786
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28368 9574 28488 9602
rect 28368 9518 28396 9574
rect 28356 9512 28408 9518
rect 28356 9454 28408 9460
rect 28264 9444 28316 9450
rect 28264 9386 28316 9392
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27540 8634 27568 8774
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27540 6798 27568 8366
rect 27620 7812 27672 7818
rect 27620 7754 27672 7760
rect 27632 7546 27660 7754
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 27160 6656 27212 6662
rect 27160 6598 27212 6604
rect 27908 6322 27936 6734
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27068 5296 27120 5302
rect 27068 5238 27120 5244
rect 27620 4752 27672 4758
rect 27620 4694 27672 4700
rect 27344 4208 27396 4214
rect 27344 4150 27396 4156
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 27068 4004 27120 4010
rect 27068 3946 27120 3952
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26620 3466 26648 3674
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 26608 3460 26660 3466
rect 26608 3402 26660 3408
rect 26896 3194 26924 3470
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 26896 800 26924 2926
rect 26988 2774 27016 3878
rect 27080 3602 27108 3946
rect 27264 3738 27292 4082
rect 27356 4049 27384 4150
rect 27436 4072 27488 4078
rect 27342 4040 27398 4049
rect 27436 4014 27488 4020
rect 27342 3975 27398 3984
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 27356 3097 27384 3878
rect 27342 3088 27398 3097
rect 27342 3023 27398 3032
rect 26988 2746 27108 2774
rect 27080 2650 27108 2746
rect 27448 2650 27476 4014
rect 27632 2774 27660 4694
rect 27724 4690 27752 5714
rect 27712 4684 27764 4690
rect 27712 4626 27764 4632
rect 27908 4010 27936 6258
rect 28276 5914 28304 9386
rect 29012 9382 29040 11018
rect 29196 10690 29224 12786
rect 29276 12776 29328 12782
rect 29276 12718 29328 12724
rect 29288 12374 29316 12718
rect 29276 12368 29328 12374
rect 29276 12310 29328 12316
rect 29276 11552 29328 11558
rect 29276 11494 29328 11500
rect 29104 10674 29224 10690
rect 29092 10668 29224 10674
rect 29144 10662 29224 10668
rect 29092 10610 29144 10616
rect 29104 9722 29132 10610
rect 29288 9926 29316 11494
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 28816 9104 28868 9110
rect 28816 9046 28868 9052
rect 28828 8974 28856 9046
rect 28816 8968 28868 8974
rect 28816 8910 28868 8916
rect 28908 8968 28960 8974
rect 28908 8910 28960 8916
rect 28920 8809 28948 8910
rect 29104 8906 29132 9658
rect 29368 9580 29420 9586
rect 29368 9522 29420 9528
rect 29380 9178 29408 9522
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29092 8900 29144 8906
rect 29092 8842 29144 8848
rect 28906 8800 28962 8809
rect 28906 8735 28962 8744
rect 29472 8634 29500 16646
rect 29564 10810 29592 16934
rect 30484 16590 30512 18022
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 29838 16348 30146 16357
rect 29838 16346 29844 16348
rect 29900 16346 29924 16348
rect 29980 16346 30004 16348
rect 30060 16346 30084 16348
rect 30140 16346 30146 16348
rect 29900 16294 29902 16346
rect 30082 16294 30084 16346
rect 29838 16292 29844 16294
rect 29900 16292 29924 16294
rect 29980 16292 30004 16294
rect 30060 16292 30084 16294
rect 30140 16292 30146 16294
rect 29838 16283 30146 16292
rect 30392 16250 30420 16390
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29656 15638 29684 16050
rect 30196 15904 30248 15910
rect 30196 15846 30248 15852
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 29644 15632 29696 15638
rect 29644 15574 29696 15580
rect 30208 15502 30236 15846
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 29838 15260 30146 15269
rect 29838 15258 29844 15260
rect 29900 15258 29924 15260
rect 29980 15258 30004 15260
rect 30060 15258 30084 15260
rect 30140 15258 30146 15260
rect 29900 15206 29902 15258
rect 30082 15206 30084 15258
rect 29838 15204 29844 15206
rect 29900 15204 29924 15206
rect 29980 15204 30004 15206
rect 30060 15204 30084 15206
rect 30140 15204 30146 15206
rect 29838 15195 30146 15204
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29748 11898 29776 14350
rect 29838 14172 30146 14181
rect 29838 14170 29844 14172
rect 29900 14170 29924 14172
rect 29980 14170 30004 14172
rect 30060 14170 30084 14172
rect 30140 14170 30146 14172
rect 29900 14118 29902 14170
rect 30082 14118 30084 14170
rect 29838 14116 29844 14118
rect 29900 14116 29924 14118
rect 29980 14116 30004 14118
rect 30060 14116 30084 14118
rect 30140 14116 30146 14118
rect 29838 14107 30146 14116
rect 29838 13084 30146 13093
rect 29838 13082 29844 13084
rect 29900 13082 29924 13084
rect 29980 13082 30004 13084
rect 30060 13082 30084 13084
rect 30140 13082 30146 13084
rect 29900 13030 29902 13082
rect 30082 13030 30084 13082
rect 29838 13028 29844 13030
rect 29900 13028 29924 13030
rect 29980 13028 30004 13030
rect 30060 13028 30084 13030
rect 30140 13028 30146 13030
rect 29838 13019 30146 13028
rect 30196 12844 30248 12850
rect 30196 12786 30248 12792
rect 29838 11996 30146 12005
rect 29838 11994 29844 11996
rect 29900 11994 29924 11996
rect 29980 11994 30004 11996
rect 30060 11994 30084 11996
rect 30140 11994 30146 11996
rect 29900 11942 29902 11994
rect 30082 11942 30084 11994
rect 29838 11940 29844 11942
rect 29900 11940 29924 11942
rect 29980 11940 30004 11942
rect 30060 11940 30084 11942
rect 30140 11940 30146 11942
rect 29838 11931 30146 11940
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29748 10690 29776 11290
rect 29838 10908 30146 10917
rect 29838 10906 29844 10908
rect 29900 10906 29924 10908
rect 29980 10906 30004 10908
rect 30060 10906 30084 10908
rect 30140 10906 30146 10908
rect 29900 10854 29902 10906
rect 30082 10854 30084 10906
rect 29838 10852 29844 10854
rect 29900 10852 29924 10854
rect 29980 10852 30004 10854
rect 30060 10852 30084 10854
rect 30140 10852 30146 10854
rect 29838 10843 30146 10852
rect 29748 10662 30052 10690
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29736 10056 29788 10062
rect 29932 10033 29960 10542
rect 30024 10198 30052 10662
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 29736 9998 29788 10004
rect 29918 10024 29974 10033
rect 29564 9722 29592 9998
rect 29552 9716 29604 9722
rect 29748 9704 29776 9998
rect 29918 9959 29974 9968
rect 29838 9820 30146 9829
rect 29838 9818 29844 9820
rect 29900 9818 29924 9820
rect 29980 9818 30004 9820
rect 30060 9818 30084 9820
rect 30140 9818 30146 9820
rect 29900 9766 29902 9818
rect 30082 9766 30084 9818
rect 29838 9764 29844 9766
rect 29900 9764 29924 9766
rect 29980 9764 30004 9766
rect 30060 9764 30084 9766
rect 30140 9764 30146 9766
rect 29838 9755 30146 9764
rect 30104 9716 30156 9722
rect 29748 9676 30104 9704
rect 29552 9658 29604 9664
rect 30104 9658 30156 9664
rect 29460 8628 29512 8634
rect 29460 8570 29512 8576
rect 29564 8498 29592 9658
rect 29736 8900 29788 8906
rect 29736 8842 29788 8848
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28644 7546 28672 7822
rect 29000 7812 29052 7818
rect 29000 7754 29052 7760
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 28264 5908 28316 5914
rect 28264 5850 28316 5856
rect 28448 5568 28500 5574
rect 28448 5510 28500 5516
rect 28460 5234 28488 5510
rect 28920 5370 28948 6258
rect 28908 5364 28960 5370
rect 28908 5306 28960 5312
rect 28448 5228 28500 5234
rect 28448 5170 28500 5176
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 27896 4004 27948 4010
rect 27896 3946 27948 3952
rect 27804 3936 27856 3942
rect 27804 3878 27856 3884
rect 27712 3120 27764 3126
rect 27816 3097 27844 3878
rect 27712 3062 27764 3068
rect 27802 3088 27858 3097
rect 27540 2746 27660 2774
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27448 800 27476 2450
rect 27540 2446 27568 2746
rect 27724 2446 27752 3062
rect 27802 3023 27858 3032
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 28000 800 28028 4558
rect 28184 3602 28212 4966
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 28184 3398 28212 3538
rect 28356 3460 28408 3466
rect 28356 3402 28408 3408
rect 28172 3392 28224 3398
rect 28172 3334 28224 3340
rect 28368 3194 28396 3402
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 28460 2990 28488 3334
rect 28552 3194 28580 3334
rect 28920 3194 28948 3334
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28448 2984 28500 2990
rect 28448 2926 28500 2932
rect 28368 1578 28396 2926
rect 29012 2650 29040 7754
rect 29104 5370 29132 8434
rect 29656 8090 29684 8774
rect 29748 8634 29776 8842
rect 29838 8732 30146 8741
rect 29838 8730 29844 8732
rect 29900 8730 29924 8732
rect 29980 8730 30004 8732
rect 30060 8730 30084 8732
rect 30140 8730 30146 8732
rect 29900 8678 29902 8730
rect 30082 8678 30084 8730
rect 29838 8676 29844 8678
rect 29900 8676 29924 8678
rect 29980 8676 30004 8678
rect 30060 8676 30084 8678
rect 30140 8676 30146 8678
rect 29838 8667 30146 8676
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29196 6798 29224 7686
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 29288 5710 29316 7482
rect 29380 6458 29408 7686
rect 29644 7336 29696 7342
rect 29644 7278 29696 7284
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29564 6458 29592 7142
rect 29656 6730 29684 7278
rect 29748 7206 29776 7822
rect 29838 7644 30146 7653
rect 29838 7642 29844 7644
rect 29900 7642 29924 7644
rect 29980 7642 30004 7644
rect 30060 7642 30084 7644
rect 30140 7642 30146 7644
rect 29900 7590 29902 7642
rect 30082 7590 30084 7642
rect 29838 7588 29844 7590
rect 29900 7588 29924 7590
rect 29980 7588 30004 7590
rect 30060 7588 30084 7590
rect 30140 7588 30146 7590
rect 29838 7579 30146 7588
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29644 6724 29696 6730
rect 29644 6666 29696 6672
rect 29368 6452 29420 6458
rect 29368 6394 29420 6400
rect 29552 6452 29604 6458
rect 29552 6394 29604 6400
rect 29564 5914 29592 6394
rect 29748 6322 29776 7142
rect 29838 6556 30146 6565
rect 29838 6554 29844 6556
rect 29900 6554 29924 6556
rect 29980 6554 30004 6556
rect 30060 6554 30084 6556
rect 30140 6554 30146 6556
rect 29900 6502 29902 6554
rect 30082 6502 30084 6554
rect 29838 6500 29844 6502
rect 29900 6500 29924 6502
rect 29980 6500 30004 6502
rect 30060 6500 30084 6502
rect 30140 6500 30146 6502
rect 29838 6491 30146 6500
rect 29736 6316 29788 6322
rect 29736 6258 29788 6264
rect 29644 6180 29696 6186
rect 29644 6122 29696 6128
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29276 5704 29328 5710
rect 29196 5664 29276 5692
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29196 4706 29224 5664
rect 29276 5646 29328 5652
rect 29552 5636 29604 5642
rect 29552 5578 29604 5584
rect 29564 5370 29592 5578
rect 29552 5364 29604 5370
rect 29552 5306 29604 5312
rect 29656 5234 29684 6122
rect 30012 6112 30064 6118
rect 30010 6080 30012 6089
rect 30064 6080 30066 6089
rect 30010 6015 30066 6024
rect 29838 5468 30146 5477
rect 29838 5466 29844 5468
rect 29900 5466 29924 5468
rect 29980 5466 30004 5468
rect 30060 5466 30084 5468
rect 30140 5466 30146 5468
rect 29900 5414 29902 5466
rect 30082 5414 30084 5466
rect 29838 5412 29844 5414
rect 29900 5412 29924 5414
rect 29980 5412 30004 5414
rect 30060 5412 30084 5414
rect 30140 5412 30146 5414
rect 29838 5403 30146 5412
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 29104 4678 29224 4706
rect 29104 3398 29132 4678
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29196 3738 29224 4558
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 28368 1550 28580 1578
rect 28552 800 28580 1550
rect 29104 800 29132 2926
rect 29288 2922 29316 5170
rect 29736 5160 29788 5166
rect 29736 5102 29788 5108
rect 29644 5024 29696 5030
rect 29644 4966 29696 4972
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29368 4480 29420 4486
rect 29368 4422 29420 4428
rect 29380 4214 29408 4422
rect 29564 4282 29592 4558
rect 29552 4276 29604 4282
rect 29552 4218 29604 4224
rect 29368 4208 29420 4214
rect 29368 4150 29420 4156
rect 29656 4128 29684 4966
rect 29748 4826 29776 5102
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 29748 4282 29776 4762
rect 29838 4380 30146 4389
rect 29838 4378 29844 4380
rect 29900 4378 29924 4380
rect 29980 4378 30004 4380
rect 30060 4378 30084 4380
rect 30140 4378 30146 4380
rect 29900 4326 29902 4378
rect 30082 4326 30084 4378
rect 29838 4324 29844 4326
rect 29900 4324 29924 4326
rect 29980 4324 30004 4326
rect 30060 4324 30084 4326
rect 30140 4324 30146 4326
rect 29838 4315 30146 4324
rect 29736 4276 29788 4282
rect 29736 4218 29788 4224
rect 29736 4140 29788 4146
rect 29656 4100 29736 4128
rect 29736 4082 29788 4088
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29564 3194 29592 3878
rect 30208 3505 30236 12786
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30300 12186 30328 12718
rect 30392 12434 30420 15846
rect 30668 14278 30696 18770
rect 30944 16250 30972 19858
rect 31208 19712 31260 19718
rect 31208 19654 31260 19660
rect 31220 19514 31248 19654
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31128 16454 31156 17614
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 30932 16244 30984 16250
rect 30932 16186 30984 16192
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 31036 14618 31064 15302
rect 31024 14612 31076 14618
rect 31024 14554 31076 14560
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30656 14272 30708 14278
rect 30656 14214 30708 14220
rect 31392 14272 31444 14278
rect 31392 14214 31444 14220
rect 30576 14074 30604 14214
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 30668 13734 30696 14214
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 30748 13932 30800 13938
rect 30748 13874 30800 13880
rect 30656 13728 30708 13734
rect 30656 13670 30708 13676
rect 30760 13326 30788 13874
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30944 13530 30972 13738
rect 30932 13524 30984 13530
rect 30932 13466 30984 13472
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30748 13320 30800 13326
rect 30800 13280 30880 13308
rect 30748 13262 30800 13268
rect 30484 12986 30512 13262
rect 30576 12986 30604 13262
rect 30748 13184 30800 13190
rect 30748 13126 30800 13132
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30760 12442 30788 13126
rect 30656 12436 30708 12442
rect 30392 12406 30512 12434
rect 30300 12158 30420 12186
rect 30392 12102 30420 12158
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30392 11898 30420 12038
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 30300 10674 30328 10950
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 30288 10532 30340 10538
rect 30288 10474 30340 10480
rect 30300 10130 30328 10474
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 30288 9920 30340 9926
rect 30288 9862 30340 9868
rect 30300 9382 30328 9862
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 30300 8430 30328 9318
rect 30392 8974 30420 9318
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30392 8430 30420 8774
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30300 7342 30328 8366
rect 30288 7336 30340 7342
rect 30288 7278 30340 7284
rect 30300 6934 30328 7278
rect 30288 6928 30340 6934
rect 30484 6914 30512 12406
rect 30656 12378 30708 12384
rect 30748 12436 30800 12442
rect 30748 12378 30800 12384
rect 30668 10810 30696 12378
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30852 10674 30880 13280
rect 31036 11898 31064 14010
rect 31404 13394 31432 14214
rect 31588 13734 31616 20556
rect 31668 20538 31720 20544
rect 32864 20596 32916 20602
rect 32864 20538 32916 20544
rect 31852 20256 31904 20262
rect 31852 20198 31904 20204
rect 33324 20256 33376 20262
rect 33324 20198 33376 20204
rect 31864 20058 31892 20198
rect 33336 20058 33364 20198
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 33324 20052 33376 20058
rect 33324 19994 33376 20000
rect 31864 17338 31892 19994
rect 33428 19378 33456 20742
rect 33600 19984 33652 19990
rect 33600 19926 33652 19932
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31956 18766 31984 19110
rect 33612 18834 33640 19926
rect 33704 19514 33732 20878
rect 34244 20800 34296 20806
rect 34244 20742 34296 20748
rect 34256 20602 34284 20742
rect 34244 20596 34296 20602
rect 34244 20538 34296 20544
rect 34152 20528 34204 20534
rect 34152 20470 34204 20476
rect 33968 20460 34020 20466
rect 33968 20402 34020 20408
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 33796 20058 33824 20334
rect 33784 20052 33836 20058
rect 33784 19994 33836 20000
rect 33980 19718 34008 20402
rect 34164 20074 34192 20470
rect 34336 20324 34388 20330
rect 34336 20266 34388 20272
rect 34164 20046 34284 20074
rect 34152 19916 34204 19922
rect 34152 19858 34204 19864
rect 33876 19712 33928 19718
rect 33876 19654 33928 19660
rect 33968 19712 34020 19718
rect 33968 19654 34020 19660
rect 33692 19508 33744 19514
rect 33692 19450 33744 19456
rect 33888 18902 33916 19654
rect 33876 18896 33928 18902
rect 33876 18838 33928 18844
rect 33600 18828 33652 18834
rect 33600 18770 33652 18776
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 33968 18216 34020 18222
rect 33968 18158 34020 18164
rect 33140 18080 33192 18086
rect 33140 18022 33192 18028
rect 33152 17746 33180 18022
rect 33140 17740 33192 17746
rect 33140 17682 33192 17688
rect 32772 17536 32824 17542
rect 32772 17478 32824 17484
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 31852 17332 31904 17338
rect 31852 17274 31904 17280
rect 31864 16794 31892 17274
rect 32784 17202 32812 17478
rect 33152 17338 33180 17478
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 32772 17196 32824 17202
rect 32772 17138 32824 17144
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 31852 16788 31904 16794
rect 31852 16730 31904 16736
rect 31680 14618 31708 16730
rect 32128 16584 32180 16590
rect 32128 16526 32180 16532
rect 32140 16250 32168 16526
rect 32680 16448 32732 16454
rect 32680 16390 32732 16396
rect 32128 16244 32180 16250
rect 32128 16186 32180 16192
rect 32692 15706 32720 16390
rect 32784 16250 32812 17138
rect 33324 17128 33376 17134
rect 33324 17070 33376 17076
rect 33336 16250 33364 17070
rect 33520 16998 33548 18158
rect 33980 17338 34008 18158
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 33508 16992 33560 16998
rect 33508 16934 33560 16940
rect 33508 16516 33560 16522
rect 33508 16458 33560 16464
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 33324 16244 33376 16250
rect 33324 16186 33376 16192
rect 33140 16108 33192 16114
rect 33140 16050 33192 16056
rect 33152 15706 33180 16050
rect 32680 15700 32732 15706
rect 32680 15642 32732 15648
rect 33140 15700 33192 15706
rect 33140 15642 33192 15648
rect 33336 15502 33364 16186
rect 33520 16046 33548 16458
rect 33508 16040 33560 16046
rect 33508 15982 33560 15988
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 33520 15162 33548 15982
rect 34060 15972 34112 15978
rect 34060 15914 34112 15920
rect 34072 15366 34100 15914
rect 34060 15360 34112 15366
rect 34060 15302 34112 15308
rect 33508 15156 33560 15162
rect 33508 15098 33560 15104
rect 33324 14816 33376 14822
rect 33324 14758 33376 14764
rect 31668 14612 31720 14618
rect 31668 14554 31720 14560
rect 31680 13938 31708 14554
rect 31852 14544 31904 14550
rect 31852 14486 31904 14492
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31576 13728 31628 13734
rect 31576 13670 31628 13676
rect 31864 13462 31892 14486
rect 33336 13734 33364 14758
rect 33324 13728 33376 13734
rect 33324 13670 33376 13676
rect 31852 13456 31904 13462
rect 31852 13398 31904 13404
rect 31392 13388 31444 13394
rect 31392 13330 31444 13336
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31484 13184 31536 13190
rect 31484 13126 31536 13132
rect 31576 13184 31628 13190
rect 31576 13126 31628 13132
rect 31496 12986 31524 13126
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 31588 12866 31616 13126
rect 31404 12838 31616 12866
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31128 11898 31156 12174
rect 31404 12102 31432 12838
rect 31484 12640 31536 12646
rect 31484 12582 31536 12588
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31024 11892 31076 11898
rect 31024 11834 31076 11840
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31496 10742 31524 12582
rect 31576 10804 31628 10810
rect 31576 10746 31628 10752
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30576 10130 30604 10406
rect 30564 10124 30616 10130
rect 30564 10066 30616 10072
rect 30748 10124 30800 10130
rect 30852 10112 30880 10610
rect 31588 10130 31616 10746
rect 30800 10084 30880 10112
rect 31576 10124 31628 10130
rect 30748 10066 30800 10072
rect 31576 10066 31628 10072
rect 31680 9926 31708 13194
rect 31852 13184 31904 13190
rect 31852 13126 31904 13132
rect 31864 12442 31892 13126
rect 31852 12436 31904 12442
rect 31852 12378 31904 12384
rect 32324 11898 32352 13262
rect 33520 12714 33548 15098
rect 34072 14618 34100 15302
rect 34060 14612 34112 14618
rect 34060 14554 34112 14560
rect 34060 13864 34112 13870
rect 34060 13806 34112 13812
rect 33600 13252 33652 13258
rect 33600 13194 33652 13200
rect 33508 12708 33560 12714
rect 33508 12650 33560 12656
rect 32772 12640 32824 12646
rect 32772 12582 32824 12588
rect 33140 12640 33192 12646
rect 33140 12582 33192 12588
rect 32784 12374 32812 12582
rect 32772 12368 32824 12374
rect 32772 12310 32824 12316
rect 33152 12306 33180 12582
rect 33612 12442 33640 13194
rect 33876 13184 33928 13190
rect 33876 13126 33928 13132
rect 33600 12436 33652 12442
rect 33600 12378 33652 12384
rect 33888 12306 33916 13126
rect 34072 12986 34100 13806
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33980 12442 34008 12786
rect 33968 12436 34020 12442
rect 33968 12378 34020 12384
rect 33140 12300 33192 12306
rect 33140 12242 33192 12248
rect 33876 12300 33928 12306
rect 33876 12242 33928 12248
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 34164 11694 34192 19858
rect 34256 18034 34284 20046
rect 34348 19786 34376 20266
rect 35360 19922 35388 20878
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 35820 19938 35848 20742
rect 35912 20262 35940 20878
rect 36728 20800 36780 20806
rect 36728 20742 36780 20748
rect 37464 20800 37516 20806
rect 37464 20742 37516 20748
rect 35992 20392 36044 20398
rect 35992 20334 36044 20340
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35912 20058 35940 20198
rect 35900 20052 35952 20058
rect 35900 19994 35952 20000
rect 35348 19916 35400 19922
rect 35820 19910 35940 19938
rect 35348 19858 35400 19864
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34336 19780 34388 19786
rect 34336 19722 34388 19728
rect 34348 19378 34376 19722
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34336 19372 34388 19378
rect 34336 19314 34388 19320
rect 34348 18970 34376 19314
rect 34440 19122 34468 19654
rect 34716 19514 34744 19790
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34520 19168 34572 19174
rect 34440 19116 34520 19122
rect 34440 19110 34572 19116
rect 34440 19094 34560 19110
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 34440 18630 34468 19094
rect 34428 18624 34480 18630
rect 34428 18566 34480 18572
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34612 18080 34664 18086
rect 34256 18006 34468 18034
rect 34612 18022 34664 18028
rect 34244 17740 34296 17746
rect 34244 17682 34296 17688
rect 34256 12850 34284 17682
rect 34336 16992 34388 16998
rect 34336 16934 34388 16940
rect 34348 16114 34376 16934
rect 34440 16130 34468 18006
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34532 16726 34560 17614
rect 34520 16720 34572 16726
rect 34520 16662 34572 16668
rect 34532 16250 34560 16662
rect 34624 16590 34652 18022
rect 34900 17134 34928 18566
rect 35360 17626 35388 19858
rect 35912 19854 35940 19910
rect 35624 19848 35676 19854
rect 35624 19790 35676 19796
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 35636 19446 35664 19790
rect 35624 19440 35676 19446
rect 35912 19394 35940 19790
rect 36004 19514 36032 20334
rect 36544 19712 36596 19718
rect 36544 19654 36596 19660
rect 35992 19508 36044 19514
rect 35992 19450 36044 19456
rect 35624 19382 35676 19388
rect 35820 19366 35940 19394
rect 36268 19440 36320 19446
rect 36268 19382 36320 19388
rect 36176 19372 36228 19378
rect 35820 19258 35848 19366
rect 36176 19314 36228 19320
rect 35544 19230 35848 19258
rect 35440 18080 35492 18086
rect 35440 18022 35492 18028
rect 35268 17598 35388 17626
rect 35268 17270 35296 17598
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 35360 17338 35388 17478
rect 35348 17332 35400 17338
rect 35348 17274 35400 17280
rect 35256 17264 35308 17270
rect 35256 17206 35308 17212
rect 34888 17128 34940 17134
rect 34888 17070 34940 17076
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 34612 16448 34664 16454
rect 34612 16390 34664 16396
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34336 16108 34388 16114
rect 34440 16102 34560 16130
rect 34336 16050 34388 16056
rect 34428 16040 34480 16046
rect 34428 15982 34480 15988
rect 34440 15706 34468 15982
rect 34428 15700 34480 15706
rect 34428 15642 34480 15648
rect 34532 15586 34560 16102
rect 34624 15910 34652 16390
rect 34612 15904 34664 15910
rect 34612 15846 34664 15852
rect 34716 15706 34744 16594
rect 34796 15904 34848 15910
rect 34796 15846 34848 15852
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 34440 15558 34560 15586
rect 34336 12912 34388 12918
rect 34336 12854 34388 12860
rect 34244 12844 34296 12850
rect 34244 12786 34296 12792
rect 34348 12374 34376 12854
rect 34440 12646 34468 15558
rect 34808 14600 34836 15846
rect 34716 14572 34836 14600
rect 34612 13864 34664 13870
rect 34612 13806 34664 13812
rect 34624 13326 34652 13806
rect 34612 13320 34664 13326
rect 34612 13262 34664 13268
rect 34428 12640 34480 12646
rect 34428 12582 34480 12588
rect 34336 12368 34388 12374
rect 34336 12310 34388 12316
rect 34348 11762 34376 12310
rect 34336 11756 34388 11762
rect 34336 11698 34388 11704
rect 34440 11694 34468 12582
rect 34716 12434 34744 14572
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34808 14074 34836 14418
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34716 12406 34836 12434
rect 34612 12232 34664 12238
rect 34612 12174 34664 12180
rect 34152 11688 34204 11694
rect 34152 11630 34204 11636
rect 34428 11688 34480 11694
rect 34428 11630 34480 11636
rect 32956 11552 33008 11558
rect 32956 11494 33008 11500
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 32968 11150 32996 11494
rect 33796 11354 33824 11494
rect 33888 11354 33916 11494
rect 33784 11348 33836 11354
rect 33784 11290 33836 11296
rect 33876 11348 33928 11354
rect 33876 11290 33928 11296
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32956 11144 33008 11150
rect 32956 11086 33008 11092
rect 32508 10470 32536 11086
rect 33600 11076 33652 11082
rect 33600 11018 33652 11024
rect 33612 10674 33640 11018
rect 33600 10668 33652 10674
rect 33600 10610 33652 10616
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31668 9920 31720 9926
rect 31668 9862 31720 9868
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30668 8634 30696 9522
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30944 7750 30972 8978
rect 30932 7744 30984 7750
rect 30932 7686 30984 7692
rect 30288 6870 30340 6876
rect 30392 6886 30512 6914
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 30300 6458 30328 6598
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 30288 5024 30340 5030
rect 30392 5012 30420 6886
rect 30656 6792 30708 6798
rect 30656 6734 30708 6740
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 6225 30512 6598
rect 30470 6216 30526 6225
rect 30470 6151 30526 6160
rect 30564 6180 30616 6186
rect 30564 6122 30616 6128
rect 30576 5953 30604 6122
rect 30562 5944 30618 5953
rect 30562 5879 30618 5888
rect 30576 5642 30604 5879
rect 30668 5778 30696 6734
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30852 6322 30880 6598
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30564 5636 30616 5642
rect 30564 5578 30616 5584
rect 30668 5370 30696 5714
rect 30748 5636 30800 5642
rect 30748 5578 30800 5584
rect 30656 5364 30708 5370
rect 30656 5306 30708 5312
rect 30340 4984 30420 5012
rect 30656 5024 30708 5030
rect 30288 4966 30340 4972
rect 30656 4966 30708 4972
rect 30564 4616 30616 4622
rect 30564 4558 30616 4564
rect 30288 4480 30340 4486
rect 30288 4422 30340 4428
rect 30300 3602 30328 4422
rect 30576 4282 30604 4558
rect 30564 4276 30616 4282
rect 30564 4218 30616 4224
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30194 3496 30250 3505
rect 30194 3431 30250 3440
rect 29838 3292 30146 3301
rect 29838 3290 29844 3292
rect 29900 3290 29924 3292
rect 29980 3290 30004 3292
rect 30060 3290 30084 3292
rect 30140 3290 30146 3292
rect 29900 3238 29902 3290
rect 30082 3238 30084 3290
rect 29838 3236 29844 3238
rect 29900 3236 29924 3238
rect 29980 3236 30004 3238
rect 30060 3236 30084 3238
rect 30140 3236 30146 3238
rect 29838 3227 30146 3236
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29276 2916 29328 2922
rect 29276 2858 29328 2864
rect 30668 2446 30696 4966
rect 30760 4010 30788 5578
rect 31036 5234 31064 9862
rect 31484 9716 31536 9722
rect 31484 9658 31536 9664
rect 31496 9042 31524 9658
rect 31772 9382 31800 9998
rect 32508 9722 32536 10406
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 32692 9722 32720 9998
rect 33232 9920 33284 9926
rect 33232 9862 33284 9868
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31484 9036 31536 9042
rect 31484 8978 31536 8984
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 31220 5574 31248 6598
rect 31312 5642 31340 7686
rect 31772 6914 31800 9318
rect 32220 8968 32272 8974
rect 32220 8910 32272 8916
rect 32128 8424 32180 8430
rect 32128 8366 32180 8372
rect 32140 7886 32168 8366
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32128 7336 32180 7342
rect 32128 7278 32180 7284
rect 32140 7002 32168 7278
rect 32128 6996 32180 7002
rect 32128 6938 32180 6944
rect 31588 6886 31800 6914
rect 31484 6248 31536 6254
rect 31588 6236 31616 6886
rect 31852 6860 31904 6866
rect 31852 6802 31904 6808
rect 31668 6452 31720 6458
rect 31668 6394 31720 6400
rect 31536 6208 31616 6236
rect 31484 6190 31536 6196
rect 31496 5642 31524 6190
rect 31300 5636 31352 5642
rect 31300 5578 31352 5584
rect 31484 5636 31536 5642
rect 31484 5578 31536 5584
rect 31116 5568 31168 5574
rect 31208 5568 31260 5574
rect 31168 5528 31208 5556
rect 31116 5510 31168 5516
rect 31208 5510 31260 5516
rect 31128 5370 31156 5510
rect 31496 5386 31524 5578
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 31312 5358 31524 5386
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 31208 4752 31260 4758
rect 31206 4720 31208 4729
rect 31260 4720 31262 4729
rect 31206 4655 31262 4664
rect 31116 4480 31168 4486
rect 31116 4422 31168 4428
rect 30748 4004 30800 4010
rect 30748 3946 30800 3952
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30840 3392 30892 3398
rect 30840 3334 30892 3340
rect 30760 3074 30788 3334
rect 30852 3194 30880 3334
rect 31128 3194 31156 4422
rect 31312 4146 31340 5358
rect 31576 5228 31628 5234
rect 31576 5170 31628 5176
rect 31392 4616 31444 4622
rect 31392 4558 31444 4564
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31208 4072 31260 4078
rect 31208 4014 31260 4020
rect 31220 3618 31248 4014
rect 31404 3670 31432 4558
rect 31484 4548 31536 4554
rect 31484 4490 31536 4496
rect 31496 4078 31524 4490
rect 31484 4072 31536 4078
rect 31484 4014 31536 4020
rect 31392 3664 31444 3670
rect 31220 3590 31340 3618
rect 31392 3606 31444 3612
rect 31312 3466 31340 3590
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31220 3233 31248 3402
rect 31206 3224 31262 3233
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31116 3188 31168 3194
rect 31206 3159 31262 3168
rect 31484 3188 31536 3194
rect 31116 3130 31168 3136
rect 31484 3130 31536 3136
rect 30760 3058 30972 3074
rect 30760 3052 30984 3058
rect 30760 3046 30932 3052
rect 30932 2994 30984 3000
rect 31496 2990 31524 3130
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31588 2650 31616 5170
rect 31680 3738 31708 6394
rect 31760 6112 31812 6118
rect 31864 6089 31892 6802
rect 31944 6656 31996 6662
rect 31944 6598 31996 6604
rect 31956 6254 31984 6598
rect 31944 6248 31996 6254
rect 31944 6190 31996 6196
rect 31760 6054 31812 6060
rect 31850 6080 31906 6089
rect 31772 4554 31800 6054
rect 31850 6015 31906 6024
rect 31864 5710 31892 6015
rect 32232 5778 32260 8910
rect 33244 8566 33272 9862
rect 33324 9444 33376 9450
rect 33324 9386 33376 9392
rect 33232 8560 33284 8566
rect 33232 8502 33284 8508
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 33060 7274 33088 7822
rect 33336 7750 33364 9386
rect 33416 8492 33468 8498
rect 33416 8434 33468 8440
rect 33324 7744 33376 7750
rect 33324 7686 33376 7692
rect 33336 7410 33364 7686
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33324 7404 33376 7410
rect 33324 7346 33376 7352
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 32772 7200 32824 7206
rect 32772 7142 32824 7148
rect 32784 6798 32812 7142
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 32416 6390 32444 6598
rect 32404 6384 32456 6390
rect 32404 6326 32456 6332
rect 32770 6216 32826 6225
rect 32770 6151 32826 6160
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 32036 5296 32088 5302
rect 32036 5238 32088 5244
rect 32048 4758 32076 5238
rect 32036 4752 32088 4758
rect 32036 4694 32088 4700
rect 31760 4548 31812 4554
rect 31760 4490 31812 4496
rect 31944 4480 31996 4486
rect 31944 4422 31996 4428
rect 31956 4282 31984 4422
rect 31944 4276 31996 4282
rect 31944 4218 31996 4224
rect 32232 4146 32260 5714
rect 32680 5024 32732 5030
rect 32680 4966 32732 4972
rect 32692 4622 32720 4966
rect 32680 4616 32732 4622
rect 32680 4558 32732 4564
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 31852 4072 31904 4078
rect 31852 4014 31904 4020
rect 31668 3732 31720 3738
rect 31668 3674 31720 3680
rect 31864 3194 31892 4014
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31668 3052 31720 3058
rect 31668 2994 31720 3000
rect 31576 2644 31628 2650
rect 31576 2586 31628 2592
rect 30748 2508 30800 2514
rect 30748 2450 30800 2456
rect 29736 2440 29788 2446
rect 29656 2400 29736 2428
rect 29656 800 29684 2400
rect 29736 2382 29788 2388
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 29838 2204 30146 2213
rect 29838 2202 29844 2204
rect 29900 2202 29924 2204
rect 29980 2202 30004 2204
rect 30060 2202 30084 2204
rect 30140 2202 30146 2204
rect 29900 2150 29902 2202
rect 30082 2150 30084 2202
rect 29838 2148 29844 2150
rect 29900 2148 29924 2150
rect 29980 2148 30004 2150
rect 30060 2148 30084 2150
rect 30140 2148 30146 2150
rect 29838 2139 30146 2148
rect 30208 800 30236 2382
rect 30760 800 30788 2450
rect 31312 870 31432 898
rect 31312 800 31340 870
rect 23124 734 23428 762
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25226 0 25282 800
rect 25778 0 25834 800
rect 26330 0 26386 800
rect 26882 0 26938 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31404 762 31432 870
rect 31680 762 31708 2994
rect 31760 2848 31812 2854
rect 31760 2790 31812 2796
rect 31772 2514 31800 2790
rect 31760 2508 31812 2514
rect 31760 2450 31812 2456
rect 32048 2106 32076 3470
rect 32312 3188 32364 3194
rect 32312 3130 32364 3136
rect 32324 2961 32352 3130
rect 32784 2972 32812 6151
rect 32876 5914 32904 6734
rect 32956 6112 33008 6118
rect 32956 6054 33008 6060
rect 32968 5953 32996 6054
rect 32954 5944 33010 5953
rect 32864 5908 32916 5914
rect 32954 5879 32956 5888
rect 32864 5850 32916 5856
rect 33008 5879 33010 5888
rect 32956 5850 33008 5856
rect 33060 5234 33088 7210
rect 33152 7002 33180 7346
rect 33140 6996 33192 7002
rect 33140 6938 33192 6944
rect 33336 6390 33364 7346
rect 33324 6384 33376 6390
rect 33428 6361 33456 8434
rect 33520 8294 33548 9998
rect 33968 9920 34020 9926
rect 33968 9862 34020 9868
rect 33980 9722 34008 9862
rect 33968 9716 34020 9722
rect 33968 9658 34020 9664
rect 34164 9654 34192 11630
rect 34440 11234 34468 11630
rect 34520 11552 34572 11558
rect 34520 11494 34572 11500
rect 34348 11206 34468 11234
rect 34348 10470 34376 11206
rect 34532 11098 34560 11494
rect 34440 11070 34560 11098
rect 34624 11082 34652 12174
rect 34612 11076 34664 11082
rect 34440 11014 34468 11070
rect 34612 11018 34664 11024
rect 34428 11008 34480 11014
rect 34428 10950 34480 10956
rect 34624 10810 34652 11018
rect 34612 10804 34664 10810
rect 34612 10746 34664 10752
rect 34244 10464 34296 10470
rect 34244 10406 34296 10412
rect 34336 10464 34388 10470
rect 34336 10406 34388 10412
rect 34152 9648 34204 9654
rect 34152 9590 34204 9596
rect 34164 9518 34192 9590
rect 34152 9512 34204 9518
rect 34152 9454 34204 9460
rect 34256 8838 34284 10406
rect 34348 9518 34376 10406
rect 34428 9648 34480 9654
rect 34428 9590 34480 9596
rect 34336 9512 34388 9518
rect 34336 9454 34388 9460
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34256 8566 34284 8774
rect 34244 8560 34296 8566
rect 34244 8502 34296 8508
rect 33508 8288 33560 8294
rect 33508 8230 33560 8236
rect 33520 8090 33548 8230
rect 33508 8084 33560 8090
rect 33508 8026 33560 8032
rect 33784 8016 33836 8022
rect 33784 7958 33836 7964
rect 33600 7336 33652 7342
rect 33600 7278 33652 7284
rect 33612 7002 33640 7278
rect 33600 6996 33652 7002
rect 33600 6938 33652 6944
rect 33796 6866 33824 7958
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 33888 7546 33916 7822
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 34348 7410 34376 9454
rect 34440 8430 34468 9590
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34428 8424 34480 8430
rect 34428 8366 34480 8372
rect 34532 7478 34560 8774
rect 34704 7880 34756 7886
rect 34704 7822 34756 7828
rect 34716 7546 34744 7822
rect 34704 7540 34756 7546
rect 34704 7482 34756 7488
rect 34520 7472 34572 7478
rect 34520 7414 34572 7420
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 34428 6452 34480 6458
rect 34428 6394 34480 6400
rect 34060 6384 34112 6390
rect 33324 6326 33376 6332
rect 33414 6352 33470 6361
rect 34060 6326 34112 6332
rect 33414 6287 33470 6296
rect 33508 6316 33560 6322
rect 33508 6258 33560 6264
rect 33048 5228 33100 5234
rect 33048 5170 33100 5176
rect 33232 4820 33284 4826
rect 33232 4762 33284 4768
rect 33244 4146 33272 4762
rect 33322 4584 33378 4593
rect 33322 4519 33324 4528
rect 33376 4519 33378 4528
rect 33324 4490 33376 4496
rect 33416 4480 33468 4486
rect 33416 4422 33468 4428
rect 33428 4185 33456 4422
rect 33414 4176 33470 4185
rect 33232 4140 33284 4146
rect 33414 4111 33470 4120
rect 33232 4082 33284 4088
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32968 3913 32996 4014
rect 33140 3936 33192 3942
rect 32954 3904 33010 3913
rect 33140 3878 33192 3884
rect 32954 3839 33010 3848
rect 33152 2990 33180 3878
rect 33520 3398 33548 6258
rect 33600 5704 33652 5710
rect 33600 5646 33652 5652
rect 33612 4826 33640 5646
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 34072 4690 34100 6326
rect 34152 5568 34204 5574
rect 34152 5510 34204 5516
rect 34164 5302 34192 5510
rect 34152 5296 34204 5302
rect 34152 5238 34204 5244
rect 34152 5024 34204 5030
rect 34152 4966 34204 4972
rect 34336 5024 34388 5030
rect 34336 4966 34388 4972
rect 34060 4684 34112 4690
rect 34060 4626 34112 4632
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 33600 3936 33652 3942
rect 33600 3878 33652 3884
rect 33612 3738 33640 3878
rect 33980 3738 34008 4422
rect 34072 4282 34100 4626
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 33600 3732 33652 3738
rect 33600 3674 33652 3680
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 34058 3224 34114 3233
rect 34058 3159 34114 3168
rect 34072 3058 34100 3159
rect 34060 3052 34112 3058
rect 34060 2994 34112 3000
rect 32864 2984 32916 2990
rect 32310 2952 32366 2961
rect 32784 2944 32864 2972
rect 32864 2926 32916 2932
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 32310 2887 32366 2896
rect 32956 2916 33008 2922
rect 32956 2858 33008 2864
rect 33508 2916 33560 2922
rect 33508 2858 33560 2864
rect 32680 2508 32732 2514
rect 32680 2450 32732 2456
rect 32036 2100 32088 2106
rect 32036 2042 32088 2048
rect 31852 1556 31904 1562
rect 31852 1498 31904 1504
rect 31864 800 31892 1498
rect 32416 870 32536 898
rect 32416 800 32444 870
rect 31404 734 31708 762
rect 31850 0 31906 800
rect 32402 0 32458 800
rect 32508 762 32536 870
rect 32692 762 32720 2450
rect 32968 800 32996 2858
rect 33520 800 33548 2858
rect 34164 2446 34192 4966
rect 34348 3602 34376 4966
rect 34440 4690 34468 6394
rect 34624 5914 34652 7142
rect 34716 6662 34744 7346
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34704 6112 34756 6118
rect 34704 6054 34756 6060
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34716 5817 34744 6054
rect 34702 5808 34758 5817
rect 34702 5743 34758 5752
rect 34716 5710 34744 5743
rect 34704 5704 34756 5710
rect 34704 5646 34756 5652
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 34624 4758 34652 5578
rect 34808 5234 34836 12406
rect 34900 10810 34928 17070
rect 34980 16040 35032 16046
rect 34980 15982 35032 15988
rect 34992 14822 35020 15982
rect 35268 15366 35296 17206
rect 35452 17134 35480 18022
rect 35440 17128 35492 17134
rect 35440 17070 35492 17076
rect 35452 15570 35480 17070
rect 35440 15564 35492 15570
rect 35440 15506 35492 15512
rect 35072 15360 35124 15366
rect 35072 15302 35124 15308
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 34980 14816 35032 14822
rect 34980 14758 35032 14764
rect 34992 14074 35020 14758
rect 34980 14068 35032 14074
rect 34980 14010 35032 14016
rect 35084 13394 35112 15302
rect 35256 14408 35308 14414
rect 35256 14350 35308 14356
rect 35268 13870 35296 14350
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 35256 13864 35308 13870
rect 35256 13806 35308 13812
rect 35072 13388 35124 13394
rect 35072 13330 35124 13336
rect 35084 12918 35112 13330
rect 35360 12986 35388 14214
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 35072 12912 35124 12918
rect 35072 12854 35124 12860
rect 35084 12434 35112 12854
rect 35164 12708 35216 12714
rect 35164 12650 35216 12656
rect 34992 12406 35112 12434
rect 34992 11218 35020 12406
rect 35072 11620 35124 11626
rect 35072 11562 35124 11568
rect 35084 11286 35112 11562
rect 35072 11280 35124 11286
rect 35072 11222 35124 11228
rect 34980 11212 35032 11218
rect 34980 11154 35032 11160
rect 34888 10804 34940 10810
rect 34888 10746 34940 10752
rect 34992 9926 35020 11154
rect 35072 11144 35124 11150
rect 35072 11086 35124 11092
rect 35084 10810 35112 11086
rect 35072 10804 35124 10810
rect 35072 10746 35124 10752
rect 34980 9920 35032 9926
rect 34980 9862 35032 9868
rect 34888 8628 34940 8634
rect 34888 8570 34940 8576
rect 34900 7954 34928 8570
rect 34992 7954 35020 9862
rect 34888 7948 34940 7954
rect 34888 7890 34940 7896
rect 34980 7948 35032 7954
rect 34980 7890 35032 7896
rect 34888 6316 34940 6322
rect 34888 6258 34940 6264
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 34704 5160 34756 5166
rect 34704 5102 34756 5108
rect 34716 4826 34744 5102
rect 34900 4865 34928 6258
rect 34992 6254 35020 7890
rect 35072 6384 35124 6390
rect 35072 6326 35124 6332
rect 34980 6248 35032 6254
rect 34980 6190 35032 6196
rect 34886 4856 34942 4865
rect 34704 4820 34756 4826
rect 34886 4791 34942 4800
rect 34704 4762 34756 4768
rect 34612 4752 34664 4758
rect 34612 4694 34664 4700
rect 34428 4684 34480 4690
rect 34428 4626 34480 4632
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34336 3596 34388 3602
rect 34336 3538 34388 3544
rect 34244 3460 34296 3466
rect 34244 3402 34296 3408
rect 34256 3194 34284 3402
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34440 2854 34468 4014
rect 34716 3516 34744 4762
rect 35084 4078 35112 6326
rect 35176 6118 35204 12650
rect 35544 12434 35572 19230
rect 36188 18970 36216 19314
rect 36176 18964 36228 18970
rect 36176 18906 36228 18912
rect 36280 18834 36308 19382
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 36268 18828 36320 18834
rect 36268 18770 36320 18776
rect 35912 18086 35940 18770
rect 35900 18080 35952 18086
rect 35900 18022 35952 18028
rect 35624 17128 35676 17134
rect 35624 17070 35676 17076
rect 35636 16454 35664 17070
rect 35992 16992 36044 16998
rect 35992 16934 36044 16940
rect 36004 16590 36032 16934
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 35624 16448 35676 16454
rect 35624 16390 35676 16396
rect 36556 16250 36584 19654
rect 36740 19514 36768 20742
rect 37476 20398 37504 20742
rect 37568 20602 37596 20878
rect 37556 20596 37608 20602
rect 37556 20538 37608 20544
rect 37844 20534 37872 22066
rect 38304 22030 38332 22578
rect 38568 22432 38620 22438
rect 38568 22374 38620 22380
rect 38660 22432 38712 22438
rect 38660 22374 38712 22380
rect 38580 22166 38608 22374
rect 38568 22160 38620 22166
rect 38568 22102 38620 22108
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38384 21344 38436 21350
rect 38384 21286 38436 21292
rect 38396 21146 38424 21286
rect 38384 21140 38436 21146
rect 38384 21082 38436 21088
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 38108 20800 38160 20806
rect 38108 20742 38160 20748
rect 37832 20528 37884 20534
rect 37832 20470 37884 20476
rect 37464 20392 37516 20398
rect 37464 20334 37516 20340
rect 36912 20256 36964 20262
rect 36912 20198 36964 20204
rect 36924 19854 36952 20198
rect 37060 20156 37368 20165
rect 37060 20154 37066 20156
rect 37122 20154 37146 20156
rect 37202 20154 37226 20156
rect 37282 20154 37306 20156
rect 37362 20154 37368 20156
rect 37122 20102 37124 20154
rect 37304 20102 37306 20154
rect 37060 20100 37066 20102
rect 37122 20100 37146 20102
rect 37202 20100 37226 20102
rect 37282 20100 37306 20102
rect 37362 20100 37368 20102
rect 37060 20091 37368 20100
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 36924 19514 36952 19790
rect 37476 19718 37504 20334
rect 38120 19786 38148 20742
rect 38304 20398 38332 20878
rect 38672 20398 38700 22374
rect 38752 21888 38804 21894
rect 38752 21830 38804 21836
rect 38764 21554 38792 21830
rect 38856 21690 38884 23054
rect 39396 22976 39448 22982
rect 39396 22918 39448 22924
rect 40040 22976 40092 22982
rect 40040 22918 40092 22924
rect 39408 22642 39436 22918
rect 40052 22710 40080 22918
rect 44282 22876 44590 22885
rect 44282 22874 44288 22876
rect 44344 22874 44368 22876
rect 44424 22874 44448 22876
rect 44504 22874 44528 22876
rect 44584 22874 44590 22876
rect 44344 22822 44346 22874
rect 44526 22822 44528 22874
rect 44282 22820 44288 22822
rect 44344 22820 44368 22822
rect 44424 22820 44448 22822
rect 44504 22820 44528 22822
rect 44584 22820 44590 22822
rect 44282 22811 44590 22820
rect 40040 22704 40092 22710
rect 40040 22646 40092 22652
rect 47584 22704 47636 22710
rect 47584 22646 47636 22652
rect 39396 22636 39448 22642
rect 39396 22578 39448 22584
rect 40052 22094 40080 22646
rect 40408 22432 40460 22438
rect 40408 22374 40460 22380
rect 39960 22066 40080 22094
rect 39212 21888 39264 21894
rect 39212 21830 39264 21836
rect 39396 21888 39448 21894
rect 39396 21830 39448 21836
rect 38844 21684 38896 21690
rect 38844 21626 38896 21632
rect 39224 21554 39252 21830
rect 39408 21690 39436 21830
rect 39396 21684 39448 21690
rect 39396 21626 39448 21632
rect 38752 21548 38804 21554
rect 38752 21490 38804 21496
rect 38936 21548 38988 21554
rect 38936 21490 38988 21496
rect 39212 21548 39264 21554
rect 39212 21490 39264 21496
rect 38844 20800 38896 20806
rect 38844 20742 38896 20748
rect 38856 20602 38884 20742
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38948 20482 38976 21490
rect 39304 21480 39356 21486
rect 39304 21422 39356 21428
rect 39028 21412 39080 21418
rect 39028 21354 39080 21360
rect 38856 20454 38976 20482
rect 38200 20392 38252 20398
rect 38200 20334 38252 20340
rect 38292 20392 38344 20398
rect 38292 20334 38344 20340
rect 38568 20392 38620 20398
rect 38568 20334 38620 20340
rect 38660 20392 38712 20398
rect 38660 20334 38712 20340
rect 38212 19922 38240 20334
rect 38304 20058 38332 20334
rect 38580 20210 38608 20334
rect 38856 20262 38884 20454
rect 39040 20330 39068 21354
rect 39212 21344 39264 21350
rect 39212 21286 39264 21292
rect 39224 20806 39252 21286
rect 39212 20800 39264 20806
rect 39212 20742 39264 20748
rect 39028 20324 39080 20330
rect 39028 20266 39080 20272
rect 38844 20256 38896 20262
rect 38580 20182 38700 20210
rect 38844 20198 38896 20204
rect 38292 20052 38344 20058
rect 38292 19994 38344 20000
rect 38200 19916 38252 19922
rect 38200 19858 38252 19864
rect 38108 19780 38160 19786
rect 38108 19722 38160 19728
rect 37464 19712 37516 19718
rect 37464 19654 37516 19660
rect 36728 19508 36780 19514
rect 36728 19450 36780 19456
rect 36912 19508 36964 19514
rect 36912 19450 36964 19456
rect 36924 18834 36952 19450
rect 38672 19378 38700 20182
rect 38856 19718 38884 20198
rect 39028 19916 39080 19922
rect 39028 19858 39080 19864
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38660 19372 38712 19378
rect 38660 19314 38712 19320
rect 38292 19168 38344 19174
rect 38292 19110 38344 19116
rect 38384 19168 38436 19174
rect 38384 19110 38436 19116
rect 37060 19068 37368 19077
rect 37060 19066 37066 19068
rect 37122 19066 37146 19068
rect 37202 19066 37226 19068
rect 37282 19066 37306 19068
rect 37362 19066 37368 19068
rect 37122 19014 37124 19066
rect 37304 19014 37306 19066
rect 37060 19012 37066 19014
rect 37122 19012 37146 19014
rect 37202 19012 37226 19014
rect 37282 19012 37306 19014
rect 37362 19012 37368 19014
rect 37060 19003 37368 19012
rect 38304 18834 38332 19110
rect 36912 18828 36964 18834
rect 36912 18770 36964 18776
rect 38292 18828 38344 18834
rect 38292 18770 38344 18776
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36728 17536 36780 17542
rect 36728 17478 36780 17484
rect 36648 16658 36676 17478
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36648 16250 36676 16594
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 36636 16244 36688 16250
rect 36636 16186 36688 16192
rect 36740 16114 36768 17478
rect 36728 16108 36780 16114
rect 36728 16050 36780 16056
rect 36360 15904 36412 15910
rect 36360 15846 36412 15852
rect 36372 15366 36400 15846
rect 36728 15564 36780 15570
rect 36728 15506 36780 15512
rect 36360 15360 36412 15366
rect 36360 15302 36412 15308
rect 36268 14816 36320 14822
rect 36268 14758 36320 14764
rect 35624 14476 35676 14482
rect 35624 14418 35676 14424
rect 35636 13394 35664 14418
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 36096 13394 36124 14010
rect 36280 13938 36308 14758
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36176 13728 36228 13734
rect 36176 13670 36228 13676
rect 35624 13388 35676 13394
rect 35624 13330 35676 13336
rect 35716 13388 35768 13394
rect 36084 13388 36136 13394
rect 35768 13348 35848 13376
rect 35716 13330 35768 13336
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35452 12406 35572 12434
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 35360 11898 35388 12038
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 35452 11558 35480 12406
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 35256 10668 35308 10674
rect 35256 10610 35308 10616
rect 35164 6112 35216 6118
rect 35164 6054 35216 6060
rect 35072 4072 35124 4078
rect 35072 4014 35124 4020
rect 35162 4040 35218 4049
rect 35162 3975 35218 3984
rect 35176 3738 35204 3975
rect 35268 3942 35296 10610
rect 35452 9586 35480 11494
rect 35624 11144 35676 11150
rect 35624 11086 35676 11092
rect 35636 11014 35664 11086
rect 35728 11014 35756 12786
rect 35820 12306 35848 13348
rect 36084 13330 36136 13336
rect 35808 12300 35860 12306
rect 35808 12242 35860 12248
rect 35992 12232 36044 12238
rect 35992 12174 36044 12180
rect 36004 11898 36032 12174
rect 35992 11892 36044 11898
rect 35992 11834 36044 11840
rect 36096 11218 36124 13330
rect 36188 13190 36216 13670
rect 36176 13184 36228 13190
rect 36176 13126 36228 13132
rect 36372 12238 36400 15302
rect 36544 14952 36596 14958
rect 36544 14894 36596 14900
rect 36556 14074 36584 14894
rect 36636 14408 36688 14414
rect 36636 14350 36688 14356
rect 36544 14068 36596 14074
rect 36544 14010 36596 14016
rect 36648 13734 36676 14350
rect 36636 13728 36688 13734
rect 36636 13670 36688 13676
rect 36740 13394 36768 15506
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 36544 13184 36596 13190
rect 36544 13126 36596 13132
rect 36360 12232 36412 12238
rect 36360 12174 36412 12180
rect 36360 11756 36412 11762
rect 36360 11698 36412 11704
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 35900 11212 35952 11218
rect 35900 11154 35952 11160
rect 36084 11212 36136 11218
rect 36084 11154 36136 11160
rect 35624 11008 35676 11014
rect 35624 10950 35676 10956
rect 35716 11008 35768 11014
rect 35716 10950 35768 10956
rect 35912 10266 35940 11154
rect 36280 10266 36308 11290
rect 36372 10470 36400 11698
rect 36556 11218 36584 13126
rect 36740 12714 36768 13330
rect 36820 13320 36872 13326
rect 36820 13262 36872 13268
rect 36728 12708 36780 12714
rect 36728 12650 36780 12656
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36648 10674 36676 12038
rect 36636 10668 36688 10674
rect 36636 10610 36688 10616
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 35900 10260 35952 10266
rect 35900 10202 35952 10208
rect 36268 10260 36320 10266
rect 36268 10202 36320 10208
rect 35532 9920 35584 9926
rect 35532 9862 35584 9868
rect 35440 9580 35492 9586
rect 35440 9522 35492 9528
rect 35544 9450 35572 9862
rect 35532 9444 35584 9450
rect 35532 9386 35584 9392
rect 35348 8288 35400 8294
rect 35348 8230 35400 8236
rect 35360 7206 35388 8230
rect 35716 8084 35768 8090
rect 35716 8026 35768 8032
rect 35728 7954 35756 8026
rect 35912 7954 35940 10202
rect 35992 9512 36044 9518
rect 35992 9454 36044 9460
rect 35716 7948 35768 7954
rect 35716 7890 35768 7896
rect 35900 7948 35952 7954
rect 35900 7890 35952 7896
rect 36004 7546 36032 9454
rect 36084 8968 36136 8974
rect 36084 8910 36136 8916
rect 35992 7540 36044 7546
rect 35992 7482 36044 7488
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 35348 7200 35400 7206
rect 35348 7142 35400 7148
rect 35360 7002 35388 7142
rect 35912 7002 35940 7346
rect 35348 6996 35400 7002
rect 35348 6938 35400 6944
rect 35900 6996 35952 7002
rect 35900 6938 35952 6944
rect 36096 6934 36124 8910
rect 36268 7948 36320 7954
rect 36268 7890 36320 7896
rect 36084 6928 36136 6934
rect 36084 6870 36136 6876
rect 35808 6724 35860 6730
rect 35808 6666 35860 6672
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35532 6112 35584 6118
rect 35532 6054 35584 6060
rect 35544 5642 35572 6054
rect 35532 5636 35584 5642
rect 35532 5578 35584 5584
rect 35440 5228 35492 5234
rect 35492 5188 35572 5216
rect 35440 5170 35492 5176
rect 35544 4078 35572 5188
rect 35636 5098 35664 6190
rect 35820 5914 35848 6666
rect 35808 5908 35860 5914
rect 35808 5850 35860 5856
rect 36280 5574 36308 7890
rect 36372 6798 36400 10406
rect 36544 9376 36596 9382
rect 36544 9318 36596 9324
rect 36556 8498 36584 9318
rect 36740 8922 36768 12650
rect 36832 12374 36860 13262
rect 36924 12434 36952 18022
rect 37060 17980 37368 17989
rect 37060 17978 37066 17980
rect 37122 17978 37146 17980
rect 37202 17978 37226 17980
rect 37282 17978 37306 17980
rect 37362 17978 37368 17980
rect 37122 17926 37124 17978
rect 37304 17926 37306 17978
rect 37060 17924 37066 17926
rect 37122 17924 37146 17926
rect 37202 17924 37226 17926
rect 37282 17924 37306 17926
rect 37362 17924 37368 17926
rect 37060 17915 37368 17924
rect 38304 17882 38332 18770
rect 38292 17876 38344 17882
rect 38292 17818 38344 17824
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 38120 17202 38148 17614
rect 38200 17536 38252 17542
rect 38200 17478 38252 17484
rect 38108 17196 38160 17202
rect 38108 17138 38160 17144
rect 37060 16892 37368 16901
rect 37060 16890 37066 16892
rect 37122 16890 37146 16892
rect 37202 16890 37226 16892
rect 37282 16890 37306 16892
rect 37362 16890 37368 16892
rect 37122 16838 37124 16890
rect 37304 16838 37306 16890
rect 37060 16836 37066 16838
rect 37122 16836 37146 16838
rect 37202 16836 37226 16838
rect 37282 16836 37306 16838
rect 37362 16836 37368 16838
rect 37060 16827 37368 16836
rect 38212 16658 38240 17478
rect 38200 16652 38252 16658
rect 38200 16594 38252 16600
rect 38200 16516 38252 16522
rect 38200 16458 38252 16464
rect 38108 16448 38160 16454
rect 38108 16390 38160 16396
rect 37060 15804 37368 15813
rect 37060 15802 37066 15804
rect 37122 15802 37146 15804
rect 37202 15802 37226 15804
rect 37282 15802 37306 15804
rect 37362 15802 37368 15804
rect 37122 15750 37124 15802
rect 37304 15750 37306 15802
rect 37060 15748 37066 15750
rect 37122 15748 37146 15750
rect 37202 15748 37226 15750
rect 37282 15748 37306 15750
rect 37362 15748 37368 15750
rect 37060 15739 37368 15748
rect 38120 15706 38148 16390
rect 38212 15706 38240 16458
rect 38108 15700 38160 15706
rect 38108 15642 38160 15648
rect 38200 15700 38252 15706
rect 38200 15642 38252 15648
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 37464 14816 37516 14822
rect 37464 14758 37516 14764
rect 37060 14716 37368 14725
rect 37060 14714 37066 14716
rect 37122 14714 37146 14716
rect 37202 14714 37226 14716
rect 37282 14714 37306 14716
rect 37362 14714 37368 14716
rect 37122 14662 37124 14714
rect 37304 14662 37306 14714
rect 37060 14660 37066 14662
rect 37122 14660 37146 14662
rect 37202 14660 37226 14662
rect 37282 14660 37306 14662
rect 37362 14660 37368 14662
rect 37060 14651 37368 14660
rect 37476 14006 37504 14758
rect 37556 14272 37608 14278
rect 37556 14214 37608 14220
rect 37464 14000 37516 14006
rect 37464 13942 37516 13948
rect 37060 13628 37368 13637
rect 37060 13626 37066 13628
rect 37122 13626 37146 13628
rect 37202 13626 37226 13628
rect 37282 13626 37306 13628
rect 37362 13626 37368 13628
rect 37122 13574 37124 13626
rect 37304 13574 37306 13626
rect 37060 13572 37066 13574
rect 37122 13572 37146 13574
rect 37202 13572 37226 13574
rect 37282 13572 37306 13574
rect 37362 13572 37368 13574
rect 37060 13563 37368 13572
rect 37568 13530 37596 14214
rect 37648 13932 37700 13938
rect 37648 13874 37700 13880
rect 37556 13524 37608 13530
rect 37556 13466 37608 13472
rect 37004 13184 37056 13190
rect 37004 13126 37056 13132
rect 37016 12986 37044 13126
rect 37004 12980 37056 12986
rect 37004 12922 37056 12928
rect 37568 12850 37596 13466
rect 37660 13394 37688 13874
rect 37844 13870 37872 15438
rect 38396 15094 38424 19110
rect 38660 18896 38712 18902
rect 38660 18838 38712 18844
rect 38568 18692 38620 18698
rect 38568 18634 38620 18640
rect 38476 18624 38528 18630
rect 38476 18566 38528 18572
rect 38488 18426 38516 18566
rect 38580 18426 38608 18634
rect 38476 18420 38528 18426
rect 38476 18362 38528 18368
rect 38568 18420 38620 18426
rect 38568 18362 38620 18368
rect 38672 18290 38700 18838
rect 38856 18630 38884 19654
rect 39040 19174 39068 19858
rect 39224 19825 39252 20742
rect 39316 20466 39344 21422
rect 39960 21146 39988 22066
rect 40420 21690 40448 22374
rect 40776 22160 40828 22166
rect 40776 22102 40828 22108
rect 40408 21684 40460 21690
rect 40408 21626 40460 21632
rect 39488 21140 39540 21146
rect 39488 21082 39540 21088
rect 39948 21140 40000 21146
rect 39948 21082 40000 21088
rect 39304 20460 39356 20466
rect 39304 20402 39356 20408
rect 39500 20448 39528 21082
rect 39580 20460 39632 20466
rect 39500 20420 39580 20448
rect 39210 19816 39266 19825
rect 39210 19751 39266 19760
rect 39304 19712 39356 19718
rect 39304 19654 39356 19660
rect 39316 19514 39344 19654
rect 39304 19508 39356 19514
rect 39304 19450 39356 19456
rect 39028 19168 39080 19174
rect 39028 19110 39080 19116
rect 38844 18624 38896 18630
rect 38844 18566 38896 18572
rect 38936 18624 38988 18630
rect 38936 18566 38988 18572
rect 38660 18284 38712 18290
rect 38660 18226 38712 18232
rect 38672 17134 38700 18226
rect 38752 17536 38804 17542
rect 38752 17478 38804 17484
rect 38660 17128 38712 17134
rect 38660 17070 38712 17076
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38476 16448 38528 16454
rect 38476 16390 38528 16396
rect 38488 15706 38516 16390
rect 38672 16250 38700 16934
rect 38660 16244 38712 16250
rect 38660 16186 38712 16192
rect 38476 15700 38528 15706
rect 38476 15642 38528 15648
rect 38672 15502 38700 16186
rect 38764 16182 38792 17478
rect 38856 16454 38884 18566
rect 38948 18426 38976 18566
rect 38936 18420 38988 18426
rect 38936 18362 38988 18368
rect 38936 17672 38988 17678
rect 38936 17614 38988 17620
rect 38948 16794 38976 17614
rect 39500 17134 39528 20420
rect 39580 20402 39632 20408
rect 39960 20398 39988 21082
rect 40788 20602 40816 22102
rect 47308 21888 47360 21894
rect 47308 21830 47360 21836
rect 44282 21788 44590 21797
rect 44282 21786 44288 21788
rect 44344 21786 44368 21788
rect 44424 21786 44448 21788
rect 44504 21786 44528 21788
rect 44584 21786 44590 21788
rect 44344 21734 44346 21786
rect 44526 21734 44528 21786
rect 44282 21732 44288 21734
rect 44344 21732 44368 21734
rect 44424 21732 44448 21734
rect 44504 21732 44528 21734
rect 44584 21732 44590 21734
rect 44282 21723 44590 21732
rect 42708 21480 42760 21486
rect 42708 21422 42760 21428
rect 46664 21480 46716 21486
rect 46664 21422 46716 21428
rect 42248 21412 42300 21418
rect 42248 21354 42300 21360
rect 41880 21344 41932 21350
rect 41880 21286 41932 21292
rect 41420 21140 41472 21146
rect 41420 21082 41472 21088
rect 40776 20596 40828 20602
rect 40776 20538 40828 20544
rect 39948 20392 40000 20398
rect 39948 20334 40000 20340
rect 39960 19786 39988 20334
rect 40788 20262 40816 20538
rect 41432 20534 41460 21082
rect 41892 20942 41920 21286
rect 42260 21146 42288 21354
rect 42248 21140 42300 21146
rect 42248 21082 42300 21088
rect 41788 20936 41840 20942
rect 41788 20878 41840 20884
rect 41880 20936 41932 20942
rect 41880 20878 41932 20884
rect 41800 20602 41828 20878
rect 41788 20596 41840 20602
rect 41788 20538 41840 20544
rect 41420 20528 41472 20534
rect 41420 20470 41472 20476
rect 40224 20256 40276 20262
rect 40224 20198 40276 20204
rect 40776 20256 40828 20262
rect 40776 20198 40828 20204
rect 40040 20052 40092 20058
rect 40040 19994 40092 20000
rect 39948 19780 40000 19786
rect 39948 19722 40000 19728
rect 39580 19712 39632 19718
rect 39580 19654 39632 19660
rect 39592 19310 39620 19654
rect 39960 19378 39988 19722
rect 39948 19372 40000 19378
rect 39948 19314 40000 19320
rect 39580 19304 39632 19310
rect 39580 19246 39632 19252
rect 40052 18834 40080 19994
rect 40040 18828 40092 18834
rect 40040 18770 40092 18776
rect 39948 18080 40000 18086
rect 39948 18022 40000 18028
rect 39028 17128 39080 17134
rect 39028 17070 39080 17076
rect 39488 17128 39540 17134
rect 39488 17070 39540 17076
rect 38936 16788 38988 16794
rect 38936 16730 38988 16736
rect 39040 16590 39068 17070
rect 39500 16776 39528 17070
rect 39764 16992 39816 16998
rect 39764 16934 39816 16940
rect 39500 16748 39620 16776
rect 39488 16652 39540 16658
rect 39488 16594 39540 16600
rect 39028 16584 39080 16590
rect 39028 16526 39080 16532
rect 38844 16448 38896 16454
rect 38844 16390 38896 16396
rect 38752 16176 38804 16182
rect 38752 16118 38804 16124
rect 39040 15706 39068 16526
rect 39304 16448 39356 16454
rect 39304 16390 39356 16396
rect 39396 16448 39448 16454
rect 39396 16390 39448 16396
rect 39028 15700 39080 15706
rect 39028 15642 39080 15648
rect 38660 15496 38712 15502
rect 38660 15438 38712 15444
rect 38200 15088 38252 15094
rect 38200 15030 38252 15036
rect 38384 15088 38436 15094
rect 38384 15030 38436 15036
rect 38108 14340 38160 14346
rect 38108 14282 38160 14288
rect 38016 14272 38068 14278
rect 38016 14214 38068 14220
rect 38028 14074 38056 14214
rect 38016 14068 38068 14074
rect 38016 14010 38068 14016
rect 37832 13864 37884 13870
rect 37832 13806 37884 13812
rect 38120 13530 38148 14282
rect 38108 13524 38160 13530
rect 38108 13466 38160 13472
rect 37648 13388 37700 13394
rect 37648 13330 37700 13336
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37060 12540 37368 12549
rect 37060 12538 37066 12540
rect 37122 12538 37146 12540
rect 37202 12538 37226 12540
rect 37282 12538 37306 12540
rect 37362 12538 37368 12540
rect 37122 12486 37124 12538
rect 37304 12486 37306 12538
rect 37060 12484 37066 12486
rect 37122 12484 37146 12486
rect 37202 12484 37226 12486
rect 37282 12484 37306 12486
rect 37362 12484 37368 12486
rect 37060 12475 37368 12484
rect 36924 12406 37044 12434
rect 36820 12368 36872 12374
rect 36820 12310 36872 12316
rect 36832 11830 36860 12310
rect 36820 11824 36872 11830
rect 36820 11766 36872 11772
rect 36912 11688 36964 11694
rect 36912 11630 36964 11636
rect 36820 11552 36872 11558
rect 36820 11494 36872 11500
rect 36832 10690 36860 11494
rect 36924 10810 36952 11630
rect 37016 11558 37044 12406
rect 37464 12232 37516 12238
rect 37464 12174 37516 12180
rect 37004 11552 37056 11558
rect 37004 11494 37056 11500
rect 37060 11452 37368 11461
rect 37060 11450 37066 11452
rect 37122 11450 37146 11452
rect 37202 11450 37226 11452
rect 37282 11450 37306 11452
rect 37362 11450 37368 11452
rect 37122 11398 37124 11450
rect 37304 11398 37306 11450
rect 37060 11396 37066 11398
rect 37122 11396 37146 11398
rect 37202 11396 37226 11398
rect 37282 11396 37306 11398
rect 37362 11396 37368 11398
rect 37060 11387 37368 11396
rect 37476 11354 37504 12174
rect 37464 11348 37516 11354
rect 37464 11290 37516 11296
rect 37556 11280 37608 11286
rect 37556 11222 37608 11228
rect 37464 11144 37516 11150
rect 37464 11086 37516 11092
rect 37476 10810 37504 11086
rect 36912 10804 36964 10810
rect 36912 10746 36964 10752
rect 37464 10804 37516 10810
rect 37464 10746 37516 10752
rect 36832 10662 36952 10690
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 36832 8974 36860 9318
rect 36648 8894 36768 8922
rect 36820 8968 36872 8974
rect 36820 8910 36872 8916
rect 36924 8906 36952 10662
rect 37060 10364 37368 10373
rect 37060 10362 37066 10364
rect 37122 10362 37146 10364
rect 37202 10362 37226 10364
rect 37282 10362 37306 10364
rect 37362 10362 37368 10364
rect 37122 10310 37124 10362
rect 37304 10310 37306 10362
rect 37060 10308 37066 10310
rect 37122 10308 37146 10310
rect 37202 10308 37226 10310
rect 37282 10308 37306 10310
rect 37362 10308 37368 10310
rect 37060 10299 37368 10308
rect 37464 9920 37516 9926
rect 37464 9862 37516 9868
rect 37060 9276 37368 9285
rect 37060 9274 37066 9276
rect 37122 9274 37146 9276
rect 37202 9274 37226 9276
rect 37282 9274 37306 9276
rect 37362 9274 37368 9276
rect 37122 9222 37124 9274
rect 37304 9222 37306 9274
rect 37060 9220 37066 9222
rect 37122 9220 37146 9222
rect 37202 9220 37226 9222
rect 37282 9220 37306 9222
rect 37362 9220 37368 9222
rect 37060 9211 37368 9220
rect 37476 8906 37504 9862
rect 36912 8900 36964 8906
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36648 7834 36676 8894
rect 36912 8842 36964 8848
rect 37464 8900 37516 8906
rect 37464 8842 37516 8848
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 36740 8634 36768 8774
rect 36728 8628 36780 8634
rect 36728 8570 36780 8576
rect 36820 8288 36872 8294
rect 36820 8230 36872 8236
rect 36832 7954 36860 8230
rect 36924 7954 36952 8842
rect 37060 8188 37368 8197
rect 37060 8186 37066 8188
rect 37122 8186 37146 8188
rect 37202 8186 37226 8188
rect 37282 8186 37306 8188
rect 37362 8186 37368 8188
rect 37122 8134 37124 8186
rect 37304 8134 37306 8186
rect 37060 8132 37066 8134
rect 37122 8132 37146 8134
rect 37202 8132 37226 8134
rect 37282 8132 37306 8134
rect 37362 8132 37368 8134
rect 37060 8123 37368 8132
rect 36820 7948 36872 7954
rect 36820 7890 36872 7896
rect 36912 7948 36964 7954
rect 36912 7890 36964 7896
rect 36648 7806 36768 7834
rect 36452 7744 36504 7750
rect 36452 7686 36504 7692
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36636 7744 36688 7750
rect 36636 7686 36688 7692
rect 36464 7546 36492 7686
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 36268 5568 36320 5574
rect 36268 5510 36320 5516
rect 36280 5234 36308 5510
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 35624 5092 35676 5098
rect 35624 5034 35676 5040
rect 36004 4826 36032 5170
rect 36452 5160 36504 5166
rect 36452 5102 36504 5108
rect 35992 4820 36044 4826
rect 35992 4762 36044 4768
rect 35808 4616 35860 4622
rect 35808 4558 35860 4564
rect 35820 4162 35848 4558
rect 35900 4548 35952 4554
rect 35900 4490 35952 4496
rect 35912 4282 35940 4490
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 35820 4134 35940 4162
rect 36004 4146 36032 4762
rect 36464 4758 36492 5102
rect 36452 4752 36504 4758
rect 36452 4694 36504 4700
rect 36556 4622 36584 7686
rect 36648 6866 36676 7686
rect 36740 7206 36768 7806
rect 36728 7200 36780 7206
rect 36728 7142 36780 7148
rect 36636 6860 36688 6866
rect 36636 6802 36688 6808
rect 36740 6202 36768 7142
rect 36924 6934 36952 7890
rect 37096 7744 37148 7750
rect 37096 7686 37148 7692
rect 37108 7546 37136 7686
rect 37096 7540 37148 7546
rect 37096 7482 37148 7488
rect 37188 7336 37240 7342
rect 37476 7290 37504 8842
rect 37240 7284 37504 7290
rect 37188 7278 37504 7284
rect 37200 7262 37504 7278
rect 37060 7100 37368 7109
rect 37060 7098 37066 7100
rect 37122 7098 37146 7100
rect 37202 7098 37226 7100
rect 37282 7098 37306 7100
rect 37362 7098 37368 7100
rect 37122 7046 37124 7098
rect 37304 7046 37306 7098
rect 37060 7044 37066 7046
rect 37122 7044 37146 7046
rect 37202 7044 37226 7046
rect 37282 7044 37306 7046
rect 37362 7044 37368 7046
rect 37060 7035 37368 7044
rect 36912 6928 36964 6934
rect 37476 6905 37504 7262
rect 36912 6870 36964 6876
rect 37462 6896 37518 6905
rect 37462 6831 37518 6840
rect 37476 6798 37504 6831
rect 37464 6792 37516 6798
rect 37464 6734 37516 6740
rect 36648 6174 36768 6202
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 36084 4480 36136 4486
rect 36084 4422 36136 4428
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 35532 4072 35584 4078
rect 35532 4014 35584 4020
rect 35256 3936 35308 3942
rect 35256 3878 35308 3884
rect 35164 3732 35216 3738
rect 35164 3674 35216 3680
rect 34796 3528 34848 3534
rect 34716 3488 34796 3516
rect 34796 3470 34848 3476
rect 34888 3528 34940 3534
rect 34888 3470 34940 3476
rect 34980 3528 35032 3534
rect 34980 3470 35032 3476
rect 35544 3482 35572 4014
rect 35912 3738 35940 4134
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 35900 3732 35952 3738
rect 35900 3674 35952 3680
rect 35992 3528 36044 3534
rect 34612 3052 34664 3058
rect 34612 2994 34664 3000
rect 34624 2961 34652 2994
rect 34610 2952 34666 2961
rect 34610 2887 34666 2896
rect 34428 2848 34480 2854
rect 34428 2790 34480 2796
rect 34808 2650 34836 3470
rect 34900 3233 34928 3470
rect 34886 3224 34942 3233
rect 34886 3159 34942 3168
rect 34992 2650 35020 3470
rect 35544 3454 35756 3482
rect 36096 3516 36124 4422
rect 36280 4214 36308 4422
rect 36268 4208 36320 4214
rect 36268 4150 36320 4156
rect 36044 3488 36124 3516
rect 35992 3470 36044 3476
rect 35728 3398 35756 3454
rect 35624 3392 35676 3398
rect 35624 3334 35676 3340
rect 35716 3392 35768 3398
rect 35716 3334 35768 3340
rect 35348 2984 35400 2990
rect 35162 2952 35218 2961
rect 35348 2926 35400 2932
rect 35162 2887 35218 2896
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 34980 2644 35032 2650
rect 34980 2586 35032 2592
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34348 2378 34468 2394
rect 34348 2372 34480 2378
rect 34348 2366 34428 2372
rect 34060 2304 34112 2310
rect 34060 2246 34112 2252
rect 34072 2106 34100 2246
rect 34060 2100 34112 2106
rect 34060 2042 34112 2048
rect 34072 870 34192 898
rect 34072 800 34100 870
rect 32508 734 32720 762
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34164 762 34192 870
rect 34348 762 34376 2366
rect 34428 2314 34480 2320
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 34808 1170 34836 2246
rect 34624 1142 34836 1170
rect 34624 800 34652 1142
rect 35176 800 35204 2887
rect 35360 1562 35388 2926
rect 35636 2514 35664 3334
rect 36280 3126 36308 4150
rect 36268 3120 36320 3126
rect 36268 3062 36320 3068
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 2582 36032 2790
rect 35992 2576 36044 2582
rect 35992 2518 36044 2524
rect 35624 2508 35676 2514
rect 35624 2450 35676 2456
rect 35716 2508 35768 2514
rect 35716 2450 35768 2456
rect 35348 1556 35400 1562
rect 35348 1498 35400 1504
rect 35728 800 35756 2450
rect 36188 2446 36216 2994
rect 36648 2922 36676 6174
rect 36728 6112 36780 6118
rect 36728 6054 36780 6060
rect 36740 5098 36768 6054
rect 37060 6012 37368 6021
rect 37060 6010 37066 6012
rect 37122 6010 37146 6012
rect 37202 6010 37226 6012
rect 37282 6010 37306 6012
rect 37362 6010 37368 6012
rect 37122 5958 37124 6010
rect 37304 5958 37306 6010
rect 37060 5956 37066 5958
rect 37122 5956 37146 5958
rect 37202 5956 37226 5958
rect 37282 5956 37306 5958
rect 37362 5956 37368 5958
rect 37060 5947 37368 5956
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 37464 5704 37516 5710
rect 37464 5646 37516 5652
rect 36924 5114 36952 5646
rect 37476 5370 37504 5646
rect 37568 5370 37596 11222
rect 38108 11008 38160 11014
rect 38108 10950 38160 10956
rect 37648 10668 37700 10674
rect 37648 10610 37700 10616
rect 37660 10266 37688 10610
rect 37648 10260 37700 10266
rect 37648 10202 37700 10208
rect 38120 10062 38148 10950
rect 38212 10470 38240 15030
rect 38660 14816 38712 14822
rect 38660 14758 38712 14764
rect 38292 14000 38344 14006
rect 38292 13942 38344 13948
rect 38304 13394 38332 13942
rect 38384 13864 38436 13870
rect 38384 13806 38436 13812
rect 38292 13388 38344 13394
rect 38292 13330 38344 13336
rect 38304 11218 38332 13330
rect 38292 11212 38344 11218
rect 38292 11154 38344 11160
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38212 9926 38240 10406
rect 38304 10130 38332 11154
rect 38292 10124 38344 10130
rect 38292 10066 38344 10072
rect 38200 9920 38252 9926
rect 38200 9862 38252 9868
rect 37740 9376 37792 9382
rect 37740 9318 37792 9324
rect 37752 8498 37780 9318
rect 38292 8832 38344 8838
rect 38292 8774 38344 8780
rect 37740 8492 37792 8498
rect 37740 8434 37792 8440
rect 37752 7954 37780 8434
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 37752 7546 37780 7890
rect 38304 7546 38332 8774
rect 37740 7540 37792 7546
rect 37740 7482 37792 7488
rect 38292 7540 38344 7546
rect 38292 7482 38344 7488
rect 37752 7002 37780 7482
rect 37740 6996 37792 7002
rect 37740 6938 37792 6944
rect 37752 6458 37780 6938
rect 38200 6656 38252 6662
rect 38200 6598 38252 6604
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 38212 6186 38240 6598
rect 38200 6180 38252 6186
rect 38200 6122 38252 6128
rect 38396 6118 38424 13806
rect 38672 12434 38700 14758
rect 39120 13184 39172 13190
rect 39120 13126 39172 13132
rect 39132 12646 39160 13126
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 38672 12406 38792 12434
rect 38764 11830 38792 12406
rect 39028 12096 39080 12102
rect 39028 12038 39080 12044
rect 38752 11824 38804 11830
rect 38752 11766 38804 11772
rect 38764 9654 38792 11766
rect 39040 11694 39068 12038
rect 39028 11688 39080 11694
rect 39028 11630 39080 11636
rect 38844 11008 38896 11014
rect 38844 10950 38896 10956
rect 38856 10810 38884 10950
rect 38844 10804 38896 10810
rect 38844 10746 38896 10752
rect 38752 9648 38804 9654
rect 38752 9590 38804 9596
rect 38660 8832 38712 8838
rect 38660 8774 38712 8780
rect 38672 8498 38700 8774
rect 38660 8492 38712 8498
rect 38660 8434 38712 8440
rect 38476 7200 38528 7206
rect 38476 7142 38528 7148
rect 38488 6866 38516 7142
rect 38476 6860 38528 6866
rect 38476 6802 38528 6808
rect 38764 6730 38792 9590
rect 38844 8968 38896 8974
rect 38844 8910 38896 8916
rect 38856 7546 38884 8910
rect 38936 7812 38988 7818
rect 38936 7754 38988 7760
rect 38844 7540 38896 7546
rect 38844 7482 38896 7488
rect 38844 7404 38896 7410
rect 38844 7346 38896 7352
rect 38856 7002 38884 7346
rect 38844 6996 38896 7002
rect 38844 6938 38896 6944
rect 38948 6866 38976 7754
rect 39040 7342 39068 11630
rect 39120 11552 39172 11558
rect 39120 11494 39172 11500
rect 39132 10062 39160 11494
rect 39120 10056 39172 10062
rect 39120 9998 39172 10004
rect 39316 9654 39344 16390
rect 39408 15706 39436 16390
rect 39500 16250 39528 16594
rect 39488 16244 39540 16250
rect 39488 16186 39540 16192
rect 39488 15904 39540 15910
rect 39488 15846 39540 15852
rect 39396 15700 39448 15706
rect 39396 15642 39448 15648
rect 39304 9648 39356 9654
rect 39304 9590 39356 9596
rect 39396 8560 39448 8566
rect 39396 8502 39448 8508
rect 39408 8090 39436 8502
rect 39396 8084 39448 8090
rect 39396 8026 39448 8032
rect 39120 7744 39172 7750
rect 39120 7686 39172 7692
rect 39028 7336 39080 7342
rect 39028 7278 39080 7284
rect 38936 6860 38988 6866
rect 38936 6802 38988 6808
rect 38752 6724 38804 6730
rect 38752 6666 38804 6672
rect 39040 6662 39068 7278
rect 39132 6866 39160 7686
rect 39120 6860 39172 6866
rect 39120 6802 39172 6808
rect 39396 6724 39448 6730
rect 39396 6666 39448 6672
rect 39028 6656 39080 6662
rect 39028 6598 39080 6604
rect 38568 6248 38620 6254
rect 38568 6190 38620 6196
rect 38384 6112 38436 6118
rect 38384 6054 38436 6060
rect 37464 5364 37516 5370
rect 37464 5306 37516 5312
rect 37556 5364 37608 5370
rect 37556 5306 37608 5312
rect 36728 5092 36780 5098
rect 36728 5034 36780 5040
rect 36832 5086 36952 5114
rect 36740 4604 36768 5034
rect 36832 4758 36860 5086
rect 36912 5024 36964 5030
rect 36912 4966 36964 4972
rect 36924 4826 36952 4966
rect 37060 4924 37368 4933
rect 37060 4922 37066 4924
rect 37122 4922 37146 4924
rect 37202 4922 37226 4924
rect 37282 4922 37306 4924
rect 37362 4922 37368 4924
rect 37122 4870 37124 4922
rect 37304 4870 37306 4922
rect 37060 4868 37066 4870
rect 37122 4868 37146 4870
rect 37202 4868 37226 4870
rect 37282 4868 37306 4870
rect 37362 4868 37368 4870
rect 37060 4859 37368 4868
rect 36912 4820 36964 4826
rect 36912 4762 36964 4768
rect 36820 4752 36872 4758
rect 36820 4694 36872 4700
rect 37280 4684 37332 4690
rect 37280 4626 37332 4632
rect 36820 4616 36872 4622
rect 36740 4576 36820 4604
rect 36820 4558 36872 4564
rect 36832 4282 36860 4558
rect 36820 4276 36872 4282
rect 36820 4218 36872 4224
rect 37292 4049 37320 4626
rect 37476 4570 37504 5306
rect 37556 5160 37608 5166
rect 37556 5102 37608 5108
rect 37384 4542 37504 4570
rect 37568 4554 37596 5102
rect 37648 5092 37700 5098
rect 37648 5034 37700 5040
rect 37556 4548 37608 4554
rect 37384 4078 37412 4542
rect 37556 4490 37608 4496
rect 37464 4480 37516 4486
rect 37464 4422 37516 4428
rect 37476 4282 37504 4422
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37372 4072 37424 4078
rect 37278 4040 37334 4049
rect 37372 4014 37424 4020
rect 37278 3975 37334 3984
rect 37060 3836 37368 3845
rect 37060 3834 37066 3836
rect 37122 3834 37146 3836
rect 37202 3834 37226 3836
rect 37282 3834 37306 3836
rect 37362 3834 37368 3836
rect 37122 3782 37124 3834
rect 37304 3782 37306 3834
rect 37060 3780 37066 3782
rect 37122 3780 37146 3782
rect 37202 3780 37226 3782
rect 37282 3780 37306 3782
rect 37362 3780 37368 3782
rect 37060 3771 37368 3780
rect 37568 3738 37596 4490
rect 37556 3732 37608 3738
rect 37556 3674 37608 3680
rect 37660 3618 37688 5034
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37740 3936 37792 3942
rect 37740 3878 37792 3884
rect 37568 3590 37688 3618
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37384 3194 37412 3470
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 36636 2916 36688 2922
rect 36636 2858 36688 2864
rect 36820 2916 36872 2922
rect 36820 2858 36872 2864
rect 36268 2848 36320 2854
rect 36268 2790 36320 2796
rect 36176 2440 36228 2446
rect 36176 2382 36228 2388
rect 35808 2304 35860 2310
rect 35808 2246 35860 2252
rect 35820 2038 35848 2246
rect 35808 2032 35860 2038
rect 35808 1974 35860 1980
rect 36280 800 36308 2790
rect 36832 800 36860 2858
rect 37476 2854 37504 3130
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37060 2748 37368 2757
rect 37060 2746 37066 2748
rect 37122 2746 37146 2748
rect 37202 2746 37226 2748
rect 37282 2746 37306 2748
rect 37362 2746 37368 2748
rect 37122 2694 37124 2746
rect 37304 2694 37306 2746
rect 37060 2692 37066 2694
rect 37122 2692 37146 2694
rect 37202 2692 37226 2694
rect 37282 2692 37306 2694
rect 37362 2692 37368 2694
rect 37060 2683 37368 2692
rect 37568 2446 37596 3590
rect 37752 3126 37780 3878
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 37844 3058 37872 4966
rect 38396 4842 38424 6054
rect 38580 5914 38608 6190
rect 38568 5908 38620 5914
rect 38568 5850 38620 5856
rect 39040 5681 39068 6598
rect 39120 6112 39172 6118
rect 39120 6054 39172 6060
rect 39026 5672 39082 5681
rect 39026 5607 39082 5616
rect 39132 5302 39160 6054
rect 39408 5778 39436 6666
rect 39396 5772 39448 5778
rect 39396 5714 39448 5720
rect 39120 5296 39172 5302
rect 39120 5238 39172 5244
rect 39396 5160 39448 5166
rect 39396 5102 39448 5108
rect 38304 4814 38424 4842
rect 38304 4758 38332 4814
rect 38292 4752 38344 4758
rect 38014 4720 38070 4729
rect 38292 4694 38344 4700
rect 38014 4655 38070 4664
rect 38028 4622 38056 4655
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 39212 4548 39264 4554
rect 39212 4490 39264 4496
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 37832 3052 37884 3058
rect 37832 2994 37884 3000
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37384 870 37504 898
rect 37384 800 37412 870
rect 34164 734 34376 762
rect 34610 0 34666 800
rect 35162 0 35218 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37476 762 37504 870
rect 37660 762 37688 2926
rect 38016 2372 38068 2378
rect 38016 2314 38068 2320
rect 38028 1306 38056 2314
rect 38212 2106 38240 4422
rect 39224 4282 39252 4490
rect 39212 4276 39264 4282
rect 39212 4218 39264 4224
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 39028 4140 39080 4146
rect 39028 4082 39080 4088
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 38200 2100 38252 2106
rect 38200 2042 38252 2048
rect 38396 1850 38424 3334
rect 38672 2650 38700 4082
rect 39040 3738 39068 4082
rect 39028 3732 39080 3738
rect 39028 3674 39080 3680
rect 39408 3670 39436 5102
rect 39500 4010 39528 15846
rect 39592 15162 39620 16748
rect 39776 16250 39804 16934
rect 39960 16561 39988 18022
rect 40132 17672 40184 17678
rect 40132 17614 40184 17620
rect 40040 17536 40092 17542
rect 40040 17478 40092 17484
rect 40052 17338 40080 17478
rect 40040 17332 40092 17338
rect 40040 17274 40092 17280
rect 40052 16658 40080 17274
rect 40144 16794 40172 17614
rect 40132 16788 40184 16794
rect 40132 16730 40184 16736
rect 40040 16652 40092 16658
rect 40040 16594 40092 16600
rect 39946 16552 40002 16561
rect 39946 16487 40002 16496
rect 40052 16250 40080 16594
rect 39764 16244 39816 16250
rect 39764 16186 39816 16192
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 40236 16182 40264 20198
rect 41052 19780 41104 19786
rect 41052 19722 41104 19728
rect 41064 18970 41092 19722
rect 41512 19712 41564 19718
rect 41512 19654 41564 19660
rect 41788 19712 41840 19718
rect 41788 19654 41840 19660
rect 41326 19408 41382 19417
rect 41326 19343 41382 19352
rect 41052 18964 41104 18970
rect 41052 18906 41104 18912
rect 41236 18624 41288 18630
rect 41236 18566 41288 18572
rect 40776 17740 40828 17746
rect 40776 17682 40828 17688
rect 40684 17536 40736 17542
rect 40684 17478 40736 17484
rect 40696 17338 40724 17478
rect 40788 17338 40816 17682
rect 40684 17332 40736 17338
rect 40684 17274 40736 17280
rect 40776 17332 40828 17338
rect 40776 17274 40828 17280
rect 40408 16652 40460 16658
rect 40408 16594 40460 16600
rect 40224 16176 40276 16182
rect 40224 16118 40276 16124
rect 40316 16176 40368 16182
rect 40316 16118 40368 16124
rect 40328 15706 40356 16118
rect 40316 15700 40368 15706
rect 40316 15642 40368 15648
rect 40420 15366 40448 16594
rect 40960 16448 41012 16454
rect 40960 16390 41012 16396
rect 41248 16402 41276 18566
rect 41340 18154 41368 19343
rect 41524 18834 41552 19654
rect 41800 19514 41828 19654
rect 41788 19508 41840 19514
rect 41788 19450 41840 19456
rect 41512 18828 41564 18834
rect 41512 18770 41564 18776
rect 41328 18148 41380 18154
rect 41328 18090 41380 18096
rect 41512 18148 41564 18154
rect 41564 18108 41644 18136
rect 41512 18090 41564 18096
rect 41512 17672 41564 17678
rect 41512 17614 41564 17620
rect 41420 17536 41472 17542
rect 41420 17478 41472 17484
rect 41432 16522 41460 17478
rect 41524 17338 41552 17614
rect 41512 17332 41564 17338
rect 41512 17274 41564 17280
rect 41616 16561 41644 18108
rect 41788 16652 41840 16658
rect 41788 16594 41840 16600
rect 41602 16552 41658 16561
rect 41420 16516 41472 16522
rect 41658 16510 41736 16538
rect 41602 16487 41658 16496
rect 41420 16458 41472 16464
rect 40972 16114 41000 16390
rect 41248 16374 41460 16402
rect 40960 16108 41012 16114
rect 40960 16050 41012 16056
rect 41432 15706 41460 16374
rect 41420 15700 41472 15706
rect 41420 15642 41472 15648
rect 41144 15496 41196 15502
rect 41144 15438 41196 15444
rect 40408 15360 40460 15366
rect 40408 15302 40460 15308
rect 39580 15156 39632 15162
rect 39580 15098 39632 15104
rect 41052 14884 41104 14890
rect 41052 14826 41104 14832
rect 39672 14816 39724 14822
rect 39672 14758 39724 14764
rect 39684 14482 39712 14758
rect 39672 14476 39724 14482
rect 39672 14418 39724 14424
rect 40684 14408 40736 14414
rect 40684 14350 40736 14356
rect 39672 14272 39724 14278
rect 39672 14214 39724 14220
rect 40132 14272 40184 14278
rect 40132 14214 40184 14220
rect 40592 14272 40644 14278
rect 40592 14214 40644 14220
rect 39684 13326 39712 14214
rect 39948 13932 40000 13938
rect 39948 13874 40000 13880
rect 39672 13320 39724 13326
rect 39672 13262 39724 13268
rect 39856 13184 39908 13190
rect 39856 13126 39908 13132
rect 39868 12986 39896 13126
rect 39960 12986 39988 13874
rect 40144 13190 40172 14214
rect 40604 13938 40632 14214
rect 40592 13932 40644 13938
rect 40592 13874 40644 13880
rect 40224 13864 40276 13870
rect 40224 13806 40276 13812
rect 40132 13184 40184 13190
rect 40132 13126 40184 13132
rect 39856 12980 39908 12986
rect 39856 12922 39908 12928
rect 39948 12980 40000 12986
rect 39948 12922 40000 12928
rect 40144 12434 40172 13126
rect 40236 12850 40264 13806
rect 40592 13728 40644 13734
rect 40592 13670 40644 13676
rect 40604 13376 40632 13670
rect 40696 13530 40724 14350
rect 41064 13802 41092 14826
rect 41052 13796 41104 13802
rect 41052 13738 41104 13744
rect 41064 13682 41092 13738
rect 40972 13654 41092 13682
rect 40684 13524 40736 13530
rect 40684 13466 40736 13472
rect 40684 13388 40736 13394
rect 40604 13348 40684 13376
rect 40684 13330 40736 13336
rect 40316 13184 40368 13190
rect 40316 13126 40368 13132
rect 40328 12986 40356 13126
rect 40696 12986 40724 13330
rect 40316 12980 40368 12986
rect 40316 12922 40368 12928
rect 40684 12980 40736 12986
rect 40684 12922 40736 12928
rect 40224 12844 40276 12850
rect 40224 12786 40276 12792
rect 40696 12442 40724 12922
rect 40684 12436 40736 12442
rect 40144 12406 40264 12434
rect 40236 11830 40264 12406
rect 40684 12378 40736 12384
rect 40224 11824 40276 11830
rect 40224 11766 40276 11772
rect 40040 11688 40092 11694
rect 40040 11630 40092 11636
rect 39672 11552 39724 11558
rect 39672 11494 39724 11500
rect 39684 11354 39712 11494
rect 40052 11354 40080 11630
rect 39672 11348 39724 11354
rect 39672 11290 39724 11296
rect 40040 11348 40092 11354
rect 40040 11290 40092 11296
rect 40236 11082 40264 11766
rect 40500 11756 40552 11762
rect 40500 11698 40552 11704
rect 40316 11620 40368 11626
rect 40316 11562 40368 11568
rect 40328 11354 40356 11562
rect 40316 11348 40368 11354
rect 40316 11290 40368 11296
rect 40408 11212 40460 11218
rect 40408 11154 40460 11160
rect 40224 11076 40276 11082
rect 40224 11018 40276 11024
rect 40420 11014 40448 11154
rect 39856 11008 39908 11014
rect 39856 10950 39908 10956
rect 40408 11008 40460 11014
rect 40408 10950 40460 10956
rect 39764 9580 39816 9586
rect 39764 9522 39816 9528
rect 39580 5160 39632 5166
rect 39580 5102 39632 5108
rect 39592 4826 39620 5102
rect 39580 4820 39632 4826
rect 39580 4762 39632 4768
rect 39776 4078 39804 9522
rect 39868 7342 39896 10950
rect 40316 10464 40368 10470
rect 40316 10406 40368 10412
rect 40132 9376 40184 9382
rect 40132 9318 40184 9324
rect 40040 8628 40092 8634
rect 40040 8570 40092 8576
rect 40052 7970 40080 8570
rect 40144 8498 40172 9318
rect 40328 9042 40356 10406
rect 40512 10266 40540 11698
rect 40684 11552 40736 11558
rect 40684 11494 40736 11500
rect 40696 11354 40724 11494
rect 40972 11354 41000 13654
rect 40684 11348 40736 11354
rect 40684 11290 40736 11296
rect 40960 11348 41012 11354
rect 40960 11290 41012 11296
rect 40972 10810 41000 11290
rect 40960 10804 41012 10810
rect 40960 10746 41012 10752
rect 40500 10260 40552 10266
rect 40500 10202 40552 10208
rect 40972 9722 41000 10746
rect 41156 10266 41184 15438
rect 41604 15156 41656 15162
rect 41604 15098 41656 15104
rect 41616 13870 41644 15098
rect 41708 14618 41736 16510
rect 41696 14612 41748 14618
rect 41696 14554 41748 14560
rect 41800 14464 41828 16594
rect 41708 14436 41828 14464
rect 41420 13864 41472 13870
rect 41340 13812 41420 13818
rect 41340 13806 41472 13812
rect 41604 13864 41656 13870
rect 41604 13806 41656 13812
rect 41340 13790 41460 13806
rect 41340 13530 41368 13790
rect 41616 13682 41644 13806
rect 41432 13654 41644 13682
rect 41328 13524 41380 13530
rect 41328 13466 41380 13472
rect 41432 12434 41460 13654
rect 41708 13546 41736 14436
rect 41788 14272 41840 14278
rect 41788 14214 41840 14220
rect 41616 13518 41736 13546
rect 41616 12866 41644 13518
rect 41696 13252 41748 13258
rect 41696 13194 41748 13200
rect 41708 12986 41736 13194
rect 41696 12980 41748 12986
rect 41696 12922 41748 12928
rect 41616 12838 41736 12866
rect 41800 12850 41828 14214
rect 41892 13326 41920 20878
rect 42340 20800 42392 20806
rect 42340 20742 42392 20748
rect 42064 20528 42116 20534
rect 42064 20470 42116 20476
rect 42076 19718 42104 20470
rect 42352 20466 42380 20742
rect 42340 20460 42392 20466
rect 42340 20402 42392 20408
rect 42720 20262 42748 21422
rect 43260 21344 43312 21350
rect 43260 21286 43312 21292
rect 43904 21344 43956 21350
rect 43904 21286 43956 21292
rect 46112 21344 46164 21350
rect 46112 21286 46164 21292
rect 46480 21344 46532 21350
rect 46480 21286 46532 21292
rect 43272 20602 43300 21286
rect 43916 21078 43944 21286
rect 46124 21078 46152 21286
rect 43904 21072 43956 21078
rect 43904 21014 43956 21020
rect 46112 21072 46164 21078
rect 46112 21014 46164 21020
rect 43260 20596 43312 20602
rect 43260 20538 43312 20544
rect 43916 20534 43944 21014
rect 44732 20936 44784 20942
rect 44732 20878 44784 20884
rect 45008 20936 45060 20942
rect 45008 20878 45060 20884
rect 44640 20800 44692 20806
rect 44640 20742 44692 20748
rect 44282 20700 44590 20709
rect 44282 20698 44288 20700
rect 44344 20698 44368 20700
rect 44424 20698 44448 20700
rect 44504 20698 44528 20700
rect 44584 20698 44590 20700
rect 44344 20646 44346 20698
rect 44526 20646 44528 20698
rect 44282 20644 44288 20646
rect 44344 20644 44368 20646
rect 44424 20644 44448 20646
rect 44504 20644 44528 20646
rect 44584 20644 44590 20646
rect 44282 20635 44590 20644
rect 43904 20528 43956 20534
rect 43074 20496 43130 20505
rect 43904 20470 43956 20476
rect 43074 20431 43130 20440
rect 43168 20460 43220 20466
rect 43088 20398 43116 20431
rect 43168 20402 43220 20408
rect 43076 20392 43128 20398
rect 43076 20334 43128 20340
rect 42708 20256 42760 20262
rect 42708 20198 42760 20204
rect 42616 19916 42668 19922
rect 42616 19858 42668 19864
rect 42064 19712 42116 19718
rect 42064 19654 42116 19660
rect 42076 19514 42104 19654
rect 42064 19508 42116 19514
rect 42064 19450 42116 19456
rect 41972 19372 42024 19378
rect 41972 19314 42024 19320
rect 41984 18970 42012 19314
rect 41972 18964 42024 18970
rect 41972 18906 42024 18912
rect 42076 18850 42104 19450
rect 42628 19378 42656 19858
rect 43180 19378 43208 20402
rect 43628 20256 43680 20262
rect 43628 20198 43680 20204
rect 43260 19916 43312 19922
rect 43260 19858 43312 19864
rect 42616 19372 42668 19378
rect 42616 19314 42668 19320
rect 43168 19372 43220 19378
rect 43168 19314 43220 19320
rect 43180 18970 43208 19314
rect 43168 18964 43220 18970
rect 43168 18906 43220 18912
rect 43272 18902 43300 19858
rect 43640 19854 43668 20198
rect 44652 19922 44680 20742
rect 44744 20262 44772 20878
rect 44916 20392 44968 20398
rect 44916 20334 44968 20340
rect 44732 20256 44784 20262
rect 44732 20198 44784 20204
rect 44744 20058 44772 20198
rect 44928 20058 44956 20334
rect 44732 20052 44784 20058
rect 44732 19994 44784 20000
rect 44916 20052 44968 20058
rect 44916 19994 44968 20000
rect 44088 19916 44140 19922
rect 44088 19858 44140 19864
rect 44640 19916 44692 19922
rect 44640 19858 44692 19864
rect 43628 19848 43680 19854
rect 43628 19790 43680 19796
rect 43996 19712 44048 19718
rect 43996 19654 44048 19660
rect 44008 19514 44036 19654
rect 43996 19508 44048 19514
rect 43996 19450 44048 19456
rect 41984 18822 42104 18850
rect 43260 18896 43312 18902
rect 43260 18838 43312 18844
rect 41984 17134 42012 18822
rect 42064 18080 42116 18086
rect 42064 18022 42116 18028
rect 42076 17134 42104 18022
rect 42156 17536 42208 17542
rect 42156 17478 42208 17484
rect 41972 17128 42024 17134
rect 41972 17070 42024 17076
rect 42064 17128 42116 17134
rect 42064 17070 42116 17076
rect 42064 16992 42116 16998
rect 42064 16934 42116 16940
rect 42076 15434 42104 16934
rect 42168 16590 42196 17478
rect 42708 17264 42760 17270
rect 42708 17206 42760 17212
rect 42432 17128 42484 17134
rect 42432 17070 42484 17076
rect 42444 16794 42472 17070
rect 42432 16788 42484 16794
rect 42432 16730 42484 16736
rect 42720 16658 42748 17206
rect 43272 16658 43300 18838
rect 43352 17740 43404 17746
rect 43352 17682 43404 17688
rect 42708 16652 42760 16658
rect 42708 16594 42760 16600
rect 43260 16652 43312 16658
rect 43260 16594 43312 16600
rect 42156 16584 42208 16590
rect 42156 16526 42208 16532
rect 42524 16448 42576 16454
rect 42524 16390 42576 16396
rect 42536 16046 42564 16390
rect 42800 16244 42852 16250
rect 42800 16186 42852 16192
rect 42432 16040 42484 16046
rect 42432 15982 42484 15988
rect 42524 16040 42576 16046
rect 42524 15982 42576 15988
rect 42444 15706 42472 15982
rect 42432 15700 42484 15706
rect 42432 15642 42484 15648
rect 42812 15570 42840 16186
rect 43364 15910 43392 17682
rect 43904 17536 43956 17542
rect 43904 17478 43956 17484
rect 43444 17128 43496 17134
rect 43444 17070 43496 17076
rect 43456 16998 43484 17070
rect 43444 16992 43496 16998
rect 43444 16934 43496 16940
rect 43456 15910 43484 16934
rect 43628 16584 43680 16590
rect 43628 16526 43680 16532
rect 43640 16250 43668 16526
rect 43628 16244 43680 16250
rect 43628 16186 43680 16192
rect 43352 15904 43404 15910
rect 43352 15846 43404 15852
rect 43444 15904 43496 15910
rect 43444 15846 43496 15852
rect 42800 15564 42852 15570
rect 42800 15506 42852 15512
rect 42064 15428 42116 15434
rect 42064 15370 42116 15376
rect 43352 15156 43404 15162
rect 43352 15098 43404 15104
rect 42064 14816 42116 14822
rect 42064 14758 42116 14764
rect 42076 14346 42104 14758
rect 43364 14482 43392 15098
rect 43352 14476 43404 14482
rect 43352 14418 43404 14424
rect 42064 14340 42116 14346
rect 42064 14282 42116 14288
rect 42076 14226 42104 14282
rect 43076 14272 43128 14278
rect 42076 14198 42196 14226
rect 43076 14214 43128 14220
rect 42168 14074 42196 14198
rect 42064 14068 42116 14074
rect 42064 14010 42116 14016
rect 42156 14068 42208 14074
rect 42156 14010 42208 14016
rect 42800 14068 42852 14074
rect 42800 14010 42852 14016
rect 42076 13530 42104 14010
rect 42432 13728 42484 13734
rect 42432 13670 42484 13676
rect 42064 13524 42116 13530
rect 42064 13466 42116 13472
rect 41880 13320 41932 13326
rect 41880 13262 41932 13268
rect 41432 12406 41552 12434
rect 41420 12300 41472 12306
rect 41420 12242 41472 12248
rect 41432 11234 41460 12242
rect 41340 11206 41460 11234
rect 41340 11150 41368 11206
rect 41328 11144 41380 11150
rect 41328 11086 41380 11092
rect 41432 10690 41460 11206
rect 41524 10810 41552 12406
rect 41708 12374 41736 12838
rect 41788 12844 41840 12850
rect 41788 12786 41840 12792
rect 41892 12434 41920 13262
rect 42076 12850 42104 13466
rect 42444 12986 42472 13670
rect 42432 12980 42484 12986
rect 42432 12922 42484 12928
rect 42064 12844 42116 12850
rect 42064 12786 42116 12792
rect 41892 12406 42104 12434
rect 41696 12368 41748 12374
rect 41696 12310 41748 12316
rect 42076 12102 42104 12406
rect 42340 12368 42392 12374
rect 42340 12310 42392 12316
rect 42248 12232 42300 12238
rect 42248 12174 42300 12180
rect 42064 12096 42116 12102
rect 42064 12038 42116 12044
rect 42156 12096 42208 12102
rect 42156 12038 42208 12044
rect 41880 11552 41932 11558
rect 41880 11494 41932 11500
rect 41892 11218 41920 11494
rect 41880 11212 41932 11218
rect 41880 11154 41932 11160
rect 41972 11144 42024 11150
rect 41972 11086 42024 11092
rect 41512 10804 41564 10810
rect 41512 10746 41564 10752
rect 41432 10662 41552 10690
rect 41144 10260 41196 10266
rect 41144 10202 41196 10208
rect 41524 9926 41552 10662
rect 41788 10260 41840 10266
rect 41788 10202 41840 10208
rect 41512 9920 41564 9926
rect 41512 9862 41564 9868
rect 40500 9716 40552 9722
rect 40500 9658 40552 9664
rect 40960 9716 41012 9722
rect 40960 9658 41012 9664
rect 40408 9512 40460 9518
rect 40408 9454 40460 9460
rect 40420 9178 40448 9454
rect 40408 9172 40460 9178
rect 40408 9114 40460 9120
rect 40316 9036 40368 9042
rect 40316 8978 40368 8984
rect 40224 8832 40276 8838
rect 40224 8774 40276 8780
rect 40132 8492 40184 8498
rect 40132 8434 40184 8440
rect 40132 8016 40184 8022
rect 40052 7964 40132 7970
rect 40052 7958 40184 7964
rect 40052 7942 40172 7958
rect 40052 7342 40080 7942
rect 40236 7546 40264 8774
rect 40408 8628 40460 8634
rect 40408 8570 40460 8576
rect 40420 7954 40448 8570
rect 40512 7954 40540 9658
rect 41144 9512 41196 9518
rect 41144 9454 41196 9460
rect 40776 9104 40828 9110
rect 40776 9046 40828 9052
rect 40788 8906 40816 9046
rect 40776 8900 40828 8906
rect 40776 8842 40828 8848
rect 41156 8634 41184 9454
rect 41328 9444 41380 9450
rect 41328 9386 41380 9392
rect 41236 9376 41288 9382
rect 41236 9318 41288 9324
rect 41248 9178 41276 9318
rect 41340 9178 41368 9386
rect 41236 9172 41288 9178
rect 41236 9114 41288 9120
rect 41328 9172 41380 9178
rect 41328 9114 41380 9120
rect 41800 9042 41828 10202
rect 41984 10130 42012 11086
rect 42076 10538 42104 12038
rect 42168 11898 42196 12038
rect 42156 11892 42208 11898
rect 42156 11834 42208 11840
rect 42260 11558 42288 12174
rect 42248 11552 42300 11558
rect 42248 11494 42300 11500
rect 42156 11144 42208 11150
rect 42156 11086 42208 11092
rect 42168 10810 42196 11086
rect 42156 10804 42208 10810
rect 42156 10746 42208 10752
rect 42064 10532 42116 10538
rect 42064 10474 42116 10480
rect 41972 10124 42024 10130
rect 41972 10066 42024 10072
rect 41880 9920 41932 9926
rect 41880 9862 41932 9868
rect 41788 9036 41840 9042
rect 41788 8978 41840 8984
rect 41144 8628 41196 8634
rect 41144 8570 41196 8576
rect 41420 8560 41472 8566
rect 41420 8502 41472 8508
rect 40776 8288 40828 8294
rect 40776 8230 40828 8236
rect 40788 8090 40816 8230
rect 40776 8084 40828 8090
rect 40776 8026 40828 8032
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 40408 7948 40460 7954
rect 40408 7890 40460 7896
rect 40500 7948 40552 7954
rect 40500 7890 40552 7896
rect 40224 7540 40276 7546
rect 40224 7482 40276 7488
rect 40132 7472 40184 7478
rect 40132 7414 40184 7420
rect 39856 7336 39908 7342
rect 39856 7278 39908 7284
rect 40040 7336 40092 7342
rect 40040 7278 40092 7284
rect 39868 6866 39896 7278
rect 40040 7200 40092 7206
rect 40040 7142 40092 7148
rect 39856 6860 39908 6866
rect 39856 6802 39908 6808
rect 39868 6458 39896 6802
rect 40052 6662 40080 7142
rect 40040 6656 40092 6662
rect 40040 6598 40092 6604
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 40144 6254 40172 7414
rect 40236 6458 40264 7482
rect 40512 7002 40540 7890
rect 40868 7880 40920 7886
rect 40868 7822 40920 7828
rect 40880 7750 40908 7822
rect 40868 7744 40920 7750
rect 40868 7686 40920 7692
rect 40972 7002 41000 8026
rect 41432 7954 41460 8502
rect 41420 7948 41472 7954
rect 41420 7890 41472 7896
rect 41052 7880 41104 7886
rect 41052 7822 41104 7828
rect 41064 7478 41092 7822
rect 41432 7546 41460 7890
rect 41696 7744 41748 7750
rect 41696 7686 41748 7692
rect 41420 7540 41472 7546
rect 41420 7482 41472 7488
rect 41052 7472 41104 7478
rect 41052 7414 41104 7420
rect 40500 6996 40552 7002
rect 40500 6938 40552 6944
rect 40684 6996 40736 7002
rect 40684 6938 40736 6944
rect 40960 6996 41012 7002
rect 40960 6938 41012 6944
rect 40500 6792 40552 6798
rect 40500 6734 40552 6740
rect 40224 6452 40276 6458
rect 40224 6394 40276 6400
rect 40132 6248 40184 6254
rect 40132 6190 40184 6196
rect 39948 6112 40000 6118
rect 39948 6054 40000 6060
rect 39960 5710 39988 6054
rect 39856 5704 39908 5710
rect 39856 5646 39908 5652
rect 39948 5704 40000 5710
rect 39948 5646 40000 5652
rect 39868 5370 39896 5646
rect 39856 5364 39908 5370
rect 39856 5306 39908 5312
rect 39960 4690 39988 5646
rect 40144 5574 40172 6190
rect 40236 5914 40264 6394
rect 40512 6390 40540 6734
rect 40500 6384 40552 6390
rect 40500 6326 40552 6332
rect 40224 5908 40276 5914
rect 40224 5850 40276 5856
rect 40132 5568 40184 5574
rect 40132 5510 40184 5516
rect 40144 5166 40172 5510
rect 40132 5160 40184 5166
rect 40132 5102 40184 5108
rect 40040 4820 40092 4826
rect 40040 4762 40092 4768
rect 39948 4684 40000 4690
rect 39948 4626 40000 4632
rect 39856 4480 39908 4486
rect 39856 4422 39908 4428
rect 39868 4146 39896 4422
rect 40052 4146 40080 4762
rect 40236 4554 40264 5850
rect 40408 5364 40460 5370
rect 40408 5306 40460 5312
rect 40420 5234 40448 5306
rect 40316 5228 40368 5234
rect 40316 5170 40368 5176
rect 40408 5228 40460 5234
rect 40408 5170 40460 5176
rect 40328 4826 40356 5170
rect 40316 4820 40368 4826
rect 40316 4762 40368 4768
rect 40512 4690 40540 6326
rect 40696 6322 40724 6938
rect 40684 6316 40736 6322
rect 40684 6258 40736 6264
rect 40592 5772 40644 5778
rect 40592 5714 40644 5720
rect 40500 4684 40552 4690
rect 40500 4626 40552 4632
rect 40224 4548 40276 4554
rect 40224 4490 40276 4496
rect 39856 4140 39908 4146
rect 39856 4082 39908 4088
rect 40040 4140 40092 4146
rect 40040 4082 40092 4088
rect 39764 4072 39816 4078
rect 39764 4014 39816 4020
rect 39488 4004 39540 4010
rect 39488 3946 39540 3952
rect 40040 3936 40092 3942
rect 40040 3878 40092 3884
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 38936 3528 38988 3534
rect 38936 3470 38988 3476
rect 38948 3194 38976 3470
rect 39212 3460 39264 3466
rect 39212 3402 39264 3408
rect 39224 3194 39252 3402
rect 39856 3392 39908 3398
rect 39856 3334 39908 3340
rect 39486 3224 39542 3233
rect 38936 3188 38988 3194
rect 38936 3130 38988 3136
rect 39212 3188 39264 3194
rect 39868 3194 39896 3334
rect 39486 3159 39542 3168
rect 39856 3188 39908 3194
rect 39212 3130 39264 3136
rect 38750 2952 38806 2961
rect 38750 2887 38806 2896
rect 38660 2644 38712 2650
rect 38660 2586 38712 2592
rect 38764 2514 38792 2887
rect 39500 2650 39528 3159
rect 39856 3130 39908 3136
rect 39948 3120 40000 3126
rect 39948 3062 40000 3068
rect 39960 2774 39988 3062
rect 39592 2746 39988 2774
rect 39488 2644 39540 2650
rect 39488 2586 39540 2592
rect 38752 2508 38804 2514
rect 38752 2450 38804 2456
rect 39028 2508 39080 2514
rect 39028 2450 39080 2456
rect 38396 1822 38516 1850
rect 37936 1278 38056 1306
rect 37936 800 37964 1278
rect 38488 800 38516 1822
rect 39040 800 39068 2450
rect 39592 800 39620 2746
rect 40052 2446 40080 3878
rect 40236 3466 40264 4490
rect 40316 4480 40368 4486
rect 40316 4422 40368 4428
rect 40328 4282 40356 4422
rect 40316 4276 40368 4282
rect 40316 4218 40368 4224
rect 40224 3460 40276 3466
rect 40224 3402 40276 3408
rect 40604 3194 40632 5714
rect 40696 5710 40724 6258
rect 40684 5704 40736 5710
rect 40684 5646 40736 5652
rect 40696 5030 40724 5646
rect 40776 5568 40828 5574
rect 40776 5510 40828 5516
rect 40684 5024 40736 5030
rect 40684 4966 40736 4972
rect 40788 4690 40816 5510
rect 40776 4684 40828 4690
rect 40776 4626 40828 4632
rect 40868 4616 40920 4622
rect 40868 4558 40920 4564
rect 40592 3188 40644 3194
rect 40592 3130 40644 3136
rect 40684 2984 40736 2990
rect 40684 2926 40736 2932
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 40144 800 40172 2382
rect 40696 800 40724 2926
rect 37476 734 37688 762
rect 37922 0 37978 800
rect 38474 0 38530 800
rect 39026 0 39082 800
rect 39578 0 39634 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 40880 762 40908 4558
rect 40972 3602 41000 6938
rect 41512 6860 41564 6866
rect 41512 6802 41564 6808
rect 41144 6656 41196 6662
rect 41144 6598 41196 6604
rect 40960 3596 41012 3602
rect 40960 3538 41012 3544
rect 41156 2854 41184 6598
rect 41524 6458 41552 6802
rect 41604 6792 41656 6798
rect 41604 6734 41656 6740
rect 41236 6452 41288 6458
rect 41236 6394 41288 6400
rect 41512 6452 41564 6458
rect 41512 6394 41564 6400
rect 41248 6186 41276 6394
rect 41616 6390 41644 6734
rect 41604 6384 41656 6390
rect 41604 6326 41656 6332
rect 41512 6316 41564 6322
rect 41512 6258 41564 6264
rect 41236 6180 41288 6186
rect 41236 6122 41288 6128
rect 41328 6112 41380 6118
rect 41328 6054 41380 6060
rect 41340 4078 41368 6054
rect 41420 5636 41472 5642
rect 41420 5578 41472 5584
rect 41432 5166 41460 5578
rect 41420 5160 41472 5166
rect 41420 5102 41472 5108
rect 41420 5024 41472 5030
rect 41420 4966 41472 4972
rect 41432 4146 41460 4966
rect 41420 4140 41472 4146
rect 41420 4082 41472 4088
rect 41328 4072 41380 4078
rect 41326 4040 41328 4049
rect 41380 4040 41382 4049
rect 41326 3975 41382 3984
rect 41144 2848 41196 2854
rect 41144 2790 41196 2796
rect 41524 2650 41552 6258
rect 41708 5370 41736 7686
rect 41892 6866 41920 9862
rect 42352 8838 42380 12310
rect 42812 11898 42840 14010
rect 43088 12986 43116 14214
rect 43456 13734 43484 15846
rect 43444 13728 43496 13734
rect 43444 13670 43496 13676
rect 43076 12980 43128 12986
rect 43076 12922 43128 12928
rect 43916 12434 43944 17478
rect 44100 16794 44128 19858
rect 44180 19712 44232 19718
rect 44180 19654 44232 19660
rect 44916 19712 44968 19718
rect 44916 19654 44968 19660
rect 44192 17678 44220 19654
rect 44282 19612 44590 19621
rect 44282 19610 44288 19612
rect 44344 19610 44368 19612
rect 44424 19610 44448 19612
rect 44504 19610 44528 19612
rect 44584 19610 44590 19612
rect 44344 19558 44346 19610
rect 44526 19558 44528 19610
rect 44282 19556 44288 19558
rect 44344 19556 44368 19558
rect 44424 19556 44448 19558
rect 44504 19556 44528 19558
rect 44584 19556 44590 19558
rect 44282 19547 44590 19556
rect 44548 19508 44600 19514
rect 44548 19450 44600 19456
rect 44560 19310 44588 19450
rect 44928 19378 44956 19654
rect 45020 19514 45048 20878
rect 45376 20868 45428 20874
rect 45376 20810 45428 20816
rect 45100 20256 45152 20262
rect 45100 20198 45152 20204
rect 45112 19514 45140 20198
rect 45388 19514 45416 20810
rect 45652 20800 45704 20806
rect 45652 20742 45704 20748
rect 45664 20534 45692 20742
rect 45652 20528 45704 20534
rect 45652 20470 45704 20476
rect 46124 20466 46152 21014
rect 46492 21010 46520 21286
rect 46676 21146 46704 21422
rect 47216 21344 47268 21350
rect 47216 21286 47268 21292
rect 46664 21140 46716 21146
rect 46664 21082 46716 21088
rect 46480 21004 46532 21010
rect 46480 20946 46532 20952
rect 46492 20505 46520 20946
rect 47228 20534 47256 21286
rect 47320 20874 47348 21830
rect 47308 20868 47360 20874
rect 47308 20810 47360 20816
rect 47216 20528 47268 20534
rect 46478 20496 46534 20505
rect 46112 20460 46164 20466
rect 47216 20470 47268 20476
rect 46478 20431 46534 20440
rect 46112 20402 46164 20408
rect 45468 20392 45520 20398
rect 45468 20334 45520 20340
rect 45480 19922 45508 20334
rect 45468 19916 45520 19922
rect 45468 19858 45520 19864
rect 45480 19825 45508 19858
rect 45466 19816 45522 19825
rect 45466 19751 45522 19760
rect 46124 19718 46152 20402
rect 46940 19916 46992 19922
rect 46940 19858 46992 19864
rect 45468 19712 45520 19718
rect 45468 19654 45520 19660
rect 46112 19712 46164 19718
rect 46112 19654 46164 19660
rect 45480 19514 45508 19654
rect 46124 19514 46152 19654
rect 45008 19508 45060 19514
rect 45008 19450 45060 19456
rect 45100 19508 45152 19514
rect 45100 19450 45152 19456
rect 45376 19508 45428 19514
rect 45376 19450 45428 19456
rect 45468 19508 45520 19514
rect 45468 19450 45520 19456
rect 46112 19508 46164 19514
rect 46112 19450 46164 19456
rect 44916 19372 44968 19378
rect 44916 19314 44968 19320
rect 44548 19304 44600 19310
rect 44548 19246 44600 19252
rect 45192 19304 45244 19310
rect 45192 19246 45244 19252
rect 45204 19174 45232 19246
rect 46952 19174 46980 19858
rect 47320 19854 47348 20810
rect 47596 20466 47624 22646
rect 47872 22234 47900 23054
rect 48504 22976 48556 22982
rect 48504 22918 48556 22924
rect 48516 22778 48544 22918
rect 58726 22876 59034 22885
rect 58726 22874 58732 22876
rect 58788 22874 58812 22876
rect 58868 22874 58892 22876
rect 58948 22874 58972 22876
rect 59028 22874 59034 22876
rect 58788 22822 58790 22874
rect 58970 22822 58972 22874
rect 58726 22820 58732 22822
rect 58788 22820 58812 22822
rect 58868 22820 58892 22822
rect 58948 22820 58972 22822
rect 59028 22820 59034 22822
rect 58726 22811 59034 22820
rect 48504 22772 48556 22778
rect 48504 22714 48556 22720
rect 50712 22568 50764 22574
rect 50712 22510 50764 22516
rect 51356 22568 51408 22574
rect 51356 22510 51408 22516
rect 52920 22568 52972 22574
rect 52920 22510 52972 22516
rect 55312 22568 55364 22574
rect 55312 22510 55364 22516
rect 55956 22568 56008 22574
rect 55956 22510 56008 22516
rect 48504 22432 48556 22438
rect 48504 22374 48556 22380
rect 49700 22432 49752 22438
rect 49700 22374 49752 22380
rect 47860 22228 47912 22234
rect 47860 22170 47912 22176
rect 48228 22160 48280 22166
rect 48228 22102 48280 22108
rect 48240 21350 48268 22102
rect 48516 22030 48544 22374
rect 49712 22098 49740 22374
rect 49700 22092 49752 22098
rect 49700 22034 49752 22040
rect 48504 22024 48556 22030
rect 48504 21966 48556 21972
rect 47860 21344 47912 21350
rect 47860 21286 47912 21292
rect 48228 21344 48280 21350
rect 48228 21286 48280 21292
rect 47676 20936 47728 20942
rect 47676 20878 47728 20884
rect 47688 20466 47716 20878
rect 47584 20460 47636 20466
rect 47584 20402 47636 20408
rect 47676 20460 47728 20466
rect 47676 20402 47728 20408
rect 47872 20369 47900 21286
rect 48240 20602 48268 21286
rect 48228 20596 48280 20602
rect 48228 20538 48280 20544
rect 47858 20360 47914 20369
rect 47858 20295 47860 20304
rect 47912 20295 47914 20304
rect 48320 20324 48372 20330
rect 47860 20266 47912 20272
rect 48320 20266 48372 20272
rect 47308 19848 47360 19854
rect 47308 19790 47360 19796
rect 47216 19780 47268 19786
rect 47216 19722 47268 19728
rect 47228 19446 47256 19722
rect 47216 19440 47268 19446
rect 47216 19382 47268 19388
rect 45192 19168 45244 19174
rect 45112 19128 45192 19156
rect 45112 18970 45140 19128
rect 45192 19110 45244 19116
rect 46940 19168 46992 19174
rect 46940 19110 46992 19116
rect 45100 18964 45152 18970
rect 45100 18906 45152 18912
rect 44282 18524 44590 18533
rect 44282 18522 44288 18524
rect 44344 18522 44368 18524
rect 44424 18522 44448 18524
rect 44504 18522 44528 18524
rect 44584 18522 44590 18524
rect 44344 18470 44346 18522
rect 44526 18470 44528 18522
rect 44282 18468 44288 18470
rect 44344 18468 44368 18470
rect 44424 18468 44448 18470
rect 44504 18468 44528 18470
rect 44584 18468 44590 18470
rect 44282 18459 44590 18468
rect 44180 17672 44232 17678
rect 44180 17614 44232 17620
rect 44640 17536 44692 17542
rect 44640 17478 44692 17484
rect 44916 17536 44968 17542
rect 44916 17478 44968 17484
rect 44282 17436 44590 17445
rect 44282 17434 44288 17436
rect 44344 17434 44368 17436
rect 44424 17434 44448 17436
rect 44504 17434 44528 17436
rect 44584 17434 44590 17436
rect 44344 17382 44346 17434
rect 44526 17382 44528 17434
rect 44282 17380 44288 17382
rect 44344 17380 44368 17382
rect 44424 17380 44448 17382
rect 44504 17380 44528 17382
rect 44584 17380 44590 17382
rect 44282 17371 44590 17380
rect 44652 16794 44680 17478
rect 44928 17338 44956 17478
rect 44916 17332 44968 17338
rect 44916 17274 44968 17280
rect 45008 17128 45060 17134
rect 45008 17070 45060 17076
rect 45020 16794 45048 17070
rect 44088 16788 44140 16794
rect 44088 16730 44140 16736
rect 44640 16788 44692 16794
rect 44640 16730 44692 16736
rect 45008 16788 45060 16794
rect 45008 16730 45060 16736
rect 44640 16516 44692 16522
rect 44640 16458 44692 16464
rect 44282 16348 44590 16357
rect 44282 16346 44288 16348
rect 44344 16346 44368 16348
rect 44424 16346 44448 16348
rect 44504 16346 44528 16348
rect 44584 16346 44590 16348
rect 44344 16294 44346 16346
rect 44526 16294 44528 16346
rect 44282 16292 44288 16294
rect 44344 16292 44368 16294
rect 44424 16292 44448 16294
rect 44504 16292 44528 16294
rect 44584 16292 44590 16294
rect 44282 16283 44590 16292
rect 44652 16250 44680 16458
rect 44916 16448 44968 16454
rect 44916 16390 44968 16396
rect 44928 16250 44956 16390
rect 43996 16244 44048 16250
rect 43996 16186 44048 16192
rect 44640 16244 44692 16250
rect 44640 16186 44692 16192
rect 44916 16244 44968 16250
rect 44916 16186 44968 16192
rect 44008 15366 44036 16186
rect 44928 15570 44956 16186
rect 45008 16040 45060 16046
rect 45008 15982 45060 15988
rect 45020 15706 45048 15982
rect 45008 15700 45060 15706
rect 45008 15642 45060 15648
rect 44916 15564 44968 15570
rect 44916 15506 44968 15512
rect 43996 15360 44048 15366
rect 43996 15302 44048 15308
rect 43732 12406 43944 12434
rect 42984 12300 43036 12306
rect 42984 12242 43036 12248
rect 42800 11892 42852 11898
rect 42800 11834 42852 11840
rect 42996 11778 43024 12242
rect 42628 11750 43024 11778
rect 43168 11824 43220 11830
rect 43168 11766 43220 11772
rect 42628 11558 42656 11750
rect 42996 11694 43024 11750
rect 42800 11688 42852 11694
rect 42800 11630 42852 11636
rect 42984 11688 43036 11694
rect 42984 11630 43036 11636
rect 42616 11552 42668 11558
rect 42616 11494 42668 11500
rect 42524 10668 42576 10674
rect 42524 10610 42576 10616
rect 42536 10198 42564 10610
rect 42524 10192 42576 10198
rect 42524 10134 42576 10140
rect 42536 9654 42564 10134
rect 42524 9648 42576 9654
rect 42524 9590 42576 9596
rect 42628 9602 42656 11494
rect 42812 11354 42840 11630
rect 42892 11552 42944 11558
rect 42892 11494 42944 11500
rect 42800 11348 42852 11354
rect 42800 11290 42852 11296
rect 42904 11218 42932 11494
rect 42892 11212 42944 11218
rect 42892 11154 42944 11160
rect 42708 10464 42760 10470
rect 42708 10406 42760 10412
rect 42720 9704 42748 10406
rect 42720 9676 42840 9704
rect 42432 9512 42484 9518
rect 42432 9454 42484 9460
rect 42340 8832 42392 8838
rect 42340 8774 42392 8780
rect 42156 8560 42208 8566
rect 42156 8502 42208 8508
rect 42168 8090 42196 8502
rect 42156 8084 42208 8090
rect 42156 8026 42208 8032
rect 42168 7546 42196 8026
rect 42156 7540 42208 7546
rect 42156 7482 42208 7488
rect 41972 7200 42024 7206
rect 41972 7142 42024 7148
rect 41984 6905 42012 7142
rect 41970 6896 42026 6905
rect 41880 6860 41932 6866
rect 41970 6831 42026 6840
rect 41880 6802 41932 6808
rect 41984 5794 42012 6831
rect 42248 6724 42300 6730
rect 42248 6666 42300 6672
rect 41892 5778 42012 5794
rect 41880 5772 42012 5778
rect 41932 5766 42012 5772
rect 41880 5714 41932 5720
rect 41972 5568 42024 5574
rect 41972 5510 42024 5516
rect 41696 5364 41748 5370
rect 41696 5306 41748 5312
rect 41984 4554 42012 5510
rect 41972 4548 42024 4554
rect 41972 4490 42024 4496
rect 42064 4548 42116 4554
rect 42064 4490 42116 4496
rect 41880 4480 41932 4486
rect 41880 4422 41932 4428
rect 41892 4214 41920 4422
rect 42076 4282 42104 4490
rect 42064 4276 42116 4282
rect 42064 4218 42116 4224
rect 41880 4208 41932 4214
rect 41880 4150 41932 4156
rect 41604 3936 41656 3942
rect 41604 3878 41656 3884
rect 41972 3936 42024 3942
rect 41972 3878 42024 3884
rect 41616 3194 41644 3878
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 41604 3188 41656 3194
rect 41604 3130 41656 3136
rect 41788 2984 41840 2990
rect 41788 2926 41840 2932
rect 41512 2644 41564 2650
rect 41512 2586 41564 2592
rect 41156 870 41276 898
rect 41156 762 41184 870
rect 41248 800 41276 870
rect 41800 800 41828 2926
rect 41892 2854 41920 3334
rect 41984 2854 42012 3878
rect 42260 3602 42288 6666
rect 42352 6186 42380 8774
rect 42444 8362 42472 9454
rect 42536 8498 42564 9590
rect 42628 9574 42748 9602
rect 42616 8832 42668 8838
rect 42616 8774 42668 8780
rect 42628 8634 42656 8774
rect 42616 8628 42668 8634
rect 42616 8570 42668 8576
rect 42524 8492 42576 8498
rect 42524 8434 42576 8440
rect 42720 8378 42748 9574
rect 42812 9450 42840 9676
rect 42800 9444 42852 9450
rect 42800 9386 42852 9392
rect 43076 9376 43128 9382
rect 43076 9318 43128 9324
rect 43088 9110 43116 9318
rect 43076 9104 43128 9110
rect 43076 9046 43128 9052
rect 42432 8356 42484 8362
rect 42432 8298 42484 8304
rect 42536 8350 42748 8378
rect 42432 7200 42484 7206
rect 42432 7142 42484 7148
rect 42444 6798 42472 7142
rect 42432 6792 42484 6798
rect 42432 6734 42484 6740
rect 42536 6662 42564 8350
rect 42616 7200 42668 7206
rect 42616 7142 42668 7148
rect 42524 6656 42576 6662
rect 42524 6598 42576 6604
rect 42340 6180 42392 6186
rect 42340 6122 42392 6128
rect 42536 5302 42564 6598
rect 42628 6118 42656 7142
rect 42708 6724 42760 6730
rect 42708 6666 42760 6672
rect 42720 6458 42748 6666
rect 42708 6452 42760 6458
rect 42708 6394 42760 6400
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42524 5296 42576 5302
rect 42524 5238 42576 5244
rect 42720 5234 42748 6394
rect 43076 5636 43128 5642
rect 43076 5578 43128 5584
rect 42708 5228 42760 5234
rect 42708 5170 42760 5176
rect 42720 4622 42748 5170
rect 43088 4826 43116 5578
rect 43076 4820 43128 4826
rect 43076 4762 43128 4768
rect 42708 4616 42760 4622
rect 42430 4584 42486 4593
rect 42708 4558 42760 4564
rect 42430 4519 42486 4528
rect 42340 4208 42392 4214
rect 42340 4150 42392 4156
rect 42248 3596 42300 3602
rect 42248 3538 42300 3544
rect 42352 3097 42380 4150
rect 42444 3942 42472 4519
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 42720 3738 42748 4558
rect 43180 4146 43208 11766
rect 43628 11552 43680 11558
rect 43628 11494 43680 11500
rect 43640 10674 43668 11494
rect 43628 10668 43680 10674
rect 43628 10610 43680 10616
rect 43260 9444 43312 9450
rect 43260 9386 43312 9392
rect 43272 7546 43300 9386
rect 43352 8968 43404 8974
rect 43352 8910 43404 8916
rect 43260 7540 43312 7546
rect 43260 7482 43312 7488
rect 43272 4214 43300 7482
rect 43364 6866 43392 8910
rect 43352 6860 43404 6866
rect 43352 6802 43404 6808
rect 43352 5704 43404 5710
rect 43352 5646 43404 5652
rect 43364 4826 43392 5646
rect 43732 5114 43760 12406
rect 43904 12096 43956 12102
rect 43904 12038 43956 12044
rect 43916 11898 43944 12038
rect 43904 11892 43956 11898
rect 43904 11834 43956 11840
rect 43812 11688 43864 11694
rect 43812 11630 43864 11636
rect 43824 11354 43852 11630
rect 43812 11348 43864 11354
rect 43812 11290 43864 11296
rect 43824 10810 43852 11290
rect 43812 10804 43864 10810
rect 43812 10746 43864 10752
rect 43904 10600 43956 10606
rect 43904 10542 43956 10548
rect 43916 10266 43944 10542
rect 43904 10260 43956 10266
rect 43904 10202 43956 10208
rect 44008 9654 44036 15302
rect 44282 15260 44590 15269
rect 44282 15258 44288 15260
rect 44344 15258 44368 15260
rect 44424 15258 44448 15260
rect 44504 15258 44528 15260
rect 44584 15258 44590 15260
rect 44344 15206 44346 15258
rect 44526 15206 44528 15258
rect 44282 15204 44288 15206
rect 44344 15204 44368 15206
rect 44424 15204 44448 15206
rect 44504 15204 44528 15206
rect 44584 15204 44590 15206
rect 44282 15195 44590 15204
rect 45112 15162 45140 18906
rect 45928 18896 45980 18902
rect 45928 18838 45980 18844
rect 45468 17536 45520 17542
rect 45468 17478 45520 17484
rect 45480 16658 45508 17478
rect 45468 16652 45520 16658
rect 45468 16594 45520 16600
rect 45940 16250 45968 18838
rect 46952 17626 46980 19110
rect 47124 18624 47176 18630
rect 47124 18566 47176 18572
rect 46860 17598 46980 17626
rect 46388 16652 46440 16658
rect 46388 16594 46440 16600
rect 45928 16244 45980 16250
rect 45928 16186 45980 16192
rect 45940 15706 45968 16186
rect 46400 15910 46428 16594
rect 46572 16584 46624 16590
rect 46572 16526 46624 16532
rect 46584 15978 46612 16526
rect 46572 15972 46624 15978
rect 46572 15914 46624 15920
rect 46388 15904 46440 15910
rect 46388 15846 46440 15852
rect 45928 15700 45980 15706
rect 45928 15642 45980 15648
rect 45100 15156 45152 15162
rect 45100 15098 45152 15104
rect 46296 15088 46348 15094
rect 46296 15030 46348 15036
rect 46480 15088 46532 15094
rect 46480 15030 46532 15036
rect 44180 14816 44232 14822
rect 44180 14758 44232 14764
rect 44916 14816 44968 14822
rect 44916 14758 44968 14764
rect 44192 14618 44220 14758
rect 44180 14612 44232 14618
rect 44180 14554 44232 14560
rect 44180 14272 44232 14278
rect 44180 14214 44232 14220
rect 44732 14272 44784 14278
rect 44732 14214 44784 14220
rect 44192 14074 44220 14214
rect 44282 14172 44590 14181
rect 44282 14170 44288 14172
rect 44344 14170 44368 14172
rect 44424 14170 44448 14172
rect 44504 14170 44528 14172
rect 44584 14170 44590 14172
rect 44344 14118 44346 14170
rect 44526 14118 44528 14170
rect 44282 14116 44288 14118
rect 44344 14116 44368 14118
rect 44424 14116 44448 14118
rect 44504 14116 44528 14118
rect 44584 14116 44590 14118
rect 44282 14107 44590 14116
rect 44180 14068 44232 14074
rect 44180 14010 44232 14016
rect 44088 13728 44140 13734
rect 44088 13670 44140 13676
rect 44100 13258 44128 13670
rect 44088 13252 44140 13258
rect 44088 13194 44140 13200
rect 44744 13190 44772 14214
rect 44928 13394 44956 14758
rect 46308 14074 46336 15030
rect 46492 14414 46520 15030
rect 46572 14816 46624 14822
rect 46572 14758 46624 14764
rect 46756 14816 46808 14822
rect 46756 14758 46808 14764
rect 46584 14618 46612 14758
rect 46572 14612 46624 14618
rect 46572 14554 46624 14560
rect 46768 14550 46796 14758
rect 46756 14544 46808 14550
rect 46756 14486 46808 14492
rect 46480 14408 46532 14414
rect 46480 14350 46532 14356
rect 45652 14068 45704 14074
rect 45652 14010 45704 14016
rect 46296 14068 46348 14074
rect 46296 14010 46348 14016
rect 44916 13388 44968 13394
rect 44916 13330 44968 13336
rect 44732 13184 44784 13190
rect 44732 13126 44784 13132
rect 44282 13084 44590 13093
rect 44282 13082 44288 13084
rect 44344 13082 44368 13084
rect 44424 13082 44448 13084
rect 44504 13082 44528 13084
rect 44584 13082 44590 13084
rect 44344 13030 44346 13082
rect 44526 13030 44528 13082
rect 44282 13028 44288 13030
rect 44344 13028 44368 13030
rect 44424 13028 44448 13030
rect 44504 13028 44528 13030
rect 44584 13028 44590 13030
rect 44282 13019 44590 13028
rect 44282 11996 44590 12005
rect 44282 11994 44288 11996
rect 44344 11994 44368 11996
rect 44424 11994 44448 11996
rect 44504 11994 44528 11996
rect 44584 11994 44590 11996
rect 44344 11942 44346 11994
rect 44526 11942 44528 11994
rect 44282 11940 44288 11942
rect 44344 11940 44368 11942
rect 44424 11940 44448 11942
rect 44504 11940 44528 11942
rect 44584 11940 44590 11942
rect 44282 11931 44590 11940
rect 44088 11280 44140 11286
rect 44088 11222 44140 11228
rect 44100 11014 44128 11222
rect 44180 11076 44232 11082
rect 44180 11018 44232 11024
rect 44088 11008 44140 11014
rect 44088 10950 44140 10956
rect 44100 10130 44128 10950
rect 44192 10810 44220 11018
rect 44744 11014 44772 13126
rect 45664 12306 45692 14010
rect 45928 13932 45980 13938
rect 45928 13874 45980 13880
rect 45836 13728 45888 13734
rect 45836 13670 45888 13676
rect 45848 13394 45876 13670
rect 45940 13530 45968 13874
rect 46296 13864 46348 13870
rect 46296 13806 46348 13812
rect 46308 13530 46336 13806
rect 46860 13802 46888 17598
rect 46940 17536 46992 17542
rect 46940 17478 46992 17484
rect 46952 16522 46980 17478
rect 47136 17202 47164 18566
rect 47320 17542 47348 19790
rect 47400 19712 47452 19718
rect 47400 19654 47452 19660
rect 47768 19712 47820 19718
rect 47768 19654 47820 19660
rect 47412 19378 47440 19654
rect 47780 19446 47808 19654
rect 47768 19440 47820 19446
rect 47768 19382 47820 19388
rect 47400 19372 47452 19378
rect 47400 19314 47452 19320
rect 47492 18760 47544 18766
rect 47492 18702 47544 18708
rect 47400 18216 47452 18222
rect 47400 18158 47452 18164
rect 47412 17882 47440 18158
rect 47400 17876 47452 17882
rect 47400 17818 47452 17824
rect 47308 17536 47360 17542
rect 47308 17478 47360 17484
rect 47320 17202 47348 17478
rect 47412 17338 47440 17818
rect 47504 17338 47532 18702
rect 48332 18426 48360 20266
rect 48516 20058 48544 21966
rect 50724 21690 50752 22510
rect 50804 22432 50856 22438
rect 50804 22374 50856 22380
rect 50816 21962 50844 22374
rect 50804 21956 50856 21962
rect 50804 21898 50856 21904
rect 51368 21894 51396 22510
rect 52000 22432 52052 22438
rect 52000 22374 52052 22380
rect 52368 22432 52420 22438
rect 52368 22374 52420 22380
rect 51504 22332 51812 22341
rect 51504 22330 51510 22332
rect 51566 22330 51590 22332
rect 51646 22330 51670 22332
rect 51726 22330 51750 22332
rect 51806 22330 51812 22332
rect 51566 22278 51568 22330
rect 51748 22278 51750 22330
rect 51504 22276 51510 22278
rect 51566 22276 51590 22278
rect 51646 22276 51670 22278
rect 51726 22276 51750 22278
rect 51806 22276 51812 22278
rect 51504 22267 51812 22276
rect 51356 21888 51408 21894
rect 51356 21830 51408 21836
rect 52012 21690 52040 22374
rect 52380 22030 52408 22374
rect 52368 22024 52420 22030
rect 52368 21966 52420 21972
rect 52460 22024 52512 22030
rect 52460 21966 52512 21972
rect 52184 21888 52236 21894
rect 52184 21830 52236 21836
rect 50712 21684 50764 21690
rect 50712 21626 50764 21632
rect 52000 21684 52052 21690
rect 52000 21626 52052 21632
rect 51354 21584 51410 21593
rect 51354 21519 51410 21528
rect 52092 21548 52144 21554
rect 51368 21486 51396 21519
rect 52092 21490 52144 21496
rect 51356 21480 51408 21486
rect 51356 21422 51408 21428
rect 51264 21344 51316 21350
rect 51264 21286 51316 21292
rect 51080 21072 51132 21078
rect 51080 21014 51132 21020
rect 49516 20936 49568 20942
rect 49516 20878 49568 20884
rect 48688 20868 48740 20874
rect 48688 20810 48740 20816
rect 48596 20392 48648 20398
rect 48596 20334 48648 20340
rect 48504 20052 48556 20058
rect 48504 19994 48556 20000
rect 48516 19514 48544 19994
rect 48608 19718 48636 20334
rect 48596 19712 48648 19718
rect 48596 19654 48648 19660
rect 48504 19508 48556 19514
rect 48504 19450 48556 19456
rect 48412 19236 48464 19242
rect 48412 19178 48464 19184
rect 48320 18420 48372 18426
rect 48320 18362 48372 18368
rect 47584 18352 47636 18358
rect 47584 18294 47636 18300
rect 47596 18086 47624 18294
rect 48320 18216 48372 18222
rect 48320 18158 48372 18164
rect 47584 18080 47636 18086
rect 47584 18022 47636 18028
rect 47676 18080 47728 18086
rect 47676 18022 47728 18028
rect 48228 18080 48280 18086
rect 48228 18022 48280 18028
rect 47400 17332 47452 17338
rect 47400 17274 47452 17280
rect 47492 17332 47544 17338
rect 47492 17274 47544 17280
rect 47124 17196 47176 17202
rect 47124 17138 47176 17144
rect 47308 17196 47360 17202
rect 47308 17138 47360 17144
rect 47492 16788 47544 16794
rect 47492 16730 47544 16736
rect 46940 16516 46992 16522
rect 46940 16458 46992 16464
rect 47400 15972 47452 15978
rect 47400 15914 47452 15920
rect 47032 15632 47084 15638
rect 47032 15574 47084 15580
rect 47044 14482 47072 15574
rect 47412 15366 47440 15914
rect 47504 15706 47532 16730
rect 47492 15700 47544 15706
rect 47492 15642 47544 15648
rect 47400 15360 47452 15366
rect 47400 15302 47452 15308
rect 47412 14958 47440 15302
rect 47400 14952 47452 14958
rect 47400 14894 47452 14900
rect 47032 14476 47084 14482
rect 47084 14436 47164 14464
rect 47032 14418 47084 14424
rect 46848 13796 46900 13802
rect 46848 13738 46900 13744
rect 45928 13524 45980 13530
rect 45928 13466 45980 13472
rect 46296 13524 46348 13530
rect 46296 13466 46348 13472
rect 45836 13388 45888 13394
rect 45836 13330 45888 13336
rect 45652 12300 45704 12306
rect 45652 12242 45704 12248
rect 45284 12232 45336 12238
rect 45284 12174 45336 12180
rect 45008 12164 45060 12170
rect 45008 12106 45060 12112
rect 45020 11898 45048 12106
rect 45296 11898 45324 12174
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 45008 11892 45060 11898
rect 45008 11834 45060 11840
rect 45284 11892 45336 11898
rect 45284 11834 45336 11840
rect 45572 11150 45600 12038
rect 45664 11898 45692 12242
rect 46020 12232 46072 12238
rect 46020 12174 46072 12180
rect 45652 11892 45704 11898
rect 45652 11834 45704 11840
rect 46032 11558 46060 12174
rect 46664 12096 46716 12102
rect 46664 12038 46716 12044
rect 46848 12096 46900 12102
rect 46848 12038 46900 12044
rect 46388 11892 46440 11898
rect 46388 11834 46440 11840
rect 46020 11552 46072 11558
rect 46020 11494 46072 11500
rect 45560 11144 45612 11150
rect 45560 11086 45612 11092
rect 44732 11008 44784 11014
rect 44732 10950 44784 10956
rect 44282 10908 44590 10917
rect 44282 10906 44288 10908
rect 44344 10906 44368 10908
rect 44424 10906 44448 10908
rect 44504 10906 44528 10908
rect 44584 10906 44590 10908
rect 44344 10854 44346 10906
rect 44526 10854 44528 10906
rect 44282 10852 44288 10854
rect 44344 10852 44368 10854
rect 44424 10852 44448 10854
rect 44504 10852 44528 10854
rect 44584 10852 44590 10854
rect 44282 10843 44590 10852
rect 44180 10804 44232 10810
rect 44180 10746 44232 10752
rect 44744 10470 44772 10950
rect 44732 10464 44784 10470
rect 44732 10406 44784 10412
rect 44744 10266 44772 10406
rect 44732 10260 44784 10266
rect 45836 10260 45888 10266
rect 44784 10220 44864 10248
rect 44732 10202 44784 10208
rect 44088 10124 44140 10130
rect 44088 10066 44140 10072
rect 44282 9820 44590 9829
rect 44282 9818 44288 9820
rect 44344 9818 44368 9820
rect 44424 9818 44448 9820
rect 44504 9818 44528 9820
rect 44584 9818 44590 9820
rect 44344 9766 44346 9818
rect 44526 9766 44528 9818
rect 44282 9764 44288 9766
rect 44344 9764 44368 9766
rect 44424 9764 44448 9766
rect 44504 9764 44528 9766
rect 44584 9764 44590 9766
rect 44282 9755 44590 9764
rect 43996 9648 44048 9654
rect 43996 9590 44048 9596
rect 44640 9580 44692 9586
rect 44640 9522 44692 9528
rect 44180 9512 44232 9518
rect 44180 9454 44232 9460
rect 43812 9376 43864 9382
rect 43812 9318 43864 9324
rect 43824 9042 43852 9318
rect 43812 9036 43864 9042
rect 43812 8978 43864 8984
rect 43904 8832 43956 8838
rect 43904 8774 43956 8780
rect 43916 8634 43944 8774
rect 43904 8628 43956 8634
rect 43904 8570 43956 8576
rect 44192 8362 44220 9454
rect 44282 8732 44590 8741
rect 44282 8730 44288 8732
rect 44344 8730 44368 8732
rect 44424 8730 44448 8732
rect 44504 8730 44528 8732
rect 44584 8730 44590 8732
rect 44344 8678 44346 8730
rect 44526 8678 44528 8730
rect 44282 8676 44288 8678
rect 44344 8676 44368 8678
rect 44424 8676 44448 8678
rect 44504 8676 44528 8678
rect 44584 8676 44590 8678
rect 44282 8667 44590 8676
rect 44180 8356 44232 8362
rect 44180 8298 44232 8304
rect 44548 8356 44600 8362
rect 44548 8298 44600 8304
rect 44088 8084 44140 8090
rect 44088 8026 44140 8032
rect 43996 7812 44048 7818
rect 43996 7754 44048 7760
rect 43904 7744 43956 7750
rect 43904 7686 43956 7692
rect 43916 7546 43944 7686
rect 44008 7546 44036 7754
rect 44100 7546 44128 8026
rect 44560 7750 44588 8298
rect 44180 7744 44232 7750
rect 44180 7686 44232 7692
rect 44548 7744 44600 7750
rect 44548 7686 44600 7692
rect 44192 7546 44220 7686
rect 44282 7644 44590 7653
rect 44282 7642 44288 7644
rect 44344 7642 44368 7644
rect 44424 7642 44448 7644
rect 44504 7642 44528 7644
rect 44584 7642 44590 7644
rect 44344 7590 44346 7642
rect 44526 7590 44528 7642
rect 44282 7588 44288 7590
rect 44344 7588 44368 7590
rect 44424 7588 44448 7590
rect 44504 7588 44528 7590
rect 44584 7588 44590 7590
rect 44282 7579 44590 7588
rect 43904 7540 43956 7546
rect 43904 7482 43956 7488
rect 43996 7540 44048 7546
rect 43996 7482 44048 7488
rect 44088 7540 44140 7546
rect 44088 7482 44140 7488
rect 44180 7540 44232 7546
rect 44180 7482 44232 7488
rect 44456 7540 44508 7546
rect 44456 7482 44508 7488
rect 44468 7002 44496 7482
rect 44456 6996 44508 7002
rect 44456 6938 44508 6944
rect 44468 6662 44496 6938
rect 44456 6656 44508 6662
rect 44456 6598 44508 6604
rect 44282 6556 44590 6565
rect 44282 6554 44288 6556
rect 44344 6554 44368 6556
rect 44424 6554 44448 6556
rect 44504 6554 44528 6556
rect 44584 6554 44590 6556
rect 44344 6502 44346 6554
rect 44526 6502 44528 6554
rect 44282 6500 44288 6502
rect 44344 6500 44368 6502
rect 44424 6500 44448 6502
rect 44504 6500 44528 6502
rect 44584 6500 44590 6502
rect 44282 6491 44590 6500
rect 43904 6248 43956 6254
rect 43904 6190 43956 6196
rect 43916 5574 43944 6190
rect 43996 5704 44048 5710
rect 43996 5646 44048 5652
rect 44180 5704 44232 5710
rect 44180 5646 44232 5652
rect 43812 5568 43864 5574
rect 43812 5510 43864 5516
rect 43904 5568 43956 5574
rect 43904 5510 43956 5516
rect 43824 5302 43852 5510
rect 43812 5296 43864 5302
rect 43812 5238 43864 5244
rect 43732 5086 43852 5114
rect 43352 4820 43404 4826
rect 43352 4762 43404 4768
rect 43628 4480 43680 4486
rect 43628 4422 43680 4428
rect 43640 4282 43668 4422
rect 43628 4276 43680 4282
rect 43628 4218 43680 4224
rect 43260 4208 43312 4214
rect 43260 4150 43312 4156
rect 43168 4140 43220 4146
rect 43168 4082 43220 4088
rect 43536 4140 43588 4146
rect 43536 4082 43588 4088
rect 42800 4072 42852 4078
rect 42892 4072 42944 4078
rect 42800 4014 42852 4020
rect 42890 4040 42892 4049
rect 42984 4072 43036 4078
rect 42944 4040 42946 4049
rect 42708 3732 42760 3738
rect 42708 3674 42760 3680
rect 42338 3088 42394 3097
rect 42338 3023 42394 3032
rect 42812 2961 42840 4014
rect 42984 4014 43036 4020
rect 42890 3975 42946 3984
rect 42904 3097 42932 3975
rect 42890 3088 42946 3097
rect 42890 3023 42946 3032
rect 42798 2952 42854 2961
rect 42798 2887 42854 2896
rect 41880 2848 41932 2854
rect 41880 2790 41932 2796
rect 41972 2848 42024 2854
rect 41972 2790 42024 2796
rect 42996 2774 43024 4014
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 43260 3936 43312 3942
rect 43260 3878 43312 3884
rect 43352 3936 43404 3942
rect 43352 3878 43404 3884
rect 43088 3738 43116 3878
rect 43076 3732 43128 3738
rect 43076 3674 43128 3680
rect 42904 2746 43024 2774
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42352 870 42472 898
rect 42352 800 42380 870
rect 40880 734 41184 762
rect 41234 0 41290 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42444 762 42472 870
rect 42628 762 42656 2450
rect 42904 800 42932 2746
rect 43272 2446 43300 3878
rect 43364 3534 43392 3878
rect 43352 3528 43404 3534
rect 43352 3470 43404 3476
rect 43548 3194 43576 4082
rect 43720 3936 43772 3942
rect 43720 3878 43772 3884
rect 43732 3398 43760 3878
rect 43824 3505 43852 5086
rect 43916 4690 43944 5510
rect 44008 5030 44036 5646
rect 44088 5568 44140 5574
rect 44088 5510 44140 5516
rect 43996 5024 44048 5030
rect 43996 4966 44048 4972
rect 44008 4826 44036 4966
rect 43996 4820 44048 4826
rect 43996 4762 44048 4768
rect 44100 4690 44128 5510
rect 43904 4684 43956 4690
rect 43904 4626 43956 4632
rect 44088 4684 44140 4690
rect 44088 4626 44140 4632
rect 44192 4622 44220 5646
rect 44282 5468 44590 5477
rect 44282 5466 44288 5468
rect 44344 5466 44368 5468
rect 44424 5466 44448 5468
rect 44504 5466 44528 5468
rect 44584 5466 44590 5468
rect 44344 5414 44346 5466
rect 44526 5414 44528 5466
rect 44282 5412 44288 5414
rect 44344 5412 44368 5414
rect 44424 5412 44448 5414
rect 44504 5412 44528 5414
rect 44584 5412 44590 5414
rect 44282 5403 44590 5412
rect 44652 4690 44680 9522
rect 44732 8900 44784 8906
rect 44732 8842 44784 8848
rect 44744 7954 44772 8842
rect 44836 8634 44864 10220
rect 45836 10202 45888 10208
rect 44916 9648 44968 9654
rect 44916 9590 44968 9596
rect 44928 8974 44956 9590
rect 45468 9512 45520 9518
rect 45468 9454 45520 9460
rect 44916 8968 44968 8974
rect 44916 8910 44968 8916
rect 44824 8628 44876 8634
rect 44824 8570 44876 8576
rect 44732 7948 44784 7954
rect 44732 7890 44784 7896
rect 44744 6662 44772 7890
rect 44836 6866 44864 8570
rect 45480 8294 45508 9454
rect 45848 9042 45876 10202
rect 46400 9654 46428 11834
rect 46676 10674 46704 12038
rect 46860 11286 46888 12038
rect 47032 11756 47084 11762
rect 47032 11698 47084 11704
rect 46940 11552 46992 11558
rect 46940 11494 46992 11500
rect 46848 11280 46900 11286
rect 46848 11222 46900 11228
rect 46952 11150 46980 11494
rect 46940 11144 46992 11150
rect 46940 11086 46992 11092
rect 47044 10810 47072 11698
rect 47136 11506 47164 14436
rect 47412 13870 47440 14894
rect 47492 14408 47544 14414
rect 47492 14350 47544 14356
rect 47504 13938 47532 14350
rect 47492 13932 47544 13938
rect 47492 13874 47544 13880
rect 47400 13864 47452 13870
rect 47400 13806 47452 13812
rect 47216 13388 47268 13394
rect 47216 13330 47268 13336
rect 47228 11898 47256 13330
rect 47412 13190 47440 13806
rect 47400 13184 47452 13190
rect 47400 13126 47452 13132
rect 47596 12434 47624 18022
rect 47688 17746 47716 18022
rect 47676 17740 47728 17746
rect 47676 17682 47728 17688
rect 47688 13462 47716 17682
rect 48136 17672 48188 17678
rect 48136 17614 48188 17620
rect 47952 17536 48004 17542
rect 47952 17478 48004 17484
rect 48044 17536 48096 17542
rect 48044 17478 48096 17484
rect 47964 16250 47992 17478
rect 47952 16244 48004 16250
rect 47952 16186 48004 16192
rect 47860 15700 47912 15706
rect 47860 15642 47912 15648
rect 47872 14482 47900 15642
rect 47860 14476 47912 14482
rect 47860 14418 47912 14424
rect 47676 13456 47728 13462
rect 47676 13398 47728 13404
rect 47768 12980 47820 12986
rect 47768 12922 47820 12928
rect 47504 12406 47624 12434
rect 47400 12096 47452 12102
rect 47400 12038 47452 12044
rect 47412 11898 47440 12038
rect 47216 11892 47268 11898
rect 47216 11834 47268 11840
rect 47400 11892 47452 11898
rect 47400 11834 47452 11840
rect 47228 11694 47256 11834
rect 47308 11756 47360 11762
rect 47308 11698 47360 11704
rect 47216 11688 47268 11694
rect 47216 11630 47268 11636
rect 47320 11506 47348 11698
rect 47136 11478 47348 11506
rect 47124 11212 47176 11218
rect 47124 11154 47176 11160
rect 47216 11212 47268 11218
rect 47320 11200 47348 11478
rect 47504 11234 47532 12406
rect 47780 12374 47808 12922
rect 47872 12442 47900 14418
rect 48056 12986 48084 17478
rect 48148 16794 48176 17614
rect 48240 17338 48268 18022
rect 48228 17332 48280 17338
rect 48228 17274 48280 17280
rect 48332 17270 48360 18158
rect 48320 17264 48372 17270
rect 48320 17206 48372 17212
rect 48136 16788 48188 16794
rect 48136 16730 48188 16736
rect 48332 16658 48360 17206
rect 48320 16652 48372 16658
rect 48320 16594 48372 16600
rect 48320 16448 48372 16454
rect 48320 16390 48372 16396
rect 48332 16114 48360 16390
rect 48320 16108 48372 16114
rect 48320 16050 48372 16056
rect 48424 15638 48452 19178
rect 48516 18970 48544 19450
rect 48608 19378 48636 19654
rect 48700 19378 48728 20810
rect 48780 20800 48832 20806
rect 48780 20742 48832 20748
rect 48792 20398 48820 20742
rect 49528 20602 49556 20878
rect 51092 20806 51120 21014
rect 51276 20942 51304 21286
rect 51368 21010 51396 21422
rect 51504 21244 51812 21253
rect 51504 21242 51510 21244
rect 51566 21242 51590 21244
rect 51646 21242 51670 21244
rect 51726 21242 51750 21244
rect 51806 21242 51812 21244
rect 51566 21190 51568 21242
rect 51748 21190 51750 21242
rect 51504 21188 51510 21190
rect 51566 21188 51590 21190
rect 51646 21188 51670 21190
rect 51726 21188 51750 21190
rect 51806 21188 51812 21190
rect 51504 21179 51812 21188
rect 51356 21004 51408 21010
rect 51356 20946 51408 20952
rect 52000 21004 52052 21010
rect 52000 20946 52052 20952
rect 51264 20936 51316 20942
rect 52012 20913 52040 20946
rect 51264 20878 51316 20884
rect 51998 20904 52054 20913
rect 51998 20839 52054 20848
rect 49700 20800 49752 20806
rect 49700 20742 49752 20748
rect 50160 20800 50212 20806
rect 50160 20742 50212 20748
rect 51080 20800 51132 20806
rect 51080 20742 51132 20748
rect 49516 20596 49568 20602
rect 49516 20538 49568 20544
rect 48780 20392 48832 20398
rect 48780 20334 48832 20340
rect 48596 19372 48648 19378
rect 48596 19314 48648 19320
rect 48688 19372 48740 19378
rect 48688 19314 48740 19320
rect 48504 18964 48556 18970
rect 48504 18906 48556 18912
rect 48688 18420 48740 18426
rect 48688 18362 48740 18368
rect 48504 18080 48556 18086
rect 48504 18022 48556 18028
rect 48516 17746 48544 18022
rect 48700 17746 48728 18362
rect 48792 18358 48820 20334
rect 49332 20256 49384 20262
rect 49332 20198 49384 20204
rect 49344 19786 49372 20198
rect 49712 20058 49740 20742
rect 50172 20398 50200 20742
rect 49976 20392 50028 20398
rect 49976 20334 50028 20340
rect 50160 20392 50212 20398
rect 50160 20334 50212 20340
rect 50436 20392 50488 20398
rect 50436 20334 50488 20340
rect 49700 20052 49752 20058
rect 49700 19994 49752 20000
rect 49608 19848 49660 19854
rect 49608 19790 49660 19796
rect 49332 19780 49384 19786
rect 49332 19722 49384 19728
rect 48780 18352 48832 18358
rect 48780 18294 48832 18300
rect 49332 18352 49384 18358
rect 49332 18294 49384 18300
rect 49344 17746 49372 18294
rect 49620 18222 49648 19790
rect 49988 18630 50016 20334
rect 50068 20256 50120 20262
rect 50068 20198 50120 20204
rect 49976 18624 50028 18630
rect 49976 18566 50028 18572
rect 49608 18216 49660 18222
rect 49608 18158 49660 18164
rect 48504 17740 48556 17746
rect 48504 17682 48556 17688
rect 48688 17740 48740 17746
rect 48688 17682 48740 17688
rect 49332 17740 49384 17746
rect 49332 17682 49384 17688
rect 49056 17672 49108 17678
rect 49344 17649 49372 17682
rect 49056 17614 49108 17620
rect 49330 17640 49386 17649
rect 49068 16522 49096 17614
rect 49330 17575 49386 17584
rect 49988 17338 50016 18566
rect 50080 17678 50108 20198
rect 50448 19786 50476 20334
rect 50436 19780 50488 19786
rect 50436 19722 50488 19728
rect 50528 19304 50580 19310
rect 50528 19246 50580 19252
rect 50540 18970 50568 19246
rect 50528 18964 50580 18970
rect 50528 18906 50580 18912
rect 50712 18828 50764 18834
rect 50712 18770 50764 18776
rect 50068 17672 50120 17678
rect 50068 17614 50120 17620
rect 50160 17536 50212 17542
rect 50160 17478 50212 17484
rect 49516 17332 49568 17338
rect 49516 17274 49568 17280
rect 49976 17332 50028 17338
rect 49976 17274 50028 17280
rect 49148 17128 49200 17134
rect 49148 17070 49200 17076
rect 49056 16516 49108 16522
rect 49056 16458 49108 16464
rect 49160 16402 49188 17070
rect 49068 16374 49188 16402
rect 49068 15910 49096 16374
rect 49056 15904 49108 15910
rect 49056 15846 49108 15852
rect 48412 15632 48464 15638
rect 48412 15574 48464 15580
rect 48424 14482 48452 15574
rect 48412 14476 48464 14482
rect 48412 14418 48464 14424
rect 48228 14272 48280 14278
rect 48228 14214 48280 14220
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 48412 14272 48464 14278
rect 48412 14214 48464 14220
rect 48780 14272 48832 14278
rect 48780 14214 48832 14220
rect 48964 14272 49016 14278
rect 48964 14214 49016 14220
rect 48240 14074 48268 14214
rect 48228 14068 48280 14074
rect 48228 14010 48280 14016
rect 48044 12980 48096 12986
rect 48044 12922 48096 12928
rect 47952 12776 48004 12782
rect 47952 12718 48004 12724
rect 47860 12436 47912 12442
rect 47860 12378 47912 12384
rect 47768 12368 47820 12374
rect 47768 12310 47820 12316
rect 47768 12096 47820 12102
rect 47768 12038 47820 12044
rect 47584 11688 47636 11694
rect 47584 11630 47636 11636
rect 47596 11354 47624 11630
rect 47584 11348 47636 11354
rect 47584 11290 47636 11296
rect 47268 11172 47348 11200
rect 47412 11206 47532 11234
rect 47216 11154 47268 11160
rect 47136 10810 47164 11154
rect 47032 10804 47084 10810
rect 47032 10746 47084 10752
rect 47124 10804 47176 10810
rect 47124 10746 47176 10752
rect 46664 10668 46716 10674
rect 46664 10610 46716 10616
rect 47228 10266 47256 11154
rect 47216 10260 47268 10266
rect 47216 10202 47268 10208
rect 46388 9648 46440 9654
rect 46388 9590 46440 9596
rect 46296 9376 46348 9382
rect 46296 9318 46348 9324
rect 46664 9376 46716 9382
rect 46664 9318 46716 9324
rect 46308 9042 46336 9318
rect 46676 9042 46704 9318
rect 47412 9178 47440 11206
rect 47492 11144 47544 11150
rect 47492 11086 47544 11092
rect 47504 10606 47532 11086
rect 47492 10600 47544 10606
rect 47492 10542 47544 10548
rect 47400 9172 47452 9178
rect 47400 9114 47452 9120
rect 45836 9036 45888 9042
rect 45836 8978 45888 8984
rect 46296 9036 46348 9042
rect 46296 8978 46348 8984
rect 46664 9036 46716 9042
rect 46664 8978 46716 8984
rect 45468 8288 45520 8294
rect 45848 8242 45876 8978
rect 46676 8922 46704 8978
rect 46492 8906 46704 8922
rect 46492 8900 46716 8906
rect 46492 8894 46664 8900
rect 46492 8634 46520 8894
rect 46664 8842 46716 8848
rect 46572 8832 46624 8838
rect 46572 8774 46624 8780
rect 46584 8634 46612 8774
rect 47412 8634 47440 9114
rect 46480 8628 46532 8634
rect 46480 8570 46532 8576
rect 46572 8628 46624 8634
rect 46572 8570 46624 8576
rect 47400 8628 47452 8634
rect 47400 8570 47452 8576
rect 47596 8498 47624 11290
rect 47676 9580 47728 9586
rect 47676 9522 47728 9528
rect 47584 8492 47636 8498
rect 47584 8434 47636 8440
rect 47216 8424 47268 8430
rect 47216 8366 47268 8372
rect 45468 8230 45520 8236
rect 45480 8022 45508 8230
rect 45664 8214 45876 8242
rect 45664 8022 45692 8214
rect 47228 8090 47256 8366
rect 47216 8084 47268 8090
rect 47216 8026 47268 8032
rect 45468 8016 45520 8022
rect 45468 7958 45520 7964
rect 45652 8016 45704 8022
rect 45652 7958 45704 7964
rect 44916 7948 44968 7954
rect 44916 7890 44968 7896
rect 45560 7948 45612 7954
rect 45560 7890 45612 7896
rect 44928 7546 44956 7890
rect 45572 7546 45600 7890
rect 44916 7540 44968 7546
rect 44916 7482 44968 7488
rect 45560 7540 45612 7546
rect 45560 7482 45612 7488
rect 45664 7478 45692 7958
rect 46388 7948 46440 7954
rect 46388 7890 46440 7896
rect 45928 7880 45980 7886
rect 45928 7822 45980 7828
rect 45940 7750 45968 7822
rect 45928 7744 45980 7750
rect 45928 7686 45980 7692
rect 46296 7540 46348 7546
rect 46296 7482 46348 7488
rect 45652 7472 45704 7478
rect 45704 7432 45784 7460
rect 45652 7414 45704 7420
rect 45192 7404 45244 7410
rect 45192 7346 45244 7352
rect 44824 6860 44876 6866
rect 44824 6802 44876 6808
rect 45204 6730 45232 7346
rect 45192 6724 45244 6730
rect 45192 6666 45244 6672
rect 44732 6656 44784 6662
rect 44732 6598 44784 6604
rect 44916 6248 44968 6254
rect 44916 6190 44968 6196
rect 44928 5914 44956 6190
rect 44916 5908 44968 5914
rect 44916 5850 44968 5856
rect 44730 5672 44786 5681
rect 44730 5607 44786 5616
rect 44640 4684 44692 4690
rect 44640 4626 44692 4632
rect 44180 4616 44232 4622
rect 44180 4558 44232 4564
rect 44088 4072 44140 4078
rect 44088 4014 44140 4020
rect 44100 3670 44128 4014
rect 44088 3664 44140 3670
rect 44088 3606 44140 3612
rect 43810 3496 43866 3505
rect 43810 3431 43866 3440
rect 43904 3460 43956 3466
rect 43904 3402 43956 3408
rect 43720 3392 43772 3398
rect 43720 3334 43772 3340
rect 43812 3392 43864 3398
rect 43812 3334 43864 3340
rect 43824 3194 43852 3334
rect 43916 3194 43944 3402
rect 43536 3188 43588 3194
rect 43536 3130 43588 3136
rect 43812 3188 43864 3194
rect 43812 3130 43864 3136
rect 43904 3188 43956 3194
rect 43904 3130 43956 3136
rect 43996 2984 44048 2990
rect 43996 2926 44048 2932
rect 43260 2440 43312 2446
rect 43260 2382 43312 2388
rect 43904 2372 43956 2378
rect 43904 2314 43956 2320
rect 43456 870 43576 898
rect 43456 800 43484 870
rect 42444 734 42656 762
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 43548 762 43576 870
rect 43916 762 43944 2314
rect 44008 800 44036 2926
rect 44100 2514 44128 3606
rect 44192 3602 44220 4558
rect 44282 4380 44590 4389
rect 44282 4378 44288 4380
rect 44344 4378 44368 4380
rect 44424 4378 44448 4380
rect 44504 4378 44528 4380
rect 44584 4378 44590 4380
rect 44344 4326 44346 4378
rect 44526 4326 44528 4378
rect 44282 4324 44288 4326
rect 44344 4324 44368 4326
rect 44424 4324 44448 4326
rect 44504 4324 44528 4326
rect 44584 4324 44590 4326
rect 44282 4315 44590 4324
rect 44744 4060 44772 5607
rect 44916 5364 44968 5370
rect 44916 5306 44968 5312
rect 44928 4758 44956 5306
rect 45204 5030 45232 6666
rect 45468 6656 45520 6662
rect 45468 6598 45520 6604
rect 45480 6458 45508 6598
rect 45468 6452 45520 6458
rect 45388 6412 45468 6440
rect 45388 5710 45416 6412
rect 45468 6394 45520 6400
rect 45560 6316 45612 6322
rect 45560 6258 45612 6264
rect 45468 6112 45520 6118
rect 45468 6054 45520 6060
rect 45376 5704 45428 5710
rect 45376 5646 45428 5652
rect 45192 5024 45244 5030
rect 45192 4966 45244 4972
rect 44916 4752 44968 4758
rect 44916 4694 44968 4700
rect 45204 4282 45232 4966
rect 45388 4706 45416 5646
rect 45480 5302 45508 6054
rect 45572 5370 45600 6258
rect 45652 6112 45704 6118
rect 45652 6054 45704 6060
rect 45664 5914 45692 6054
rect 45652 5908 45704 5914
rect 45652 5850 45704 5856
rect 45560 5364 45612 5370
rect 45560 5306 45612 5312
rect 45652 5364 45704 5370
rect 45652 5306 45704 5312
rect 45468 5296 45520 5302
rect 45468 5238 45520 5244
rect 45664 4842 45692 5306
rect 45480 4814 45692 4842
rect 45480 4758 45508 4814
rect 45296 4678 45416 4706
rect 45468 4752 45520 4758
rect 45756 4706 45784 7432
rect 46112 6860 46164 6866
rect 46112 6802 46164 6808
rect 46124 6390 46152 6802
rect 46308 6798 46336 7482
rect 46296 6792 46348 6798
rect 46296 6734 46348 6740
rect 46112 6384 46164 6390
rect 46112 6326 46164 6332
rect 45836 5704 45888 5710
rect 45836 5646 45888 5652
rect 45848 5370 45876 5646
rect 45836 5364 45888 5370
rect 45836 5306 45888 5312
rect 46204 5160 46256 5166
rect 46204 5102 46256 5108
rect 46216 4826 46244 5102
rect 46204 4820 46256 4826
rect 46204 4762 46256 4768
rect 45468 4694 45520 4700
rect 45664 4690 45784 4706
rect 46400 4690 46428 7890
rect 47596 7886 47624 8434
rect 47584 7880 47636 7886
rect 47584 7822 47636 7828
rect 46848 7744 46900 7750
rect 46848 7686 46900 7692
rect 46572 7336 46624 7342
rect 46572 7278 46624 7284
rect 46584 7002 46612 7278
rect 46572 6996 46624 7002
rect 46572 6938 46624 6944
rect 46860 5370 46888 7686
rect 46940 6656 46992 6662
rect 46940 6598 46992 6604
rect 46952 6186 46980 6598
rect 47124 6248 47176 6254
rect 47124 6190 47176 6196
rect 46940 6180 46992 6186
rect 46940 6122 46992 6128
rect 46952 5914 46980 6122
rect 46940 5908 46992 5914
rect 46940 5850 46992 5856
rect 46848 5364 46900 5370
rect 46848 5306 46900 5312
rect 46952 4690 46980 5850
rect 47136 5098 47164 6190
rect 47124 5092 47176 5098
rect 47124 5034 47176 5040
rect 47032 5024 47084 5030
rect 47032 4966 47084 4972
rect 45560 4684 45612 4690
rect 45192 4276 45244 4282
rect 45192 4218 45244 4224
rect 44468 4032 44772 4060
rect 44468 3602 44496 4032
rect 44824 4004 44876 4010
rect 44824 3946 44876 3952
rect 44836 3738 44864 3946
rect 44824 3732 44876 3738
rect 44824 3674 44876 3680
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 44456 3596 44508 3602
rect 44456 3538 44508 3544
rect 45204 3534 45232 4218
rect 45296 4010 45324 4678
rect 45560 4626 45612 4632
rect 45652 4684 45784 4690
rect 45704 4678 45784 4684
rect 46388 4684 46440 4690
rect 45652 4626 45704 4632
rect 46388 4626 46440 4632
rect 46940 4684 46992 4690
rect 46940 4626 46992 4632
rect 45376 4616 45428 4622
rect 45428 4576 45508 4604
rect 45376 4558 45428 4564
rect 45480 4026 45508 4576
rect 45572 4146 45600 4626
rect 46020 4616 46072 4622
rect 46020 4558 46072 4564
rect 45652 4480 45704 4486
rect 45652 4422 45704 4428
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 45284 4004 45336 4010
rect 45480 3998 45600 4026
rect 45284 3946 45336 3952
rect 44824 3528 44876 3534
rect 44824 3470 44876 3476
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44192 2650 44220 3334
rect 44282 3292 44590 3301
rect 44282 3290 44288 3292
rect 44344 3290 44368 3292
rect 44424 3290 44448 3292
rect 44504 3290 44528 3292
rect 44584 3290 44590 3292
rect 44344 3238 44346 3290
rect 44526 3238 44528 3290
rect 44282 3236 44288 3238
rect 44344 3236 44368 3238
rect 44424 3236 44448 3238
rect 44504 3236 44528 3238
rect 44584 3236 44590 3238
rect 44282 3227 44590 3236
rect 44836 3058 44864 3470
rect 45572 3194 45600 3998
rect 45560 3188 45612 3194
rect 45560 3130 45612 3136
rect 45100 3120 45152 3126
rect 45284 3120 45336 3126
rect 45152 3080 45284 3108
rect 45100 3062 45152 3068
rect 45284 3062 45336 3068
rect 44824 3052 44876 3058
rect 44824 2994 44876 3000
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 44732 2916 44784 2922
rect 44732 2858 44784 2864
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 44088 2508 44140 2514
rect 44088 2450 44140 2456
rect 44282 2204 44590 2213
rect 44282 2202 44288 2204
rect 44344 2202 44368 2204
rect 44424 2202 44448 2204
rect 44504 2202 44528 2204
rect 44584 2202 44590 2204
rect 44344 2150 44346 2202
rect 44526 2150 44528 2202
rect 44282 2148 44288 2150
rect 44344 2148 44368 2150
rect 44424 2148 44448 2150
rect 44504 2148 44528 2150
rect 44584 2148 44590 2150
rect 44282 2139 44590 2148
rect 44744 1442 44772 2858
rect 44560 1414 44772 1442
rect 44560 800 44588 1414
rect 45112 800 45140 2926
rect 45664 2774 45692 4422
rect 45836 4208 45888 4214
rect 45836 4150 45888 4156
rect 45848 3738 45876 4150
rect 46032 4078 46060 4558
rect 46480 4140 46532 4146
rect 46480 4082 46532 4088
rect 46020 4072 46072 4078
rect 46020 4014 46072 4020
rect 46492 3738 46520 4082
rect 45836 3732 45888 3738
rect 45836 3674 45888 3680
rect 46480 3732 46532 3738
rect 46480 3674 46532 3680
rect 46754 3632 46810 3641
rect 46754 3567 46810 3576
rect 46478 3496 46534 3505
rect 46478 3431 46534 3440
rect 46386 3088 46442 3097
rect 46492 3058 46520 3431
rect 46768 3058 46796 3567
rect 47044 3194 47072 4966
rect 47136 4554 47164 5034
rect 47216 5024 47268 5030
rect 47216 4966 47268 4972
rect 47228 4622 47256 4966
rect 47216 4616 47268 4622
rect 47216 4558 47268 4564
rect 47124 4548 47176 4554
rect 47124 4490 47176 4496
rect 47582 4040 47638 4049
rect 47582 3975 47638 3984
rect 47400 3732 47452 3738
rect 47400 3674 47452 3680
rect 47032 3188 47084 3194
rect 47032 3130 47084 3136
rect 46386 3023 46388 3032
rect 46440 3023 46442 3032
rect 46480 3052 46532 3058
rect 46388 2994 46440 3000
rect 46480 2994 46532 3000
rect 46756 3052 46808 3058
rect 46756 2994 46808 3000
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46860 2774 46888 2926
rect 45572 2746 45692 2774
rect 46768 2746 46888 2774
rect 45572 2650 45600 2746
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 45652 2508 45704 2514
rect 45652 2450 45704 2456
rect 45664 800 45692 2450
rect 46204 2372 46256 2378
rect 46204 2314 46256 2320
rect 46216 800 46244 2314
rect 46768 800 46796 2746
rect 47136 2446 47164 2994
rect 47412 2650 47440 3674
rect 47596 3602 47624 3975
rect 47688 3942 47716 9522
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47780 3738 47808 12038
rect 47872 11200 47900 12378
rect 47964 11558 47992 12718
rect 48332 12238 48360 14214
rect 48424 13394 48452 14214
rect 48792 14074 48820 14214
rect 48780 14068 48832 14074
rect 48780 14010 48832 14016
rect 48780 13932 48832 13938
rect 48780 13874 48832 13880
rect 48792 13530 48820 13874
rect 48780 13524 48832 13530
rect 48780 13466 48832 13472
rect 48412 13388 48464 13394
rect 48412 13330 48464 13336
rect 48872 12640 48924 12646
rect 48872 12582 48924 12588
rect 48884 12238 48912 12582
rect 48320 12232 48372 12238
rect 48320 12174 48372 12180
rect 48872 12232 48924 12238
rect 48872 12174 48924 12180
rect 48976 12170 49004 14214
rect 48964 12164 49016 12170
rect 48964 12106 49016 12112
rect 48228 12096 48280 12102
rect 48228 12038 48280 12044
rect 47952 11552 48004 11558
rect 47952 11494 48004 11500
rect 48240 11286 48268 12038
rect 48228 11280 48280 11286
rect 48228 11222 48280 11228
rect 48976 11218 49004 12106
rect 49068 11218 49096 15846
rect 49240 14952 49292 14958
rect 49240 14894 49292 14900
rect 49252 14618 49280 14894
rect 49240 14612 49292 14618
rect 49240 14554 49292 14560
rect 49148 14408 49200 14414
rect 49148 14350 49200 14356
rect 49160 13530 49188 14350
rect 49148 13524 49200 13530
rect 49148 13466 49200 13472
rect 49160 11558 49188 13466
rect 49332 12436 49384 12442
rect 49332 12378 49384 12384
rect 49344 11898 49372 12378
rect 49332 11892 49384 11898
rect 49332 11834 49384 11840
rect 49148 11552 49200 11558
rect 49148 11494 49200 11500
rect 47952 11212 48004 11218
rect 47872 11172 47952 11200
rect 47872 8634 47900 11172
rect 47952 11154 48004 11160
rect 48964 11212 49016 11218
rect 48964 11154 49016 11160
rect 49056 11212 49108 11218
rect 49056 11154 49108 11160
rect 48872 11144 48924 11150
rect 48872 11086 48924 11092
rect 48884 10674 48912 11086
rect 48872 10668 48924 10674
rect 48872 10610 48924 10616
rect 49068 9926 49096 11154
rect 49528 10266 49556 17274
rect 49700 16992 49752 16998
rect 49700 16934 49752 16940
rect 49712 15706 49740 16934
rect 49792 15972 49844 15978
rect 49792 15914 49844 15920
rect 49700 15700 49752 15706
rect 49700 15642 49752 15648
rect 49804 15570 49832 15914
rect 49792 15564 49844 15570
rect 49792 15506 49844 15512
rect 49804 15314 49832 15506
rect 49712 15286 49832 15314
rect 49712 14906 49740 15286
rect 49620 14878 49740 14906
rect 49620 12850 49648 14878
rect 49700 14816 49752 14822
rect 49700 14758 49752 14764
rect 49712 14618 49740 14758
rect 49700 14612 49752 14618
rect 49700 14554 49752 14560
rect 49608 12844 49660 12850
rect 49608 12786 49660 12792
rect 49620 12306 49648 12786
rect 50172 12434 50200 17478
rect 50528 17128 50580 17134
rect 50528 17070 50580 17076
rect 50436 16992 50488 16998
rect 50436 16934 50488 16940
rect 50448 16590 50476 16934
rect 50540 16794 50568 17070
rect 50528 16788 50580 16794
rect 50528 16730 50580 16736
rect 50436 16584 50488 16590
rect 50436 16526 50488 16532
rect 50724 15978 50752 18770
rect 50988 18760 51040 18766
rect 50988 18702 51040 18708
rect 51000 18086 51028 18702
rect 50988 18080 51040 18086
rect 50988 18022 51040 18028
rect 51092 16250 51120 20742
rect 51264 20392 51316 20398
rect 51264 20334 51316 20340
rect 51276 19514 51304 20334
rect 52000 20256 52052 20262
rect 52000 20198 52052 20204
rect 51504 20156 51812 20165
rect 51504 20154 51510 20156
rect 51566 20154 51590 20156
rect 51646 20154 51670 20156
rect 51726 20154 51750 20156
rect 51806 20154 51812 20156
rect 51566 20102 51568 20154
rect 51748 20102 51750 20154
rect 51504 20100 51510 20102
rect 51566 20100 51590 20102
rect 51646 20100 51670 20102
rect 51726 20100 51750 20102
rect 51806 20100 51812 20102
rect 51504 20091 51812 20100
rect 52012 20058 52040 20198
rect 52000 20052 52052 20058
rect 52000 19994 52052 20000
rect 51356 19712 51408 19718
rect 51356 19654 51408 19660
rect 51264 19508 51316 19514
rect 51264 19450 51316 19456
rect 51172 19168 51224 19174
rect 51172 19110 51224 19116
rect 51184 18358 51212 19110
rect 51172 18352 51224 18358
rect 51172 18294 51224 18300
rect 51368 17678 51396 19654
rect 52104 19378 52132 21490
rect 52196 21010 52224 21830
rect 52274 21720 52330 21729
rect 52274 21655 52330 21664
rect 52288 21486 52316 21655
rect 52380 21622 52408 21966
rect 52368 21616 52420 21622
rect 52368 21558 52420 21564
rect 52472 21554 52500 21966
rect 52736 21888 52788 21894
rect 52736 21830 52788 21836
rect 52460 21548 52512 21554
rect 52460 21490 52512 21496
rect 52276 21480 52328 21486
rect 52276 21422 52328 21428
rect 52644 21344 52696 21350
rect 52644 21286 52696 21292
rect 52656 21010 52684 21286
rect 52184 21004 52236 21010
rect 52184 20946 52236 20952
rect 52644 21004 52696 21010
rect 52644 20946 52696 20952
rect 52460 20936 52512 20942
rect 52460 20878 52512 20884
rect 52472 19922 52500 20878
rect 52460 19916 52512 19922
rect 52460 19858 52512 19864
rect 52092 19372 52144 19378
rect 52092 19314 52144 19320
rect 51504 19068 51812 19077
rect 51504 19066 51510 19068
rect 51566 19066 51590 19068
rect 51646 19066 51670 19068
rect 51726 19066 51750 19068
rect 51806 19066 51812 19068
rect 51566 19014 51568 19066
rect 51748 19014 51750 19066
rect 51504 19012 51510 19014
rect 51566 19012 51590 19014
rect 51646 19012 51670 19014
rect 51726 19012 51750 19014
rect 51806 19012 51812 19014
rect 51504 19003 51812 19012
rect 51504 17980 51812 17989
rect 51504 17978 51510 17980
rect 51566 17978 51590 17980
rect 51646 17978 51670 17980
rect 51726 17978 51750 17980
rect 51806 17978 51812 17980
rect 51566 17926 51568 17978
rect 51748 17926 51750 17978
rect 51504 17924 51510 17926
rect 51566 17924 51590 17926
rect 51646 17924 51670 17926
rect 51726 17924 51750 17926
rect 51806 17924 51812 17926
rect 51504 17915 51812 17924
rect 52460 17876 52512 17882
rect 52460 17818 52512 17824
rect 51356 17672 51408 17678
rect 51356 17614 51408 17620
rect 51908 17536 51960 17542
rect 51908 17478 51960 17484
rect 51504 16892 51812 16901
rect 51504 16890 51510 16892
rect 51566 16890 51590 16892
rect 51646 16890 51670 16892
rect 51726 16890 51750 16892
rect 51806 16890 51812 16892
rect 51566 16838 51568 16890
rect 51748 16838 51750 16890
rect 51504 16836 51510 16838
rect 51566 16836 51590 16838
rect 51646 16836 51670 16838
rect 51726 16836 51750 16838
rect 51806 16836 51812 16838
rect 51504 16827 51812 16836
rect 51920 16794 51948 17478
rect 51908 16788 51960 16794
rect 51908 16730 51960 16736
rect 51908 16448 51960 16454
rect 51908 16390 51960 16396
rect 51080 16244 51132 16250
rect 51080 16186 51132 16192
rect 51172 16244 51224 16250
rect 51172 16186 51224 16192
rect 50712 15972 50764 15978
rect 50712 15914 50764 15920
rect 50712 15496 50764 15502
rect 51092 15484 51120 16186
rect 51184 15638 51212 16186
rect 51920 16046 51948 16390
rect 51908 16040 51960 16046
rect 51908 15982 51960 15988
rect 51504 15804 51812 15813
rect 51504 15802 51510 15804
rect 51566 15802 51590 15804
rect 51646 15802 51670 15804
rect 51726 15802 51750 15804
rect 51806 15802 51812 15804
rect 51566 15750 51568 15802
rect 51748 15750 51750 15802
rect 51504 15748 51510 15750
rect 51566 15748 51590 15750
rect 51646 15748 51670 15750
rect 51726 15748 51750 15750
rect 51806 15748 51812 15750
rect 51504 15739 51812 15748
rect 51172 15632 51224 15638
rect 51172 15574 51224 15580
rect 51920 15570 51948 15982
rect 51448 15564 51500 15570
rect 51276 15524 51448 15552
rect 51276 15484 51304 15524
rect 51448 15506 51500 15512
rect 51908 15564 51960 15570
rect 51908 15506 51960 15512
rect 50712 15438 50764 15444
rect 51000 15456 51304 15484
rect 52276 15496 52328 15502
rect 50724 15162 50752 15438
rect 50712 15156 50764 15162
rect 50712 15098 50764 15104
rect 50252 14408 50304 14414
rect 50252 14350 50304 14356
rect 50264 14074 50292 14350
rect 50252 14068 50304 14074
rect 50252 14010 50304 14016
rect 50172 12406 50476 12434
rect 49608 12300 49660 12306
rect 49608 12242 49660 12248
rect 49884 12096 49936 12102
rect 49884 12038 49936 12044
rect 50160 12096 50212 12102
rect 50160 12038 50212 12044
rect 49896 11898 49924 12038
rect 49884 11892 49936 11898
rect 49884 11834 49936 11840
rect 49608 11552 49660 11558
rect 49608 11494 49660 11500
rect 49516 10260 49568 10266
rect 49516 10202 49568 10208
rect 48872 9920 48924 9926
rect 48872 9862 48924 9868
rect 49056 9920 49108 9926
rect 49056 9862 49108 9868
rect 48044 9512 48096 9518
rect 48044 9454 48096 9460
rect 48780 9512 48832 9518
rect 48780 9454 48832 9460
rect 48056 9178 48084 9454
rect 48136 9376 48188 9382
rect 48136 9318 48188 9324
rect 48044 9172 48096 9178
rect 48044 9114 48096 9120
rect 47952 8968 48004 8974
rect 47952 8910 48004 8916
rect 47860 8628 47912 8634
rect 47860 8570 47912 8576
rect 47964 7546 47992 8910
rect 48148 7818 48176 9318
rect 48320 8832 48372 8838
rect 48320 8774 48372 8780
rect 48412 8832 48464 8838
rect 48412 8774 48464 8780
rect 48688 8832 48740 8838
rect 48688 8774 48740 8780
rect 48136 7812 48188 7818
rect 48136 7754 48188 7760
rect 47952 7540 48004 7546
rect 47952 7482 48004 7488
rect 48332 7002 48360 8774
rect 48424 7750 48452 8774
rect 48700 8498 48728 8774
rect 48688 8492 48740 8498
rect 48688 8434 48740 8440
rect 48792 8090 48820 9454
rect 48780 8084 48832 8090
rect 48780 8026 48832 8032
rect 48412 7744 48464 7750
rect 48412 7686 48464 7692
rect 48424 7546 48452 7686
rect 48412 7540 48464 7546
rect 48412 7482 48464 7488
rect 48320 6996 48372 7002
rect 48320 6938 48372 6944
rect 48228 6656 48280 6662
rect 48228 6598 48280 6604
rect 48240 6322 48268 6598
rect 48228 6316 48280 6322
rect 48228 6258 48280 6264
rect 48240 5681 48268 6258
rect 48226 5672 48282 5681
rect 48226 5607 48282 5616
rect 48240 5166 48268 5607
rect 48424 5370 48452 7482
rect 48792 7410 48820 8026
rect 48780 7404 48832 7410
rect 48780 7346 48832 7352
rect 48504 7336 48556 7342
rect 48504 7278 48556 7284
rect 48516 6866 48544 7278
rect 48596 7268 48648 7274
rect 48596 7210 48648 7216
rect 48608 7002 48636 7210
rect 48596 6996 48648 7002
rect 48596 6938 48648 6944
rect 48504 6860 48556 6866
rect 48504 6802 48556 6808
rect 48608 6458 48636 6938
rect 48596 6452 48648 6458
rect 48596 6394 48648 6400
rect 48884 6118 48912 9862
rect 49332 9376 49384 9382
rect 49332 9318 49384 9324
rect 49344 9178 49372 9318
rect 49332 9172 49384 9178
rect 49332 9114 49384 9120
rect 49424 8492 49476 8498
rect 49424 8434 49476 8440
rect 49148 8016 49200 8022
rect 49148 7958 49200 7964
rect 49056 7812 49108 7818
rect 49056 7754 49108 7760
rect 49068 7410 49096 7754
rect 49056 7404 49108 7410
rect 49056 7346 49108 7352
rect 49160 6934 49188 7958
rect 49436 7954 49464 8434
rect 49620 8022 49648 11494
rect 50172 11354 50200 12038
rect 50160 11348 50212 11354
rect 50160 11290 50212 11296
rect 49700 11076 49752 11082
rect 49700 11018 49752 11024
rect 49712 10810 49740 11018
rect 49700 10804 49752 10810
rect 49700 10746 49752 10752
rect 49884 9512 49936 9518
rect 49884 9454 49936 9460
rect 49896 8634 49924 9454
rect 50068 9376 50120 9382
rect 50068 9318 50120 9324
rect 49884 8628 49936 8634
rect 49884 8570 49936 8576
rect 49608 8016 49660 8022
rect 49608 7958 49660 7964
rect 49424 7948 49476 7954
rect 49424 7890 49476 7896
rect 49896 7410 49924 8570
rect 49976 7744 50028 7750
rect 49976 7686 50028 7692
rect 49884 7404 49936 7410
rect 49884 7346 49936 7352
rect 49514 7304 49570 7313
rect 49514 7239 49516 7248
rect 49568 7239 49570 7248
rect 49516 7210 49568 7216
rect 49988 7018 50016 7686
rect 50080 7206 50108 9318
rect 50160 8968 50212 8974
rect 50160 8910 50212 8916
rect 50172 8090 50200 8910
rect 50252 8288 50304 8294
rect 50252 8230 50304 8236
rect 50160 8084 50212 8090
rect 50160 8026 50212 8032
rect 50264 7342 50292 8230
rect 50252 7336 50304 7342
rect 50252 7278 50304 7284
rect 50068 7200 50120 7206
rect 50068 7142 50120 7148
rect 50160 7200 50212 7206
rect 50160 7142 50212 7148
rect 50172 7018 50200 7142
rect 49608 6996 49660 7002
rect 49988 6990 50200 7018
rect 50264 7002 50292 7278
rect 49608 6938 49660 6944
rect 49148 6928 49200 6934
rect 49148 6870 49200 6876
rect 49160 6633 49188 6870
rect 49146 6624 49202 6633
rect 49146 6559 49202 6568
rect 49148 6452 49200 6458
rect 49148 6394 49200 6400
rect 48872 6112 48924 6118
rect 48872 6054 48924 6060
rect 48688 5704 48740 5710
rect 48688 5646 48740 5652
rect 48504 5568 48556 5574
rect 48504 5510 48556 5516
rect 48412 5364 48464 5370
rect 48412 5306 48464 5312
rect 48228 5160 48280 5166
rect 48148 5108 48228 5114
rect 48148 5102 48280 5108
rect 48148 5086 48268 5102
rect 47860 4140 47912 4146
rect 47860 4082 47912 4088
rect 47768 3732 47820 3738
rect 47768 3674 47820 3680
rect 47676 3664 47728 3670
rect 47676 3606 47728 3612
rect 47584 3596 47636 3602
rect 47584 3538 47636 3544
rect 47688 2854 47716 3606
rect 47872 3194 47900 4082
rect 48148 3777 48176 5086
rect 48228 4752 48280 4758
rect 48228 4694 48280 4700
rect 48240 4146 48268 4694
rect 48424 4622 48452 5306
rect 48516 4690 48544 5510
rect 48596 5092 48648 5098
rect 48596 5034 48648 5040
rect 48504 4684 48556 4690
rect 48504 4626 48556 4632
rect 48412 4616 48464 4622
rect 48412 4558 48464 4564
rect 48608 4282 48636 5034
rect 48700 4826 48728 5646
rect 48780 5160 48832 5166
rect 48780 5102 48832 5108
rect 48792 4826 48820 5102
rect 49160 5098 49188 6394
rect 49620 6254 49648 6938
rect 49884 6928 49936 6934
rect 49884 6870 49936 6876
rect 49896 6390 49924 6870
rect 49884 6384 49936 6390
rect 49884 6326 49936 6332
rect 50068 6316 50120 6322
rect 50068 6258 50120 6264
rect 49608 6248 49660 6254
rect 49608 6190 49660 6196
rect 49620 5914 49648 6190
rect 49608 5908 49660 5914
rect 49608 5850 49660 5856
rect 49620 5794 49648 5850
rect 49620 5766 49740 5794
rect 49424 5568 49476 5574
rect 49424 5510 49476 5516
rect 49436 5234 49464 5510
rect 49712 5234 49740 5766
rect 49424 5228 49476 5234
rect 49424 5170 49476 5176
rect 49700 5228 49752 5234
rect 49700 5170 49752 5176
rect 49148 5092 49200 5098
rect 49148 5034 49200 5040
rect 48688 4820 48740 4826
rect 48688 4762 48740 4768
rect 48780 4820 48832 4826
rect 48780 4762 48832 4768
rect 49436 4690 49464 5170
rect 49792 5024 49844 5030
rect 49792 4966 49844 4972
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49240 4616 49292 4622
rect 49240 4558 49292 4564
rect 49252 4282 49280 4558
rect 48596 4276 48648 4282
rect 48596 4218 48648 4224
rect 49240 4276 49292 4282
rect 49240 4218 49292 4224
rect 49424 4276 49476 4282
rect 49424 4218 49476 4224
rect 48228 4140 48280 4146
rect 48228 4082 48280 4088
rect 49332 4072 49384 4078
rect 49332 4014 49384 4020
rect 49344 3913 49372 4014
rect 49330 3904 49386 3913
rect 49330 3839 49386 3848
rect 48134 3768 48190 3777
rect 49436 3738 49464 4218
rect 49804 4060 49832 4966
rect 50080 4826 50108 6258
rect 50172 5710 50200 6990
rect 50252 6996 50304 7002
rect 50252 6938 50304 6944
rect 50344 6112 50396 6118
rect 50344 6054 50396 6060
rect 50356 5778 50384 6054
rect 50344 5772 50396 5778
rect 50344 5714 50396 5720
rect 50160 5704 50212 5710
rect 50160 5646 50212 5652
rect 50344 5024 50396 5030
rect 50344 4966 50396 4972
rect 50356 4826 50384 4966
rect 50068 4820 50120 4826
rect 50068 4762 50120 4768
rect 50344 4820 50396 4826
rect 50344 4762 50396 4768
rect 50160 4480 50212 4486
rect 50160 4422 50212 4428
rect 49884 4072 49936 4078
rect 49804 4032 49884 4060
rect 49516 3936 49568 3942
rect 49516 3878 49568 3884
rect 48134 3703 48190 3712
rect 49424 3732 49476 3738
rect 49424 3674 49476 3680
rect 48044 3528 48096 3534
rect 48044 3470 48096 3476
rect 47860 3188 47912 3194
rect 47860 3130 47912 3136
rect 48056 3126 48084 3470
rect 49528 3466 49556 3878
rect 49804 3738 49832 4032
rect 49884 4014 49936 4020
rect 49792 3732 49844 3738
rect 49792 3674 49844 3680
rect 49516 3460 49568 3466
rect 49516 3402 49568 3408
rect 48320 3392 48372 3398
rect 48320 3334 48372 3340
rect 49700 3392 49752 3398
rect 49700 3334 49752 3340
rect 48044 3120 48096 3126
rect 48042 3088 48044 3097
rect 48096 3088 48098 3097
rect 48042 3023 48098 3032
rect 47860 2984 47912 2990
rect 47860 2926 47912 2932
rect 47676 2848 47728 2854
rect 47676 2790 47728 2796
rect 47400 2644 47452 2650
rect 47400 2586 47452 2592
rect 47492 2508 47544 2514
rect 47320 2468 47492 2496
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47320 800 47348 2468
rect 47492 2450 47544 2456
rect 47872 800 47900 2926
rect 48332 2446 48360 3334
rect 49240 2984 49292 2990
rect 49240 2926 49292 2932
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 48424 800 48452 2382
rect 48976 870 49096 898
rect 48976 800 49004 870
rect 43548 734 43944 762
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46202 0 46258 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47858 0 47914 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49068 762 49096 870
rect 49252 762 49280 2926
rect 49712 2650 49740 3334
rect 50172 3126 50200 4422
rect 50448 3466 50476 12406
rect 51000 11898 51028 15456
rect 52276 15438 52328 15444
rect 52368 15496 52420 15502
rect 52368 15438 52420 15444
rect 51356 15428 51408 15434
rect 51356 15370 51408 15376
rect 51264 15360 51316 15366
rect 51264 15302 51316 15308
rect 51276 14346 51304 15302
rect 51368 14958 51396 15370
rect 51356 14952 51408 14958
rect 51356 14894 51408 14900
rect 51908 14952 51960 14958
rect 51908 14894 51960 14900
rect 51368 14482 51396 14894
rect 51504 14716 51812 14725
rect 51504 14714 51510 14716
rect 51566 14714 51590 14716
rect 51646 14714 51670 14716
rect 51726 14714 51750 14716
rect 51806 14714 51812 14716
rect 51566 14662 51568 14714
rect 51748 14662 51750 14714
rect 51504 14660 51510 14662
rect 51566 14660 51590 14662
rect 51646 14660 51670 14662
rect 51726 14660 51750 14662
rect 51806 14660 51812 14662
rect 51504 14651 51812 14660
rect 51920 14618 51948 14894
rect 52000 14816 52052 14822
rect 52000 14758 52052 14764
rect 51908 14612 51960 14618
rect 51908 14554 51960 14560
rect 51356 14476 51408 14482
rect 51356 14418 51408 14424
rect 51264 14340 51316 14346
rect 51264 14282 51316 14288
rect 51724 14340 51776 14346
rect 51724 14282 51776 14288
rect 51632 14272 51684 14278
rect 51632 14214 51684 14220
rect 51644 14074 51672 14214
rect 51632 14068 51684 14074
rect 51632 14010 51684 14016
rect 51736 13802 51764 14282
rect 52012 14278 52040 14758
rect 52092 14476 52144 14482
rect 52092 14418 52144 14424
rect 52184 14476 52236 14482
rect 52184 14418 52236 14424
rect 52000 14272 52052 14278
rect 52000 14214 52052 14220
rect 52012 14074 52040 14214
rect 52000 14068 52052 14074
rect 52000 14010 52052 14016
rect 52104 14006 52132 14418
rect 52092 14000 52144 14006
rect 52092 13942 52144 13948
rect 51724 13796 51776 13802
rect 51724 13738 51776 13744
rect 51504 13628 51812 13637
rect 51504 13626 51510 13628
rect 51566 13626 51590 13628
rect 51646 13626 51670 13628
rect 51726 13626 51750 13628
rect 51806 13626 51812 13628
rect 51566 13574 51568 13626
rect 51748 13574 51750 13626
rect 51504 13572 51510 13574
rect 51566 13572 51590 13574
rect 51646 13572 51670 13574
rect 51726 13572 51750 13574
rect 51806 13572 51812 13574
rect 51504 13563 51812 13572
rect 52196 13530 52224 14418
rect 52288 14346 52316 15438
rect 52380 15026 52408 15438
rect 52472 15162 52500 17818
rect 52656 16250 52684 20946
rect 52748 20806 52776 21830
rect 52736 20800 52788 20806
rect 52736 20742 52788 20748
rect 52932 20602 52960 22510
rect 53564 22432 53616 22438
rect 53564 22374 53616 22380
rect 54852 22432 54904 22438
rect 54852 22374 54904 22380
rect 53576 21554 53604 22374
rect 54484 21888 54536 21894
rect 54484 21830 54536 21836
rect 54760 21888 54812 21894
rect 54760 21830 54812 21836
rect 54496 21690 54524 21830
rect 54772 21690 54800 21830
rect 54484 21684 54536 21690
rect 54484 21626 54536 21632
rect 54760 21684 54812 21690
rect 54760 21626 54812 21632
rect 53564 21548 53616 21554
rect 53564 21490 53616 21496
rect 53748 21344 53800 21350
rect 53748 21286 53800 21292
rect 53760 21078 53788 21286
rect 54772 21146 54800 21626
rect 54864 21622 54892 22374
rect 55324 22234 55352 22510
rect 55772 22432 55824 22438
rect 55772 22374 55824 22380
rect 55312 22228 55364 22234
rect 55312 22170 55364 22176
rect 55784 22098 55812 22374
rect 55772 22092 55824 22098
rect 55772 22034 55824 22040
rect 55864 22092 55916 22098
rect 55864 22034 55916 22040
rect 54852 21616 54904 21622
rect 55876 21593 55904 22034
rect 55968 21690 55996 22510
rect 56692 22432 56744 22438
rect 56692 22374 56744 22380
rect 56704 22166 56732 22374
rect 56692 22160 56744 22166
rect 56692 22102 56744 22108
rect 56704 21729 56732 22102
rect 58532 21956 58584 21962
rect 58532 21898 58584 21904
rect 57796 21888 57848 21894
rect 57796 21830 57848 21836
rect 57980 21888 58032 21894
rect 57980 21830 58032 21836
rect 56690 21720 56746 21729
rect 55956 21684 56008 21690
rect 55956 21626 56008 21632
rect 56508 21684 56560 21690
rect 56690 21655 56746 21664
rect 56508 21626 56560 21632
rect 54852 21558 54904 21564
rect 55862 21584 55918 21593
rect 55862 21519 55918 21528
rect 56048 21548 56100 21554
rect 56048 21490 56100 21496
rect 54760 21140 54812 21146
rect 54760 21082 54812 21088
rect 53748 21072 53800 21078
rect 53748 21014 53800 21020
rect 53564 20936 53616 20942
rect 53194 20904 53250 20913
rect 53564 20878 53616 20884
rect 53194 20839 53196 20848
rect 53248 20839 53250 20848
rect 53196 20810 53248 20816
rect 53288 20800 53340 20806
rect 53288 20742 53340 20748
rect 52920 20596 52972 20602
rect 52920 20538 52972 20544
rect 53196 20392 53248 20398
rect 53196 20334 53248 20340
rect 53012 19712 53064 19718
rect 53012 19654 53064 19660
rect 53024 19514 53052 19654
rect 53012 19508 53064 19514
rect 53012 19450 53064 19456
rect 53208 19378 53236 20334
rect 53012 19372 53064 19378
rect 53012 19314 53064 19320
rect 53196 19372 53248 19378
rect 53196 19314 53248 19320
rect 52828 18760 52880 18766
rect 52828 18702 52880 18708
rect 52736 18080 52788 18086
rect 52736 18022 52788 18028
rect 52748 17610 52776 18022
rect 52736 17604 52788 17610
rect 52736 17546 52788 17552
rect 52644 16244 52696 16250
rect 52644 16186 52696 16192
rect 52656 16130 52684 16186
rect 52564 16102 52684 16130
rect 52564 15570 52592 16102
rect 52552 15564 52604 15570
rect 52552 15506 52604 15512
rect 52644 15360 52696 15366
rect 52644 15302 52696 15308
rect 52460 15156 52512 15162
rect 52460 15098 52512 15104
rect 52368 15020 52420 15026
rect 52368 14962 52420 14968
rect 52276 14340 52328 14346
rect 52276 14282 52328 14288
rect 52184 13524 52236 13530
rect 52184 13466 52236 13472
rect 51172 12776 51224 12782
rect 51172 12718 51224 12724
rect 51356 12776 51408 12782
rect 51356 12718 51408 12724
rect 51080 12640 51132 12646
rect 51080 12582 51132 12588
rect 51092 12170 51120 12582
rect 51080 12164 51132 12170
rect 51080 12106 51132 12112
rect 51184 11898 51212 12718
rect 51368 12434 51396 12718
rect 52368 12640 52420 12646
rect 52368 12582 52420 12588
rect 51504 12540 51812 12549
rect 51504 12538 51510 12540
rect 51566 12538 51590 12540
rect 51646 12538 51670 12540
rect 51726 12538 51750 12540
rect 51806 12538 51812 12540
rect 51566 12486 51568 12538
rect 51748 12486 51750 12538
rect 51504 12484 51510 12486
rect 51566 12484 51590 12486
rect 51646 12484 51670 12486
rect 51726 12484 51750 12486
rect 51806 12484 51812 12486
rect 51504 12475 51812 12484
rect 51448 12436 51500 12442
rect 51368 12406 51448 12434
rect 50988 11892 51040 11898
rect 51172 11892 51224 11898
rect 51040 11852 51120 11880
rect 50988 11834 51040 11840
rect 51092 11540 51120 11852
rect 51172 11834 51224 11840
rect 51264 11756 51316 11762
rect 51264 11698 51316 11704
rect 51172 11552 51224 11558
rect 51092 11512 51172 11540
rect 51172 11494 51224 11500
rect 51276 10810 51304 11698
rect 51368 11218 51396 12406
rect 51448 12378 51500 12384
rect 52184 12096 52236 12102
rect 52184 12038 52236 12044
rect 52000 11688 52052 11694
rect 52000 11630 52052 11636
rect 52092 11688 52144 11694
rect 52092 11630 52144 11636
rect 51504 11452 51812 11461
rect 51504 11450 51510 11452
rect 51566 11450 51590 11452
rect 51646 11450 51670 11452
rect 51726 11450 51750 11452
rect 51806 11450 51812 11452
rect 51566 11398 51568 11450
rect 51748 11398 51750 11450
rect 51504 11396 51510 11398
rect 51566 11396 51590 11398
rect 51646 11396 51670 11398
rect 51726 11396 51750 11398
rect 51806 11396 51812 11398
rect 51504 11387 51812 11396
rect 51356 11212 51408 11218
rect 51356 11154 51408 11160
rect 52012 10810 52040 11630
rect 51264 10804 51316 10810
rect 51264 10746 51316 10752
rect 52000 10804 52052 10810
rect 52000 10746 52052 10752
rect 52104 10742 52132 11630
rect 52196 11218 52224 12038
rect 52380 11898 52408 12582
rect 52368 11892 52420 11898
rect 52368 11834 52420 11840
rect 52656 11642 52684 15302
rect 52472 11614 52684 11642
rect 52276 11552 52328 11558
rect 52276 11494 52328 11500
rect 52288 11218 52316 11494
rect 52184 11212 52236 11218
rect 52184 11154 52236 11160
rect 52276 11212 52328 11218
rect 52276 11154 52328 11160
rect 52276 10804 52328 10810
rect 52276 10746 52328 10752
rect 51356 10736 51408 10742
rect 51356 10678 51408 10684
rect 52092 10736 52144 10742
rect 52092 10678 52144 10684
rect 51264 10668 51316 10674
rect 51264 10610 51316 10616
rect 50896 10192 50948 10198
rect 50896 10134 50948 10140
rect 50908 9926 50936 10134
rect 50896 9920 50948 9926
rect 50896 9862 50948 9868
rect 50988 9920 51040 9926
rect 50988 9862 51040 9868
rect 50804 8832 50856 8838
rect 50804 8774 50856 8780
rect 50816 8634 50844 8774
rect 50804 8628 50856 8634
rect 50804 8570 50856 8576
rect 50620 8288 50672 8294
rect 50620 8230 50672 8236
rect 50712 8288 50764 8294
rect 50712 8230 50764 8236
rect 50632 7478 50660 8230
rect 50724 7546 50752 8230
rect 50804 7880 50856 7886
rect 50804 7822 50856 7828
rect 50816 7546 50844 7822
rect 50712 7540 50764 7546
rect 50712 7482 50764 7488
rect 50804 7540 50856 7546
rect 50804 7482 50856 7488
rect 50620 7472 50672 7478
rect 50620 7414 50672 7420
rect 50712 7200 50764 7206
rect 50712 7142 50764 7148
rect 50528 6112 50580 6118
rect 50528 6054 50580 6060
rect 50540 5234 50568 6054
rect 50528 5228 50580 5234
rect 50528 5170 50580 5176
rect 50540 3602 50568 5170
rect 50724 4554 50752 7142
rect 50908 6934 50936 9862
rect 51000 9586 51028 9862
rect 51276 9722 51304 10610
rect 51368 10130 51396 10678
rect 52288 10606 52316 10746
rect 52276 10600 52328 10606
rect 52276 10542 52328 10548
rect 51504 10364 51812 10373
rect 51504 10362 51510 10364
rect 51566 10362 51590 10364
rect 51646 10362 51670 10364
rect 51726 10362 51750 10364
rect 51806 10362 51812 10364
rect 51566 10310 51568 10362
rect 51748 10310 51750 10362
rect 51504 10308 51510 10310
rect 51566 10308 51590 10310
rect 51646 10308 51670 10310
rect 51726 10308 51750 10310
rect 51806 10308 51812 10310
rect 51504 10299 51812 10308
rect 51356 10124 51408 10130
rect 51356 10066 51408 10072
rect 52288 9722 52316 10542
rect 51264 9716 51316 9722
rect 51264 9658 51316 9664
rect 52276 9716 52328 9722
rect 52276 9658 52328 9664
rect 50988 9580 51040 9586
rect 50988 9522 51040 9528
rect 51504 9276 51812 9285
rect 51504 9274 51510 9276
rect 51566 9274 51590 9276
rect 51646 9274 51670 9276
rect 51726 9274 51750 9276
rect 51806 9274 51812 9276
rect 51566 9222 51568 9274
rect 51748 9222 51750 9274
rect 51504 9220 51510 9222
rect 51566 9220 51590 9222
rect 51646 9220 51670 9222
rect 51726 9220 51750 9222
rect 51806 9220 51812 9222
rect 51504 9211 51812 9220
rect 52288 9042 52316 9658
rect 52276 9036 52328 9042
rect 52276 8978 52328 8984
rect 52288 8634 52316 8978
rect 52276 8628 52328 8634
rect 52276 8570 52328 8576
rect 51356 8424 51408 8430
rect 51356 8366 51408 8372
rect 51368 8090 51396 8366
rect 52184 8288 52236 8294
rect 52184 8230 52236 8236
rect 52276 8288 52328 8294
rect 52276 8230 52328 8236
rect 51504 8188 51812 8197
rect 51504 8186 51510 8188
rect 51566 8186 51590 8188
rect 51646 8186 51670 8188
rect 51726 8186 51750 8188
rect 51806 8186 51812 8188
rect 51566 8134 51568 8186
rect 51748 8134 51750 8186
rect 51504 8132 51510 8134
rect 51566 8132 51590 8134
rect 51646 8132 51670 8134
rect 51726 8132 51750 8134
rect 51806 8132 51812 8134
rect 51504 8123 51812 8132
rect 51356 8084 51408 8090
rect 51356 8026 51408 8032
rect 51368 7750 51396 8026
rect 51356 7744 51408 7750
rect 51356 7686 51408 7692
rect 51448 7744 51500 7750
rect 51448 7686 51500 7692
rect 51356 7336 51408 7342
rect 51460 7324 51488 7686
rect 52196 7546 52224 8230
rect 52184 7540 52236 7546
rect 52184 7482 52236 7488
rect 51408 7296 51488 7324
rect 51356 7278 51408 7284
rect 51368 7002 51396 7278
rect 52184 7200 52236 7206
rect 52184 7142 52236 7148
rect 51504 7100 51812 7109
rect 51504 7098 51510 7100
rect 51566 7098 51590 7100
rect 51646 7098 51670 7100
rect 51726 7098 51750 7100
rect 51806 7098 51812 7100
rect 51566 7046 51568 7098
rect 51748 7046 51750 7098
rect 51504 7044 51510 7046
rect 51566 7044 51590 7046
rect 51646 7044 51670 7046
rect 51726 7044 51750 7046
rect 51806 7044 51812 7046
rect 51504 7035 51812 7044
rect 51356 6996 51408 7002
rect 51356 6938 51408 6944
rect 51632 6996 51684 7002
rect 51632 6938 51684 6944
rect 50896 6928 50948 6934
rect 50896 6870 50948 6876
rect 51644 6390 51672 6938
rect 52196 6458 52224 7142
rect 52184 6452 52236 6458
rect 52184 6394 52236 6400
rect 51632 6384 51684 6390
rect 51632 6326 51684 6332
rect 52288 6254 52316 8230
rect 52276 6248 52328 6254
rect 52276 6190 52328 6196
rect 51504 6012 51812 6021
rect 51504 6010 51510 6012
rect 51566 6010 51590 6012
rect 51646 6010 51670 6012
rect 51726 6010 51750 6012
rect 51806 6010 51812 6012
rect 51566 5958 51568 6010
rect 51748 5958 51750 6010
rect 51504 5956 51510 5958
rect 51566 5956 51590 5958
rect 51646 5956 51670 5958
rect 51726 5956 51750 5958
rect 51806 5956 51812 5958
rect 51504 5947 51812 5956
rect 50988 5704 51040 5710
rect 50988 5646 51040 5652
rect 51000 5370 51028 5646
rect 52368 5568 52420 5574
rect 52368 5510 52420 5516
rect 50988 5364 51040 5370
rect 50988 5306 51040 5312
rect 52092 5296 52144 5302
rect 52092 5238 52144 5244
rect 52104 5030 52132 5238
rect 52380 5234 52408 5510
rect 52368 5228 52420 5234
rect 52368 5170 52420 5176
rect 52276 5160 52328 5166
rect 52276 5102 52328 5108
rect 51080 5024 51132 5030
rect 51080 4966 51132 4972
rect 52092 5024 52144 5030
rect 52092 4966 52144 4972
rect 50712 4548 50764 4554
rect 50712 4490 50764 4496
rect 51092 3913 51120 4966
rect 51504 4924 51812 4933
rect 51504 4922 51510 4924
rect 51566 4922 51590 4924
rect 51646 4922 51670 4924
rect 51726 4922 51750 4924
rect 51806 4922 51812 4924
rect 51566 4870 51568 4922
rect 51748 4870 51750 4922
rect 51504 4868 51510 4870
rect 51566 4868 51590 4870
rect 51646 4868 51670 4870
rect 51726 4868 51750 4870
rect 51806 4868 51812 4870
rect 51504 4859 51812 4868
rect 52288 4826 52316 5102
rect 52276 4820 52328 4826
rect 52276 4762 52328 4768
rect 51448 4616 51500 4622
rect 51448 4558 51500 4564
rect 51264 4480 51316 4486
rect 51264 4422 51316 4428
rect 51276 4049 51304 4422
rect 51262 4040 51318 4049
rect 51460 4026 51488 4558
rect 52092 4480 52144 4486
rect 52092 4422 52144 4428
rect 51262 3975 51318 3984
rect 51368 3998 51488 4026
rect 52000 4072 52052 4078
rect 52000 4014 52052 4020
rect 51078 3904 51134 3913
rect 51078 3839 51134 3848
rect 50710 3768 50766 3777
rect 50710 3703 50712 3712
rect 50764 3703 50766 3712
rect 50712 3674 50764 3680
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50988 3528 51040 3534
rect 51040 3488 51120 3516
rect 50988 3470 51040 3476
rect 50252 3460 50304 3466
rect 50252 3402 50304 3408
rect 50436 3460 50488 3466
rect 50436 3402 50488 3408
rect 50160 3120 50212 3126
rect 50160 3062 50212 3068
rect 50068 2984 50120 2990
rect 50068 2926 50120 2932
rect 49700 2644 49752 2650
rect 49700 2586 49752 2592
rect 49700 2440 49752 2446
rect 49528 2400 49700 2428
rect 49528 800 49556 2400
rect 49700 2382 49752 2388
rect 50080 800 50108 2926
rect 50264 2650 50292 3402
rect 51092 3194 51120 3488
rect 51264 3392 51316 3398
rect 51264 3334 51316 3340
rect 51080 3188 51132 3194
rect 51080 3130 51132 3136
rect 51276 3074 51304 3334
rect 51092 3046 51304 3074
rect 50252 2644 50304 2650
rect 50252 2586 50304 2592
rect 50620 2508 50672 2514
rect 50620 2450 50672 2456
rect 50632 800 50660 2450
rect 51092 2446 51120 3046
rect 51172 2848 51224 2854
rect 51172 2790 51224 2796
rect 51184 2446 51212 2790
rect 51368 2774 51396 3998
rect 51504 3836 51812 3845
rect 51504 3834 51510 3836
rect 51566 3834 51590 3836
rect 51646 3834 51670 3836
rect 51726 3834 51750 3836
rect 51806 3834 51812 3836
rect 51566 3782 51568 3834
rect 51748 3782 51750 3834
rect 51504 3780 51510 3782
rect 51566 3780 51590 3782
rect 51646 3780 51670 3782
rect 51726 3780 51750 3782
rect 51806 3780 51812 3782
rect 51504 3771 51812 3780
rect 52012 3505 52040 4014
rect 52104 3641 52132 4422
rect 52090 3632 52146 3641
rect 52090 3567 52146 3576
rect 51998 3496 52054 3505
rect 51998 3431 52054 3440
rect 52472 3058 52500 11614
rect 52552 11552 52604 11558
rect 52552 11494 52604 11500
rect 52564 11354 52592 11494
rect 52552 11348 52604 11354
rect 52552 11290 52604 11296
rect 52552 11212 52604 11218
rect 52552 11154 52604 11160
rect 52564 10606 52592 11154
rect 52644 11144 52696 11150
rect 52644 11086 52696 11092
rect 52552 10600 52604 10606
rect 52552 10542 52604 10548
rect 52656 10538 52684 11086
rect 52644 10532 52696 10538
rect 52644 10474 52696 10480
rect 52656 10130 52684 10474
rect 52644 10124 52696 10130
rect 52644 10066 52696 10072
rect 52644 9920 52696 9926
rect 52644 9862 52696 9868
rect 52552 8968 52604 8974
rect 52552 8910 52604 8916
rect 52564 7886 52592 8910
rect 52552 7880 52604 7886
rect 52552 7822 52604 7828
rect 52564 6322 52592 7822
rect 52552 6316 52604 6322
rect 52552 6258 52604 6264
rect 52564 5778 52592 6258
rect 52552 5772 52604 5778
rect 52552 5714 52604 5720
rect 52552 3936 52604 3942
rect 52550 3904 52552 3913
rect 52604 3904 52606 3913
rect 52550 3839 52606 3848
rect 52552 3460 52604 3466
rect 52552 3402 52604 3408
rect 52564 3194 52592 3402
rect 52552 3188 52604 3194
rect 52552 3130 52604 3136
rect 52460 3052 52512 3058
rect 52460 2994 52512 3000
rect 51908 2984 51960 2990
rect 51908 2926 51960 2932
rect 51276 2746 51396 2774
rect 51504 2748 51812 2757
rect 51504 2746 51510 2748
rect 51566 2746 51590 2748
rect 51646 2746 51670 2748
rect 51726 2746 51750 2748
rect 51806 2746 51812 2748
rect 51080 2440 51132 2446
rect 51080 2382 51132 2388
rect 51172 2440 51224 2446
rect 51172 2382 51224 2388
rect 51276 2258 51304 2746
rect 51566 2694 51568 2746
rect 51748 2694 51750 2746
rect 51504 2692 51510 2694
rect 51566 2692 51590 2694
rect 51646 2692 51670 2694
rect 51726 2692 51750 2694
rect 51806 2692 51812 2694
rect 51504 2683 51812 2692
rect 51184 2230 51304 2258
rect 51184 800 51212 2230
rect 51920 1578 51948 2926
rect 52460 2848 52512 2854
rect 52460 2790 52512 2796
rect 52368 2508 52420 2514
rect 51736 1550 51948 1578
rect 52288 2468 52368 2496
rect 51736 800 51764 1550
rect 52288 800 52316 2468
rect 52368 2450 52420 2456
rect 52472 2446 52500 2790
rect 52656 2774 52684 9862
rect 52748 9654 52776 17546
rect 52840 17338 52868 18702
rect 52828 17332 52880 17338
rect 52828 17274 52880 17280
rect 53024 17202 53052 19314
rect 53104 18216 53156 18222
rect 53104 18158 53156 18164
rect 53116 17542 53144 18158
rect 53104 17536 53156 17542
rect 53104 17478 53156 17484
rect 53012 17196 53064 17202
rect 53012 17138 53064 17144
rect 53024 16046 53052 17138
rect 53012 16040 53064 16046
rect 53012 15982 53064 15988
rect 53116 15706 53144 17478
rect 53196 16584 53248 16590
rect 53196 16526 53248 16532
rect 53208 16250 53236 16526
rect 53196 16244 53248 16250
rect 53196 16186 53248 16192
rect 53196 16040 53248 16046
rect 53196 15982 53248 15988
rect 53104 15700 53156 15706
rect 53104 15642 53156 15648
rect 53104 15564 53156 15570
rect 53104 15506 53156 15512
rect 53116 15162 53144 15506
rect 53208 15314 53236 15982
rect 53300 15502 53328 20742
rect 53472 18624 53524 18630
rect 53472 18566 53524 18572
rect 53380 18080 53432 18086
rect 53380 18022 53432 18028
rect 53392 17338 53420 18022
rect 53484 17678 53512 18566
rect 53576 18290 53604 20878
rect 53760 20398 53788 21014
rect 56060 21010 56088 21490
rect 56520 21434 56548 21626
rect 56876 21548 56928 21554
rect 56876 21490 56928 21496
rect 56520 21406 56640 21434
rect 56508 21344 56560 21350
rect 56508 21286 56560 21292
rect 55588 21004 55640 21010
rect 55588 20946 55640 20952
rect 56048 21004 56100 21010
rect 56048 20946 56100 20952
rect 56232 21004 56284 21010
rect 56232 20946 56284 20952
rect 56416 21004 56468 21010
rect 56416 20946 56468 20952
rect 55036 20868 55088 20874
rect 55036 20810 55088 20816
rect 53748 20392 53800 20398
rect 53748 20334 53800 20340
rect 54852 20392 54904 20398
rect 54852 20334 54904 20340
rect 54668 20256 54720 20262
rect 54668 20198 54720 20204
rect 54680 20058 54708 20198
rect 54668 20052 54720 20058
rect 54668 19994 54720 20000
rect 53932 19712 53984 19718
rect 53932 19654 53984 19660
rect 53944 19310 53972 19654
rect 53932 19304 53984 19310
rect 53932 19246 53984 19252
rect 54024 19304 54076 19310
rect 54024 19246 54076 19252
rect 53564 18284 53616 18290
rect 53564 18226 53616 18232
rect 53472 17672 53524 17678
rect 53472 17614 53524 17620
rect 53576 17542 53604 18226
rect 53564 17536 53616 17542
rect 53564 17478 53616 17484
rect 53380 17332 53432 17338
rect 53380 17274 53432 17280
rect 53576 17134 53604 17478
rect 53380 17128 53432 17134
rect 53380 17070 53432 17076
rect 53564 17128 53616 17134
rect 53564 17070 53616 17076
rect 53288 15496 53340 15502
rect 53288 15438 53340 15444
rect 53208 15286 53328 15314
rect 53104 15156 53156 15162
rect 53104 15098 53156 15104
rect 53300 14074 53328 15286
rect 53288 14068 53340 14074
rect 53288 14010 53340 14016
rect 53300 12986 53328 14010
rect 53392 12986 53420 17070
rect 53840 16992 53892 16998
rect 53840 16934 53892 16940
rect 53852 16658 53880 16934
rect 53840 16652 53892 16658
rect 53840 16594 53892 16600
rect 53472 16040 53524 16046
rect 53472 15982 53524 15988
rect 53484 15910 53512 15982
rect 53472 15904 53524 15910
rect 53472 15846 53524 15852
rect 53288 12980 53340 12986
rect 53288 12922 53340 12928
rect 53380 12980 53432 12986
rect 53380 12922 53432 12928
rect 53196 12844 53248 12850
rect 53196 12786 53248 12792
rect 53012 12776 53064 12782
rect 53012 12718 53064 12724
rect 52920 12436 52972 12442
rect 52920 12378 52972 12384
rect 52932 12322 52960 12378
rect 52840 12294 52960 12322
rect 52840 11218 52868 12294
rect 53024 11898 53052 12718
rect 53012 11892 53064 11898
rect 53012 11834 53064 11840
rect 52828 11212 52880 11218
rect 52828 11154 52880 11160
rect 52736 9648 52788 9654
rect 52736 9590 52788 9596
rect 53012 8288 53064 8294
rect 53012 8230 53064 8236
rect 52736 7540 52788 7546
rect 52736 7482 52788 7488
rect 52748 6186 52776 7482
rect 53024 7410 53052 8230
rect 53012 7404 53064 7410
rect 53012 7346 53064 7352
rect 53104 6996 53156 7002
rect 53104 6938 53156 6944
rect 52828 6928 52880 6934
rect 52828 6870 52880 6876
rect 52840 6390 52868 6870
rect 52828 6384 52880 6390
rect 52828 6326 52880 6332
rect 52736 6180 52788 6186
rect 52736 6122 52788 6128
rect 52920 5024 52972 5030
rect 52920 4966 52972 4972
rect 52932 4690 52960 4966
rect 53116 4690 53144 6938
rect 52920 4684 52972 4690
rect 52920 4626 52972 4632
rect 53104 4684 53156 4690
rect 53104 4626 53156 4632
rect 52736 4140 52788 4146
rect 52736 4082 52788 4088
rect 52748 3602 52776 4082
rect 53104 3936 53156 3942
rect 53104 3878 53156 3884
rect 52736 3596 52788 3602
rect 52736 3538 52788 3544
rect 52828 3392 52880 3398
rect 52828 3334 52880 3340
rect 52840 3194 52868 3334
rect 52828 3188 52880 3194
rect 52828 3130 52880 3136
rect 52656 2746 52776 2774
rect 52748 2650 52776 2746
rect 52736 2644 52788 2650
rect 52736 2586 52788 2592
rect 52460 2440 52512 2446
rect 52460 2382 52512 2388
rect 52840 870 52960 898
rect 52840 800 52868 870
rect 49068 734 49280 762
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 52932 762 52960 870
rect 53116 762 53144 3878
rect 53208 2310 53236 12786
rect 53484 12434 53512 15846
rect 53852 14958 53880 16594
rect 53840 14952 53892 14958
rect 53840 14894 53892 14900
rect 53852 14414 53880 14894
rect 53840 14408 53892 14414
rect 53840 14350 53892 14356
rect 53944 13870 53972 19246
rect 54036 18970 54064 19246
rect 54576 19168 54628 19174
rect 54576 19110 54628 19116
rect 54024 18964 54076 18970
rect 54024 18906 54076 18912
rect 54024 18624 54076 18630
rect 54024 18566 54076 18572
rect 54036 13938 54064 18566
rect 54588 18358 54616 19110
rect 54864 18630 54892 20334
rect 55048 20058 55076 20810
rect 55600 20398 55628 20946
rect 56244 20890 56272 20946
rect 55784 20862 56272 20890
rect 55784 20806 55812 20862
rect 55772 20800 55824 20806
rect 55772 20742 55824 20748
rect 56428 20466 56456 20946
rect 56416 20460 56468 20466
rect 56416 20402 56468 20408
rect 55220 20392 55272 20398
rect 55140 20340 55220 20346
rect 55140 20334 55272 20340
rect 55588 20392 55640 20398
rect 55588 20334 55640 20340
rect 55140 20318 55260 20334
rect 55036 20052 55088 20058
rect 55036 19994 55088 20000
rect 55140 19718 55168 20318
rect 56520 19854 56548 21286
rect 56612 20942 56640 21406
rect 56888 21010 56916 21490
rect 57520 21344 57572 21350
rect 57520 21286 57572 21292
rect 57532 21146 57560 21286
rect 57520 21140 57572 21146
rect 57520 21082 57572 21088
rect 56876 21004 56928 21010
rect 56876 20946 56928 20952
rect 56600 20936 56652 20942
rect 56600 20878 56652 20884
rect 57808 20874 57836 21830
rect 57992 21690 58020 21830
rect 58544 21690 58572 21898
rect 58726 21788 59034 21797
rect 58726 21786 58732 21788
rect 58788 21786 58812 21788
rect 58868 21786 58892 21788
rect 58948 21786 58972 21788
rect 59028 21786 59034 21788
rect 58788 21734 58790 21786
rect 58970 21734 58972 21786
rect 58726 21732 58732 21734
rect 58788 21732 58812 21734
rect 58868 21732 58892 21734
rect 58948 21732 58972 21734
rect 59028 21732 59034 21734
rect 58726 21723 59034 21732
rect 57980 21684 58032 21690
rect 57980 21626 58032 21632
rect 58532 21684 58584 21690
rect 58532 21626 58584 21632
rect 58164 21004 58216 21010
rect 58164 20946 58216 20952
rect 57796 20868 57848 20874
rect 57796 20810 57848 20816
rect 56968 20800 57020 20806
rect 56968 20742 57020 20748
rect 57520 20800 57572 20806
rect 57520 20742 57572 20748
rect 57612 20800 57664 20806
rect 57612 20742 57664 20748
rect 57704 20800 57756 20806
rect 57704 20742 57756 20748
rect 56980 20466 57008 20742
rect 56968 20460 57020 20466
rect 56968 20402 57020 20408
rect 56980 20074 57008 20402
rect 56980 20058 57100 20074
rect 56980 20052 57112 20058
rect 56980 20046 57060 20052
rect 57060 19994 57112 20000
rect 56508 19848 56560 19854
rect 56508 19790 56560 19796
rect 55128 19712 55180 19718
rect 55128 19654 55180 19660
rect 55680 18896 55732 18902
rect 55680 18838 55732 18844
rect 54852 18624 54904 18630
rect 54852 18566 54904 18572
rect 54576 18352 54628 18358
rect 54576 18294 54628 18300
rect 54760 16652 54812 16658
rect 54760 16594 54812 16600
rect 54772 16250 54800 16594
rect 54864 16590 54892 18566
rect 55692 18290 55720 18838
rect 56520 18766 56548 19790
rect 57532 19514 57560 20742
rect 57624 20466 57652 20742
rect 57716 20602 57744 20742
rect 57704 20596 57756 20602
rect 57704 20538 57756 20544
rect 57612 20460 57664 20466
rect 57612 20402 57664 20408
rect 56600 19508 56652 19514
rect 56600 19450 56652 19456
rect 57520 19508 57572 19514
rect 57520 19450 57572 19456
rect 56048 18760 56100 18766
rect 56048 18702 56100 18708
rect 56508 18760 56560 18766
rect 56508 18702 56560 18708
rect 55680 18284 55732 18290
rect 55680 18226 55732 18232
rect 56060 17678 56088 18702
rect 56508 18624 56560 18630
rect 56508 18566 56560 18572
rect 56520 18426 56548 18566
rect 56508 18420 56560 18426
rect 56508 18362 56560 18368
rect 56520 18290 56548 18362
rect 56508 18284 56560 18290
rect 56508 18226 56560 18232
rect 56140 18216 56192 18222
rect 56140 18158 56192 18164
rect 56416 18216 56468 18222
rect 56416 18158 56468 18164
rect 56048 17672 56100 17678
rect 55494 17640 55550 17649
rect 56048 17614 56100 17620
rect 55494 17575 55496 17584
rect 55548 17575 55550 17584
rect 55496 17546 55548 17552
rect 55404 17332 55456 17338
rect 55404 17274 55456 17280
rect 55128 17128 55180 17134
rect 55128 17070 55180 17076
rect 55140 16794 55168 17070
rect 55128 16788 55180 16794
rect 55128 16730 55180 16736
rect 55416 16658 55444 17274
rect 55404 16652 55456 16658
rect 55404 16594 55456 16600
rect 54852 16584 54904 16590
rect 54852 16526 54904 16532
rect 54760 16244 54812 16250
rect 54760 16186 54812 16192
rect 54772 15450 54800 16186
rect 55220 15904 55272 15910
rect 55220 15846 55272 15852
rect 55232 15502 55260 15846
rect 54496 15422 54800 15450
rect 55220 15496 55272 15502
rect 55220 15438 55272 15444
rect 54496 14618 54524 15422
rect 54576 15360 54628 15366
rect 54576 15302 54628 15308
rect 54484 14612 54536 14618
rect 54484 14554 54536 14560
rect 54024 13932 54076 13938
rect 54024 13874 54076 13880
rect 53932 13864 53984 13870
rect 53932 13806 53984 13812
rect 53748 12436 53800 12442
rect 53484 12406 53604 12434
rect 53472 11756 53524 11762
rect 53472 11698 53524 11704
rect 53380 11688 53432 11694
rect 53380 11630 53432 11636
rect 53392 7750 53420 11630
rect 53484 8634 53512 11698
rect 53576 10062 53604 12406
rect 53748 12378 53800 12384
rect 53760 11762 53788 12378
rect 53840 12368 53892 12374
rect 53840 12310 53892 12316
rect 53852 11762 53880 12310
rect 53748 11756 53800 11762
rect 53748 11698 53800 11704
rect 53840 11756 53892 11762
rect 53840 11698 53892 11704
rect 53852 10674 53880 11698
rect 53840 10668 53892 10674
rect 53840 10610 53892 10616
rect 53564 10056 53616 10062
rect 53564 9998 53616 10004
rect 53852 9722 53880 10610
rect 53944 10266 53972 13806
rect 54036 11150 54064 13874
rect 54116 12640 54168 12646
rect 54116 12582 54168 12588
rect 54128 12306 54156 12582
rect 54496 12434 54524 14554
rect 54588 14346 54616 15302
rect 54760 14476 54812 14482
rect 54760 14418 54812 14424
rect 54576 14340 54628 14346
rect 54576 14282 54628 14288
rect 54772 13870 54800 14418
rect 54760 13864 54812 13870
rect 54760 13806 54812 13812
rect 54496 12406 54616 12434
rect 54588 12374 54616 12406
rect 54576 12368 54628 12374
rect 54576 12310 54628 12316
rect 54116 12300 54168 12306
rect 54116 12242 54168 12248
rect 54484 12232 54536 12238
rect 54484 12174 54536 12180
rect 54392 12096 54444 12102
rect 54392 12038 54444 12044
rect 54404 11898 54432 12038
rect 54392 11892 54444 11898
rect 54392 11834 54444 11840
rect 54496 11354 54524 12174
rect 55128 12096 55180 12102
rect 55128 12038 55180 12044
rect 55140 11898 55168 12038
rect 55128 11892 55180 11898
rect 55128 11834 55180 11840
rect 54484 11348 54536 11354
rect 54484 11290 54536 11296
rect 54024 11144 54076 11150
rect 54024 11086 54076 11092
rect 53932 10260 53984 10266
rect 53932 10202 53984 10208
rect 54036 10146 54064 11086
rect 54668 11076 54720 11082
rect 54668 11018 54720 11024
rect 53944 10118 54064 10146
rect 53840 9716 53892 9722
rect 53840 9658 53892 9664
rect 53852 9042 53880 9658
rect 53840 9036 53892 9042
rect 53840 8978 53892 8984
rect 53852 8634 53880 8978
rect 53472 8628 53524 8634
rect 53472 8570 53524 8576
rect 53840 8628 53892 8634
rect 53840 8570 53892 8576
rect 53484 7886 53512 8570
rect 53944 8430 53972 10118
rect 54576 9376 54628 9382
rect 54576 9318 54628 9324
rect 54024 8900 54076 8906
rect 54024 8842 54076 8848
rect 53932 8424 53984 8430
rect 53932 8366 53984 8372
rect 53472 7880 53524 7886
rect 53472 7822 53524 7828
rect 53380 7744 53432 7750
rect 53380 7686 53432 7692
rect 53484 7546 53512 7822
rect 53564 7812 53616 7818
rect 53564 7754 53616 7760
rect 53576 7546 53604 7754
rect 53932 7744 53984 7750
rect 53932 7686 53984 7692
rect 53944 7546 53972 7686
rect 54036 7546 54064 8842
rect 54588 8838 54616 9318
rect 54680 8974 54708 11018
rect 55232 10810 55260 15438
rect 55508 15162 55536 17546
rect 55680 16040 55732 16046
rect 55680 15982 55732 15988
rect 55588 15360 55640 15366
rect 55588 15302 55640 15308
rect 55496 15156 55548 15162
rect 55496 15098 55548 15104
rect 55404 15020 55456 15026
rect 55404 14962 55456 14968
rect 55312 14272 55364 14278
rect 55312 14214 55364 14220
rect 55324 14074 55352 14214
rect 55416 14074 55444 14962
rect 55600 14482 55628 15302
rect 55692 14822 55720 15982
rect 55864 15904 55916 15910
rect 55864 15846 55916 15852
rect 55772 15360 55824 15366
rect 55772 15302 55824 15308
rect 55680 14816 55732 14822
rect 55680 14758 55732 14764
rect 55588 14476 55640 14482
rect 55588 14418 55640 14424
rect 55312 14068 55364 14074
rect 55312 14010 55364 14016
rect 55404 14068 55456 14074
rect 55404 14010 55456 14016
rect 55600 13954 55628 14418
rect 55784 14074 55812 15302
rect 55876 14346 55904 15846
rect 56060 15570 56088 17614
rect 56152 15706 56180 18158
rect 56428 17338 56456 18158
rect 56416 17332 56468 17338
rect 56416 17274 56468 17280
rect 56324 16992 56376 16998
rect 56324 16934 56376 16940
rect 56416 16992 56468 16998
rect 56416 16934 56468 16940
rect 56140 15700 56192 15706
rect 56140 15642 56192 15648
rect 56048 15564 56100 15570
rect 56048 15506 56100 15512
rect 56152 15314 56180 15642
rect 56336 15484 56364 16934
rect 56428 16794 56456 16934
rect 56416 16788 56468 16794
rect 56416 16730 56468 16736
rect 56336 15456 56456 15484
rect 56152 15286 56364 15314
rect 55956 14952 56008 14958
rect 55956 14894 56008 14900
rect 55968 14618 55996 14894
rect 56336 14890 56364 15286
rect 56140 14884 56192 14890
rect 56140 14826 56192 14832
rect 56324 14884 56376 14890
rect 56324 14826 56376 14832
rect 56152 14618 56180 14826
rect 55956 14612 56008 14618
rect 55956 14554 56008 14560
rect 56140 14612 56192 14618
rect 56140 14554 56192 14560
rect 55864 14340 55916 14346
rect 55864 14282 55916 14288
rect 55772 14068 55824 14074
rect 55772 14010 55824 14016
rect 55968 14006 55996 14554
rect 55956 14000 56008 14006
rect 55600 13926 55720 13954
rect 55956 13942 56008 13948
rect 55692 13870 55720 13926
rect 55680 13864 55732 13870
rect 55680 13806 55732 13812
rect 56324 13728 56376 13734
rect 56324 13670 56376 13676
rect 56336 13190 56364 13670
rect 55680 13184 55732 13190
rect 55680 13126 55732 13132
rect 56324 13184 56376 13190
rect 56324 13126 56376 13132
rect 55312 12232 55364 12238
rect 55312 12174 55364 12180
rect 55324 11801 55352 12174
rect 55310 11792 55366 11801
rect 55310 11727 55312 11736
rect 55364 11727 55366 11736
rect 55312 11698 55364 11704
rect 55692 11694 55720 13126
rect 56232 12980 56284 12986
rect 56232 12922 56284 12928
rect 55864 12368 55916 12374
rect 55864 12310 55916 12316
rect 55680 11688 55732 11694
rect 55586 11656 55642 11665
rect 55680 11630 55732 11636
rect 55586 11591 55642 11600
rect 55600 11558 55628 11591
rect 55588 11552 55640 11558
rect 55588 11494 55640 11500
rect 55876 11218 55904 12310
rect 55956 12096 56008 12102
rect 55956 12038 56008 12044
rect 56048 12096 56100 12102
rect 56048 12038 56100 12044
rect 55968 11354 55996 12038
rect 55956 11348 56008 11354
rect 55956 11290 56008 11296
rect 55496 11212 55548 11218
rect 55496 11154 55548 11160
rect 55864 11212 55916 11218
rect 55864 11154 55916 11160
rect 55220 10804 55272 10810
rect 55220 10746 55272 10752
rect 55312 10464 55364 10470
rect 55312 10406 55364 10412
rect 55220 9376 55272 9382
rect 55220 9318 55272 9324
rect 54668 8968 54720 8974
rect 54668 8910 54720 8916
rect 54116 8832 54168 8838
rect 54116 8774 54168 8780
rect 54300 8832 54352 8838
rect 54300 8774 54352 8780
rect 54576 8832 54628 8838
rect 54576 8774 54628 8780
rect 54128 8430 54156 8774
rect 54208 8560 54260 8566
rect 54208 8502 54260 8508
rect 54116 8424 54168 8430
rect 54116 8366 54168 8372
rect 53472 7540 53524 7546
rect 53472 7482 53524 7488
rect 53564 7540 53616 7546
rect 53564 7482 53616 7488
rect 53932 7540 53984 7546
rect 53932 7482 53984 7488
rect 54024 7540 54076 7546
rect 54024 7482 54076 7488
rect 54220 6866 54248 8502
rect 54208 6860 54260 6866
rect 54208 6802 54260 6808
rect 53288 6792 53340 6798
rect 53288 6734 53340 6740
rect 53300 4622 53328 6734
rect 54220 6662 54248 6802
rect 53932 6656 53984 6662
rect 53932 6598 53984 6604
rect 54116 6656 54168 6662
rect 54116 6598 54168 6604
rect 54208 6656 54260 6662
rect 54208 6598 54260 6604
rect 53748 6452 53800 6458
rect 53748 6394 53800 6400
rect 53760 5370 53788 6394
rect 53944 5710 53972 6598
rect 54024 6112 54076 6118
rect 54024 6054 54076 6060
rect 53932 5704 53984 5710
rect 53932 5646 53984 5652
rect 53748 5364 53800 5370
rect 53748 5306 53800 5312
rect 53656 5160 53708 5166
rect 53656 5102 53708 5108
rect 53288 4616 53340 4622
rect 53288 4558 53340 4564
rect 53300 3398 53328 4558
rect 53668 4049 53696 5102
rect 53760 4282 53788 5306
rect 53840 5024 53892 5030
rect 53840 4966 53892 4972
rect 53748 4276 53800 4282
rect 53748 4218 53800 4224
rect 53654 4040 53710 4049
rect 53654 3975 53710 3984
rect 53288 3392 53340 3398
rect 53288 3334 53340 3340
rect 53300 2650 53328 3334
rect 53668 3058 53696 3975
rect 53852 3602 53880 4966
rect 54036 4826 54064 6054
rect 54128 5370 54156 6598
rect 54208 5908 54260 5914
rect 54208 5850 54260 5856
rect 54116 5364 54168 5370
rect 54116 5306 54168 5312
rect 54220 5166 54248 5850
rect 54208 5160 54260 5166
rect 54208 5102 54260 5108
rect 54024 4820 54076 4826
rect 54024 4762 54076 4768
rect 54024 4616 54076 4622
rect 54024 4558 54076 4564
rect 54116 4616 54168 4622
rect 54116 4558 54168 4564
rect 54036 4214 54064 4558
rect 54024 4208 54076 4214
rect 54024 4150 54076 4156
rect 54128 4010 54156 4558
rect 54312 4026 54340 8774
rect 54392 8492 54444 8498
rect 54392 8434 54444 8440
rect 54404 7546 54432 8434
rect 54588 8430 54616 8774
rect 54576 8424 54628 8430
rect 54576 8366 54628 8372
rect 55036 8424 55088 8430
rect 55036 8366 55088 8372
rect 54668 8356 54720 8362
rect 54668 8298 54720 8304
rect 54484 8084 54536 8090
rect 54484 8026 54536 8032
rect 54392 7540 54444 7546
rect 54392 7482 54444 7488
rect 54496 7410 54524 8026
rect 54576 7948 54628 7954
rect 54576 7890 54628 7896
rect 54484 7404 54536 7410
rect 54484 7346 54536 7352
rect 54588 7002 54616 7890
rect 54680 7750 54708 8298
rect 55048 8090 55076 8366
rect 55036 8084 55088 8090
rect 55036 8026 55088 8032
rect 55232 7886 55260 9318
rect 55324 7954 55352 10406
rect 55508 9042 55536 11154
rect 55772 11008 55824 11014
rect 55772 10950 55824 10956
rect 55784 10266 55812 10950
rect 55876 10470 55904 11154
rect 55864 10464 55916 10470
rect 55864 10406 55916 10412
rect 55772 10260 55824 10266
rect 55772 10202 55824 10208
rect 55864 9444 55916 9450
rect 55864 9386 55916 9392
rect 55496 9036 55548 9042
rect 55496 8978 55548 8984
rect 55508 8838 55536 8978
rect 55772 8900 55824 8906
rect 55772 8842 55824 8848
rect 55496 8832 55548 8838
rect 55496 8774 55548 8780
rect 55588 8832 55640 8838
rect 55588 8774 55640 8780
rect 55404 8424 55456 8430
rect 55404 8366 55456 8372
rect 55416 8090 55444 8366
rect 55404 8084 55456 8090
rect 55404 8026 55456 8032
rect 55312 7948 55364 7954
rect 55312 7890 55364 7896
rect 55220 7880 55272 7886
rect 55220 7822 55272 7828
rect 54668 7744 54720 7750
rect 54668 7686 54720 7692
rect 54944 7744 54996 7750
rect 54944 7686 54996 7692
rect 54956 7313 54984 7686
rect 55324 7546 55352 7890
rect 55416 7546 55444 8026
rect 55508 7834 55536 8774
rect 55600 8022 55628 8774
rect 55784 8566 55812 8842
rect 55772 8560 55824 8566
rect 55772 8502 55824 8508
rect 55588 8016 55640 8022
rect 55588 7958 55640 7964
rect 55508 7806 55628 7834
rect 55600 7750 55628 7806
rect 55588 7744 55640 7750
rect 55588 7686 55640 7692
rect 55312 7540 55364 7546
rect 55312 7482 55364 7488
rect 55404 7540 55456 7546
rect 55404 7482 55456 7488
rect 55496 7472 55548 7478
rect 55496 7414 55548 7420
rect 54942 7304 54998 7313
rect 54942 7239 54998 7248
rect 54956 7018 54984 7239
rect 55508 7206 55536 7414
rect 55496 7200 55548 7206
rect 55496 7142 55548 7148
rect 54864 7002 54984 7018
rect 54576 6996 54628 7002
rect 54576 6938 54628 6944
rect 54864 6996 54996 7002
rect 54864 6990 54944 6996
rect 54484 5228 54536 5234
rect 54484 5170 54536 5176
rect 54116 4004 54168 4010
rect 54312 3998 54432 4026
rect 54116 3946 54168 3952
rect 54208 3936 54260 3942
rect 54208 3878 54260 3884
rect 54300 3936 54352 3942
rect 54300 3878 54352 3884
rect 54220 3738 54248 3878
rect 54208 3732 54260 3738
rect 54208 3674 54260 3680
rect 54312 3618 54340 3878
rect 54128 3602 54340 3618
rect 53840 3596 53892 3602
rect 53840 3538 53892 3544
rect 54116 3596 54340 3602
rect 54168 3590 54340 3596
rect 54116 3538 54168 3544
rect 54404 3194 54432 3998
rect 54392 3188 54444 3194
rect 54392 3130 54444 3136
rect 53656 3052 53708 3058
rect 53656 2994 53708 3000
rect 54208 2984 54260 2990
rect 54208 2926 54260 2932
rect 53378 2816 53434 2825
rect 53378 2751 53434 2760
rect 53288 2644 53340 2650
rect 53288 2586 53340 2592
rect 53196 2304 53248 2310
rect 53196 2246 53248 2252
rect 53392 800 53420 2751
rect 53944 870 54064 898
rect 53944 800 53972 870
rect 52932 734 53144 762
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54036 762 54064 870
rect 54220 762 54248 2926
rect 54496 800 54524 5170
rect 54576 4072 54628 4078
rect 54576 4014 54628 4020
rect 54588 3398 54616 4014
rect 54864 4010 54892 6990
rect 54944 6938 54996 6944
rect 55404 6996 55456 7002
rect 55404 6938 55456 6944
rect 54944 6860 54996 6866
rect 54944 6802 54996 6808
rect 54956 6322 54984 6802
rect 54944 6316 54996 6322
rect 54944 6258 54996 6264
rect 55036 6248 55088 6254
rect 55036 6190 55088 6196
rect 55048 5914 55076 6190
rect 55416 6186 55444 6938
rect 55312 6180 55364 6186
rect 55312 6122 55364 6128
rect 55404 6180 55456 6186
rect 55404 6122 55456 6128
rect 55324 5914 55352 6122
rect 55036 5908 55088 5914
rect 55036 5850 55088 5856
rect 55312 5908 55364 5914
rect 55312 5850 55364 5856
rect 55508 5710 55536 7142
rect 55128 5704 55180 5710
rect 55126 5672 55128 5681
rect 55496 5704 55548 5710
rect 55180 5672 55182 5681
rect 55036 5636 55088 5642
rect 55126 5607 55182 5616
rect 55416 5664 55496 5692
rect 55036 5578 55088 5584
rect 54944 5568 54996 5574
rect 54944 5510 54996 5516
rect 54852 4004 54904 4010
rect 54852 3946 54904 3952
rect 54576 3392 54628 3398
rect 54576 3334 54628 3340
rect 54588 3194 54616 3334
rect 54576 3188 54628 3194
rect 54576 3130 54628 3136
rect 54956 2446 54984 5510
rect 55048 3534 55076 5578
rect 55312 4480 55364 4486
rect 55312 4422 55364 4428
rect 55324 4321 55352 4422
rect 55310 4312 55366 4321
rect 55310 4247 55366 4256
rect 55416 4049 55444 5664
rect 55496 5646 55548 5652
rect 55600 5030 55628 7686
rect 55876 7478 55904 9386
rect 56060 8498 56088 12038
rect 56138 11656 56194 11665
rect 56138 11591 56140 11600
rect 56192 11591 56194 11600
rect 56140 11562 56192 11568
rect 56140 9512 56192 9518
rect 56140 9454 56192 9460
rect 56152 9178 56180 9454
rect 56140 9172 56192 9178
rect 56140 9114 56192 9120
rect 56244 9042 56272 12922
rect 56428 12434 56456 15456
rect 56508 13728 56560 13734
rect 56508 13670 56560 13676
rect 56520 13394 56548 13670
rect 56508 13388 56560 13394
rect 56508 13330 56560 13336
rect 56428 12406 56548 12434
rect 56232 9036 56284 9042
rect 56232 8978 56284 8984
rect 55956 8492 56008 8498
rect 55956 8434 56008 8440
rect 56048 8492 56100 8498
rect 56048 8434 56100 8440
rect 55968 7954 55996 8434
rect 56244 8090 56272 8978
rect 56324 8288 56376 8294
rect 56324 8230 56376 8236
rect 56336 8090 56364 8230
rect 56048 8084 56100 8090
rect 56048 8026 56100 8032
rect 56232 8084 56284 8090
rect 56232 8026 56284 8032
rect 56324 8084 56376 8090
rect 56324 8026 56376 8032
rect 55956 7948 56008 7954
rect 55956 7890 56008 7896
rect 55864 7472 55916 7478
rect 55864 7414 55916 7420
rect 55772 6656 55824 6662
rect 55772 6598 55824 6604
rect 55784 6322 55812 6598
rect 55772 6316 55824 6322
rect 55772 6258 55824 6264
rect 55784 6118 55812 6258
rect 55772 6112 55824 6118
rect 55772 6054 55824 6060
rect 55864 6112 55916 6118
rect 55864 6054 55916 6060
rect 55876 5710 55904 6054
rect 55864 5704 55916 5710
rect 55864 5646 55916 5652
rect 55680 5160 55732 5166
rect 55680 5102 55732 5108
rect 55588 5024 55640 5030
rect 55588 4966 55640 4972
rect 55496 4072 55548 4078
rect 55402 4040 55458 4049
rect 55496 4014 55548 4020
rect 55402 3975 55458 3984
rect 55508 3942 55536 4014
rect 55600 3942 55628 4966
rect 55692 4282 55720 5102
rect 56060 4622 56088 8026
rect 56416 7948 56468 7954
rect 56416 7890 56468 7896
rect 56232 7540 56284 7546
rect 56232 7482 56284 7488
rect 56244 6934 56272 7482
rect 56232 6928 56284 6934
rect 56152 6888 56232 6916
rect 56152 6254 56180 6888
rect 56232 6870 56284 6876
rect 56428 6866 56456 7890
rect 56416 6860 56468 6866
rect 56416 6802 56468 6808
rect 56140 6248 56192 6254
rect 56140 6190 56192 6196
rect 56048 4616 56100 4622
rect 56048 4558 56100 4564
rect 55772 4480 55824 4486
rect 55772 4422 55824 4428
rect 55680 4276 55732 4282
rect 55680 4218 55732 4224
rect 55496 3936 55548 3942
rect 55496 3878 55548 3884
rect 55588 3936 55640 3942
rect 55588 3878 55640 3884
rect 55036 3528 55088 3534
rect 55036 3470 55088 3476
rect 55312 3528 55364 3534
rect 55312 3470 55364 3476
rect 55128 3392 55180 3398
rect 55128 3334 55180 3340
rect 55140 2961 55168 3334
rect 55126 2952 55182 2961
rect 55036 2916 55088 2922
rect 55126 2887 55182 2896
rect 55036 2858 55088 2864
rect 54944 2440 54996 2446
rect 54944 2382 54996 2388
rect 55048 800 55076 2858
rect 55324 2650 55352 3470
rect 55784 3194 55812 4422
rect 56152 4010 56180 6190
rect 56520 5658 56548 12406
rect 56612 6254 56640 19450
rect 57428 19304 57480 19310
rect 57428 19246 57480 19252
rect 56784 19168 56836 19174
rect 56784 19110 56836 19116
rect 56692 18216 56744 18222
rect 56692 18158 56744 18164
rect 56704 17678 56732 18158
rect 56692 17672 56744 17678
rect 56692 17614 56744 17620
rect 56692 17332 56744 17338
rect 56692 17274 56744 17280
rect 56704 16794 56732 17274
rect 56692 16788 56744 16794
rect 56692 16730 56744 16736
rect 56796 16182 56824 19110
rect 57440 18426 57468 19246
rect 57428 18420 57480 18426
rect 57428 18362 57480 18368
rect 57428 18080 57480 18086
rect 57428 18022 57480 18028
rect 57440 17882 57468 18022
rect 57428 17876 57480 17882
rect 57428 17818 57480 17824
rect 56876 17672 56928 17678
rect 56876 17614 56928 17620
rect 56784 16176 56836 16182
rect 56784 16118 56836 16124
rect 56888 15026 56916 17614
rect 57060 17604 57112 17610
rect 57060 17546 57112 17552
rect 57072 16794 57100 17546
rect 57440 17134 57468 17818
rect 57520 17740 57572 17746
rect 57520 17682 57572 17688
rect 57428 17128 57480 17134
rect 57428 17070 57480 17076
rect 57428 16992 57480 16998
rect 57532 16946 57560 17682
rect 57808 17542 57836 20810
rect 58176 20602 58204 20946
rect 58726 20700 59034 20709
rect 58726 20698 58732 20700
rect 58788 20698 58812 20700
rect 58868 20698 58892 20700
rect 58948 20698 58972 20700
rect 59028 20698 59034 20700
rect 58788 20646 58790 20698
rect 58970 20646 58972 20698
rect 58726 20644 58732 20646
rect 58788 20644 58812 20646
rect 58868 20644 58892 20646
rect 58948 20644 58972 20646
rect 59028 20644 59034 20646
rect 58726 20635 59034 20644
rect 58164 20596 58216 20602
rect 58164 20538 58216 20544
rect 58726 19612 59034 19621
rect 58726 19610 58732 19612
rect 58788 19610 58812 19612
rect 58868 19610 58892 19612
rect 58948 19610 58972 19612
rect 59028 19610 59034 19612
rect 58788 19558 58790 19610
rect 58970 19558 58972 19610
rect 58726 19556 58732 19558
rect 58788 19556 58812 19558
rect 58868 19556 58892 19558
rect 58948 19556 58972 19558
rect 59028 19556 59034 19558
rect 58726 19547 59034 19556
rect 58164 19372 58216 19378
rect 58164 19314 58216 19320
rect 57888 19168 57940 19174
rect 57888 19110 57940 19116
rect 57900 18970 57928 19110
rect 57888 18964 57940 18970
rect 57888 18906 57940 18912
rect 57888 18216 57940 18222
rect 57888 18158 57940 18164
rect 57900 17882 57928 18158
rect 57888 17876 57940 17882
rect 57888 17818 57940 17824
rect 58176 17678 58204 19314
rect 58532 18692 58584 18698
rect 58532 18634 58584 18640
rect 58544 18426 58572 18634
rect 58726 18524 59034 18533
rect 58726 18522 58732 18524
rect 58788 18522 58812 18524
rect 58868 18522 58892 18524
rect 58948 18522 58972 18524
rect 59028 18522 59034 18524
rect 58788 18470 58790 18522
rect 58970 18470 58972 18522
rect 58726 18468 58732 18470
rect 58788 18468 58812 18470
rect 58868 18468 58892 18470
rect 58948 18468 58972 18470
rect 59028 18468 59034 18470
rect 58726 18459 59034 18468
rect 58532 18420 58584 18426
rect 58532 18362 58584 18368
rect 58164 17672 58216 17678
rect 58164 17614 58216 17620
rect 57796 17536 57848 17542
rect 57796 17478 57848 17484
rect 58440 17536 58492 17542
rect 58440 17478 58492 17484
rect 58452 17338 58480 17478
rect 58726 17436 59034 17445
rect 58726 17434 58732 17436
rect 58788 17434 58812 17436
rect 58868 17434 58892 17436
rect 58948 17434 58972 17436
rect 59028 17434 59034 17436
rect 58788 17382 58790 17434
rect 58970 17382 58972 17434
rect 58726 17380 58732 17382
rect 58788 17380 58812 17382
rect 58868 17380 58892 17382
rect 58948 17380 58972 17382
rect 59028 17380 59034 17382
rect 58726 17371 59034 17380
rect 58440 17332 58492 17338
rect 58440 17274 58492 17280
rect 57480 16940 57560 16946
rect 57428 16934 57560 16940
rect 57440 16918 57560 16934
rect 57060 16788 57112 16794
rect 57060 16730 57112 16736
rect 57336 15360 57388 15366
rect 57336 15302 57388 15308
rect 57348 15162 57376 15302
rect 57336 15156 57388 15162
rect 57336 15098 57388 15104
rect 56876 15020 56928 15026
rect 56876 14962 56928 14968
rect 56692 14952 56744 14958
rect 56692 14894 56744 14900
rect 56704 14822 56732 14894
rect 56692 14816 56744 14822
rect 56692 14758 56744 14764
rect 57336 14476 57388 14482
rect 57336 14418 57388 14424
rect 57152 14340 57204 14346
rect 57152 14282 57204 14288
rect 56876 14272 56928 14278
rect 56876 14214 56928 14220
rect 56888 14074 56916 14214
rect 56876 14068 56928 14074
rect 56876 14010 56928 14016
rect 56692 13864 56744 13870
rect 56692 13806 56744 13812
rect 56704 12986 56732 13806
rect 57164 13530 57192 14282
rect 57348 13870 57376 14418
rect 57336 13864 57388 13870
rect 57336 13806 57388 13812
rect 57152 13524 57204 13530
rect 57152 13466 57204 13472
rect 56692 12980 56744 12986
rect 56692 12922 56744 12928
rect 56704 12866 56732 12922
rect 56704 12838 56916 12866
rect 56692 12640 56744 12646
rect 56692 12582 56744 12588
rect 56704 12238 56732 12582
rect 56888 12434 56916 12838
rect 57348 12442 57376 13806
rect 57336 12436 57388 12442
rect 56888 12406 57008 12434
rect 56692 12232 56744 12238
rect 56692 12174 56744 12180
rect 56782 11792 56838 11801
rect 56692 11756 56744 11762
rect 56782 11727 56784 11736
rect 56692 11698 56744 11704
rect 56836 11727 56838 11736
rect 56784 11698 56836 11704
rect 56704 10810 56732 11698
rect 56876 11280 56928 11286
rect 56876 11222 56928 11228
rect 56888 11121 56916 11222
rect 56874 11112 56930 11121
rect 56874 11047 56930 11056
rect 56980 11014 57008 12406
rect 57336 12378 57388 12384
rect 57336 12164 57388 12170
rect 57336 12106 57388 12112
rect 57152 12096 57204 12102
rect 57152 12038 57204 12044
rect 57164 11558 57192 12038
rect 57348 11694 57376 12106
rect 57336 11688 57388 11694
rect 57336 11630 57388 11636
rect 57152 11552 57204 11558
rect 57152 11494 57204 11500
rect 56784 11008 56836 11014
rect 56784 10950 56836 10956
rect 56968 11008 57020 11014
rect 56968 10950 57020 10956
rect 56692 10804 56744 10810
rect 56692 10746 56744 10752
rect 56704 10130 56732 10746
rect 56796 10742 56824 10950
rect 56784 10736 56836 10742
rect 56784 10678 56836 10684
rect 56692 10124 56744 10130
rect 56692 10066 56744 10072
rect 56980 9926 57008 10950
rect 56876 9920 56928 9926
rect 56876 9862 56928 9868
rect 56968 9920 57020 9926
rect 56968 9862 57020 9868
rect 56888 9382 56916 9862
rect 57440 9466 57468 16918
rect 57888 16040 57940 16046
rect 57888 15982 57940 15988
rect 57900 15366 57928 15982
rect 57980 15904 58032 15910
rect 57980 15846 58032 15852
rect 57888 15360 57940 15366
rect 57888 15302 57940 15308
rect 57888 14952 57940 14958
rect 57888 14894 57940 14900
rect 57520 14816 57572 14822
rect 57520 14758 57572 14764
rect 57532 11150 57560 14758
rect 57900 14618 57928 14894
rect 57888 14612 57940 14618
rect 57888 14554 57940 14560
rect 57704 14544 57756 14550
rect 57704 14486 57756 14492
rect 57716 13870 57744 14486
rect 57992 14414 58020 15846
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 57704 13864 57756 13870
rect 57704 13806 57756 13812
rect 57796 12776 57848 12782
rect 57796 12718 57848 12724
rect 57808 12102 57836 12718
rect 58452 12442 58480 17274
rect 58726 16348 59034 16357
rect 58726 16346 58732 16348
rect 58788 16346 58812 16348
rect 58868 16346 58892 16348
rect 58948 16346 58972 16348
rect 59028 16346 59034 16348
rect 58788 16294 58790 16346
rect 58970 16294 58972 16346
rect 58726 16292 58732 16294
rect 58788 16292 58812 16294
rect 58868 16292 58892 16294
rect 58948 16292 58972 16294
rect 59028 16292 59034 16294
rect 58726 16283 59034 16292
rect 58532 15428 58584 15434
rect 58532 15370 58584 15376
rect 58544 15162 58572 15370
rect 58726 15260 59034 15269
rect 58726 15258 58732 15260
rect 58788 15258 58812 15260
rect 58868 15258 58892 15260
rect 58948 15258 58972 15260
rect 59028 15258 59034 15260
rect 58788 15206 58790 15258
rect 58970 15206 58972 15258
rect 58726 15204 58732 15206
rect 58788 15204 58812 15206
rect 58868 15204 58892 15206
rect 58948 15204 58972 15206
rect 59028 15204 59034 15206
rect 58726 15195 59034 15204
rect 58532 15156 58584 15162
rect 58532 15098 58584 15104
rect 58726 14172 59034 14181
rect 58726 14170 58732 14172
rect 58788 14170 58812 14172
rect 58868 14170 58892 14172
rect 58948 14170 58972 14172
rect 59028 14170 59034 14172
rect 58788 14118 58790 14170
rect 58970 14118 58972 14170
rect 58726 14116 58732 14118
rect 58788 14116 58812 14118
rect 58868 14116 58892 14118
rect 58948 14116 58972 14118
rect 59028 14116 59034 14118
rect 58726 14107 59034 14116
rect 58726 13084 59034 13093
rect 58726 13082 58732 13084
rect 58788 13082 58812 13084
rect 58868 13082 58892 13084
rect 58948 13082 58972 13084
rect 59028 13082 59034 13084
rect 58788 13030 58790 13082
rect 58970 13030 58972 13082
rect 58726 13028 58732 13030
rect 58788 13028 58812 13030
rect 58868 13028 58892 13030
rect 58948 13028 58972 13030
rect 59028 13028 59034 13030
rect 58726 13019 59034 13028
rect 58440 12436 58492 12442
rect 58440 12378 58492 12384
rect 57888 12368 57940 12374
rect 57888 12310 57940 12316
rect 57796 12096 57848 12102
rect 57796 12038 57848 12044
rect 57704 11892 57756 11898
rect 57704 11834 57756 11840
rect 57612 11552 57664 11558
rect 57612 11494 57664 11500
rect 57624 11150 57652 11494
rect 57520 11144 57572 11150
rect 57520 11086 57572 11092
rect 57612 11144 57664 11150
rect 57612 11086 57664 11092
rect 57716 10810 57744 11834
rect 57900 10826 57928 12310
rect 58256 12164 58308 12170
rect 58256 12106 58308 12112
rect 57704 10804 57756 10810
rect 57900 10798 58020 10826
rect 57704 10746 57756 10752
rect 57716 10130 57744 10746
rect 57888 10600 57940 10606
rect 57888 10542 57940 10548
rect 57900 10266 57928 10542
rect 57888 10260 57940 10266
rect 57888 10202 57940 10208
rect 57704 10124 57756 10130
rect 57704 10066 57756 10072
rect 57704 9920 57756 9926
rect 57704 9862 57756 9868
rect 56980 9438 57468 9466
rect 56784 9376 56836 9382
rect 56784 9318 56836 9324
rect 56876 9376 56928 9382
rect 56876 9318 56928 9324
rect 56796 8634 56824 9318
rect 56876 9172 56928 9178
rect 56876 9114 56928 9120
rect 56888 8634 56916 9114
rect 56784 8628 56836 8634
rect 56784 8570 56836 8576
rect 56876 8628 56928 8634
rect 56876 8570 56928 8576
rect 56876 7540 56928 7546
rect 56876 7482 56928 7488
rect 56692 7336 56744 7342
rect 56692 7278 56744 7284
rect 56704 6798 56732 7278
rect 56784 7200 56836 7206
rect 56784 7142 56836 7148
rect 56692 6792 56744 6798
rect 56692 6734 56744 6740
rect 56796 6610 56824 7142
rect 56704 6582 56824 6610
rect 56600 6248 56652 6254
rect 56600 6190 56652 6196
rect 56600 6112 56652 6118
rect 56600 6054 56652 6060
rect 56428 5630 56548 5658
rect 56324 5160 56376 5166
rect 56428 5137 56456 5630
rect 56508 5568 56560 5574
rect 56508 5510 56560 5516
rect 56324 5102 56376 5108
rect 56414 5128 56470 5137
rect 56232 5024 56284 5030
rect 56232 4966 56284 4972
rect 56244 4622 56272 4966
rect 56336 4826 56364 5102
rect 56414 5063 56470 5072
rect 56520 4826 56548 5510
rect 56324 4820 56376 4826
rect 56324 4762 56376 4768
rect 56508 4820 56560 4826
rect 56508 4762 56560 4768
rect 56232 4616 56284 4622
rect 56232 4558 56284 4564
rect 56612 4282 56640 6054
rect 56704 5234 56732 6582
rect 56888 6458 56916 7482
rect 56876 6452 56928 6458
rect 56876 6394 56928 6400
rect 56784 6316 56836 6322
rect 56784 6258 56836 6264
rect 56796 5574 56824 6258
rect 56784 5568 56836 5574
rect 56784 5510 56836 5516
rect 56692 5228 56744 5234
rect 56692 5170 56744 5176
rect 56692 5092 56744 5098
rect 56692 5034 56744 5040
rect 56600 4276 56652 4282
rect 56600 4218 56652 4224
rect 56416 4140 56468 4146
rect 56416 4082 56468 4088
rect 56428 4026 56456 4082
rect 56140 4004 56192 4010
rect 56140 3946 56192 3952
rect 56336 3998 56456 4026
rect 56598 4040 56654 4049
rect 56336 3942 56364 3998
rect 56598 3975 56654 3984
rect 56612 3942 56640 3975
rect 56324 3936 56376 3942
rect 56324 3878 56376 3884
rect 56416 3936 56468 3942
rect 56416 3878 56468 3884
rect 56600 3936 56652 3942
rect 56600 3878 56652 3884
rect 55772 3188 55824 3194
rect 55772 3130 55824 3136
rect 56324 3188 56376 3194
rect 56324 3130 56376 3136
rect 55404 2848 55456 2854
rect 55404 2790 55456 2796
rect 55312 2644 55364 2650
rect 55312 2586 55364 2592
rect 55416 2446 55444 2790
rect 55588 2508 55640 2514
rect 55588 2450 55640 2456
rect 55404 2440 55456 2446
rect 55404 2382 55456 2388
rect 55600 800 55628 2450
rect 56336 1850 56364 3130
rect 56428 2650 56456 3878
rect 56416 2644 56468 2650
rect 56416 2586 56468 2592
rect 56152 1822 56364 1850
rect 56152 800 56180 1822
rect 56704 800 56732 5034
rect 56796 4690 56824 5510
rect 56784 4684 56836 4690
rect 56784 4626 56836 4632
rect 56888 3602 56916 6394
rect 56980 5273 57008 9438
rect 57060 9376 57112 9382
rect 57060 9318 57112 9324
rect 57428 9376 57480 9382
rect 57428 9318 57480 9324
rect 57072 9042 57100 9318
rect 57336 9104 57388 9110
rect 57336 9046 57388 9052
rect 57060 9036 57112 9042
rect 57060 8978 57112 8984
rect 57072 7206 57100 8978
rect 57348 8634 57376 9046
rect 57336 8628 57388 8634
rect 57336 8570 57388 8576
rect 57440 7546 57468 9318
rect 57612 8968 57664 8974
rect 57612 8910 57664 8916
rect 57520 8356 57572 8362
rect 57520 8298 57572 8304
rect 57532 7886 57560 8298
rect 57624 8090 57652 8910
rect 57612 8084 57664 8090
rect 57612 8026 57664 8032
rect 57520 7880 57572 7886
rect 57520 7822 57572 7828
rect 57716 7546 57744 9862
rect 57992 9654 58020 10798
rect 57980 9648 58032 9654
rect 57980 9590 58032 9596
rect 57428 7540 57480 7546
rect 57428 7482 57480 7488
rect 57704 7540 57756 7546
rect 57704 7482 57756 7488
rect 57060 7200 57112 7206
rect 57060 7142 57112 7148
rect 57704 7200 57756 7206
rect 57704 7142 57756 7148
rect 57336 6792 57388 6798
rect 57336 6734 57388 6740
rect 57242 6624 57298 6633
rect 57348 6610 57376 6734
rect 57298 6582 57376 6610
rect 57242 6559 57298 6568
rect 57256 6254 57284 6559
rect 57152 6248 57204 6254
rect 57152 6190 57204 6196
rect 57244 6248 57296 6254
rect 57244 6190 57296 6196
rect 57060 5908 57112 5914
rect 57060 5850 57112 5856
rect 56966 5264 57022 5273
rect 57072 5234 57100 5850
rect 57164 5370 57192 6190
rect 57520 6112 57572 6118
rect 57520 6054 57572 6060
rect 57428 5908 57480 5914
rect 57428 5850 57480 5856
rect 57152 5364 57204 5370
rect 57152 5306 57204 5312
rect 57440 5234 57468 5850
rect 57532 5778 57560 6054
rect 57520 5772 57572 5778
rect 57520 5714 57572 5720
rect 57716 5710 57744 7142
rect 57796 6316 57848 6322
rect 57796 6258 57848 6264
rect 57704 5704 57756 5710
rect 57704 5646 57756 5652
rect 56966 5199 57022 5208
rect 57060 5228 57112 5234
rect 57060 5170 57112 5176
rect 57428 5228 57480 5234
rect 57428 5170 57480 5176
rect 57060 5092 57112 5098
rect 57060 5034 57112 5040
rect 56968 5024 57020 5030
rect 56968 4966 57020 4972
rect 56876 3596 56928 3602
rect 56876 3538 56928 3544
rect 56980 3534 57008 4966
rect 57072 4690 57100 5034
rect 57060 4684 57112 4690
rect 57060 4626 57112 4632
rect 57152 4072 57204 4078
rect 57150 4040 57152 4049
rect 57244 4072 57296 4078
rect 57204 4040 57206 4049
rect 57244 4014 57296 4020
rect 57150 3975 57206 3984
rect 57256 3942 57284 4014
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 57612 3936 57664 3942
rect 57612 3878 57664 3884
rect 57256 3584 57284 3878
rect 57164 3556 57284 3584
rect 56968 3528 57020 3534
rect 56968 3470 57020 3476
rect 57164 2446 57192 3556
rect 57428 3528 57480 3534
rect 57428 3470 57480 3476
rect 57440 3194 57468 3470
rect 57624 3194 57652 3878
rect 57428 3188 57480 3194
rect 57428 3130 57480 3136
rect 57612 3188 57664 3194
rect 57612 3130 57664 3136
rect 57244 2984 57296 2990
rect 57244 2926 57296 2932
rect 57152 2440 57204 2446
rect 57152 2382 57204 2388
rect 57256 800 57284 2926
rect 57808 800 57836 6258
rect 57992 5778 58020 9590
rect 58072 9376 58124 9382
rect 58072 9318 58124 9324
rect 58084 8634 58112 9318
rect 58072 8628 58124 8634
rect 58072 8570 58124 8576
rect 58072 7200 58124 7206
rect 58072 7142 58124 7148
rect 58084 6798 58112 7142
rect 58072 6792 58124 6798
rect 58072 6734 58124 6740
rect 58268 6662 58296 12106
rect 58726 11996 59034 12005
rect 58726 11994 58732 11996
rect 58788 11994 58812 11996
rect 58868 11994 58892 11996
rect 58948 11994 58972 11996
rect 59028 11994 59034 11996
rect 58788 11942 58790 11994
rect 58970 11942 58972 11994
rect 58726 11940 58732 11942
rect 58788 11940 58812 11942
rect 58868 11940 58892 11942
rect 58948 11940 58972 11942
rect 59028 11940 59034 11942
rect 58726 11931 59034 11940
rect 58726 10908 59034 10917
rect 58726 10906 58732 10908
rect 58788 10906 58812 10908
rect 58868 10906 58892 10908
rect 58948 10906 58972 10908
rect 59028 10906 59034 10908
rect 58788 10854 58790 10906
rect 58970 10854 58972 10906
rect 58726 10852 58732 10854
rect 58788 10852 58812 10854
rect 58868 10852 58892 10854
rect 58948 10852 58972 10854
rect 59028 10852 59034 10854
rect 58726 10843 59034 10852
rect 58726 9820 59034 9829
rect 58726 9818 58732 9820
rect 58788 9818 58812 9820
rect 58868 9818 58892 9820
rect 58948 9818 58972 9820
rect 59028 9818 59034 9820
rect 58788 9766 58790 9818
rect 58970 9766 58972 9818
rect 58726 9764 58732 9766
rect 58788 9764 58812 9766
rect 58868 9764 58892 9766
rect 58948 9764 58972 9766
rect 59028 9764 59034 9766
rect 58726 9755 59034 9764
rect 58726 8732 59034 8741
rect 58726 8730 58732 8732
rect 58788 8730 58812 8732
rect 58868 8730 58892 8732
rect 58948 8730 58972 8732
rect 59028 8730 59034 8732
rect 58788 8678 58790 8730
rect 58970 8678 58972 8730
rect 58726 8676 58732 8678
rect 58788 8676 58812 8678
rect 58868 8676 58892 8678
rect 58948 8676 58972 8678
rect 59028 8676 59034 8678
rect 58726 8667 59034 8676
rect 58726 7644 59034 7653
rect 58726 7642 58732 7644
rect 58788 7642 58812 7644
rect 58868 7642 58892 7644
rect 58948 7642 58972 7644
rect 59028 7642 59034 7644
rect 58788 7590 58790 7642
rect 58970 7590 58972 7642
rect 58726 7588 58732 7590
rect 58788 7588 58812 7590
rect 58868 7588 58892 7590
rect 58948 7588 58972 7590
rect 59028 7588 59034 7590
rect 58726 7579 59034 7588
rect 58348 7404 58400 7410
rect 58348 7346 58400 7352
rect 58256 6656 58308 6662
rect 58256 6598 58308 6604
rect 58360 5914 58388 7346
rect 58440 6792 58492 6798
rect 58440 6734 58492 6740
rect 58348 5908 58400 5914
rect 58348 5850 58400 5856
rect 57980 5772 58032 5778
rect 57980 5714 58032 5720
rect 57888 5704 57940 5710
rect 57888 5646 57940 5652
rect 57978 5672 58034 5681
rect 57900 5370 57928 5646
rect 57978 5607 58034 5616
rect 57888 5364 57940 5370
rect 57888 5306 57940 5312
rect 57886 4312 57942 4321
rect 57886 4247 57942 4256
rect 57900 4146 57928 4247
rect 57888 4140 57940 4146
rect 57888 4082 57940 4088
rect 57992 3194 58020 5607
rect 58256 3936 58308 3942
rect 58452 3913 58480 6734
rect 58532 6724 58584 6730
rect 58532 6666 58584 6672
rect 58544 5370 58572 6666
rect 58726 6556 59034 6565
rect 58726 6554 58732 6556
rect 58788 6554 58812 6556
rect 58868 6554 58892 6556
rect 58948 6554 58972 6556
rect 59028 6554 59034 6556
rect 58788 6502 58790 6554
rect 58970 6502 58972 6554
rect 58726 6500 58732 6502
rect 58788 6500 58812 6502
rect 58868 6500 58892 6502
rect 58948 6500 58972 6502
rect 59028 6500 59034 6502
rect 58726 6491 59034 6500
rect 58726 5468 59034 5477
rect 58726 5466 58732 5468
rect 58788 5466 58812 5468
rect 58868 5466 58892 5468
rect 58948 5466 58972 5468
rect 59028 5466 59034 5468
rect 58788 5414 58790 5466
rect 58970 5414 58972 5466
rect 58726 5412 58732 5414
rect 58788 5412 58812 5414
rect 58868 5412 58892 5414
rect 58948 5412 58972 5414
rect 59028 5412 59034 5414
rect 58726 5403 59034 5412
rect 58532 5364 58584 5370
rect 58532 5306 58584 5312
rect 59084 4548 59136 4554
rect 59084 4490 59136 4496
rect 58532 4480 58584 4486
rect 58532 4422 58584 4428
rect 58256 3878 58308 3884
rect 58438 3904 58494 3913
rect 58268 3670 58296 3878
rect 58438 3839 58494 3848
rect 58256 3664 58308 3670
rect 58256 3606 58308 3612
rect 58346 3496 58402 3505
rect 58346 3431 58402 3440
rect 57980 3188 58032 3194
rect 57980 3130 58032 3136
rect 57886 2816 57942 2825
rect 57886 2751 57942 2760
rect 57900 2514 57928 2751
rect 57888 2508 57940 2514
rect 57888 2450 57940 2456
rect 58360 800 58388 3431
rect 58544 2650 58572 4422
rect 58726 4380 59034 4389
rect 58726 4378 58732 4380
rect 58788 4378 58812 4380
rect 58868 4378 58892 4380
rect 58948 4378 58972 4380
rect 59028 4378 59034 4380
rect 58788 4326 58790 4378
rect 58970 4326 58972 4378
rect 58726 4324 58732 4326
rect 58788 4324 58812 4326
rect 58868 4324 58892 4326
rect 58948 4324 58972 4326
rect 59028 4324 59034 4326
rect 58726 4315 59034 4324
rect 58726 3292 59034 3301
rect 58726 3290 58732 3292
rect 58788 3290 58812 3292
rect 58868 3290 58892 3292
rect 58948 3290 58972 3292
rect 59028 3290 59034 3292
rect 58788 3238 58790 3290
rect 58970 3238 58972 3290
rect 58726 3236 58732 3238
rect 58788 3236 58812 3238
rect 58868 3236 58892 3238
rect 58948 3236 58972 3238
rect 59028 3236 59034 3238
rect 58726 3227 59034 3236
rect 58532 2644 58584 2650
rect 58532 2586 58584 2592
rect 58726 2204 59034 2213
rect 58726 2202 58732 2204
rect 58788 2202 58812 2204
rect 58868 2202 58892 2204
rect 58948 2202 58972 2204
rect 59028 2202 59034 2204
rect 58788 2150 58790 2202
rect 58970 2150 58972 2202
rect 58726 2148 58732 2150
rect 58788 2148 58812 2150
rect 58868 2148 58892 2150
rect 58948 2148 58972 2150
rect 59028 2148 59034 2150
rect 58726 2139 59034 2148
rect 59096 1986 59124 4490
rect 58912 1958 59124 1986
rect 58912 800 58940 1958
rect 54036 734 54248 762
rect 54482 0 54538 800
rect 55034 0 55090 800
rect 55586 0 55642 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58898 0 58954 800
<< via2 >>
rect 8178 27770 8234 27772
rect 8258 27770 8314 27772
rect 8338 27770 8394 27772
rect 8418 27770 8474 27772
rect 8178 27718 8224 27770
rect 8224 27718 8234 27770
rect 8258 27718 8288 27770
rect 8288 27718 8300 27770
rect 8300 27718 8314 27770
rect 8338 27718 8352 27770
rect 8352 27718 8364 27770
rect 8364 27718 8394 27770
rect 8418 27718 8428 27770
rect 8428 27718 8474 27770
rect 8178 27716 8234 27718
rect 8258 27716 8314 27718
rect 8338 27716 8394 27718
rect 8418 27716 8474 27718
rect 22622 27770 22678 27772
rect 22702 27770 22758 27772
rect 22782 27770 22838 27772
rect 22862 27770 22918 27772
rect 22622 27718 22668 27770
rect 22668 27718 22678 27770
rect 22702 27718 22732 27770
rect 22732 27718 22744 27770
rect 22744 27718 22758 27770
rect 22782 27718 22796 27770
rect 22796 27718 22808 27770
rect 22808 27718 22838 27770
rect 22862 27718 22872 27770
rect 22872 27718 22918 27770
rect 22622 27716 22678 27718
rect 22702 27716 22758 27718
rect 22782 27716 22838 27718
rect 22862 27716 22918 27718
rect 37066 27770 37122 27772
rect 37146 27770 37202 27772
rect 37226 27770 37282 27772
rect 37306 27770 37362 27772
rect 37066 27718 37112 27770
rect 37112 27718 37122 27770
rect 37146 27718 37176 27770
rect 37176 27718 37188 27770
rect 37188 27718 37202 27770
rect 37226 27718 37240 27770
rect 37240 27718 37252 27770
rect 37252 27718 37282 27770
rect 37306 27718 37316 27770
rect 37316 27718 37362 27770
rect 37066 27716 37122 27718
rect 37146 27716 37202 27718
rect 37226 27716 37282 27718
rect 37306 27716 37362 27718
rect 51510 27770 51566 27772
rect 51590 27770 51646 27772
rect 51670 27770 51726 27772
rect 51750 27770 51806 27772
rect 51510 27718 51556 27770
rect 51556 27718 51566 27770
rect 51590 27718 51620 27770
rect 51620 27718 51632 27770
rect 51632 27718 51646 27770
rect 51670 27718 51684 27770
rect 51684 27718 51696 27770
rect 51696 27718 51726 27770
rect 51750 27718 51760 27770
rect 51760 27718 51806 27770
rect 51510 27716 51566 27718
rect 51590 27716 51646 27718
rect 51670 27716 51726 27718
rect 51750 27716 51806 27718
rect 15400 27226 15456 27228
rect 15480 27226 15536 27228
rect 15560 27226 15616 27228
rect 15640 27226 15696 27228
rect 15400 27174 15446 27226
rect 15446 27174 15456 27226
rect 15480 27174 15510 27226
rect 15510 27174 15522 27226
rect 15522 27174 15536 27226
rect 15560 27174 15574 27226
rect 15574 27174 15586 27226
rect 15586 27174 15616 27226
rect 15640 27174 15650 27226
rect 15650 27174 15696 27226
rect 15400 27172 15456 27174
rect 15480 27172 15536 27174
rect 15560 27172 15616 27174
rect 15640 27172 15696 27174
rect 29844 27226 29900 27228
rect 29924 27226 29980 27228
rect 30004 27226 30060 27228
rect 30084 27226 30140 27228
rect 29844 27174 29890 27226
rect 29890 27174 29900 27226
rect 29924 27174 29954 27226
rect 29954 27174 29966 27226
rect 29966 27174 29980 27226
rect 30004 27174 30018 27226
rect 30018 27174 30030 27226
rect 30030 27174 30060 27226
rect 30084 27174 30094 27226
rect 30094 27174 30140 27226
rect 29844 27172 29900 27174
rect 29924 27172 29980 27174
rect 30004 27172 30060 27174
rect 30084 27172 30140 27174
rect 44288 27226 44344 27228
rect 44368 27226 44424 27228
rect 44448 27226 44504 27228
rect 44528 27226 44584 27228
rect 44288 27174 44334 27226
rect 44334 27174 44344 27226
rect 44368 27174 44398 27226
rect 44398 27174 44410 27226
rect 44410 27174 44424 27226
rect 44448 27174 44462 27226
rect 44462 27174 44474 27226
rect 44474 27174 44504 27226
rect 44528 27174 44538 27226
rect 44538 27174 44584 27226
rect 44288 27172 44344 27174
rect 44368 27172 44424 27174
rect 44448 27172 44504 27174
rect 44528 27172 44584 27174
rect 58732 27226 58788 27228
rect 58812 27226 58868 27228
rect 58892 27226 58948 27228
rect 58972 27226 59028 27228
rect 58732 27174 58778 27226
rect 58778 27174 58788 27226
rect 58812 27174 58842 27226
rect 58842 27174 58854 27226
rect 58854 27174 58868 27226
rect 58892 27174 58906 27226
rect 58906 27174 58918 27226
rect 58918 27174 58948 27226
rect 58972 27174 58982 27226
rect 58982 27174 59028 27226
rect 58732 27172 58788 27174
rect 58812 27172 58868 27174
rect 58892 27172 58948 27174
rect 58972 27172 59028 27174
rect 8178 26682 8234 26684
rect 8258 26682 8314 26684
rect 8338 26682 8394 26684
rect 8418 26682 8474 26684
rect 8178 26630 8224 26682
rect 8224 26630 8234 26682
rect 8258 26630 8288 26682
rect 8288 26630 8300 26682
rect 8300 26630 8314 26682
rect 8338 26630 8352 26682
rect 8352 26630 8364 26682
rect 8364 26630 8394 26682
rect 8418 26630 8428 26682
rect 8428 26630 8474 26682
rect 8178 26628 8234 26630
rect 8258 26628 8314 26630
rect 8338 26628 8394 26630
rect 8418 26628 8474 26630
rect 22622 26682 22678 26684
rect 22702 26682 22758 26684
rect 22782 26682 22838 26684
rect 22862 26682 22918 26684
rect 22622 26630 22668 26682
rect 22668 26630 22678 26682
rect 22702 26630 22732 26682
rect 22732 26630 22744 26682
rect 22744 26630 22758 26682
rect 22782 26630 22796 26682
rect 22796 26630 22808 26682
rect 22808 26630 22838 26682
rect 22862 26630 22872 26682
rect 22872 26630 22918 26682
rect 22622 26628 22678 26630
rect 22702 26628 22758 26630
rect 22782 26628 22838 26630
rect 22862 26628 22918 26630
rect 37066 26682 37122 26684
rect 37146 26682 37202 26684
rect 37226 26682 37282 26684
rect 37306 26682 37362 26684
rect 37066 26630 37112 26682
rect 37112 26630 37122 26682
rect 37146 26630 37176 26682
rect 37176 26630 37188 26682
rect 37188 26630 37202 26682
rect 37226 26630 37240 26682
rect 37240 26630 37252 26682
rect 37252 26630 37282 26682
rect 37306 26630 37316 26682
rect 37316 26630 37362 26682
rect 37066 26628 37122 26630
rect 37146 26628 37202 26630
rect 37226 26628 37282 26630
rect 37306 26628 37362 26630
rect 51510 26682 51566 26684
rect 51590 26682 51646 26684
rect 51670 26682 51726 26684
rect 51750 26682 51806 26684
rect 51510 26630 51556 26682
rect 51556 26630 51566 26682
rect 51590 26630 51620 26682
rect 51620 26630 51632 26682
rect 51632 26630 51646 26682
rect 51670 26630 51684 26682
rect 51684 26630 51696 26682
rect 51696 26630 51726 26682
rect 51750 26630 51760 26682
rect 51760 26630 51806 26682
rect 51510 26628 51566 26630
rect 51590 26628 51646 26630
rect 51670 26628 51726 26630
rect 51750 26628 51806 26630
rect 15400 26138 15456 26140
rect 15480 26138 15536 26140
rect 15560 26138 15616 26140
rect 15640 26138 15696 26140
rect 15400 26086 15446 26138
rect 15446 26086 15456 26138
rect 15480 26086 15510 26138
rect 15510 26086 15522 26138
rect 15522 26086 15536 26138
rect 15560 26086 15574 26138
rect 15574 26086 15586 26138
rect 15586 26086 15616 26138
rect 15640 26086 15650 26138
rect 15650 26086 15696 26138
rect 15400 26084 15456 26086
rect 15480 26084 15536 26086
rect 15560 26084 15616 26086
rect 15640 26084 15696 26086
rect 29844 26138 29900 26140
rect 29924 26138 29980 26140
rect 30004 26138 30060 26140
rect 30084 26138 30140 26140
rect 29844 26086 29890 26138
rect 29890 26086 29900 26138
rect 29924 26086 29954 26138
rect 29954 26086 29966 26138
rect 29966 26086 29980 26138
rect 30004 26086 30018 26138
rect 30018 26086 30030 26138
rect 30030 26086 30060 26138
rect 30084 26086 30094 26138
rect 30094 26086 30140 26138
rect 29844 26084 29900 26086
rect 29924 26084 29980 26086
rect 30004 26084 30060 26086
rect 30084 26084 30140 26086
rect 44288 26138 44344 26140
rect 44368 26138 44424 26140
rect 44448 26138 44504 26140
rect 44528 26138 44584 26140
rect 44288 26086 44334 26138
rect 44334 26086 44344 26138
rect 44368 26086 44398 26138
rect 44398 26086 44410 26138
rect 44410 26086 44424 26138
rect 44448 26086 44462 26138
rect 44462 26086 44474 26138
rect 44474 26086 44504 26138
rect 44528 26086 44538 26138
rect 44538 26086 44584 26138
rect 44288 26084 44344 26086
rect 44368 26084 44424 26086
rect 44448 26084 44504 26086
rect 44528 26084 44584 26086
rect 58732 26138 58788 26140
rect 58812 26138 58868 26140
rect 58892 26138 58948 26140
rect 58972 26138 59028 26140
rect 58732 26086 58778 26138
rect 58778 26086 58788 26138
rect 58812 26086 58842 26138
rect 58842 26086 58854 26138
rect 58854 26086 58868 26138
rect 58892 26086 58906 26138
rect 58906 26086 58918 26138
rect 58918 26086 58948 26138
rect 58972 26086 58982 26138
rect 58982 26086 59028 26138
rect 58732 26084 58788 26086
rect 58812 26084 58868 26086
rect 58892 26084 58948 26086
rect 58972 26084 59028 26086
rect 8178 25594 8234 25596
rect 8258 25594 8314 25596
rect 8338 25594 8394 25596
rect 8418 25594 8474 25596
rect 8178 25542 8224 25594
rect 8224 25542 8234 25594
rect 8258 25542 8288 25594
rect 8288 25542 8300 25594
rect 8300 25542 8314 25594
rect 8338 25542 8352 25594
rect 8352 25542 8364 25594
rect 8364 25542 8394 25594
rect 8418 25542 8428 25594
rect 8428 25542 8474 25594
rect 8178 25540 8234 25542
rect 8258 25540 8314 25542
rect 8338 25540 8394 25542
rect 8418 25540 8474 25542
rect 22622 25594 22678 25596
rect 22702 25594 22758 25596
rect 22782 25594 22838 25596
rect 22862 25594 22918 25596
rect 22622 25542 22668 25594
rect 22668 25542 22678 25594
rect 22702 25542 22732 25594
rect 22732 25542 22744 25594
rect 22744 25542 22758 25594
rect 22782 25542 22796 25594
rect 22796 25542 22808 25594
rect 22808 25542 22838 25594
rect 22862 25542 22872 25594
rect 22872 25542 22918 25594
rect 22622 25540 22678 25542
rect 22702 25540 22758 25542
rect 22782 25540 22838 25542
rect 22862 25540 22918 25542
rect 37066 25594 37122 25596
rect 37146 25594 37202 25596
rect 37226 25594 37282 25596
rect 37306 25594 37362 25596
rect 37066 25542 37112 25594
rect 37112 25542 37122 25594
rect 37146 25542 37176 25594
rect 37176 25542 37188 25594
rect 37188 25542 37202 25594
rect 37226 25542 37240 25594
rect 37240 25542 37252 25594
rect 37252 25542 37282 25594
rect 37306 25542 37316 25594
rect 37316 25542 37362 25594
rect 37066 25540 37122 25542
rect 37146 25540 37202 25542
rect 37226 25540 37282 25542
rect 37306 25540 37362 25542
rect 51510 25594 51566 25596
rect 51590 25594 51646 25596
rect 51670 25594 51726 25596
rect 51750 25594 51806 25596
rect 51510 25542 51556 25594
rect 51556 25542 51566 25594
rect 51590 25542 51620 25594
rect 51620 25542 51632 25594
rect 51632 25542 51646 25594
rect 51670 25542 51684 25594
rect 51684 25542 51696 25594
rect 51696 25542 51726 25594
rect 51750 25542 51760 25594
rect 51760 25542 51806 25594
rect 51510 25540 51566 25542
rect 51590 25540 51646 25542
rect 51670 25540 51726 25542
rect 51750 25540 51806 25542
rect 15400 25050 15456 25052
rect 15480 25050 15536 25052
rect 15560 25050 15616 25052
rect 15640 25050 15696 25052
rect 15400 24998 15446 25050
rect 15446 24998 15456 25050
rect 15480 24998 15510 25050
rect 15510 24998 15522 25050
rect 15522 24998 15536 25050
rect 15560 24998 15574 25050
rect 15574 24998 15586 25050
rect 15586 24998 15616 25050
rect 15640 24998 15650 25050
rect 15650 24998 15696 25050
rect 15400 24996 15456 24998
rect 15480 24996 15536 24998
rect 15560 24996 15616 24998
rect 15640 24996 15696 24998
rect 29844 25050 29900 25052
rect 29924 25050 29980 25052
rect 30004 25050 30060 25052
rect 30084 25050 30140 25052
rect 29844 24998 29890 25050
rect 29890 24998 29900 25050
rect 29924 24998 29954 25050
rect 29954 24998 29966 25050
rect 29966 24998 29980 25050
rect 30004 24998 30018 25050
rect 30018 24998 30030 25050
rect 30030 24998 30060 25050
rect 30084 24998 30094 25050
rect 30094 24998 30140 25050
rect 29844 24996 29900 24998
rect 29924 24996 29980 24998
rect 30004 24996 30060 24998
rect 30084 24996 30140 24998
rect 44288 25050 44344 25052
rect 44368 25050 44424 25052
rect 44448 25050 44504 25052
rect 44528 25050 44584 25052
rect 44288 24998 44334 25050
rect 44334 24998 44344 25050
rect 44368 24998 44398 25050
rect 44398 24998 44410 25050
rect 44410 24998 44424 25050
rect 44448 24998 44462 25050
rect 44462 24998 44474 25050
rect 44474 24998 44504 25050
rect 44528 24998 44538 25050
rect 44538 24998 44584 25050
rect 44288 24996 44344 24998
rect 44368 24996 44424 24998
rect 44448 24996 44504 24998
rect 44528 24996 44584 24998
rect 58732 25050 58788 25052
rect 58812 25050 58868 25052
rect 58892 25050 58948 25052
rect 58972 25050 59028 25052
rect 58732 24998 58778 25050
rect 58778 24998 58788 25050
rect 58812 24998 58842 25050
rect 58842 24998 58854 25050
rect 58854 24998 58868 25050
rect 58892 24998 58906 25050
rect 58906 24998 58918 25050
rect 58918 24998 58948 25050
rect 58972 24998 58982 25050
rect 58982 24998 59028 25050
rect 58732 24996 58788 24998
rect 58812 24996 58868 24998
rect 58892 24996 58948 24998
rect 58972 24996 59028 24998
rect 8178 24506 8234 24508
rect 8258 24506 8314 24508
rect 8338 24506 8394 24508
rect 8418 24506 8474 24508
rect 8178 24454 8224 24506
rect 8224 24454 8234 24506
rect 8258 24454 8288 24506
rect 8288 24454 8300 24506
rect 8300 24454 8314 24506
rect 8338 24454 8352 24506
rect 8352 24454 8364 24506
rect 8364 24454 8394 24506
rect 8418 24454 8428 24506
rect 8428 24454 8474 24506
rect 8178 24452 8234 24454
rect 8258 24452 8314 24454
rect 8338 24452 8394 24454
rect 8418 24452 8474 24454
rect 22622 24506 22678 24508
rect 22702 24506 22758 24508
rect 22782 24506 22838 24508
rect 22862 24506 22918 24508
rect 22622 24454 22668 24506
rect 22668 24454 22678 24506
rect 22702 24454 22732 24506
rect 22732 24454 22744 24506
rect 22744 24454 22758 24506
rect 22782 24454 22796 24506
rect 22796 24454 22808 24506
rect 22808 24454 22838 24506
rect 22862 24454 22872 24506
rect 22872 24454 22918 24506
rect 22622 24452 22678 24454
rect 22702 24452 22758 24454
rect 22782 24452 22838 24454
rect 22862 24452 22918 24454
rect 37066 24506 37122 24508
rect 37146 24506 37202 24508
rect 37226 24506 37282 24508
rect 37306 24506 37362 24508
rect 37066 24454 37112 24506
rect 37112 24454 37122 24506
rect 37146 24454 37176 24506
rect 37176 24454 37188 24506
rect 37188 24454 37202 24506
rect 37226 24454 37240 24506
rect 37240 24454 37252 24506
rect 37252 24454 37282 24506
rect 37306 24454 37316 24506
rect 37316 24454 37362 24506
rect 37066 24452 37122 24454
rect 37146 24452 37202 24454
rect 37226 24452 37282 24454
rect 37306 24452 37362 24454
rect 51510 24506 51566 24508
rect 51590 24506 51646 24508
rect 51670 24506 51726 24508
rect 51750 24506 51806 24508
rect 51510 24454 51556 24506
rect 51556 24454 51566 24506
rect 51590 24454 51620 24506
rect 51620 24454 51632 24506
rect 51632 24454 51646 24506
rect 51670 24454 51684 24506
rect 51684 24454 51696 24506
rect 51696 24454 51726 24506
rect 51750 24454 51760 24506
rect 51760 24454 51806 24506
rect 51510 24452 51566 24454
rect 51590 24452 51646 24454
rect 51670 24452 51726 24454
rect 51750 24452 51806 24454
rect 15400 23962 15456 23964
rect 15480 23962 15536 23964
rect 15560 23962 15616 23964
rect 15640 23962 15696 23964
rect 15400 23910 15446 23962
rect 15446 23910 15456 23962
rect 15480 23910 15510 23962
rect 15510 23910 15522 23962
rect 15522 23910 15536 23962
rect 15560 23910 15574 23962
rect 15574 23910 15586 23962
rect 15586 23910 15616 23962
rect 15640 23910 15650 23962
rect 15650 23910 15696 23962
rect 15400 23908 15456 23910
rect 15480 23908 15536 23910
rect 15560 23908 15616 23910
rect 15640 23908 15696 23910
rect 29844 23962 29900 23964
rect 29924 23962 29980 23964
rect 30004 23962 30060 23964
rect 30084 23962 30140 23964
rect 29844 23910 29890 23962
rect 29890 23910 29900 23962
rect 29924 23910 29954 23962
rect 29954 23910 29966 23962
rect 29966 23910 29980 23962
rect 30004 23910 30018 23962
rect 30018 23910 30030 23962
rect 30030 23910 30060 23962
rect 30084 23910 30094 23962
rect 30094 23910 30140 23962
rect 29844 23908 29900 23910
rect 29924 23908 29980 23910
rect 30004 23908 30060 23910
rect 30084 23908 30140 23910
rect 44288 23962 44344 23964
rect 44368 23962 44424 23964
rect 44448 23962 44504 23964
rect 44528 23962 44584 23964
rect 44288 23910 44334 23962
rect 44334 23910 44344 23962
rect 44368 23910 44398 23962
rect 44398 23910 44410 23962
rect 44410 23910 44424 23962
rect 44448 23910 44462 23962
rect 44462 23910 44474 23962
rect 44474 23910 44504 23962
rect 44528 23910 44538 23962
rect 44538 23910 44584 23962
rect 44288 23908 44344 23910
rect 44368 23908 44424 23910
rect 44448 23908 44504 23910
rect 44528 23908 44584 23910
rect 58732 23962 58788 23964
rect 58812 23962 58868 23964
rect 58892 23962 58948 23964
rect 58972 23962 59028 23964
rect 58732 23910 58778 23962
rect 58778 23910 58788 23962
rect 58812 23910 58842 23962
rect 58842 23910 58854 23962
rect 58854 23910 58868 23962
rect 58892 23910 58906 23962
rect 58906 23910 58918 23962
rect 58918 23910 58948 23962
rect 58972 23910 58982 23962
rect 58982 23910 59028 23962
rect 58732 23908 58788 23910
rect 58812 23908 58868 23910
rect 58892 23908 58948 23910
rect 58972 23908 59028 23910
rect 8178 23418 8234 23420
rect 8258 23418 8314 23420
rect 8338 23418 8394 23420
rect 8418 23418 8474 23420
rect 8178 23366 8224 23418
rect 8224 23366 8234 23418
rect 8258 23366 8288 23418
rect 8288 23366 8300 23418
rect 8300 23366 8314 23418
rect 8338 23366 8352 23418
rect 8352 23366 8364 23418
rect 8364 23366 8394 23418
rect 8418 23366 8428 23418
rect 8428 23366 8474 23418
rect 8178 23364 8234 23366
rect 8258 23364 8314 23366
rect 8338 23364 8394 23366
rect 8418 23364 8474 23366
rect 22622 23418 22678 23420
rect 22702 23418 22758 23420
rect 22782 23418 22838 23420
rect 22862 23418 22918 23420
rect 22622 23366 22668 23418
rect 22668 23366 22678 23418
rect 22702 23366 22732 23418
rect 22732 23366 22744 23418
rect 22744 23366 22758 23418
rect 22782 23366 22796 23418
rect 22796 23366 22808 23418
rect 22808 23366 22838 23418
rect 22862 23366 22872 23418
rect 22872 23366 22918 23418
rect 22622 23364 22678 23366
rect 22702 23364 22758 23366
rect 22782 23364 22838 23366
rect 22862 23364 22918 23366
rect 37066 23418 37122 23420
rect 37146 23418 37202 23420
rect 37226 23418 37282 23420
rect 37306 23418 37362 23420
rect 37066 23366 37112 23418
rect 37112 23366 37122 23418
rect 37146 23366 37176 23418
rect 37176 23366 37188 23418
rect 37188 23366 37202 23418
rect 37226 23366 37240 23418
rect 37240 23366 37252 23418
rect 37252 23366 37282 23418
rect 37306 23366 37316 23418
rect 37316 23366 37362 23418
rect 37066 23364 37122 23366
rect 37146 23364 37202 23366
rect 37226 23364 37282 23366
rect 37306 23364 37362 23366
rect 51510 23418 51566 23420
rect 51590 23418 51646 23420
rect 51670 23418 51726 23420
rect 51750 23418 51806 23420
rect 51510 23366 51556 23418
rect 51556 23366 51566 23418
rect 51590 23366 51620 23418
rect 51620 23366 51632 23418
rect 51632 23366 51646 23418
rect 51670 23366 51684 23418
rect 51684 23366 51696 23418
rect 51696 23366 51726 23418
rect 51750 23366 51760 23418
rect 51760 23366 51806 23418
rect 51510 23364 51566 23366
rect 51590 23364 51646 23366
rect 51670 23364 51726 23366
rect 51750 23364 51806 23366
rect 15400 22874 15456 22876
rect 15480 22874 15536 22876
rect 15560 22874 15616 22876
rect 15640 22874 15696 22876
rect 15400 22822 15446 22874
rect 15446 22822 15456 22874
rect 15480 22822 15510 22874
rect 15510 22822 15522 22874
rect 15522 22822 15536 22874
rect 15560 22822 15574 22874
rect 15574 22822 15586 22874
rect 15586 22822 15616 22874
rect 15640 22822 15650 22874
rect 15650 22822 15696 22874
rect 15400 22820 15456 22822
rect 15480 22820 15536 22822
rect 15560 22820 15616 22822
rect 15640 22820 15696 22822
rect 29844 22874 29900 22876
rect 29924 22874 29980 22876
rect 30004 22874 30060 22876
rect 30084 22874 30140 22876
rect 29844 22822 29890 22874
rect 29890 22822 29900 22874
rect 29924 22822 29954 22874
rect 29954 22822 29966 22874
rect 29966 22822 29980 22874
rect 30004 22822 30018 22874
rect 30018 22822 30030 22874
rect 30030 22822 30060 22874
rect 30084 22822 30094 22874
rect 30094 22822 30140 22874
rect 29844 22820 29900 22822
rect 29924 22820 29980 22822
rect 30004 22820 30060 22822
rect 30084 22820 30140 22822
rect 8178 22330 8234 22332
rect 8258 22330 8314 22332
rect 8338 22330 8394 22332
rect 8418 22330 8474 22332
rect 8178 22278 8224 22330
rect 8224 22278 8234 22330
rect 8258 22278 8288 22330
rect 8288 22278 8300 22330
rect 8300 22278 8314 22330
rect 8338 22278 8352 22330
rect 8352 22278 8364 22330
rect 8364 22278 8394 22330
rect 8418 22278 8428 22330
rect 8428 22278 8474 22330
rect 8178 22276 8234 22278
rect 8258 22276 8314 22278
rect 8338 22276 8394 22278
rect 8418 22276 8474 22278
rect 22622 22330 22678 22332
rect 22702 22330 22758 22332
rect 22782 22330 22838 22332
rect 22862 22330 22918 22332
rect 22622 22278 22668 22330
rect 22668 22278 22678 22330
rect 22702 22278 22732 22330
rect 22732 22278 22744 22330
rect 22744 22278 22758 22330
rect 22782 22278 22796 22330
rect 22796 22278 22808 22330
rect 22808 22278 22838 22330
rect 22862 22278 22872 22330
rect 22872 22278 22918 22330
rect 22622 22276 22678 22278
rect 22702 22276 22758 22278
rect 22782 22276 22838 22278
rect 22862 22276 22918 22278
rect 938 3440 994 3496
rect 8178 21242 8234 21244
rect 8258 21242 8314 21244
rect 8338 21242 8394 21244
rect 8418 21242 8474 21244
rect 8178 21190 8224 21242
rect 8224 21190 8234 21242
rect 8258 21190 8288 21242
rect 8288 21190 8300 21242
rect 8300 21190 8314 21242
rect 8338 21190 8352 21242
rect 8352 21190 8364 21242
rect 8364 21190 8394 21242
rect 8418 21190 8428 21242
rect 8428 21190 8474 21242
rect 8178 21188 8234 21190
rect 8258 21188 8314 21190
rect 8338 21188 8394 21190
rect 8418 21188 8474 21190
rect 6826 9988 6882 10024
rect 6826 9968 6828 9988
rect 6828 9968 6880 9988
rect 6880 9968 6882 9988
rect 8178 20154 8234 20156
rect 8258 20154 8314 20156
rect 8338 20154 8394 20156
rect 8418 20154 8474 20156
rect 8178 20102 8224 20154
rect 8224 20102 8234 20154
rect 8258 20102 8288 20154
rect 8288 20102 8300 20154
rect 8300 20102 8314 20154
rect 8338 20102 8352 20154
rect 8352 20102 8364 20154
rect 8364 20102 8394 20154
rect 8418 20102 8428 20154
rect 8428 20102 8474 20154
rect 8178 20100 8234 20102
rect 8258 20100 8314 20102
rect 8338 20100 8394 20102
rect 8418 20100 8474 20102
rect 11518 20340 11520 20360
rect 11520 20340 11572 20360
rect 11572 20340 11574 20360
rect 11518 20304 11574 20340
rect 8178 19066 8234 19068
rect 8258 19066 8314 19068
rect 8338 19066 8394 19068
rect 8418 19066 8474 19068
rect 8178 19014 8224 19066
rect 8224 19014 8234 19066
rect 8258 19014 8288 19066
rect 8288 19014 8300 19066
rect 8300 19014 8314 19066
rect 8338 19014 8352 19066
rect 8352 19014 8364 19066
rect 8364 19014 8394 19066
rect 8418 19014 8428 19066
rect 8428 19014 8474 19066
rect 8178 19012 8234 19014
rect 8258 19012 8314 19014
rect 8338 19012 8394 19014
rect 8418 19012 8474 19014
rect 8178 17978 8234 17980
rect 8258 17978 8314 17980
rect 8338 17978 8394 17980
rect 8418 17978 8474 17980
rect 8178 17926 8224 17978
rect 8224 17926 8234 17978
rect 8258 17926 8288 17978
rect 8288 17926 8300 17978
rect 8300 17926 8314 17978
rect 8338 17926 8352 17978
rect 8352 17926 8364 17978
rect 8364 17926 8394 17978
rect 8418 17926 8428 17978
rect 8428 17926 8474 17978
rect 8178 17924 8234 17926
rect 8258 17924 8314 17926
rect 8338 17924 8394 17926
rect 8418 17924 8474 17926
rect 8178 16890 8234 16892
rect 8258 16890 8314 16892
rect 8338 16890 8394 16892
rect 8418 16890 8474 16892
rect 8178 16838 8224 16890
rect 8224 16838 8234 16890
rect 8258 16838 8288 16890
rect 8288 16838 8300 16890
rect 8300 16838 8314 16890
rect 8338 16838 8352 16890
rect 8352 16838 8364 16890
rect 8364 16838 8394 16890
rect 8418 16838 8428 16890
rect 8428 16838 8474 16890
rect 8178 16836 8234 16838
rect 8258 16836 8314 16838
rect 8338 16836 8394 16838
rect 8418 16836 8474 16838
rect 8178 15802 8234 15804
rect 8258 15802 8314 15804
rect 8338 15802 8394 15804
rect 8418 15802 8474 15804
rect 8178 15750 8224 15802
rect 8224 15750 8234 15802
rect 8258 15750 8288 15802
rect 8288 15750 8300 15802
rect 8300 15750 8314 15802
rect 8338 15750 8352 15802
rect 8352 15750 8364 15802
rect 8364 15750 8394 15802
rect 8418 15750 8428 15802
rect 8428 15750 8474 15802
rect 8178 15748 8234 15750
rect 8258 15748 8314 15750
rect 8338 15748 8394 15750
rect 8418 15748 8474 15750
rect 8178 14714 8234 14716
rect 8258 14714 8314 14716
rect 8338 14714 8394 14716
rect 8418 14714 8474 14716
rect 8178 14662 8224 14714
rect 8224 14662 8234 14714
rect 8258 14662 8288 14714
rect 8288 14662 8300 14714
rect 8300 14662 8314 14714
rect 8338 14662 8352 14714
rect 8352 14662 8364 14714
rect 8364 14662 8394 14714
rect 8418 14662 8428 14714
rect 8428 14662 8474 14714
rect 8178 14660 8234 14662
rect 8258 14660 8314 14662
rect 8338 14660 8394 14662
rect 8418 14660 8474 14662
rect 5446 4140 5502 4176
rect 5446 4120 5448 4140
rect 5448 4120 5500 4140
rect 5500 4120 5502 4140
rect 5998 3576 6054 3632
rect 8178 13626 8234 13628
rect 8258 13626 8314 13628
rect 8338 13626 8394 13628
rect 8418 13626 8474 13628
rect 8178 13574 8224 13626
rect 8224 13574 8234 13626
rect 8258 13574 8288 13626
rect 8288 13574 8300 13626
rect 8300 13574 8314 13626
rect 8338 13574 8352 13626
rect 8352 13574 8364 13626
rect 8364 13574 8394 13626
rect 8418 13574 8428 13626
rect 8428 13574 8474 13626
rect 8178 13572 8234 13574
rect 8258 13572 8314 13574
rect 8338 13572 8394 13574
rect 8418 13572 8474 13574
rect 8178 12538 8234 12540
rect 8258 12538 8314 12540
rect 8338 12538 8394 12540
rect 8418 12538 8474 12540
rect 8178 12486 8224 12538
rect 8224 12486 8234 12538
rect 8258 12486 8288 12538
rect 8288 12486 8300 12538
rect 8300 12486 8314 12538
rect 8338 12486 8352 12538
rect 8352 12486 8364 12538
rect 8364 12486 8394 12538
rect 8418 12486 8428 12538
rect 8428 12486 8474 12538
rect 8178 12484 8234 12486
rect 8258 12484 8314 12486
rect 8338 12484 8394 12486
rect 8418 12484 8474 12486
rect 8390 11620 8446 11656
rect 8390 11600 8392 11620
rect 8392 11600 8444 11620
rect 8444 11600 8446 11620
rect 8178 11450 8234 11452
rect 8258 11450 8314 11452
rect 8338 11450 8394 11452
rect 8418 11450 8474 11452
rect 8178 11398 8224 11450
rect 8224 11398 8234 11450
rect 8258 11398 8288 11450
rect 8288 11398 8300 11450
rect 8300 11398 8314 11450
rect 8338 11398 8352 11450
rect 8352 11398 8364 11450
rect 8364 11398 8394 11450
rect 8418 11398 8428 11450
rect 8428 11398 8474 11450
rect 8178 11396 8234 11398
rect 8258 11396 8314 11398
rect 8338 11396 8394 11398
rect 8418 11396 8474 11398
rect 8178 10362 8234 10364
rect 8258 10362 8314 10364
rect 8338 10362 8394 10364
rect 8418 10362 8474 10364
rect 8178 10310 8224 10362
rect 8224 10310 8234 10362
rect 8258 10310 8288 10362
rect 8288 10310 8300 10362
rect 8300 10310 8314 10362
rect 8338 10310 8352 10362
rect 8352 10310 8364 10362
rect 8364 10310 8394 10362
rect 8418 10310 8428 10362
rect 8428 10310 8474 10362
rect 8178 10308 8234 10310
rect 8258 10308 8314 10310
rect 8338 10308 8394 10310
rect 8418 10308 8474 10310
rect 8178 9274 8234 9276
rect 8258 9274 8314 9276
rect 8338 9274 8394 9276
rect 8418 9274 8474 9276
rect 8178 9222 8224 9274
rect 8224 9222 8234 9274
rect 8258 9222 8288 9274
rect 8288 9222 8300 9274
rect 8300 9222 8314 9274
rect 8338 9222 8352 9274
rect 8352 9222 8364 9274
rect 8364 9222 8394 9274
rect 8418 9222 8428 9274
rect 8428 9222 8474 9274
rect 8178 9220 8234 9222
rect 8258 9220 8314 9222
rect 8338 9220 8394 9222
rect 8418 9220 8474 9222
rect 8178 8186 8234 8188
rect 8258 8186 8314 8188
rect 8338 8186 8394 8188
rect 8418 8186 8474 8188
rect 8178 8134 8224 8186
rect 8224 8134 8234 8186
rect 8258 8134 8288 8186
rect 8288 8134 8300 8186
rect 8300 8134 8314 8186
rect 8338 8134 8352 8186
rect 8352 8134 8364 8186
rect 8364 8134 8394 8186
rect 8418 8134 8428 8186
rect 8428 8134 8474 8186
rect 8178 8132 8234 8134
rect 8258 8132 8314 8134
rect 8338 8132 8394 8134
rect 8418 8132 8474 8134
rect 8178 7098 8234 7100
rect 8258 7098 8314 7100
rect 8338 7098 8394 7100
rect 8418 7098 8474 7100
rect 8178 7046 8224 7098
rect 8224 7046 8234 7098
rect 8258 7046 8288 7098
rect 8288 7046 8300 7098
rect 8300 7046 8314 7098
rect 8338 7046 8352 7098
rect 8352 7046 8364 7098
rect 8364 7046 8394 7098
rect 8418 7046 8428 7098
rect 8428 7046 8474 7098
rect 8178 7044 8234 7046
rect 8258 7044 8314 7046
rect 8338 7044 8394 7046
rect 8418 7044 8474 7046
rect 8178 6010 8234 6012
rect 8258 6010 8314 6012
rect 8338 6010 8394 6012
rect 8418 6010 8474 6012
rect 8178 5958 8224 6010
rect 8224 5958 8234 6010
rect 8258 5958 8288 6010
rect 8288 5958 8300 6010
rect 8300 5958 8314 6010
rect 8338 5958 8352 6010
rect 8352 5958 8364 6010
rect 8364 5958 8394 6010
rect 8418 5958 8428 6010
rect 8428 5958 8474 6010
rect 8178 5956 8234 5958
rect 8258 5956 8314 5958
rect 8338 5956 8394 5958
rect 8418 5956 8474 5958
rect 8666 6316 8722 6352
rect 8666 6296 8668 6316
rect 8668 6296 8720 6316
rect 8720 6296 8722 6316
rect 8942 5752 8998 5808
rect 8178 4922 8234 4924
rect 8258 4922 8314 4924
rect 8338 4922 8394 4924
rect 8418 4922 8474 4924
rect 8178 4870 8224 4922
rect 8224 4870 8234 4922
rect 8258 4870 8288 4922
rect 8288 4870 8300 4922
rect 8300 4870 8314 4922
rect 8338 4870 8352 4922
rect 8352 4870 8364 4922
rect 8364 4870 8394 4922
rect 8418 4870 8428 4922
rect 8428 4870 8474 4922
rect 8178 4868 8234 4870
rect 8258 4868 8314 4870
rect 8338 4868 8394 4870
rect 8418 4868 8474 4870
rect 8178 3834 8234 3836
rect 8258 3834 8314 3836
rect 8338 3834 8394 3836
rect 8418 3834 8474 3836
rect 8178 3782 8224 3834
rect 8224 3782 8234 3834
rect 8258 3782 8288 3834
rect 8288 3782 8300 3834
rect 8300 3782 8314 3834
rect 8338 3782 8352 3834
rect 8352 3782 8364 3834
rect 8364 3782 8394 3834
rect 8418 3782 8428 3834
rect 8428 3782 8474 3834
rect 8178 3780 8234 3782
rect 8258 3780 8314 3782
rect 8338 3780 8394 3782
rect 8418 3780 8474 3782
rect 9126 4664 9182 4720
rect 8178 2746 8234 2748
rect 8258 2746 8314 2748
rect 8338 2746 8394 2748
rect 8418 2746 8474 2748
rect 8178 2694 8224 2746
rect 8224 2694 8234 2746
rect 8258 2694 8288 2746
rect 8288 2694 8300 2746
rect 8300 2694 8314 2746
rect 8338 2694 8352 2746
rect 8352 2694 8364 2746
rect 8364 2694 8394 2746
rect 8418 2694 8428 2746
rect 8428 2694 8474 2746
rect 8178 2692 8234 2694
rect 8258 2692 8314 2694
rect 8338 2692 8394 2694
rect 8418 2692 8474 2694
rect 9586 11600 9642 11656
rect 9494 10648 9550 10704
rect 9770 9596 9772 9616
rect 9772 9596 9824 9616
rect 9824 9596 9826 9616
rect 9770 9560 9826 9596
rect 12898 17756 12900 17776
rect 12900 17756 12952 17776
rect 12952 17756 12954 17776
rect 12898 17720 12954 17756
rect 15400 21786 15456 21788
rect 15480 21786 15536 21788
rect 15560 21786 15616 21788
rect 15640 21786 15696 21788
rect 15400 21734 15446 21786
rect 15446 21734 15456 21786
rect 15480 21734 15510 21786
rect 15510 21734 15522 21786
rect 15522 21734 15536 21786
rect 15560 21734 15574 21786
rect 15574 21734 15586 21786
rect 15586 21734 15616 21786
rect 15640 21734 15650 21786
rect 15650 21734 15696 21786
rect 15400 21732 15456 21734
rect 15480 21732 15536 21734
rect 15560 21732 15616 21734
rect 15640 21732 15696 21734
rect 9494 3052 9550 3088
rect 9494 3032 9496 3052
rect 9496 3032 9548 3052
rect 9548 3032 9550 3052
rect 11150 5092 11206 5128
rect 11150 5072 11152 5092
rect 11152 5072 11204 5092
rect 11204 5072 11206 5092
rect 15400 20698 15456 20700
rect 15480 20698 15536 20700
rect 15560 20698 15616 20700
rect 15640 20698 15696 20700
rect 15400 20646 15446 20698
rect 15446 20646 15456 20698
rect 15480 20646 15510 20698
rect 15510 20646 15522 20698
rect 15522 20646 15536 20698
rect 15560 20646 15574 20698
rect 15574 20646 15586 20698
rect 15586 20646 15616 20698
rect 15640 20646 15650 20698
rect 15650 20646 15696 20698
rect 15400 20644 15456 20646
rect 15480 20644 15536 20646
rect 15560 20644 15616 20646
rect 15640 20644 15696 20646
rect 18142 20324 18198 20360
rect 18142 20304 18144 20324
rect 18144 20304 18196 20324
rect 18196 20304 18198 20324
rect 15400 19610 15456 19612
rect 15480 19610 15536 19612
rect 15560 19610 15616 19612
rect 15640 19610 15696 19612
rect 15400 19558 15446 19610
rect 15446 19558 15456 19610
rect 15480 19558 15510 19610
rect 15510 19558 15522 19610
rect 15522 19558 15536 19610
rect 15560 19558 15574 19610
rect 15574 19558 15586 19610
rect 15586 19558 15616 19610
rect 15640 19558 15650 19610
rect 15650 19558 15696 19610
rect 15400 19556 15456 19558
rect 15480 19556 15536 19558
rect 15560 19556 15616 19558
rect 15640 19556 15696 19558
rect 15400 18522 15456 18524
rect 15480 18522 15536 18524
rect 15560 18522 15616 18524
rect 15640 18522 15696 18524
rect 15400 18470 15446 18522
rect 15446 18470 15456 18522
rect 15480 18470 15510 18522
rect 15510 18470 15522 18522
rect 15522 18470 15536 18522
rect 15560 18470 15574 18522
rect 15574 18470 15586 18522
rect 15586 18470 15616 18522
rect 15640 18470 15650 18522
rect 15650 18470 15696 18522
rect 15400 18468 15456 18470
rect 15480 18468 15536 18470
rect 15560 18468 15616 18470
rect 15640 18468 15696 18470
rect 15934 17720 15990 17776
rect 15400 17434 15456 17436
rect 15480 17434 15536 17436
rect 15560 17434 15616 17436
rect 15640 17434 15696 17436
rect 15400 17382 15446 17434
rect 15446 17382 15456 17434
rect 15480 17382 15510 17434
rect 15510 17382 15522 17434
rect 15522 17382 15536 17434
rect 15560 17382 15574 17434
rect 15574 17382 15586 17434
rect 15586 17382 15616 17434
rect 15640 17382 15650 17434
rect 15650 17382 15696 17434
rect 15400 17380 15456 17382
rect 15480 17380 15536 17382
rect 15560 17380 15616 17382
rect 15640 17380 15696 17382
rect 11610 3032 11666 3088
rect 13726 5228 13782 5264
rect 13726 5208 13728 5228
rect 13728 5208 13780 5228
rect 13780 5208 13782 5228
rect 12346 3032 12402 3088
rect 15400 16346 15456 16348
rect 15480 16346 15536 16348
rect 15560 16346 15616 16348
rect 15640 16346 15696 16348
rect 15400 16294 15446 16346
rect 15446 16294 15456 16346
rect 15480 16294 15510 16346
rect 15510 16294 15522 16346
rect 15522 16294 15536 16346
rect 15560 16294 15574 16346
rect 15574 16294 15586 16346
rect 15586 16294 15616 16346
rect 15640 16294 15650 16346
rect 15650 16294 15696 16346
rect 15400 16292 15456 16294
rect 15480 16292 15536 16294
rect 15560 16292 15616 16294
rect 15640 16292 15696 16294
rect 15400 15258 15456 15260
rect 15480 15258 15536 15260
rect 15560 15258 15616 15260
rect 15640 15258 15696 15260
rect 15400 15206 15446 15258
rect 15446 15206 15456 15258
rect 15480 15206 15510 15258
rect 15510 15206 15522 15258
rect 15522 15206 15536 15258
rect 15560 15206 15574 15258
rect 15574 15206 15586 15258
rect 15586 15206 15616 15258
rect 15640 15206 15650 15258
rect 15650 15206 15696 15258
rect 15400 15204 15456 15206
rect 15480 15204 15536 15206
rect 15560 15204 15616 15206
rect 15640 15204 15696 15206
rect 15400 14170 15456 14172
rect 15480 14170 15536 14172
rect 15560 14170 15616 14172
rect 15640 14170 15696 14172
rect 15400 14118 15446 14170
rect 15446 14118 15456 14170
rect 15480 14118 15510 14170
rect 15510 14118 15522 14170
rect 15522 14118 15536 14170
rect 15560 14118 15574 14170
rect 15574 14118 15586 14170
rect 15586 14118 15616 14170
rect 15640 14118 15650 14170
rect 15650 14118 15696 14170
rect 15400 14116 15456 14118
rect 15480 14116 15536 14118
rect 15560 14116 15616 14118
rect 15640 14116 15696 14118
rect 15400 13082 15456 13084
rect 15480 13082 15536 13084
rect 15560 13082 15616 13084
rect 15640 13082 15696 13084
rect 15400 13030 15446 13082
rect 15446 13030 15456 13082
rect 15480 13030 15510 13082
rect 15510 13030 15522 13082
rect 15522 13030 15536 13082
rect 15560 13030 15574 13082
rect 15574 13030 15586 13082
rect 15586 13030 15616 13082
rect 15640 13030 15650 13082
rect 15650 13030 15696 13082
rect 15400 13028 15456 13030
rect 15480 13028 15536 13030
rect 15560 13028 15616 13030
rect 15640 13028 15696 13030
rect 15400 11994 15456 11996
rect 15480 11994 15536 11996
rect 15560 11994 15616 11996
rect 15640 11994 15696 11996
rect 15400 11942 15446 11994
rect 15446 11942 15456 11994
rect 15480 11942 15510 11994
rect 15510 11942 15522 11994
rect 15522 11942 15536 11994
rect 15560 11942 15574 11994
rect 15574 11942 15586 11994
rect 15586 11942 15616 11994
rect 15640 11942 15650 11994
rect 15650 11942 15696 11994
rect 15400 11940 15456 11942
rect 15480 11940 15536 11942
rect 15560 11940 15616 11942
rect 15640 11940 15696 11942
rect 15400 10906 15456 10908
rect 15480 10906 15536 10908
rect 15560 10906 15616 10908
rect 15640 10906 15696 10908
rect 15400 10854 15446 10906
rect 15446 10854 15456 10906
rect 15480 10854 15510 10906
rect 15510 10854 15522 10906
rect 15522 10854 15536 10906
rect 15560 10854 15574 10906
rect 15574 10854 15586 10906
rect 15586 10854 15616 10906
rect 15640 10854 15650 10906
rect 15650 10854 15696 10906
rect 15400 10852 15456 10854
rect 15480 10852 15536 10854
rect 15560 10852 15616 10854
rect 15640 10852 15696 10854
rect 15400 9818 15456 9820
rect 15480 9818 15536 9820
rect 15560 9818 15616 9820
rect 15640 9818 15696 9820
rect 15400 9766 15446 9818
rect 15446 9766 15456 9818
rect 15480 9766 15510 9818
rect 15510 9766 15522 9818
rect 15522 9766 15536 9818
rect 15560 9766 15574 9818
rect 15574 9766 15586 9818
rect 15586 9766 15616 9818
rect 15640 9766 15650 9818
rect 15650 9766 15696 9818
rect 15400 9764 15456 9766
rect 15480 9764 15536 9766
rect 15560 9764 15616 9766
rect 15640 9764 15696 9766
rect 15400 8730 15456 8732
rect 15480 8730 15536 8732
rect 15560 8730 15616 8732
rect 15640 8730 15696 8732
rect 15400 8678 15446 8730
rect 15446 8678 15456 8730
rect 15480 8678 15510 8730
rect 15510 8678 15522 8730
rect 15522 8678 15536 8730
rect 15560 8678 15574 8730
rect 15574 8678 15586 8730
rect 15586 8678 15616 8730
rect 15640 8678 15650 8730
rect 15650 8678 15696 8730
rect 15400 8676 15456 8678
rect 15480 8676 15536 8678
rect 15560 8676 15616 8678
rect 15640 8676 15696 8678
rect 15400 7642 15456 7644
rect 15480 7642 15536 7644
rect 15560 7642 15616 7644
rect 15640 7642 15696 7644
rect 15400 7590 15446 7642
rect 15446 7590 15456 7642
rect 15480 7590 15510 7642
rect 15510 7590 15522 7642
rect 15522 7590 15536 7642
rect 15560 7590 15574 7642
rect 15574 7590 15586 7642
rect 15586 7590 15616 7642
rect 15640 7590 15650 7642
rect 15650 7590 15696 7642
rect 15400 7588 15456 7590
rect 15480 7588 15536 7590
rect 15560 7588 15616 7590
rect 15640 7588 15696 7590
rect 15400 6554 15456 6556
rect 15480 6554 15536 6556
rect 15560 6554 15616 6556
rect 15640 6554 15696 6556
rect 15400 6502 15446 6554
rect 15446 6502 15456 6554
rect 15480 6502 15510 6554
rect 15510 6502 15522 6554
rect 15522 6502 15536 6554
rect 15560 6502 15574 6554
rect 15574 6502 15586 6554
rect 15586 6502 15616 6554
rect 15640 6502 15650 6554
rect 15650 6502 15696 6554
rect 15400 6500 15456 6502
rect 15480 6500 15536 6502
rect 15560 6500 15616 6502
rect 15640 6500 15696 6502
rect 15400 5466 15456 5468
rect 15480 5466 15536 5468
rect 15560 5466 15616 5468
rect 15640 5466 15696 5468
rect 15400 5414 15446 5466
rect 15446 5414 15456 5466
rect 15480 5414 15510 5466
rect 15510 5414 15522 5466
rect 15522 5414 15536 5466
rect 15560 5414 15574 5466
rect 15574 5414 15586 5466
rect 15586 5414 15616 5466
rect 15640 5414 15650 5466
rect 15650 5414 15696 5466
rect 15400 5412 15456 5414
rect 15480 5412 15536 5414
rect 15560 5412 15616 5414
rect 15640 5412 15696 5414
rect 16026 9596 16028 9616
rect 16028 9596 16080 9616
rect 16080 9596 16082 9616
rect 16026 9560 16082 9596
rect 17682 10512 17738 10568
rect 17038 10260 17094 10296
rect 17038 10240 17040 10260
rect 17040 10240 17092 10260
rect 17092 10240 17094 10260
rect 15400 4378 15456 4380
rect 15480 4378 15536 4380
rect 15560 4378 15616 4380
rect 15640 4378 15696 4380
rect 15400 4326 15446 4378
rect 15446 4326 15456 4378
rect 15480 4326 15510 4378
rect 15510 4326 15522 4378
rect 15522 4326 15536 4378
rect 15560 4326 15574 4378
rect 15574 4326 15586 4378
rect 15586 4326 15616 4378
rect 15640 4326 15650 4378
rect 15650 4326 15696 4378
rect 15400 4324 15456 4326
rect 15480 4324 15536 4326
rect 15560 4324 15616 4326
rect 15640 4324 15696 4326
rect 15106 2896 15162 2952
rect 15400 3290 15456 3292
rect 15480 3290 15536 3292
rect 15560 3290 15616 3292
rect 15640 3290 15696 3292
rect 15400 3238 15446 3290
rect 15446 3238 15456 3290
rect 15480 3238 15510 3290
rect 15510 3238 15522 3290
rect 15522 3238 15536 3290
rect 15560 3238 15574 3290
rect 15574 3238 15586 3290
rect 15586 3238 15616 3290
rect 15640 3238 15650 3290
rect 15650 3238 15696 3290
rect 15400 3236 15456 3238
rect 15480 3236 15536 3238
rect 15560 3236 15616 3238
rect 15640 3236 15696 3238
rect 16302 3032 16358 3088
rect 15400 2202 15456 2204
rect 15480 2202 15536 2204
rect 15560 2202 15616 2204
rect 15640 2202 15696 2204
rect 15400 2150 15446 2202
rect 15446 2150 15456 2202
rect 15480 2150 15510 2202
rect 15510 2150 15522 2202
rect 15522 2150 15536 2202
rect 15560 2150 15574 2202
rect 15574 2150 15586 2202
rect 15586 2150 15616 2202
rect 15640 2150 15650 2202
rect 15650 2150 15696 2202
rect 15400 2148 15456 2150
rect 15480 2148 15536 2150
rect 15560 2148 15616 2150
rect 15640 2148 15696 2150
rect 18418 10648 18474 10704
rect 18602 10240 18658 10296
rect 22622 21242 22678 21244
rect 22702 21242 22758 21244
rect 22782 21242 22838 21244
rect 22862 21242 22918 21244
rect 22622 21190 22668 21242
rect 22668 21190 22678 21242
rect 22702 21190 22732 21242
rect 22732 21190 22744 21242
rect 22744 21190 22758 21242
rect 22782 21190 22796 21242
rect 22796 21190 22808 21242
rect 22808 21190 22838 21242
rect 22862 21190 22872 21242
rect 22872 21190 22918 21242
rect 22622 21188 22678 21190
rect 22702 21188 22758 21190
rect 22782 21188 22838 21190
rect 22862 21188 22918 21190
rect 20534 17740 20590 17776
rect 20534 17720 20536 17740
rect 20536 17720 20588 17740
rect 20588 17720 20590 17740
rect 19062 10548 19064 10568
rect 19064 10548 19116 10568
rect 19116 10548 19118 10568
rect 19062 10512 19118 10548
rect 18970 2916 19026 2952
rect 18970 2896 18972 2916
rect 18972 2896 19024 2916
rect 19024 2896 19026 2916
rect 22622 20154 22678 20156
rect 22702 20154 22758 20156
rect 22782 20154 22838 20156
rect 22862 20154 22918 20156
rect 22622 20102 22668 20154
rect 22668 20102 22678 20154
rect 22702 20102 22732 20154
rect 22732 20102 22744 20154
rect 22744 20102 22758 20154
rect 22782 20102 22796 20154
rect 22796 20102 22808 20154
rect 22808 20102 22838 20154
rect 22862 20102 22872 20154
rect 22872 20102 22918 20154
rect 22622 20100 22678 20102
rect 22702 20100 22758 20102
rect 22782 20100 22838 20102
rect 22862 20100 22918 20102
rect 37066 22330 37122 22332
rect 37146 22330 37202 22332
rect 37226 22330 37282 22332
rect 37306 22330 37362 22332
rect 37066 22278 37112 22330
rect 37112 22278 37122 22330
rect 37146 22278 37176 22330
rect 37176 22278 37188 22330
rect 37188 22278 37202 22330
rect 37226 22278 37240 22330
rect 37240 22278 37252 22330
rect 37252 22278 37282 22330
rect 37306 22278 37316 22330
rect 37316 22278 37362 22330
rect 37066 22276 37122 22278
rect 37146 22276 37202 22278
rect 37226 22276 37282 22278
rect 37306 22276 37362 22278
rect 29844 21786 29900 21788
rect 29924 21786 29980 21788
rect 30004 21786 30060 21788
rect 30084 21786 30140 21788
rect 29844 21734 29890 21786
rect 29890 21734 29900 21786
rect 29924 21734 29954 21786
rect 29954 21734 29966 21786
rect 29966 21734 29980 21786
rect 30004 21734 30018 21786
rect 30018 21734 30030 21786
rect 30030 21734 30060 21786
rect 30084 21734 30094 21786
rect 30094 21734 30140 21786
rect 29844 21732 29900 21734
rect 29924 21732 29980 21734
rect 30004 21732 30060 21734
rect 30084 21732 30140 21734
rect 24306 20868 24362 20904
rect 24306 20848 24308 20868
rect 24308 20848 24360 20868
rect 24360 20848 24362 20868
rect 22622 19066 22678 19068
rect 22702 19066 22758 19068
rect 22782 19066 22838 19068
rect 22862 19066 22918 19068
rect 22622 19014 22668 19066
rect 22668 19014 22678 19066
rect 22702 19014 22732 19066
rect 22732 19014 22744 19066
rect 22744 19014 22758 19066
rect 22782 19014 22796 19066
rect 22796 19014 22808 19066
rect 22808 19014 22838 19066
rect 22862 19014 22872 19066
rect 22872 19014 22918 19066
rect 22622 19012 22678 19014
rect 22702 19012 22758 19014
rect 22782 19012 22838 19014
rect 22862 19012 22918 19014
rect 22622 17978 22678 17980
rect 22702 17978 22758 17980
rect 22782 17978 22838 17980
rect 22862 17978 22918 17980
rect 22622 17926 22668 17978
rect 22668 17926 22678 17978
rect 22702 17926 22732 17978
rect 22732 17926 22744 17978
rect 22744 17926 22758 17978
rect 22782 17926 22796 17978
rect 22796 17926 22808 17978
rect 22808 17926 22838 17978
rect 22862 17926 22872 17978
rect 22872 17926 22918 17978
rect 22622 17924 22678 17926
rect 22702 17924 22758 17926
rect 22782 17924 22838 17926
rect 22862 17924 22918 17926
rect 22622 16890 22678 16892
rect 22702 16890 22758 16892
rect 22782 16890 22838 16892
rect 22862 16890 22918 16892
rect 22622 16838 22668 16890
rect 22668 16838 22678 16890
rect 22702 16838 22732 16890
rect 22732 16838 22744 16890
rect 22744 16838 22758 16890
rect 22782 16838 22796 16890
rect 22796 16838 22808 16890
rect 22808 16838 22838 16890
rect 22862 16838 22872 16890
rect 22872 16838 22918 16890
rect 22622 16836 22678 16838
rect 22702 16836 22758 16838
rect 22782 16836 22838 16838
rect 22862 16836 22918 16838
rect 22622 15802 22678 15804
rect 22702 15802 22758 15804
rect 22782 15802 22838 15804
rect 22862 15802 22918 15804
rect 22622 15750 22668 15802
rect 22668 15750 22678 15802
rect 22702 15750 22732 15802
rect 22732 15750 22744 15802
rect 22744 15750 22758 15802
rect 22782 15750 22796 15802
rect 22796 15750 22808 15802
rect 22808 15750 22838 15802
rect 22862 15750 22872 15802
rect 22872 15750 22918 15802
rect 22622 15748 22678 15750
rect 22702 15748 22758 15750
rect 22782 15748 22838 15750
rect 22862 15748 22918 15750
rect 22622 14714 22678 14716
rect 22702 14714 22758 14716
rect 22782 14714 22838 14716
rect 22862 14714 22918 14716
rect 22622 14662 22668 14714
rect 22668 14662 22678 14714
rect 22702 14662 22732 14714
rect 22732 14662 22744 14714
rect 22744 14662 22758 14714
rect 22782 14662 22796 14714
rect 22796 14662 22808 14714
rect 22808 14662 22838 14714
rect 22862 14662 22872 14714
rect 22872 14662 22918 14714
rect 22622 14660 22678 14662
rect 22702 14660 22758 14662
rect 22782 14660 22838 14662
rect 22862 14660 22918 14662
rect 22622 13626 22678 13628
rect 22702 13626 22758 13628
rect 22782 13626 22838 13628
rect 22862 13626 22918 13628
rect 22622 13574 22668 13626
rect 22668 13574 22678 13626
rect 22702 13574 22732 13626
rect 22732 13574 22744 13626
rect 22744 13574 22758 13626
rect 22782 13574 22796 13626
rect 22796 13574 22808 13626
rect 22808 13574 22838 13626
rect 22862 13574 22872 13626
rect 22872 13574 22918 13626
rect 22622 13572 22678 13574
rect 22702 13572 22758 13574
rect 22782 13572 22838 13574
rect 22862 13572 22918 13574
rect 22622 12538 22678 12540
rect 22702 12538 22758 12540
rect 22782 12538 22838 12540
rect 22862 12538 22918 12540
rect 22622 12486 22668 12538
rect 22668 12486 22678 12538
rect 22702 12486 22732 12538
rect 22732 12486 22744 12538
rect 22744 12486 22758 12538
rect 22782 12486 22796 12538
rect 22796 12486 22808 12538
rect 22808 12486 22838 12538
rect 22862 12486 22872 12538
rect 22872 12486 22918 12538
rect 22622 12484 22678 12486
rect 22702 12484 22758 12486
rect 22782 12484 22838 12486
rect 22862 12484 22918 12486
rect 22622 11450 22678 11452
rect 22702 11450 22758 11452
rect 22782 11450 22838 11452
rect 22862 11450 22918 11452
rect 22622 11398 22668 11450
rect 22668 11398 22678 11450
rect 22702 11398 22732 11450
rect 22732 11398 22744 11450
rect 22744 11398 22758 11450
rect 22782 11398 22796 11450
rect 22796 11398 22808 11450
rect 22808 11398 22838 11450
rect 22862 11398 22872 11450
rect 22872 11398 22918 11450
rect 22622 11396 22678 11398
rect 22702 11396 22758 11398
rect 22782 11396 22838 11398
rect 22862 11396 22918 11398
rect 20258 5616 20314 5672
rect 22622 10362 22678 10364
rect 22702 10362 22758 10364
rect 22782 10362 22838 10364
rect 22862 10362 22918 10364
rect 22622 10310 22668 10362
rect 22668 10310 22678 10362
rect 22702 10310 22732 10362
rect 22732 10310 22744 10362
rect 22744 10310 22758 10362
rect 22782 10310 22796 10362
rect 22796 10310 22808 10362
rect 22808 10310 22838 10362
rect 22862 10310 22872 10362
rect 22872 10310 22918 10362
rect 22622 10308 22678 10310
rect 22702 10308 22758 10310
rect 22782 10308 22838 10310
rect 22862 10308 22918 10310
rect 24858 20324 24914 20360
rect 25502 20848 25558 20904
rect 24858 20304 24860 20324
rect 24860 20304 24912 20324
rect 24912 20304 24914 20324
rect 29844 20698 29900 20700
rect 29924 20698 29980 20700
rect 30004 20698 30060 20700
rect 30084 20698 30140 20700
rect 29844 20646 29890 20698
rect 29890 20646 29900 20698
rect 29924 20646 29954 20698
rect 29954 20646 29966 20698
rect 29966 20646 29980 20698
rect 30004 20646 30018 20698
rect 30018 20646 30030 20698
rect 30030 20646 30060 20698
rect 30084 20646 30094 20698
rect 30094 20646 30140 20698
rect 29844 20644 29900 20646
rect 29924 20644 29980 20646
rect 30004 20644 30060 20646
rect 30084 20644 30140 20646
rect 22622 9274 22678 9276
rect 22702 9274 22758 9276
rect 22782 9274 22838 9276
rect 22862 9274 22918 9276
rect 22622 9222 22668 9274
rect 22668 9222 22678 9274
rect 22702 9222 22732 9274
rect 22732 9222 22744 9274
rect 22744 9222 22758 9274
rect 22782 9222 22796 9274
rect 22796 9222 22808 9274
rect 22808 9222 22838 9274
rect 22862 9222 22872 9274
rect 22872 9222 22918 9274
rect 22622 9220 22678 9222
rect 22702 9220 22758 9222
rect 22782 9220 22838 9222
rect 22862 9220 22918 9222
rect 23294 8744 23350 8800
rect 22622 8186 22678 8188
rect 22702 8186 22758 8188
rect 22782 8186 22838 8188
rect 22862 8186 22918 8188
rect 22622 8134 22668 8186
rect 22668 8134 22678 8186
rect 22702 8134 22732 8186
rect 22732 8134 22744 8186
rect 22744 8134 22758 8186
rect 22782 8134 22796 8186
rect 22796 8134 22808 8186
rect 22808 8134 22838 8186
rect 22862 8134 22872 8186
rect 22872 8134 22918 8186
rect 22622 8132 22678 8134
rect 22702 8132 22758 8134
rect 22782 8132 22838 8134
rect 22862 8132 22918 8134
rect 22622 7098 22678 7100
rect 22702 7098 22758 7100
rect 22782 7098 22838 7100
rect 22862 7098 22918 7100
rect 22622 7046 22668 7098
rect 22668 7046 22678 7098
rect 22702 7046 22732 7098
rect 22732 7046 22744 7098
rect 22744 7046 22758 7098
rect 22782 7046 22796 7098
rect 22796 7046 22808 7098
rect 22808 7046 22838 7098
rect 22862 7046 22872 7098
rect 22872 7046 22918 7098
rect 22622 7044 22678 7046
rect 22702 7044 22758 7046
rect 22782 7044 22838 7046
rect 22862 7044 22918 7046
rect 22622 6010 22678 6012
rect 22702 6010 22758 6012
rect 22782 6010 22838 6012
rect 22862 6010 22918 6012
rect 22622 5958 22668 6010
rect 22668 5958 22678 6010
rect 22702 5958 22732 6010
rect 22732 5958 22744 6010
rect 22744 5958 22758 6010
rect 22782 5958 22796 6010
rect 22796 5958 22808 6010
rect 22808 5958 22838 6010
rect 22862 5958 22872 6010
rect 22872 5958 22918 6010
rect 22622 5956 22678 5958
rect 22702 5956 22758 5958
rect 22782 5956 22838 5958
rect 22862 5956 22918 5958
rect 22622 4922 22678 4924
rect 22702 4922 22758 4924
rect 22782 4922 22838 4924
rect 22862 4922 22918 4924
rect 22622 4870 22668 4922
rect 22668 4870 22678 4922
rect 22702 4870 22732 4922
rect 22732 4870 22744 4922
rect 22744 4870 22758 4922
rect 22782 4870 22796 4922
rect 22796 4870 22808 4922
rect 22808 4870 22838 4922
rect 22862 4870 22872 4922
rect 22872 4870 22918 4922
rect 22622 4868 22678 4870
rect 22702 4868 22758 4870
rect 22782 4868 22838 4870
rect 22862 4868 22918 4870
rect 22622 3834 22678 3836
rect 22702 3834 22758 3836
rect 22782 3834 22838 3836
rect 22862 3834 22918 3836
rect 22622 3782 22668 3834
rect 22668 3782 22678 3834
rect 22702 3782 22732 3834
rect 22732 3782 22744 3834
rect 22744 3782 22758 3834
rect 22782 3782 22796 3834
rect 22796 3782 22808 3834
rect 22808 3782 22838 3834
rect 22862 3782 22872 3834
rect 22872 3782 22918 3834
rect 22622 3780 22678 3782
rect 22702 3780 22758 3782
rect 22782 3780 22838 3782
rect 22862 3780 22918 3782
rect 23386 5652 23388 5672
rect 23388 5652 23440 5672
rect 23440 5652 23442 5672
rect 23386 5616 23442 5652
rect 24766 5616 24822 5672
rect 22622 2746 22678 2748
rect 22702 2746 22758 2748
rect 22782 2746 22838 2748
rect 22862 2746 22918 2748
rect 22622 2694 22668 2746
rect 22668 2694 22678 2746
rect 22702 2694 22732 2746
rect 22732 2694 22744 2746
rect 22744 2694 22758 2746
rect 22782 2694 22796 2746
rect 22796 2694 22808 2746
rect 22808 2694 22838 2746
rect 22862 2694 22872 2746
rect 22872 2694 22918 2746
rect 22622 2692 22678 2694
rect 22702 2692 22758 2694
rect 22782 2692 22838 2694
rect 22862 2692 22918 2694
rect 26974 17740 27030 17776
rect 26974 17720 26976 17740
rect 26976 17720 27028 17740
rect 27028 17720 27030 17740
rect 37066 21242 37122 21244
rect 37146 21242 37202 21244
rect 37226 21242 37282 21244
rect 37306 21242 37362 21244
rect 37066 21190 37112 21242
rect 37112 21190 37122 21242
rect 37146 21190 37176 21242
rect 37176 21190 37188 21242
rect 37188 21190 37202 21242
rect 37226 21190 37240 21242
rect 37240 21190 37252 21242
rect 37252 21190 37282 21242
rect 37306 21190 37316 21242
rect 37316 21190 37362 21242
rect 37066 21188 37122 21190
rect 37146 21188 37202 21190
rect 37226 21188 37282 21190
rect 37306 21188 37362 21190
rect 29844 19610 29900 19612
rect 29924 19610 29980 19612
rect 30004 19610 30060 19612
rect 30084 19610 30140 19612
rect 29844 19558 29890 19610
rect 29890 19558 29900 19610
rect 29924 19558 29954 19610
rect 29954 19558 29966 19610
rect 29966 19558 29980 19610
rect 30004 19558 30018 19610
rect 30018 19558 30030 19610
rect 30030 19558 30060 19610
rect 30084 19558 30094 19610
rect 30094 19558 30140 19610
rect 29844 19556 29900 19558
rect 29924 19556 29980 19558
rect 30004 19556 30060 19558
rect 30084 19556 30140 19558
rect 29844 18522 29900 18524
rect 29924 18522 29980 18524
rect 30004 18522 30060 18524
rect 30084 18522 30140 18524
rect 29844 18470 29890 18522
rect 29890 18470 29900 18522
rect 29924 18470 29954 18522
rect 29954 18470 29966 18522
rect 29966 18470 29980 18522
rect 30004 18470 30018 18522
rect 30018 18470 30030 18522
rect 30030 18470 30060 18522
rect 30084 18470 30094 18522
rect 30094 18470 30140 18522
rect 29844 18468 29900 18470
rect 29924 18468 29980 18470
rect 30004 18468 30060 18470
rect 30084 18468 30140 18470
rect 29844 17434 29900 17436
rect 29924 17434 29980 17436
rect 30004 17434 30060 17436
rect 30084 17434 30140 17436
rect 29844 17382 29890 17434
rect 29890 17382 29900 17434
rect 29924 17382 29954 17434
rect 29954 17382 29966 17434
rect 29966 17382 29980 17434
rect 30004 17382 30018 17434
rect 30018 17382 30030 17434
rect 30030 17382 30060 17434
rect 30084 17382 30094 17434
rect 30094 17382 30140 17434
rect 29844 17380 29900 17382
rect 29924 17380 29980 17382
rect 30004 17380 30060 17382
rect 30084 17380 30140 17382
rect 27342 3984 27398 4040
rect 27342 3032 27398 3088
rect 28906 8744 28962 8800
rect 29844 16346 29900 16348
rect 29924 16346 29980 16348
rect 30004 16346 30060 16348
rect 30084 16346 30140 16348
rect 29844 16294 29890 16346
rect 29890 16294 29900 16346
rect 29924 16294 29954 16346
rect 29954 16294 29966 16346
rect 29966 16294 29980 16346
rect 30004 16294 30018 16346
rect 30018 16294 30030 16346
rect 30030 16294 30060 16346
rect 30084 16294 30094 16346
rect 30094 16294 30140 16346
rect 29844 16292 29900 16294
rect 29924 16292 29980 16294
rect 30004 16292 30060 16294
rect 30084 16292 30140 16294
rect 29844 15258 29900 15260
rect 29924 15258 29980 15260
rect 30004 15258 30060 15260
rect 30084 15258 30140 15260
rect 29844 15206 29890 15258
rect 29890 15206 29900 15258
rect 29924 15206 29954 15258
rect 29954 15206 29966 15258
rect 29966 15206 29980 15258
rect 30004 15206 30018 15258
rect 30018 15206 30030 15258
rect 30030 15206 30060 15258
rect 30084 15206 30094 15258
rect 30094 15206 30140 15258
rect 29844 15204 29900 15206
rect 29924 15204 29980 15206
rect 30004 15204 30060 15206
rect 30084 15204 30140 15206
rect 29844 14170 29900 14172
rect 29924 14170 29980 14172
rect 30004 14170 30060 14172
rect 30084 14170 30140 14172
rect 29844 14118 29890 14170
rect 29890 14118 29900 14170
rect 29924 14118 29954 14170
rect 29954 14118 29966 14170
rect 29966 14118 29980 14170
rect 30004 14118 30018 14170
rect 30018 14118 30030 14170
rect 30030 14118 30060 14170
rect 30084 14118 30094 14170
rect 30094 14118 30140 14170
rect 29844 14116 29900 14118
rect 29924 14116 29980 14118
rect 30004 14116 30060 14118
rect 30084 14116 30140 14118
rect 29844 13082 29900 13084
rect 29924 13082 29980 13084
rect 30004 13082 30060 13084
rect 30084 13082 30140 13084
rect 29844 13030 29890 13082
rect 29890 13030 29900 13082
rect 29924 13030 29954 13082
rect 29954 13030 29966 13082
rect 29966 13030 29980 13082
rect 30004 13030 30018 13082
rect 30018 13030 30030 13082
rect 30030 13030 30060 13082
rect 30084 13030 30094 13082
rect 30094 13030 30140 13082
rect 29844 13028 29900 13030
rect 29924 13028 29980 13030
rect 30004 13028 30060 13030
rect 30084 13028 30140 13030
rect 29844 11994 29900 11996
rect 29924 11994 29980 11996
rect 30004 11994 30060 11996
rect 30084 11994 30140 11996
rect 29844 11942 29890 11994
rect 29890 11942 29900 11994
rect 29924 11942 29954 11994
rect 29954 11942 29966 11994
rect 29966 11942 29980 11994
rect 30004 11942 30018 11994
rect 30018 11942 30030 11994
rect 30030 11942 30060 11994
rect 30084 11942 30094 11994
rect 30094 11942 30140 11994
rect 29844 11940 29900 11942
rect 29924 11940 29980 11942
rect 30004 11940 30060 11942
rect 30084 11940 30140 11942
rect 29844 10906 29900 10908
rect 29924 10906 29980 10908
rect 30004 10906 30060 10908
rect 30084 10906 30140 10908
rect 29844 10854 29890 10906
rect 29890 10854 29900 10906
rect 29924 10854 29954 10906
rect 29954 10854 29966 10906
rect 29966 10854 29980 10906
rect 30004 10854 30018 10906
rect 30018 10854 30030 10906
rect 30030 10854 30060 10906
rect 30084 10854 30094 10906
rect 30094 10854 30140 10906
rect 29844 10852 29900 10854
rect 29924 10852 29980 10854
rect 30004 10852 30060 10854
rect 30084 10852 30140 10854
rect 29918 9968 29974 10024
rect 29844 9818 29900 9820
rect 29924 9818 29980 9820
rect 30004 9818 30060 9820
rect 30084 9818 30140 9820
rect 29844 9766 29890 9818
rect 29890 9766 29900 9818
rect 29924 9766 29954 9818
rect 29954 9766 29966 9818
rect 29966 9766 29980 9818
rect 30004 9766 30018 9818
rect 30018 9766 30030 9818
rect 30030 9766 30060 9818
rect 30084 9766 30094 9818
rect 30094 9766 30140 9818
rect 29844 9764 29900 9766
rect 29924 9764 29980 9766
rect 30004 9764 30060 9766
rect 30084 9764 30140 9766
rect 27802 3032 27858 3088
rect 29844 8730 29900 8732
rect 29924 8730 29980 8732
rect 30004 8730 30060 8732
rect 30084 8730 30140 8732
rect 29844 8678 29890 8730
rect 29890 8678 29900 8730
rect 29924 8678 29954 8730
rect 29954 8678 29966 8730
rect 29966 8678 29980 8730
rect 30004 8678 30018 8730
rect 30018 8678 30030 8730
rect 30030 8678 30060 8730
rect 30084 8678 30094 8730
rect 30094 8678 30140 8730
rect 29844 8676 29900 8678
rect 29924 8676 29980 8678
rect 30004 8676 30060 8678
rect 30084 8676 30140 8678
rect 29844 7642 29900 7644
rect 29924 7642 29980 7644
rect 30004 7642 30060 7644
rect 30084 7642 30140 7644
rect 29844 7590 29890 7642
rect 29890 7590 29900 7642
rect 29924 7590 29954 7642
rect 29954 7590 29966 7642
rect 29966 7590 29980 7642
rect 30004 7590 30018 7642
rect 30018 7590 30030 7642
rect 30030 7590 30060 7642
rect 30084 7590 30094 7642
rect 30094 7590 30140 7642
rect 29844 7588 29900 7590
rect 29924 7588 29980 7590
rect 30004 7588 30060 7590
rect 30084 7588 30140 7590
rect 29844 6554 29900 6556
rect 29924 6554 29980 6556
rect 30004 6554 30060 6556
rect 30084 6554 30140 6556
rect 29844 6502 29890 6554
rect 29890 6502 29900 6554
rect 29924 6502 29954 6554
rect 29954 6502 29966 6554
rect 29966 6502 29980 6554
rect 30004 6502 30018 6554
rect 30018 6502 30030 6554
rect 30030 6502 30060 6554
rect 30084 6502 30094 6554
rect 30094 6502 30140 6554
rect 29844 6500 29900 6502
rect 29924 6500 29980 6502
rect 30004 6500 30060 6502
rect 30084 6500 30140 6502
rect 30010 6060 30012 6080
rect 30012 6060 30064 6080
rect 30064 6060 30066 6080
rect 30010 6024 30066 6060
rect 29844 5466 29900 5468
rect 29924 5466 29980 5468
rect 30004 5466 30060 5468
rect 30084 5466 30140 5468
rect 29844 5414 29890 5466
rect 29890 5414 29900 5466
rect 29924 5414 29954 5466
rect 29954 5414 29966 5466
rect 29966 5414 29980 5466
rect 30004 5414 30018 5466
rect 30018 5414 30030 5466
rect 30030 5414 30060 5466
rect 30084 5414 30094 5466
rect 30094 5414 30140 5466
rect 29844 5412 29900 5414
rect 29924 5412 29980 5414
rect 30004 5412 30060 5414
rect 30084 5412 30140 5414
rect 29844 4378 29900 4380
rect 29924 4378 29980 4380
rect 30004 4378 30060 4380
rect 30084 4378 30140 4380
rect 29844 4326 29890 4378
rect 29890 4326 29900 4378
rect 29924 4326 29954 4378
rect 29954 4326 29966 4378
rect 29966 4326 29980 4378
rect 30004 4326 30018 4378
rect 30018 4326 30030 4378
rect 30030 4326 30060 4378
rect 30084 4326 30094 4378
rect 30094 4326 30140 4378
rect 29844 4324 29900 4326
rect 29924 4324 29980 4326
rect 30004 4324 30060 4326
rect 30084 4324 30140 4326
rect 30470 6160 30526 6216
rect 30562 5888 30618 5944
rect 30194 3440 30250 3496
rect 29844 3290 29900 3292
rect 29924 3290 29980 3292
rect 30004 3290 30060 3292
rect 30084 3290 30140 3292
rect 29844 3238 29890 3290
rect 29890 3238 29900 3290
rect 29924 3238 29954 3290
rect 29954 3238 29966 3290
rect 29966 3238 29980 3290
rect 30004 3238 30018 3290
rect 30018 3238 30030 3290
rect 30030 3238 30060 3290
rect 30084 3238 30094 3290
rect 30094 3238 30140 3290
rect 29844 3236 29900 3238
rect 29924 3236 29980 3238
rect 30004 3236 30060 3238
rect 30084 3236 30140 3238
rect 31206 4700 31208 4720
rect 31208 4700 31260 4720
rect 31260 4700 31262 4720
rect 31206 4664 31262 4700
rect 31206 3168 31262 3224
rect 31850 6024 31906 6080
rect 32770 6160 32826 6216
rect 29844 2202 29900 2204
rect 29924 2202 29980 2204
rect 30004 2202 30060 2204
rect 30084 2202 30140 2204
rect 29844 2150 29890 2202
rect 29890 2150 29900 2202
rect 29924 2150 29954 2202
rect 29954 2150 29966 2202
rect 29966 2150 29980 2202
rect 30004 2150 30018 2202
rect 30018 2150 30030 2202
rect 30030 2150 30060 2202
rect 30084 2150 30094 2202
rect 30094 2150 30140 2202
rect 29844 2148 29900 2150
rect 29924 2148 29980 2150
rect 30004 2148 30060 2150
rect 30084 2148 30140 2150
rect 32954 5908 33010 5944
rect 32954 5888 32956 5908
rect 32956 5888 33008 5908
rect 33008 5888 33010 5908
rect 33414 6296 33470 6352
rect 33322 4548 33378 4584
rect 33322 4528 33324 4548
rect 33324 4528 33376 4548
rect 33376 4528 33378 4548
rect 33414 4120 33470 4176
rect 32954 3848 33010 3904
rect 34058 3168 34114 3224
rect 32310 2896 32366 2952
rect 34702 5752 34758 5808
rect 34886 4800 34942 4856
rect 37066 20154 37122 20156
rect 37146 20154 37202 20156
rect 37226 20154 37282 20156
rect 37306 20154 37362 20156
rect 37066 20102 37112 20154
rect 37112 20102 37122 20154
rect 37146 20102 37176 20154
rect 37176 20102 37188 20154
rect 37188 20102 37202 20154
rect 37226 20102 37240 20154
rect 37240 20102 37252 20154
rect 37252 20102 37282 20154
rect 37306 20102 37316 20154
rect 37316 20102 37362 20154
rect 37066 20100 37122 20102
rect 37146 20100 37202 20102
rect 37226 20100 37282 20102
rect 37306 20100 37362 20102
rect 44288 22874 44344 22876
rect 44368 22874 44424 22876
rect 44448 22874 44504 22876
rect 44528 22874 44584 22876
rect 44288 22822 44334 22874
rect 44334 22822 44344 22874
rect 44368 22822 44398 22874
rect 44398 22822 44410 22874
rect 44410 22822 44424 22874
rect 44448 22822 44462 22874
rect 44462 22822 44474 22874
rect 44474 22822 44504 22874
rect 44528 22822 44538 22874
rect 44538 22822 44584 22874
rect 44288 22820 44344 22822
rect 44368 22820 44424 22822
rect 44448 22820 44504 22822
rect 44528 22820 44584 22822
rect 37066 19066 37122 19068
rect 37146 19066 37202 19068
rect 37226 19066 37282 19068
rect 37306 19066 37362 19068
rect 37066 19014 37112 19066
rect 37112 19014 37122 19066
rect 37146 19014 37176 19066
rect 37176 19014 37188 19066
rect 37188 19014 37202 19066
rect 37226 19014 37240 19066
rect 37240 19014 37252 19066
rect 37252 19014 37282 19066
rect 37306 19014 37316 19066
rect 37316 19014 37362 19066
rect 37066 19012 37122 19014
rect 37146 19012 37202 19014
rect 37226 19012 37282 19014
rect 37306 19012 37362 19014
rect 35162 3984 35218 4040
rect 37066 17978 37122 17980
rect 37146 17978 37202 17980
rect 37226 17978 37282 17980
rect 37306 17978 37362 17980
rect 37066 17926 37112 17978
rect 37112 17926 37122 17978
rect 37146 17926 37176 17978
rect 37176 17926 37188 17978
rect 37188 17926 37202 17978
rect 37226 17926 37240 17978
rect 37240 17926 37252 17978
rect 37252 17926 37282 17978
rect 37306 17926 37316 17978
rect 37316 17926 37362 17978
rect 37066 17924 37122 17926
rect 37146 17924 37202 17926
rect 37226 17924 37282 17926
rect 37306 17924 37362 17926
rect 37066 16890 37122 16892
rect 37146 16890 37202 16892
rect 37226 16890 37282 16892
rect 37306 16890 37362 16892
rect 37066 16838 37112 16890
rect 37112 16838 37122 16890
rect 37146 16838 37176 16890
rect 37176 16838 37188 16890
rect 37188 16838 37202 16890
rect 37226 16838 37240 16890
rect 37240 16838 37252 16890
rect 37252 16838 37282 16890
rect 37306 16838 37316 16890
rect 37316 16838 37362 16890
rect 37066 16836 37122 16838
rect 37146 16836 37202 16838
rect 37226 16836 37282 16838
rect 37306 16836 37362 16838
rect 37066 15802 37122 15804
rect 37146 15802 37202 15804
rect 37226 15802 37282 15804
rect 37306 15802 37362 15804
rect 37066 15750 37112 15802
rect 37112 15750 37122 15802
rect 37146 15750 37176 15802
rect 37176 15750 37188 15802
rect 37188 15750 37202 15802
rect 37226 15750 37240 15802
rect 37240 15750 37252 15802
rect 37252 15750 37282 15802
rect 37306 15750 37316 15802
rect 37316 15750 37362 15802
rect 37066 15748 37122 15750
rect 37146 15748 37202 15750
rect 37226 15748 37282 15750
rect 37306 15748 37362 15750
rect 37066 14714 37122 14716
rect 37146 14714 37202 14716
rect 37226 14714 37282 14716
rect 37306 14714 37362 14716
rect 37066 14662 37112 14714
rect 37112 14662 37122 14714
rect 37146 14662 37176 14714
rect 37176 14662 37188 14714
rect 37188 14662 37202 14714
rect 37226 14662 37240 14714
rect 37240 14662 37252 14714
rect 37252 14662 37282 14714
rect 37306 14662 37316 14714
rect 37316 14662 37362 14714
rect 37066 14660 37122 14662
rect 37146 14660 37202 14662
rect 37226 14660 37282 14662
rect 37306 14660 37362 14662
rect 37066 13626 37122 13628
rect 37146 13626 37202 13628
rect 37226 13626 37282 13628
rect 37306 13626 37362 13628
rect 37066 13574 37112 13626
rect 37112 13574 37122 13626
rect 37146 13574 37176 13626
rect 37176 13574 37188 13626
rect 37188 13574 37202 13626
rect 37226 13574 37240 13626
rect 37240 13574 37252 13626
rect 37252 13574 37282 13626
rect 37306 13574 37316 13626
rect 37316 13574 37362 13626
rect 37066 13572 37122 13574
rect 37146 13572 37202 13574
rect 37226 13572 37282 13574
rect 37306 13572 37362 13574
rect 39210 19760 39266 19816
rect 44288 21786 44344 21788
rect 44368 21786 44424 21788
rect 44448 21786 44504 21788
rect 44528 21786 44584 21788
rect 44288 21734 44334 21786
rect 44334 21734 44344 21786
rect 44368 21734 44398 21786
rect 44398 21734 44410 21786
rect 44410 21734 44424 21786
rect 44448 21734 44462 21786
rect 44462 21734 44474 21786
rect 44474 21734 44504 21786
rect 44528 21734 44538 21786
rect 44538 21734 44584 21786
rect 44288 21732 44344 21734
rect 44368 21732 44424 21734
rect 44448 21732 44504 21734
rect 44528 21732 44584 21734
rect 37066 12538 37122 12540
rect 37146 12538 37202 12540
rect 37226 12538 37282 12540
rect 37306 12538 37362 12540
rect 37066 12486 37112 12538
rect 37112 12486 37122 12538
rect 37146 12486 37176 12538
rect 37176 12486 37188 12538
rect 37188 12486 37202 12538
rect 37226 12486 37240 12538
rect 37240 12486 37252 12538
rect 37252 12486 37282 12538
rect 37306 12486 37316 12538
rect 37316 12486 37362 12538
rect 37066 12484 37122 12486
rect 37146 12484 37202 12486
rect 37226 12484 37282 12486
rect 37306 12484 37362 12486
rect 37066 11450 37122 11452
rect 37146 11450 37202 11452
rect 37226 11450 37282 11452
rect 37306 11450 37362 11452
rect 37066 11398 37112 11450
rect 37112 11398 37122 11450
rect 37146 11398 37176 11450
rect 37176 11398 37188 11450
rect 37188 11398 37202 11450
rect 37226 11398 37240 11450
rect 37240 11398 37252 11450
rect 37252 11398 37282 11450
rect 37306 11398 37316 11450
rect 37316 11398 37362 11450
rect 37066 11396 37122 11398
rect 37146 11396 37202 11398
rect 37226 11396 37282 11398
rect 37306 11396 37362 11398
rect 37066 10362 37122 10364
rect 37146 10362 37202 10364
rect 37226 10362 37282 10364
rect 37306 10362 37362 10364
rect 37066 10310 37112 10362
rect 37112 10310 37122 10362
rect 37146 10310 37176 10362
rect 37176 10310 37188 10362
rect 37188 10310 37202 10362
rect 37226 10310 37240 10362
rect 37240 10310 37252 10362
rect 37252 10310 37282 10362
rect 37306 10310 37316 10362
rect 37316 10310 37362 10362
rect 37066 10308 37122 10310
rect 37146 10308 37202 10310
rect 37226 10308 37282 10310
rect 37306 10308 37362 10310
rect 37066 9274 37122 9276
rect 37146 9274 37202 9276
rect 37226 9274 37282 9276
rect 37306 9274 37362 9276
rect 37066 9222 37112 9274
rect 37112 9222 37122 9274
rect 37146 9222 37176 9274
rect 37176 9222 37188 9274
rect 37188 9222 37202 9274
rect 37226 9222 37240 9274
rect 37240 9222 37252 9274
rect 37252 9222 37282 9274
rect 37306 9222 37316 9274
rect 37316 9222 37362 9274
rect 37066 9220 37122 9222
rect 37146 9220 37202 9222
rect 37226 9220 37282 9222
rect 37306 9220 37362 9222
rect 37066 8186 37122 8188
rect 37146 8186 37202 8188
rect 37226 8186 37282 8188
rect 37306 8186 37362 8188
rect 37066 8134 37112 8186
rect 37112 8134 37122 8186
rect 37146 8134 37176 8186
rect 37176 8134 37188 8186
rect 37188 8134 37202 8186
rect 37226 8134 37240 8186
rect 37240 8134 37252 8186
rect 37252 8134 37282 8186
rect 37306 8134 37316 8186
rect 37316 8134 37362 8186
rect 37066 8132 37122 8134
rect 37146 8132 37202 8134
rect 37226 8132 37282 8134
rect 37306 8132 37362 8134
rect 37066 7098 37122 7100
rect 37146 7098 37202 7100
rect 37226 7098 37282 7100
rect 37306 7098 37362 7100
rect 37066 7046 37112 7098
rect 37112 7046 37122 7098
rect 37146 7046 37176 7098
rect 37176 7046 37188 7098
rect 37188 7046 37202 7098
rect 37226 7046 37240 7098
rect 37240 7046 37252 7098
rect 37252 7046 37282 7098
rect 37306 7046 37316 7098
rect 37316 7046 37362 7098
rect 37066 7044 37122 7046
rect 37146 7044 37202 7046
rect 37226 7044 37282 7046
rect 37306 7044 37362 7046
rect 37462 6840 37518 6896
rect 34610 2896 34666 2952
rect 34886 3168 34942 3224
rect 35162 2896 35218 2952
rect 37066 6010 37122 6012
rect 37146 6010 37202 6012
rect 37226 6010 37282 6012
rect 37306 6010 37362 6012
rect 37066 5958 37112 6010
rect 37112 5958 37122 6010
rect 37146 5958 37176 6010
rect 37176 5958 37188 6010
rect 37188 5958 37202 6010
rect 37226 5958 37240 6010
rect 37240 5958 37252 6010
rect 37252 5958 37282 6010
rect 37306 5958 37316 6010
rect 37316 5958 37362 6010
rect 37066 5956 37122 5958
rect 37146 5956 37202 5958
rect 37226 5956 37282 5958
rect 37306 5956 37362 5958
rect 37066 4922 37122 4924
rect 37146 4922 37202 4924
rect 37226 4922 37282 4924
rect 37306 4922 37362 4924
rect 37066 4870 37112 4922
rect 37112 4870 37122 4922
rect 37146 4870 37176 4922
rect 37176 4870 37188 4922
rect 37188 4870 37202 4922
rect 37226 4870 37240 4922
rect 37240 4870 37252 4922
rect 37252 4870 37282 4922
rect 37306 4870 37316 4922
rect 37316 4870 37362 4922
rect 37066 4868 37122 4870
rect 37146 4868 37202 4870
rect 37226 4868 37282 4870
rect 37306 4868 37362 4870
rect 37278 3984 37334 4040
rect 37066 3834 37122 3836
rect 37146 3834 37202 3836
rect 37226 3834 37282 3836
rect 37306 3834 37362 3836
rect 37066 3782 37112 3834
rect 37112 3782 37122 3834
rect 37146 3782 37176 3834
rect 37176 3782 37188 3834
rect 37188 3782 37202 3834
rect 37226 3782 37240 3834
rect 37240 3782 37252 3834
rect 37252 3782 37282 3834
rect 37306 3782 37316 3834
rect 37316 3782 37362 3834
rect 37066 3780 37122 3782
rect 37146 3780 37202 3782
rect 37226 3780 37282 3782
rect 37306 3780 37362 3782
rect 37066 2746 37122 2748
rect 37146 2746 37202 2748
rect 37226 2746 37282 2748
rect 37306 2746 37362 2748
rect 37066 2694 37112 2746
rect 37112 2694 37122 2746
rect 37146 2694 37176 2746
rect 37176 2694 37188 2746
rect 37188 2694 37202 2746
rect 37226 2694 37240 2746
rect 37240 2694 37252 2746
rect 37252 2694 37282 2746
rect 37306 2694 37316 2746
rect 37316 2694 37362 2746
rect 37066 2692 37122 2694
rect 37146 2692 37202 2694
rect 37226 2692 37282 2694
rect 37306 2692 37362 2694
rect 39026 5616 39082 5672
rect 38014 4664 38070 4720
rect 39946 16496 40002 16552
rect 41326 19352 41382 19408
rect 41602 16496 41658 16552
rect 44288 20698 44344 20700
rect 44368 20698 44424 20700
rect 44448 20698 44504 20700
rect 44528 20698 44584 20700
rect 44288 20646 44334 20698
rect 44334 20646 44344 20698
rect 44368 20646 44398 20698
rect 44398 20646 44410 20698
rect 44410 20646 44424 20698
rect 44448 20646 44462 20698
rect 44462 20646 44474 20698
rect 44474 20646 44504 20698
rect 44528 20646 44538 20698
rect 44538 20646 44584 20698
rect 44288 20644 44344 20646
rect 44368 20644 44424 20646
rect 44448 20644 44504 20646
rect 44528 20644 44584 20646
rect 43074 20440 43130 20496
rect 39486 3168 39542 3224
rect 38750 2896 38806 2952
rect 41326 4020 41328 4040
rect 41328 4020 41380 4040
rect 41380 4020 41382 4040
rect 41326 3984 41382 4020
rect 44288 19610 44344 19612
rect 44368 19610 44424 19612
rect 44448 19610 44504 19612
rect 44528 19610 44584 19612
rect 44288 19558 44334 19610
rect 44334 19558 44344 19610
rect 44368 19558 44398 19610
rect 44398 19558 44410 19610
rect 44410 19558 44424 19610
rect 44448 19558 44462 19610
rect 44462 19558 44474 19610
rect 44474 19558 44504 19610
rect 44528 19558 44538 19610
rect 44538 19558 44584 19610
rect 44288 19556 44344 19558
rect 44368 19556 44424 19558
rect 44448 19556 44504 19558
rect 44528 19556 44584 19558
rect 46478 20440 46534 20496
rect 45466 19760 45522 19816
rect 58732 22874 58788 22876
rect 58812 22874 58868 22876
rect 58892 22874 58948 22876
rect 58972 22874 59028 22876
rect 58732 22822 58778 22874
rect 58778 22822 58788 22874
rect 58812 22822 58842 22874
rect 58842 22822 58854 22874
rect 58854 22822 58868 22874
rect 58892 22822 58906 22874
rect 58906 22822 58918 22874
rect 58918 22822 58948 22874
rect 58972 22822 58982 22874
rect 58982 22822 59028 22874
rect 58732 22820 58788 22822
rect 58812 22820 58868 22822
rect 58892 22820 58948 22822
rect 58972 22820 59028 22822
rect 47858 20324 47914 20360
rect 47858 20304 47860 20324
rect 47860 20304 47912 20324
rect 47912 20304 47914 20324
rect 44288 18522 44344 18524
rect 44368 18522 44424 18524
rect 44448 18522 44504 18524
rect 44528 18522 44584 18524
rect 44288 18470 44334 18522
rect 44334 18470 44344 18522
rect 44368 18470 44398 18522
rect 44398 18470 44410 18522
rect 44410 18470 44424 18522
rect 44448 18470 44462 18522
rect 44462 18470 44474 18522
rect 44474 18470 44504 18522
rect 44528 18470 44538 18522
rect 44538 18470 44584 18522
rect 44288 18468 44344 18470
rect 44368 18468 44424 18470
rect 44448 18468 44504 18470
rect 44528 18468 44584 18470
rect 44288 17434 44344 17436
rect 44368 17434 44424 17436
rect 44448 17434 44504 17436
rect 44528 17434 44584 17436
rect 44288 17382 44334 17434
rect 44334 17382 44344 17434
rect 44368 17382 44398 17434
rect 44398 17382 44410 17434
rect 44410 17382 44424 17434
rect 44448 17382 44462 17434
rect 44462 17382 44474 17434
rect 44474 17382 44504 17434
rect 44528 17382 44538 17434
rect 44538 17382 44584 17434
rect 44288 17380 44344 17382
rect 44368 17380 44424 17382
rect 44448 17380 44504 17382
rect 44528 17380 44584 17382
rect 44288 16346 44344 16348
rect 44368 16346 44424 16348
rect 44448 16346 44504 16348
rect 44528 16346 44584 16348
rect 44288 16294 44334 16346
rect 44334 16294 44344 16346
rect 44368 16294 44398 16346
rect 44398 16294 44410 16346
rect 44410 16294 44424 16346
rect 44448 16294 44462 16346
rect 44462 16294 44474 16346
rect 44474 16294 44504 16346
rect 44528 16294 44538 16346
rect 44538 16294 44584 16346
rect 44288 16292 44344 16294
rect 44368 16292 44424 16294
rect 44448 16292 44504 16294
rect 44528 16292 44584 16294
rect 41970 6840 42026 6896
rect 42430 4528 42486 4584
rect 44288 15258 44344 15260
rect 44368 15258 44424 15260
rect 44448 15258 44504 15260
rect 44528 15258 44584 15260
rect 44288 15206 44334 15258
rect 44334 15206 44344 15258
rect 44368 15206 44398 15258
rect 44398 15206 44410 15258
rect 44410 15206 44424 15258
rect 44448 15206 44462 15258
rect 44462 15206 44474 15258
rect 44474 15206 44504 15258
rect 44528 15206 44538 15258
rect 44538 15206 44584 15258
rect 44288 15204 44344 15206
rect 44368 15204 44424 15206
rect 44448 15204 44504 15206
rect 44528 15204 44584 15206
rect 44288 14170 44344 14172
rect 44368 14170 44424 14172
rect 44448 14170 44504 14172
rect 44528 14170 44584 14172
rect 44288 14118 44334 14170
rect 44334 14118 44344 14170
rect 44368 14118 44398 14170
rect 44398 14118 44410 14170
rect 44410 14118 44424 14170
rect 44448 14118 44462 14170
rect 44462 14118 44474 14170
rect 44474 14118 44504 14170
rect 44528 14118 44538 14170
rect 44538 14118 44584 14170
rect 44288 14116 44344 14118
rect 44368 14116 44424 14118
rect 44448 14116 44504 14118
rect 44528 14116 44584 14118
rect 44288 13082 44344 13084
rect 44368 13082 44424 13084
rect 44448 13082 44504 13084
rect 44528 13082 44584 13084
rect 44288 13030 44334 13082
rect 44334 13030 44344 13082
rect 44368 13030 44398 13082
rect 44398 13030 44410 13082
rect 44410 13030 44424 13082
rect 44448 13030 44462 13082
rect 44462 13030 44474 13082
rect 44474 13030 44504 13082
rect 44528 13030 44538 13082
rect 44538 13030 44584 13082
rect 44288 13028 44344 13030
rect 44368 13028 44424 13030
rect 44448 13028 44504 13030
rect 44528 13028 44584 13030
rect 44288 11994 44344 11996
rect 44368 11994 44424 11996
rect 44448 11994 44504 11996
rect 44528 11994 44584 11996
rect 44288 11942 44334 11994
rect 44334 11942 44344 11994
rect 44368 11942 44398 11994
rect 44398 11942 44410 11994
rect 44410 11942 44424 11994
rect 44448 11942 44462 11994
rect 44462 11942 44474 11994
rect 44474 11942 44504 11994
rect 44528 11942 44538 11994
rect 44538 11942 44584 11994
rect 44288 11940 44344 11942
rect 44368 11940 44424 11942
rect 44448 11940 44504 11942
rect 44528 11940 44584 11942
rect 51510 22330 51566 22332
rect 51590 22330 51646 22332
rect 51670 22330 51726 22332
rect 51750 22330 51806 22332
rect 51510 22278 51556 22330
rect 51556 22278 51566 22330
rect 51590 22278 51620 22330
rect 51620 22278 51632 22330
rect 51632 22278 51646 22330
rect 51670 22278 51684 22330
rect 51684 22278 51696 22330
rect 51696 22278 51726 22330
rect 51750 22278 51760 22330
rect 51760 22278 51806 22330
rect 51510 22276 51566 22278
rect 51590 22276 51646 22278
rect 51670 22276 51726 22278
rect 51750 22276 51806 22278
rect 51354 21528 51410 21584
rect 44288 10906 44344 10908
rect 44368 10906 44424 10908
rect 44448 10906 44504 10908
rect 44528 10906 44584 10908
rect 44288 10854 44334 10906
rect 44334 10854 44344 10906
rect 44368 10854 44398 10906
rect 44398 10854 44410 10906
rect 44410 10854 44424 10906
rect 44448 10854 44462 10906
rect 44462 10854 44474 10906
rect 44474 10854 44504 10906
rect 44528 10854 44538 10906
rect 44538 10854 44584 10906
rect 44288 10852 44344 10854
rect 44368 10852 44424 10854
rect 44448 10852 44504 10854
rect 44528 10852 44584 10854
rect 44288 9818 44344 9820
rect 44368 9818 44424 9820
rect 44448 9818 44504 9820
rect 44528 9818 44584 9820
rect 44288 9766 44334 9818
rect 44334 9766 44344 9818
rect 44368 9766 44398 9818
rect 44398 9766 44410 9818
rect 44410 9766 44424 9818
rect 44448 9766 44462 9818
rect 44462 9766 44474 9818
rect 44474 9766 44504 9818
rect 44528 9766 44538 9818
rect 44538 9766 44584 9818
rect 44288 9764 44344 9766
rect 44368 9764 44424 9766
rect 44448 9764 44504 9766
rect 44528 9764 44584 9766
rect 44288 8730 44344 8732
rect 44368 8730 44424 8732
rect 44448 8730 44504 8732
rect 44528 8730 44584 8732
rect 44288 8678 44334 8730
rect 44334 8678 44344 8730
rect 44368 8678 44398 8730
rect 44398 8678 44410 8730
rect 44410 8678 44424 8730
rect 44448 8678 44462 8730
rect 44462 8678 44474 8730
rect 44474 8678 44504 8730
rect 44528 8678 44538 8730
rect 44538 8678 44584 8730
rect 44288 8676 44344 8678
rect 44368 8676 44424 8678
rect 44448 8676 44504 8678
rect 44528 8676 44584 8678
rect 44288 7642 44344 7644
rect 44368 7642 44424 7644
rect 44448 7642 44504 7644
rect 44528 7642 44584 7644
rect 44288 7590 44334 7642
rect 44334 7590 44344 7642
rect 44368 7590 44398 7642
rect 44398 7590 44410 7642
rect 44410 7590 44424 7642
rect 44448 7590 44462 7642
rect 44462 7590 44474 7642
rect 44474 7590 44504 7642
rect 44528 7590 44538 7642
rect 44538 7590 44584 7642
rect 44288 7588 44344 7590
rect 44368 7588 44424 7590
rect 44448 7588 44504 7590
rect 44528 7588 44584 7590
rect 44288 6554 44344 6556
rect 44368 6554 44424 6556
rect 44448 6554 44504 6556
rect 44528 6554 44584 6556
rect 44288 6502 44334 6554
rect 44334 6502 44344 6554
rect 44368 6502 44398 6554
rect 44398 6502 44410 6554
rect 44410 6502 44424 6554
rect 44448 6502 44462 6554
rect 44462 6502 44474 6554
rect 44474 6502 44504 6554
rect 44528 6502 44538 6554
rect 44538 6502 44584 6554
rect 44288 6500 44344 6502
rect 44368 6500 44424 6502
rect 44448 6500 44504 6502
rect 44528 6500 44584 6502
rect 42890 4020 42892 4040
rect 42892 4020 42944 4040
rect 42944 4020 42946 4040
rect 42338 3032 42394 3088
rect 42890 3984 42946 4020
rect 42890 3032 42946 3088
rect 42798 2896 42854 2952
rect 44288 5466 44344 5468
rect 44368 5466 44424 5468
rect 44448 5466 44504 5468
rect 44528 5466 44584 5468
rect 44288 5414 44334 5466
rect 44334 5414 44344 5466
rect 44368 5414 44398 5466
rect 44398 5414 44410 5466
rect 44410 5414 44424 5466
rect 44448 5414 44462 5466
rect 44462 5414 44474 5466
rect 44474 5414 44504 5466
rect 44528 5414 44538 5466
rect 44538 5414 44584 5466
rect 44288 5412 44344 5414
rect 44368 5412 44424 5414
rect 44448 5412 44504 5414
rect 44528 5412 44584 5414
rect 51510 21242 51566 21244
rect 51590 21242 51646 21244
rect 51670 21242 51726 21244
rect 51750 21242 51806 21244
rect 51510 21190 51556 21242
rect 51556 21190 51566 21242
rect 51590 21190 51620 21242
rect 51620 21190 51632 21242
rect 51632 21190 51646 21242
rect 51670 21190 51684 21242
rect 51684 21190 51696 21242
rect 51696 21190 51726 21242
rect 51750 21190 51760 21242
rect 51760 21190 51806 21242
rect 51510 21188 51566 21190
rect 51590 21188 51646 21190
rect 51670 21188 51726 21190
rect 51750 21188 51806 21190
rect 51998 20848 52054 20904
rect 49330 17584 49386 17640
rect 44730 5616 44786 5672
rect 43810 3440 43866 3496
rect 44288 4378 44344 4380
rect 44368 4378 44424 4380
rect 44448 4378 44504 4380
rect 44528 4378 44584 4380
rect 44288 4326 44334 4378
rect 44334 4326 44344 4378
rect 44368 4326 44398 4378
rect 44398 4326 44410 4378
rect 44410 4326 44424 4378
rect 44448 4326 44462 4378
rect 44462 4326 44474 4378
rect 44474 4326 44504 4378
rect 44528 4326 44538 4378
rect 44538 4326 44584 4378
rect 44288 4324 44344 4326
rect 44368 4324 44424 4326
rect 44448 4324 44504 4326
rect 44528 4324 44584 4326
rect 44288 3290 44344 3292
rect 44368 3290 44424 3292
rect 44448 3290 44504 3292
rect 44528 3290 44584 3292
rect 44288 3238 44334 3290
rect 44334 3238 44344 3290
rect 44368 3238 44398 3290
rect 44398 3238 44410 3290
rect 44410 3238 44424 3290
rect 44448 3238 44462 3290
rect 44462 3238 44474 3290
rect 44474 3238 44504 3290
rect 44528 3238 44538 3290
rect 44538 3238 44584 3290
rect 44288 3236 44344 3238
rect 44368 3236 44424 3238
rect 44448 3236 44504 3238
rect 44528 3236 44584 3238
rect 44288 2202 44344 2204
rect 44368 2202 44424 2204
rect 44448 2202 44504 2204
rect 44528 2202 44584 2204
rect 44288 2150 44334 2202
rect 44334 2150 44344 2202
rect 44368 2150 44398 2202
rect 44398 2150 44410 2202
rect 44410 2150 44424 2202
rect 44448 2150 44462 2202
rect 44462 2150 44474 2202
rect 44474 2150 44504 2202
rect 44528 2150 44538 2202
rect 44538 2150 44584 2202
rect 44288 2148 44344 2150
rect 44368 2148 44424 2150
rect 44448 2148 44504 2150
rect 44528 2148 44584 2150
rect 46754 3576 46810 3632
rect 46478 3440 46534 3496
rect 46386 3052 46442 3088
rect 47582 3984 47638 4040
rect 46386 3032 46388 3052
rect 46388 3032 46440 3052
rect 46440 3032 46442 3052
rect 51510 20154 51566 20156
rect 51590 20154 51646 20156
rect 51670 20154 51726 20156
rect 51750 20154 51806 20156
rect 51510 20102 51556 20154
rect 51556 20102 51566 20154
rect 51590 20102 51620 20154
rect 51620 20102 51632 20154
rect 51632 20102 51646 20154
rect 51670 20102 51684 20154
rect 51684 20102 51696 20154
rect 51696 20102 51726 20154
rect 51750 20102 51760 20154
rect 51760 20102 51806 20154
rect 51510 20100 51566 20102
rect 51590 20100 51646 20102
rect 51670 20100 51726 20102
rect 51750 20100 51806 20102
rect 52274 21664 52330 21720
rect 51510 19066 51566 19068
rect 51590 19066 51646 19068
rect 51670 19066 51726 19068
rect 51750 19066 51806 19068
rect 51510 19014 51556 19066
rect 51556 19014 51566 19066
rect 51590 19014 51620 19066
rect 51620 19014 51632 19066
rect 51632 19014 51646 19066
rect 51670 19014 51684 19066
rect 51684 19014 51696 19066
rect 51696 19014 51726 19066
rect 51750 19014 51760 19066
rect 51760 19014 51806 19066
rect 51510 19012 51566 19014
rect 51590 19012 51646 19014
rect 51670 19012 51726 19014
rect 51750 19012 51806 19014
rect 51510 17978 51566 17980
rect 51590 17978 51646 17980
rect 51670 17978 51726 17980
rect 51750 17978 51806 17980
rect 51510 17926 51556 17978
rect 51556 17926 51566 17978
rect 51590 17926 51620 17978
rect 51620 17926 51632 17978
rect 51632 17926 51646 17978
rect 51670 17926 51684 17978
rect 51684 17926 51696 17978
rect 51696 17926 51726 17978
rect 51750 17926 51760 17978
rect 51760 17926 51806 17978
rect 51510 17924 51566 17926
rect 51590 17924 51646 17926
rect 51670 17924 51726 17926
rect 51750 17924 51806 17926
rect 51510 16890 51566 16892
rect 51590 16890 51646 16892
rect 51670 16890 51726 16892
rect 51750 16890 51806 16892
rect 51510 16838 51556 16890
rect 51556 16838 51566 16890
rect 51590 16838 51620 16890
rect 51620 16838 51632 16890
rect 51632 16838 51646 16890
rect 51670 16838 51684 16890
rect 51684 16838 51696 16890
rect 51696 16838 51726 16890
rect 51750 16838 51760 16890
rect 51760 16838 51806 16890
rect 51510 16836 51566 16838
rect 51590 16836 51646 16838
rect 51670 16836 51726 16838
rect 51750 16836 51806 16838
rect 51510 15802 51566 15804
rect 51590 15802 51646 15804
rect 51670 15802 51726 15804
rect 51750 15802 51806 15804
rect 51510 15750 51556 15802
rect 51556 15750 51566 15802
rect 51590 15750 51620 15802
rect 51620 15750 51632 15802
rect 51632 15750 51646 15802
rect 51670 15750 51684 15802
rect 51684 15750 51696 15802
rect 51696 15750 51726 15802
rect 51750 15750 51760 15802
rect 51760 15750 51806 15802
rect 51510 15748 51566 15750
rect 51590 15748 51646 15750
rect 51670 15748 51726 15750
rect 51750 15748 51806 15750
rect 48226 5616 48282 5672
rect 49514 7268 49570 7304
rect 49514 7248 49516 7268
rect 49516 7248 49568 7268
rect 49568 7248 49570 7268
rect 49146 6568 49202 6624
rect 49330 3848 49386 3904
rect 48134 3712 48190 3768
rect 48042 3068 48044 3088
rect 48044 3068 48096 3088
rect 48096 3068 48098 3088
rect 48042 3032 48098 3068
rect 51510 14714 51566 14716
rect 51590 14714 51646 14716
rect 51670 14714 51726 14716
rect 51750 14714 51806 14716
rect 51510 14662 51556 14714
rect 51556 14662 51566 14714
rect 51590 14662 51620 14714
rect 51620 14662 51632 14714
rect 51632 14662 51646 14714
rect 51670 14662 51684 14714
rect 51684 14662 51696 14714
rect 51696 14662 51726 14714
rect 51750 14662 51760 14714
rect 51760 14662 51806 14714
rect 51510 14660 51566 14662
rect 51590 14660 51646 14662
rect 51670 14660 51726 14662
rect 51750 14660 51806 14662
rect 51510 13626 51566 13628
rect 51590 13626 51646 13628
rect 51670 13626 51726 13628
rect 51750 13626 51806 13628
rect 51510 13574 51556 13626
rect 51556 13574 51566 13626
rect 51590 13574 51620 13626
rect 51620 13574 51632 13626
rect 51632 13574 51646 13626
rect 51670 13574 51684 13626
rect 51684 13574 51696 13626
rect 51696 13574 51726 13626
rect 51750 13574 51760 13626
rect 51760 13574 51806 13626
rect 51510 13572 51566 13574
rect 51590 13572 51646 13574
rect 51670 13572 51726 13574
rect 51750 13572 51806 13574
rect 56690 21664 56746 21720
rect 55862 21528 55918 21584
rect 53194 20868 53250 20904
rect 53194 20848 53196 20868
rect 53196 20848 53248 20868
rect 53248 20848 53250 20868
rect 51510 12538 51566 12540
rect 51590 12538 51646 12540
rect 51670 12538 51726 12540
rect 51750 12538 51806 12540
rect 51510 12486 51556 12538
rect 51556 12486 51566 12538
rect 51590 12486 51620 12538
rect 51620 12486 51632 12538
rect 51632 12486 51646 12538
rect 51670 12486 51684 12538
rect 51684 12486 51696 12538
rect 51696 12486 51726 12538
rect 51750 12486 51760 12538
rect 51760 12486 51806 12538
rect 51510 12484 51566 12486
rect 51590 12484 51646 12486
rect 51670 12484 51726 12486
rect 51750 12484 51806 12486
rect 51510 11450 51566 11452
rect 51590 11450 51646 11452
rect 51670 11450 51726 11452
rect 51750 11450 51806 11452
rect 51510 11398 51556 11450
rect 51556 11398 51566 11450
rect 51590 11398 51620 11450
rect 51620 11398 51632 11450
rect 51632 11398 51646 11450
rect 51670 11398 51684 11450
rect 51684 11398 51696 11450
rect 51696 11398 51726 11450
rect 51750 11398 51760 11450
rect 51760 11398 51806 11450
rect 51510 11396 51566 11398
rect 51590 11396 51646 11398
rect 51670 11396 51726 11398
rect 51750 11396 51806 11398
rect 51510 10362 51566 10364
rect 51590 10362 51646 10364
rect 51670 10362 51726 10364
rect 51750 10362 51806 10364
rect 51510 10310 51556 10362
rect 51556 10310 51566 10362
rect 51590 10310 51620 10362
rect 51620 10310 51632 10362
rect 51632 10310 51646 10362
rect 51670 10310 51684 10362
rect 51684 10310 51696 10362
rect 51696 10310 51726 10362
rect 51750 10310 51760 10362
rect 51760 10310 51806 10362
rect 51510 10308 51566 10310
rect 51590 10308 51646 10310
rect 51670 10308 51726 10310
rect 51750 10308 51806 10310
rect 51510 9274 51566 9276
rect 51590 9274 51646 9276
rect 51670 9274 51726 9276
rect 51750 9274 51806 9276
rect 51510 9222 51556 9274
rect 51556 9222 51566 9274
rect 51590 9222 51620 9274
rect 51620 9222 51632 9274
rect 51632 9222 51646 9274
rect 51670 9222 51684 9274
rect 51684 9222 51696 9274
rect 51696 9222 51726 9274
rect 51750 9222 51760 9274
rect 51760 9222 51806 9274
rect 51510 9220 51566 9222
rect 51590 9220 51646 9222
rect 51670 9220 51726 9222
rect 51750 9220 51806 9222
rect 51510 8186 51566 8188
rect 51590 8186 51646 8188
rect 51670 8186 51726 8188
rect 51750 8186 51806 8188
rect 51510 8134 51556 8186
rect 51556 8134 51566 8186
rect 51590 8134 51620 8186
rect 51620 8134 51632 8186
rect 51632 8134 51646 8186
rect 51670 8134 51684 8186
rect 51684 8134 51696 8186
rect 51696 8134 51726 8186
rect 51750 8134 51760 8186
rect 51760 8134 51806 8186
rect 51510 8132 51566 8134
rect 51590 8132 51646 8134
rect 51670 8132 51726 8134
rect 51750 8132 51806 8134
rect 51510 7098 51566 7100
rect 51590 7098 51646 7100
rect 51670 7098 51726 7100
rect 51750 7098 51806 7100
rect 51510 7046 51556 7098
rect 51556 7046 51566 7098
rect 51590 7046 51620 7098
rect 51620 7046 51632 7098
rect 51632 7046 51646 7098
rect 51670 7046 51684 7098
rect 51684 7046 51696 7098
rect 51696 7046 51726 7098
rect 51750 7046 51760 7098
rect 51760 7046 51806 7098
rect 51510 7044 51566 7046
rect 51590 7044 51646 7046
rect 51670 7044 51726 7046
rect 51750 7044 51806 7046
rect 51510 6010 51566 6012
rect 51590 6010 51646 6012
rect 51670 6010 51726 6012
rect 51750 6010 51806 6012
rect 51510 5958 51556 6010
rect 51556 5958 51566 6010
rect 51590 5958 51620 6010
rect 51620 5958 51632 6010
rect 51632 5958 51646 6010
rect 51670 5958 51684 6010
rect 51684 5958 51696 6010
rect 51696 5958 51726 6010
rect 51750 5958 51760 6010
rect 51760 5958 51806 6010
rect 51510 5956 51566 5958
rect 51590 5956 51646 5958
rect 51670 5956 51726 5958
rect 51750 5956 51806 5958
rect 51510 4922 51566 4924
rect 51590 4922 51646 4924
rect 51670 4922 51726 4924
rect 51750 4922 51806 4924
rect 51510 4870 51556 4922
rect 51556 4870 51566 4922
rect 51590 4870 51620 4922
rect 51620 4870 51632 4922
rect 51632 4870 51646 4922
rect 51670 4870 51684 4922
rect 51684 4870 51696 4922
rect 51696 4870 51726 4922
rect 51750 4870 51760 4922
rect 51760 4870 51806 4922
rect 51510 4868 51566 4870
rect 51590 4868 51646 4870
rect 51670 4868 51726 4870
rect 51750 4868 51806 4870
rect 51262 3984 51318 4040
rect 51078 3848 51134 3904
rect 50710 3732 50766 3768
rect 50710 3712 50712 3732
rect 50712 3712 50764 3732
rect 50764 3712 50766 3732
rect 51510 3834 51566 3836
rect 51590 3834 51646 3836
rect 51670 3834 51726 3836
rect 51750 3834 51806 3836
rect 51510 3782 51556 3834
rect 51556 3782 51566 3834
rect 51590 3782 51620 3834
rect 51620 3782 51632 3834
rect 51632 3782 51646 3834
rect 51670 3782 51684 3834
rect 51684 3782 51696 3834
rect 51696 3782 51726 3834
rect 51750 3782 51760 3834
rect 51760 3782 51806 3834
rect 51510 3780 51566 3782
rect 51590 3780 51646 3782
rect 51670 3780 51726 3782
rect 51750 3780 51806 3782
rect 52090 3576 52146 3632
rect 51998 3440 52054 3496
rect 52550 3884 52552 3904
rect 52552 3884 52604 3904
rect 52604 3884 52606 3904
rect 52550 3848 52606 3884
rect 51510 2746 51566 2748
rect 51590 2746 51646 2748
rect 51670 2746 51726 2748
rect 51750 2746 51806 2748
rect 51510 2694 51556 2746
rect 51556 2694 51566 2746
rect 51590 2694 51620 2746
rect 51620 2694 51632 2746
rect 51632 2694 51646 2746
rect 51670 2694 51684 2746
rect 51684 2694 51696 2746
rect 51696 2694 51726 2746
rect 51750 2694 51760 2746
rect 51760 2694 51806 2746
rect 51510 2692 51566 2694
rect 51590 2692 51646 2694
rect 51670 2692 51726 2694
rect 51750 2692 51806 2694
rect 58732 21786 58788 21788
rect 58812 21786 58868 21788
rect 58892 21786 58948 21788
rect 58972 21786 59028 21788
rect 58732 21734 58778 21786
rect 58778 21734 58788 21786
rect 58812 21734 58842 21786
rect 58842 21734 58854 21786
rect 58854 21734 58868 21786
rect 58892 21734 58906 21786
rect 58906 21734 58918 21786
rect 58918 21734 58948 21786
rect 58972 21734 58982 21786
rect 58982 21734 59028 21786
rect 58732 21732 58788 21734
rect 58812 21732 58868 21734
rect 58892 21732 58948 21734
rect 58972 21732 59028 21734
rect 55494 17604 55550 17640
rect 55494 17584 55496 17604
rect 55496 17584 55548 17604
rect 55548 17584 55550 17604
rect 55310 11756 55366 11792
rect 55310 11736 55312 11756
rect 55312 11736 55364 11756
rect 55364 11736 55366 11756
rect 55586 11600 55642 11656
rect 53654 3984 53710 4040
rect 54942 7248 54998 7304
rect 53378 2760 53434 2816
rect 55126 5652 55128 5672
rect 55128 5652 55180 5672
rect 55180 5652 55182 5672
rect 55126 5616 55182 5652
rect 55310 4256 55366 4312
rect 56138 11620 56194 11656
rect 56138 11600 56140 11620
rect 56140 11600 56192 11620
rect 56192 11600 56194 11620
rect 55402 3984 55458 4040
rect 55126 2896 55182 2952
rect 58732 20698 58788 20700
rect 58812 20698 58868 20700
rect 58892 20698 58948 20700
rect 58972 20698 59028 20700
rect 58732 20646 58778 20698
rect 58778 20646 58788 20698
rect 58812 20646 58842 20698
rect 58842 20646 58854 20698
rect 58854 20646 58868 20698
rect 58892 20646 58906 20698
rect 58906 20646 58918 20698
rect 58918 20646 58948 20698
rect 58972 20646 58982 20698
rect 58982 20646 59028 20698
rect 58732 20644 58788 20646
rect 58812 20644 58868 20646
rect 58892 20644 58948 20646
rect 58972 20644 59028 20646
rect 58732 19610 58788 19612
rect 58812 19610 58868 19612
rect 58892 19610 58948 19612
rect 58972 19610 59028 19612
rect 58732 19558 58778 19610
rect 58778 19558 58788 19610
rect 58812 19558 58842 19610
rect 58842 19558 58854 19610
rect 58854 19558 58868 19610
rect 58892 19558 58906 19610
rect 58906 19558 58918 19610
rect 58918 19558 58948 19610
rect 58972 19558 58982 19610
rect 58982 19558 59028 19610
rect 58732 19556 58788 19558
rect 58812 19556 58868 19558
rect 58892 19556 58948 19558
rect 58972 19556 59028 19558
rect 58732 18522 58788 18524
rect 58812 18522 58868 18524
rect 58892 18522 58948 18524
rect 58972 18522 59028 18524
rect 58732 18470 58778 18522
rect 58778 18470 58788 18522
rect 58812 18470 58842 18522
rect 58842 18470 58854 18522
rect 58854 18470 58868 18522
rect 58892 18470 58906 18522
rect 58906 18470 58918 18522
rect 58918 18470 58948 18522
rect 58972 18470 58982 18522
rect 58982 18470 59028 18522
rect 58732 18468 58788 18470
rect 58812 18468 58868 18470
rect 58892 18468 58948 18470
rect 58972 18468 59028 18470
rect 58732 17434 58788 17436
rect 58812 17434 58868 17436
rect 58892 17434 58948 17436
rect 58972 17434 59028 17436
rect 58732 17382 58778 17434
rect 58778 17382 58788 17434
rect 58812 17382 58842 17434
rect 58842 17382 58854 17434
rect 58854 17382 58868 17434
rect 58892 17382 58906 17434
rect 58906 17382 58918 17434
rect 58918 17382 58948 17434
rect 58972 17382 58982 17434
rect 58982 17382 59028 17434
rect 58732 17380 58788 17382
rect 58812 17380 58868 17382
rect 58892 17380 58948 17382
rect 58972 17380 59028 17382
rect 56782 11756 56838 11792
rect 56782 11736 56784 11756
rect 56784 11736 56836 11756
rect 56836 11736 56838 11756
rect 56874 11056 56930 11112
rect 58732 16346 58788 16348
rect 58812 16346 58868 16348
rect 58892 16346 58948 16348
rect 58972 16346 59028 16348
rect 58732 16294 58778 16346
rect 58778 16294 58788 16346
rect 58812 16294 58842 16346
rect 58842 16294 58854 16346
rect 58854 16294 58868 16346
rect 58892 16294 58906 16346
rect 58906 16294 58918 16346
rect 58918 16294 58948 16346
rect 58972 16294 58982 16346
rect 58982 16294 59028 16346
rect 58732 16292 58788 16294
rect 58812 16292 58868 16294
rect 58892 16292 58948 16294
rect 58972 16292 59028 16294
rect 58732 15258 58788 15260
rect 58812 15258 58868 15260
rect 58892 15258 58948 15260
rect 58972 15258 59028 15260
rect 58732 15206 58778 15258
rect 58778 15206 58788 15258
rect 58812 15206 58842 15258
rect 58842 15206 58854 15258
rect 58854 15206 58868 15258
rect 58892 15206 58906 15258
rect 58906 15206 58918 15258
rect 58918 15206 58948 15258
rect 58972 15206 58982 15258
rect 58982 15206 59028 15258
rect 58732 15204 58788 15206
rect 58812 15204 58868 15206
rect 58892 15204 58948 15206
rect 58972 15204 59028 15206
rect 58732 14170 58788 14172
rect 58812 14170 58868 14172
rect 58892 14170 58948 14172
rect 58972 14170 59028 14172
rect 58732 14118 58778 14170
rect 58778 14118 58788 14170
rect 58812 14118 58842 14170
rect 58842 14118 58854 14170
rect 58854 14118 58868 14170
rect 58892 14118 58906 14170
rect 58906 14118 58918 14170
rect 58918 14118 58948 14170
rect 58972 14118 58982 14170
rect 58982 14118 59028 14170
rect 58732 14116 58788 14118
rect 58812 14116 58868 14118
rect 58892 14116 58948 14118
rect 58972 14116 59028 14118
rect 58732 13082 58788 13084
rect 58812 13082 58868 13084
rect 58892 13082 58948 13084
rect 58972 13082 59028 13084
rect 58732 13030 58778 13082
rect 58778 13030 58788 13082
rect 58812 13030 58842 13082
rect 58842 13030 58854 13082
rect 58854 13030 58868 13082
rect 58892 13030 58906 13082
rect 58906 13030 58918 13082
rect 58918 13030 58948 13082
rect 58972 13030 58982 13082
rect 58982 13030 59028 13082
rect 58732 13028 58788 13030
rect 58812 13028 58868 13030
rect 58892 13028 58948 13030
rect 58972 13028 59028 13030
rect 56414 5072 56470 5128
rect 56598 3984 56654 4040
rect 57242 6568 57298 6624
rect 56966 5208 57022 5264
rect 57150 4020 57152 4040
rect 57152 4020 57204 4040
rect 57204 4020 57206 4040
rect 57150 3984 57206 4020
rect 58732 11994 58788 11996
rect 58812 11994 58868 11996
rect 58892 11994 58948 11996
rect 58972 11994 59028 11996
rect 58732 11942 58778 11994
rect 58778 11942 58788 11994
rect 58812 11942 58842 11994
rect 58842 11942 58854 11994
rect 58854 11942 58868 11994
rect 58892 11942 58906 11994
rect 58906 11942 58918 11994
rect 58918 11942 58948 11994
rect 58972 11942 58982 11994
rect 58982 11942 59028 11994
rect 58732 11940 58788 11942
rect 58812 11940 58868 11942
rect 58892 11940 58948 11942
rect 58972 11940 59028 11942
rect 58732 10906 58788 10908
rect 58812 10906 58868 10908
rect 58892 10906 58948 10908
rect 58972 10906 59028 10908
rect 58732 10854 58778 10906
rect 58778 10854 58788 10906
rect 58812 10854 58842 10906
rect 58842 10854 58854 10906
rect 58854 10854 58868 10906
rect 58892 10854 58906 10906
rect 58906 10854 58918 10906
rect 58918 10854 58948 10906
rect 58972 10854 58982 10906
rect 58982 10854 59028 10906
rect 58732 10852 58788 10854
rect 58812 10852 58868 10854
rect 58892 10852 58948 10854
rect 58972 10852 59028 10854
rect 58732 9818 58788 9820
rect 58812 9818 58868 9820
rect 58892 9818 58948 9820
rect 58972 9818 59028 9820
rect 58732 9766 58778 9818
rect 58778 9766 58788 9818
rect 58812 9766 58842 9818
rect 58842 9766 58854 9818
rect 58854 9766 58868 9818
rect 58892 9766 58906 9818
rect 58906 9766 58918 9818
rect 58918 9766 58948 9818
rect 58972 9766 58982 9818
rect 58982 9766 59028 9818
rect 58732 9764 58788 9766
rect 58812 9764 58868 9766
rect 58892 9764 58948 9766
rect 58972 9764 59028 9766
rect 58732 8730 58788 8732
rect 58812 8730 58868 8732
rect 58892 8730 58948 8732
rect 58972 8730 59028 8732
rect 58732 8678 58778 8730
rect 58778 8678 58788 8730
rect 58812 8678 58842 8730
rect 58842 8678 58854 8730
rect 58854 8678 58868 8730
rect 58892 8678 58906 8730
rect 58906 8678 58918 8730
rect 58918 8678 58948 8730
rect 58972 8678 58982 8730
rect 58982 8678 59028 8730
rect 58732 8676 58788 8678
rect 58812 8676 58868 8678
rect 58892 8676 58948 8678
rect 58972 8676 59028 8678
rect 58732 7642 58788 7644
rect 58812 7642 58868 7644
rect 58892 7642 58948 7644
rect 58972 7642 59028 7644
rect 58732 7590 58778 7642
rect 58778 7590 58788 7642
rect 58812 7590 58842 7642
rect 58842 7590 58854 7642
rect 58854 7590 58868 7642
rect 58892 7590 58906 7642
rect 58906 7590 58918 7642
rect 58918 7590 58948 7642
rect 58972 7590 58982 7642
rect 58982 7590 59028 7642
rect 58732 7588 58788 7590
rect 58812 7588 58868 7590
rect 58892 7588 58948 7590
rect 58972 7588 59028 7590
rect 57978 5616 58034 5672
rect 57886 4256 57942 4312
rect 58732 6554 58788 6556
rect 58812 6554 58868 6556
rect 58892 6554 58948 6556
rect 58972 6554 59028 6556
rect 58732 6502 58778 6554
rect 58778 6502 58788 6554
rect 58812 6502 58842 6554
rect 58842 6502 58854 6554
rect 58854 6502 58868 6554
rect 58892 6502 58906 6554
rect 58906 6502 58918 6554
rect 58918 6502 58948 6554
rect 58972 6502 58982 6554
rect 58982 6502 59028 6554
rect 58732 6500 58788 6502
rect 58812 6500 58868 6502
rect 58892 6500 58948 6502
rect 58972 6500 59028 6502
rect 58732 5466 58788 5468
rect 58812 5466 58868 5468
rect 58892 5466 58948 5468
rect 58972 5466 59028 5468
rect 58732 5414 58778 5466
rect 58778 5414 58788 5466
rect 58812 5414 58842 5466
rect 58842 5414 58854 5466
rect 58854 5414 58868 5466
rect 58892 5414 58906 5466
rect 58906 5414 58918 5466
rect 58918 5414 58948 5466
rect 58972 5414 58982 5466
rect 58982 5414 59028 5466
rect 58732 5412 58788 5414
rect 58812 5412 58868 5414
rect 58892 5412 58948 5414
rect 58972 5412 59028 5414
rect 58438 3848 58494 3904
rect 58346 3440 58402 3496
rect 57886 2760 57942 2816
rect 58732 4378 58788 4380
rect 58812 4378 58868 4380
rect 58892 4378 58948 4380
rect 58972 4378 59028 4380
rect 58732 4326 58778 4378
rect 58778 4326 58788 4378
rect 58812 4326 58842 4378
rect 58842 4326 58854 4378
rect 58854 4326 58868 4378
rect 58892 4326 58906 4378
rect 58906 4326 58918 4378
rect 58918 4326 58948 4378
rect 58972 4326 58982 4378
rect 58982 4326 59028 4378
rect 58732 4324 58788 4326
rect 58812 4324 58868 4326
rect 58892 4324 58948 4326
rect 58972 4324 59028 4326
rect 58732 3290 58788 3292
rect 58812 3290 58868 3292
rect 58892 3290 58948 3292
rect 58972 3290 59028 3292
rect 58732 3238 58778 3290
rect 58778 3238 58788 3290
rect 58812 3238 58842 3290
rect 58842 3238 58854 3290
rect 58854 3238 58868 3290
rect 58892 3238 58906 3290
rect 58906 3238 58918 3290
rect 58918 3238 58948 3290
rect 58972 3238 58982 3290
rect 58982 3238 59028 3290
rect 58732 3236 58788 3238
rect 58812 3236 58868 3238
rect 58892 3236 58948 3238
rect 58972 3236 59028 3238
rect 58732 2202 58788 2204
rect 58812 2202 58868 2204
rect 58892 2202 58948 2204
rect 58972 2202 59028 2204
rect 58732 2150 58778 2202
rect 58778 2150 58788 2202
rect 58812 2150 58842 2202
rect 58842 2150 58854 2202
rect 58854 2150 58868 2202
rect 58892 2150 58906 2202
rect 58906 2150 58918 2202
rect 58918 2150 58948 2202
rect 58972 2150 58982 2202
rect 58982 2150 59028 2202
rect 58732 2148 58788 2150
rect 58812 2148 58868 2150
rect 58892 2148 58948 2150
rect 58972 2148 59028 2150
<< metal3 >>
rect 8168 27776 8484 27777
rect 8168 27712 8174 27776
rect 8238 27712 8254 27776
rect 8318 27712 8334 27776
rect 8398 27712 8414 27776
rect 8478 27712 8484 27776
rect 8168 27711 8484 27712
rect 22612 27776 22928 27777
rect 22612 27712 22618 27776
rect 22682 27712 22698 27776
rect 22762 27712 22778 27776
rect 22842 27712 22858 27776
rect 22922 27712 22928 27776
rect 22612 27711 22928 27712
rect 37056 27776 37372 27777
rect 37056 27712 37062 27776
rect 37126 27712 37142 27776
rect 37206 27712 37222 27776
rect 37286 27712 37302 27776
rect 37366 27712 37372 27776
rect 37056 27711 37372 27712
rect 51500 27776 51816 27777
rect 51500 27712 51506 27776
rect 51570 27712 51586 27776
rect 51650 27712 51666 27776
rect 51730 27712 51746 27776
rect 51810 27712 51816 27776
rect 51500 27711 51816 27712
rect 15390 27232 15706 27233
rect 15390 27168 15396 27232
rect 15460 27168 15476 27232
rect 15540 27168 15556 27232
rect 15620 27168 15636 27232
rect 15700 27168 15706 27232
rect 15390 27167 15706 27168
rect 29834 27232 30150 27233
rect 29834 27168 29840 27232
rect 29904 27168 29920 27232
rect 29984 27168 30000 27232
rect 30064 27168 30080 27232
rect 30144 27168 30150 27232
rect 29834 27167 30150 27168
rect 44278 27232 44594 27233
rect 44278 27168 44284 27232
rect 44348 27168 44364 27232
rect 44428 27168 44444 27232
rect 44508 27168 44524 27232
rect 44588 27168 44594 27232
rect 44278 27167 44594 27168
rect 58722 27232 59038 27233
rect 58722 27168 58728 27232
rect 58792 27168 58808 27232
rect 58872 27168 58888 27232
rect 58952 27168 58968 27232
rect 59032 27168 59038 27232
rect 58722 27167 59038 27168
rect 8168 26688 8484 26689
rect 8168 26624 8174 26688
rect 8238 26624 8254 26688
rect 8318 26624 8334 26688
rect 8398 26624 8414 26688
rect 8478 26624 8484 26688
rect 8168 26623 8484 26624
rect 22612 26688 22928 26689
rect 22612 26624 22618 26688
rect 22682 26624 22698 26688
rect 22762 26624 22778 26688
rect 22842 26624 22858 26688
rect 22922 26624 22928 26688
rect 22612 26623 22928 26624
rect 37056 26688 37372 26689
rect 37056 26624 37062 26688
rect 37126 26624 37142 26688
rect 37206 26624 37222 26688
rect 37286 26624 37302 26688
rect 37366 26624 37372 26688
rect 37056 26623 37372 26624
rect 51500 26688 51816 26689
rect 51500 26624 51506 26688
rect 51570 26624 51586 26688
rect 51650 26624 51666 26688
rect 51730 26624 51746 26688
rect 51810 26624 51816 26688
rect 51500 26623 51816 26624
rect 15390 26144 15706 26145
rect 15390 26080 15396 26144
rect 15460 26080 15476 26144
rect 15540 26080 15556 26144
rect 15620 26080 15636 26144
rect 15700 26080 15706 26144
rect 15390 26079 15706 26080
rect 29834 26144 30150 26145
rect 29834 26080 29840 26144
rect 29904 26080 29920 26144
rect 29984 26080 30000 26144
rect 30064 26080 30080 26144
rect 30144 26080 30150 26144
rect 29834 26079 30150 26080
rect 44278 26144 44594 26145
rect 44278 26080 44284 26144
rect 44348 26080 44364 26144
rect 44428 26080 44444 26144
rect 44508 26080 44524 26144
rect 44588 26080 44594 26144
rect 44278 26079 44594 26080
rect 58722 26144 59038 26145
rect 58722 26080 58728 26144
rect 58792 26080 58808 26144
rect 58872 26080 58888 26144
rect 58952 26080 58968 26144
rect 59032 26080 59038 26144
rect 58722 26079 59038 26080
rect 8168 25600 8484 25601
rect 8168 25536 8174 25600
rect 8238 25536 8254 25600
rect 8318 25536 8334 25600
rect 8398 25536 8414 25600
rect 8478 25536 8484 25600
rect 8168 25535 8484 25536
rect 22612 25600 22928 25601
rect 22612 25536 22618 25600
rect 22682 25536 22698 25600
rect 22762 25536 22778 25600
rect 22842 25536 22858 25600
rect 22922 25536 22928 25600
rect 22612 25535 22928 25536
rect 37056 25600 37372 25601
rect 37056 25536 37062 25600
rect 37126 25536 37142 25600
rect 37206 25536 37222 25600
rect 37286 25536 37302 25600
rect 37366 25536 37372 25600
rect 37056 25535 37372 25536
rect 51500 25600 51816 25601
rect 51500 25536 51506 25600
rect 51570 25536 51586 25600
rect 51650 25536 51666 25600
rect 51730 25536 51746 25600
rect 51810 25536 51816 25600
rect 51500 25535 51816 25536
rect 15390 25056 15706 25057
rect 15390 24992 15396 25056
rect 15460 24992 15476 25056
rect 15540 24992 15556 25056
rect 15620 24992 15636 25056
rect 15700 24992 15706 25056
rect 15390 24991 15706 24992
rect 29834 25056 30150 25057
rect 29834 24992 29840 25056
rect 29904 24992 29920 25056
rect 29984 24992 30000 25056
rect 30064 24992 30080 25056
rect 30144 24992 30150 25056
rect 29834 24991 30150 24992
rect 44278 25056 44594 25057
rect 44278 24992 44284 25056
rect 44348 24992 44364 25056
rect 44428 24992 44444 25056
rect 44508 24992 44524 25056
rect 44588 24992 44594 25056
rect 44278 24991 44594 24992
rect 58722 25056 59038 25057
rect 58722 24992 58728 25056
rect 58792 24992 58808 25056
rect 58872 24992 58888 25056
rect 58952 24992 58968 25056
rect 59032 24992 59038 25056
rect 58722 24991 59038 24992
rect 8168 24512 8484 24513
rect 8168 24448 8174 24512
rect 8238 24448 8254 24512
rect 8318 24448 8334 24512
rect 8398 24448 8414 24512
rect 8478 24448 8484 24512
rect 8168 24447 8484 24448
rect 22612 24512 22928 24513
rect 22612 24448 22618 24512
rect 22682 24448 22698 24512
rect 22762 24448 22778 24512
rect 22842 24448 22858 24512
rect 22922 24448 22928 24512
rect 22612 24447 22928 24448
rect 37056 24512 37372 24513
rect 37056 24448 37062 24512
rect 37126 24448 37142 24512
rect 37206 24448 37222 24512
rect 37286 24448 37302 24512
rect 37366 24448 37372 24512
rect 37056 24447 37372 24448
rect 51500 24512 51816 24513
rect 51500 24448 51506 24512
rect 51570 24448 51586 24512
rect 51650 24448 51666 24512
rect 51730 24448 51746 24512
rect 51810 24448 51816 24512
rect 51500 24447 51816 24448
rect 15390 23968 15706 23969
rect 15390 23904 15396 23968
rect 15460 23904 15476 23968
rect 15540 23904 15556 23968
rect 15620 23904 15636 23968
rect 15700 23904 15706 23968
rect 15390 23903 15706 23904
rect 29834 23968 30150 23969
rect 29834 23904 29840 23968
rect 29904 23904 29920 23968
rect 29984 23904 30000 23968
rect 30064 23904 30080 23968
rect 30144 23904 30150 23968
rect 29834 23903 30150 23904
rect 44278 23968 44594 23969
rect 44278 23904 44284 23968
rect 44348 23904 44364 23968
rect 44428 23904 44444 23968
rect 44508 23904 44524 23968
rect 44588 23904 44594 23968
rect 44278 23903 44594 23904
rect 58722 23968 59038 23969
rect 58722 23904 58728 23968
rect 58792 23904 58808 23968
rect 58872 23904 58888 23968
rect 58952 23904 58968 23968
rect 59032 23904 59038 23968
rect 58722 23903 59038 23904
rect 8168 23424 8484 23425
rect 8168 23360 8174 23424
rect 8238 23360 8254 23424
rect 8318 23360 8334 23424
rect 8398 23360 8414 23424
rect 8478 23360 8484 23424
rect 8168 23359 8484 23360
rect 22612 23424 22928 23425
rect 22612 23360 22618 23424
rect 22682 23360 22698 23424
rect 22762 23360 22778 23424
rect 22842 23360 22858 23424
rect 22922 23360 22928 23424
rect 22612 23359 22928 23360
rect 37056 23424 37372 23425
rect 37056 23360 37062 23424
rect 37126 23360 37142 23424
rect 37206 23360 37222 23424
rect 37286 23360 37302 23424
rect 37366 23360 37372 23424
rect 37056 23359 37372 23360
rect 51500 23424 51816 23425
rect 51500 23360 51506 23424
rect 51570 23360 51586 23424
rect 51650 23360 51666 23424
rect 51730 23360 51746 23424
rect 51810 23360 51816 23424
rect 51500 23359 51816 23360
rect 15390 22880 15706 22881
rect 15390 22816 15396 22880
rect 15460 22816 15476 22880
rect 15540 22816 15556 22880
rect 15620 22816 15636 22880
rect 15700 22816 15706 22880
rect 15390 22815 15706 22816
rect 29834 22880 30150 22881
rect 29834 22816 29840 22880
rect 29904 22816 29920 22880
rect 29984 22816 30000 22880
rect 30064 22816 30080 22880
rect 30144 22816 30150 22880
rect 29834 22815 30150 22816
rect 44278 22880 44594 22881
rect 44278 22816 44284 22880
rect 44348 22816 44364 22880
rect 44428 22816 44444 22880
rect 44508 22816 44524 22880
rect 44588 22816 44594 22880
rect 44278 22815 44594 22816
rect 58722 22880 59038 22881
rect 58722 22816 58728 22880
rect 58792 22816 58808 22880
rect 58872 22816 58888 22880
rect 58952 22816 58968 22880
rect 59032 22816 59038 22880
rect 58722 22815 59038 22816
rect 8168 22336 8484 22337
rect 8168 22272 8174 22336
rect 8238 22272 8254 22336
rect 8318 22272 8334 22336
rect 8398 22272 8414 22336
rect 8478 22272 8484 22336
rect 8168 22271 8484 22272
rect 22612 22336 22928 22337
rect 22612 22272 22618 22336
rect 22682 22272 22698 22336
rect 22762 22272 22778 22336
rect 22842 22272 22858 22336
rect 22922 22272 22928 22336
rect 22612 22271 22928 22272
rect 37056 22336 37372 22337
rect 37056 22272 37062 22336
rect 37126 22272 37142 22336
rect 37206 22272 37222 22336
rect 37286 22272 37302 22336
rect 37366 22272 37372 22336
rect 37056 22271 37372 22272
rect 51500 22336 51816 22337
rect 51500 22272 51506 22336
rect 51570 22272 51586 22336
rect 51650 22272 51666 22336
rect 51730 22272 51746 22336
rect 51810 22272 51816 22336
rect 51500 22271 51816 22272
rect 15390 21792 15706 21793
rect 15390 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15706 21792
rect 15390 21727 15706 21728
rect 29834 21792 30150 21793
rect 29834 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30150 21792
rect 29834 21727 30150 21728
rect 44278 21792 44594 21793
rect 44278 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44594 21792
rect 44278 21727 44594 21728
rect 58722 21792 59038 21793
rect 58722 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59038 21792
rect 58722 21727 59038 21728
rect 52269 21722 52335 21725
rect 56685 21722 56751 21725
rect 52269 21720 56751 21722
rect 52269 21664 52274 21720
rect 52330 21664 56690 21720
rect 56746 21664 56751 21720
rect 52269 21662 56751 21664
rect 52269 21659 52335 21662
rect 56685 21659 56751 21662
rect 51349 21586 51415 21589
rect 55857 21586 55923 21589
rect 51349 21584 55923 21586
rect 51349 21528 51354 21584
rect 51410 21528 55862 21584
rect 55918 21528 55923 21584
rect 51349 21526 55923 21528
rect 51349 21523 51415 21526
rect 55857 21523 55923 21526
rect 8168 21248 8484 21249
rect 8168 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8484 21248
rect 8168 21183 8484 21184
rect 22612 21248 22928 21249
rect 22612 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22928 21248
rect 22612 21183 22928 21184
rect 37056 21248 37372 21249
rect 37056 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37372 21248
rect 37056 21183 37372 21184
rect 51500 21248 51816 21249
rect 51500 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51816 21248
rect 51500 21183 51816 21184
rect 24301 20906 24367 20909
rect 25497 20906 25563 20909
rect 24301 20904 25563 20906
rect 24301 20848 24306 20904
rect 24362 20848 25502 20904
rect 25558 20848 25563 20904
rect 24301 20846 25563 20848
rect 24301 20843 24367 20846
rect 25497 20843 25563 20846
rect 51993 20906 52059 20909
rect 53189 20906 53255 20909
rect 51993 20904 53255 20906
rect 51993 20848 51998 20904
rect 52054 20848 53194 20904
rect 53250 20848 53255 20904
rect 51993 20846 53255 20848
rect 51993 20843 52059 20846
rect 53189 20843 53255 20846
rect 15390 20704 15706 20705
rect 15390 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15706 20704
rect 15390 20639 15706 20640
rect 29834 20704 30150 20705
rect 29834 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30150 20704
rect 29834 20639 30150 20640
rect 44278 20704 44594 20705
rect 44278 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44594 20704
rect 44278 20639 44594 20640
rect 58722 20704 59038 20705
rect 58722 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59038 20704
rect 58722 20639 59038 20640
rect 43069 20498 43135 20501
rect 46473 20498 46539 20501
rect 43069 20496 46539 20498
rect 43069 20440 43074 20496
rect 43130 20440 46478 20496
rect 46534 20440 46539 20496
rect 43069 20438 46539 20440
rect 43069 20435 43135 20438
rect 46473 20435 46539 20438
rect 11513 20362 11579 20365
rect 18137 20362 18203 20365
rect 11513 20360 18203 20362
rect 11513 20304 11518 20360
rect 11574 20304 18142 20360
rect 18198 20304 18203 20360
rect 11513 20302 18203 20304
rect 11513 20299 11579 20302
rect 18137 20299 18203 20302
rect 24853 20362 24919 20365
rect 47853 20362 47919 20365
rect 24853 20360 47919 20362
rect 24853 20304 24858 20360
rect 24914 20304 47858 20360
rect 47914 20304 47919 20360
rect 24853 20302 47919 20304
rect 24853 20299 24919 20302
rect 47853 20299 47919 20302
rect 8168 20160 8484 20161
rect 8168 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8484 20160
rect 8168 20095 8484 20096
rect 22612 20160 22928 20161
rect 22612 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22928 20160
rect 22612 20095 22928 20096
rect 37056 20160 37372 20161
rect 37056 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37372 20160
rect 37056 20095 37372 20096
rect 51500 20160 51816 20161
rect 51500 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51816 20160
rect 51500 20095 51816 20096
rect 39205 19818 39271 19821
rect 45461 19818 45527 19821
rect 39205 19816 45527 19818
rect 39205 19760 39210 19816
rect 39266 19760 45466 19816
rect 45522 19760 45527 19816
rect 39205 19758 45527 19760
rect 39205 19755 39271 19758
rect 15390 19616 15706 19617
rect 15390 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15706 19616
rect 15390 19551 15706 19552
rect 29834 19616 30150 19617
rect 29834 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30150 19616
rect 29834 19551 30150 19552
rect 41370 19413 41430 19758
rect 45461 19755 45527 19758
rect 44278 19616 44594 19617
rect 44278 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44594 19616
rect 44278 19551 44594 19552
rect 58722 19616 59038 19617
rect 58722 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59038 19616
rect 58722 19551 59038 19552
rect 41321 19408 41430 19413
rect 41321 19352 41326 19408
rect 41382 19352 41430 19408
rect 41321 19350 41430 19352
rect 41321 19347 41387 19350
rect 8168 19072 8484 19073
rect 8168 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8484 19072
rect 8168 19007 8484 19008
rect 22612 19072 22928 19073
rect 22612 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22928 19072
rect 22612 19007 22928 19008
rect 37056 19072 37372 19073
rect 37056 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37372 19072
rect 37056 19007 37372 19008
rect 51500 19072 51816 19073
rect 51500 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51816 19072
rect 51500 19007 51816 19008
rect 15390 18528 15706 18529
rect 15390 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15706 18528
rect 15390 18463 15706 18464
rect 29834 18528 30150 18529
rect 29834 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30150 18528
rect 29834 18463 30150 18464
rect 44278 18528 44594 18529
rect 44278 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44594 18528
rect 44278 18463 44594 18464
rect 58722 18528 59038 18529
rect 58722 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59038 18528
rect 58722 18463 59038 18464
rect 8168 17984 8484 17985
rect 8168 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8484 17984
rect 8168 17919 8484 17920
rect 22612 17984 22928 17985
rect 22612 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22928 17984
rect 22612 17919 22928 17920
rect 37056 17984 37372 17985
rect 37056 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37372 17984
rect 37056 17919 37372 17920
rect 51500 17984 51816 17985
rect 51500 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51816 17984
rect 51500 17919 51816 17920
rect 12893 17778 12959 17781
rect 15929 17778 15995 17781
rect 12893 17776 15995 17778
rect 12893 17720 12898 17776
rect 12954 17720 15934 17776
rect 15990 17720 15995 17776
rect 12893 17718 15995 17720
rect 12893 17715 12959 17718
rect 15929 17715 15995 17718
rect 20529 17778 20595 17781
rect 26969 17778 27035 17781
rect 20529 17776 27035 17778
rect 20529 17720 20534 17776
rect 20590 17720 26974 17776
rect 27030 17720 27035 17776
rect 20529 17718 27035 17720
rect 20529 17715 20595 17718
rect 26969 17715 27035 17718
rect 49325 17642 49391 17645
rect 55489 17642 55555 17645
rect 49325 17640 55555 17642
rect 49325 17584 49330 17640
rect 49386 17584 55494 17640
rect 55550 17584 55555 17640
rect 49325 17582 55555 17584
rect 49325 17579 49391 17582
rect 55489 17579 55555 17582
rect 15390 17440 15706 17441
rect 15390 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15706 17440
rect 15390 17375 15706 17376
rect 29834 17440 30150 17441
rect 29834 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30150 17440
rect 29834 17375 30150 17376
rect 44278 17440 44594 17441
rect 44278 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44594 17440
rect 44278 17375 44594 17376
rect 58722 17440 59038 17441
rect 58722 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59038 17440
rect 58722 17375 59038 17376
rect 8168 16896 8484 16897
rect 8168 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8484 16896
rect 8168 16831 8484 16832
rect 22612 16896 22928 16897
rect 22612 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22928 16896
rect 22612 16831 22928 16832
rect 37056 16896 37372 16897
rect 37056 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37372 16896
rect 37056 16831 37372 16832
rect 51500 16896 51816 16897
rect 51500 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51816 16896
rect 51500 16831 51816 16832
rect 39941 16554 40007 16557
rect 41597 16554 41663 16557
rect 39941 16552 41663 16554
rect 39941 16496 39946 16552
rect 40002 16496 41602 16552
rect 41658 16496 41663 16552
rect 39941 16494 41663 16496
rect 39941 16491 40007 16494
rect 41597 16491 41663 16494
rect 15390 16352 15706 16353
rect 15390 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15706 16352
rect 15390 16287 15706 16288
rect 29834 16352 30150 16353
rect 29834 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30150 16352
rect 29834 16287 30150 16288
rect 44278 16352 44594 16353
rect 44278 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44594 16352
rect 44278 16287 44594 16288
rect 58722 16352 59038 16353
rect 58722 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59038 16352
rect 58722 16287 59038 16288
rect 8168 15808 8484 15809
rect 8168 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8484 15808
rect 8168 15743 8484 15744
rect 22612 15808 22928 15809
rect 22612 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22928 15808
rect 22612 15743 22928 15744
rect 37056 15808 37372 15809
rect 37056 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37372 15808
rect 37056 15743 37372 15744
rect 51500 15808 51816 15809
rect 51500 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51816 15808
rect 51500 15743 51816 15744
rect 15390 15264 15706 15265
rect 15390 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15706 15264
rect 15390 15199 15706 15200
rect 29834 15264 30150 15265
rect 29834 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30150 15264
rect 29834 15199 30150 15200
rect 44278 15264 44594 15265
rect 44278 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44594 15264
rect 44278 15199 44594 15200
rect 58722 15264 59038 15265
rect 58722 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59038 15264
rect 58722 15199 59038 15200
rect 8168 14720 8484 14721
rect 8168 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8484 14720
rect 8168 14655 8484 14656
rect 22612 14720 22928 14721
rect 22612 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22928 14720
rect 22612 14655 22928 14656
rect 37056 14720 37372 14721
rect 37056 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37372 14720
rect 37056 14655 37372 14656
rect 51500 14720 51816 14721
rect 51500 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51816 14720
rect 51500 14655 51816 14656
rect 15390 14176 15706 14177
rect 15390 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15706 14176
rect 15390 14111 15706 14112
rect 29834 14176 30150 14177
rect 29834 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30150 14176
rect 29834 14111 30150 14112
rect 44278 14176 44594 14177
rect 44278 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44594 14176
rect 44278 14111 44594 14112
rect 58722 14176 59038 14177
rect 58722 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59038 14176
rect 58722 14111 59038 14112
rect 8168 13632 8484 13633
rect 8168 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8484 13632
rect 8168 13567 8484 13568
rect 22612 13632 22928 13633
rect 22612 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22928 13632
rect 22612 13567 22928 13568
rect 37056 13632 37372 13633
rect 37056 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37372 13632
rect 37056 13567 37372 13568
rect 51500 13632 51816 13633
rect 51500 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51816 13632
rect 51500 13567 51816 13568
rect 15390 13088 15706 13089
rect 15390 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15706 13088
rect 15390 13023 15706 13024
rect 29834 13088 30150 13089
rect 29834 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30150 13088
rect 29834 13023 30150 13024
rect 44278 13088 44594 13089
rect 44278 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44594 13088
rect 44278 13023 44594 13024
rect 58722 13088 59038 13089
rect 58722 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59038 13088
rect 58722 13023 59038 13024
rect 8168 12544 8484 12545
rect 8168 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8484 12544
rect 8168 12479 8484 12480
rect 22612 12544 22928 12545
rect 22612 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22928 12544
rect 22612 12479 22928 12480
rect 37056 12544 37372 12545
rect 37056 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37372 12544
rect 37056 12479 37372 12480
rect 51500 12544 51816 12545
rect 51500 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51816 12544
rect 51500 12479 51816 12480
rect 15390 12000 15706 12001
rect 15390 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15706 12000
rect 15390 11935 15706 11936
rect 29834 12000 30150 12001
rect 29834 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30150 12000
rect 29834 11935 30150 11936
rect 44278 12000 44594 12001
rect 44278 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44594 12000
rect 44278 11935 44594 11936
rect 58722 12000 59038 12001
rect 58722 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59038 12000
rect 58722 11935 59038 11936
rect 55305 11794 55371 11797
rect 56777 11794 56843 11797
rect 55305 11792 56843 11794
rect 55305 11736 55310 11792
rect 55366 11736 56782 11792
rect 56838 11736 56843 11792
rect 55305 11734 56843 11736
rect 55305 11731 55371 11734
rect 56777 11731 56843 11734
rect 8385 11658 8451 11661
rect 9581 11658 9647 11661
rect 8385 11656 9647 11658
rect 8385 11600 8390 11656
rect 8446 11600 9586 11656
rect 9642 11600 9647 11656
rect 8385 11598 9647 11600
rect 8385 11595 8451 11598
rect 9581 11595 9647 11598
rect 55581 11658 55647 11661
rect 56133 11658 56199 11661
rect 55581 11656 56199 11658
rect 55581 11600 55586 11656
rect 55642 11600 56138 11656
rect 56194 11600 56199 11656
rect 55581 11598 56199 11600
rect 55581 11595 55647 11598
rect 56133 11595 56199 11598
rect 8168 11456 8484 11457
rect 8168 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8484 11456
rect 8168 11391 8484 11392
rect 22612 11456 22928 11457
rect 22612 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22928 11456
rect 22612 11391 22928 11392
rect 37056 11456 37372 11457
rect 37056 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37372 11456
rect 37056 11391 37372 11392
rect 51500 11456 51816 11457
rect 51500 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51816 11456
rect 51500 11391 51816 11392
rect 56869 11114 56935 11117
rect 57094 11114 57100 11116
rect 56869 11112 57100 11114
rect 56869 11056 56874 11112
rect 56930 11056 57100 11112
rect 56869 11054 57100 11056
rect 56869 11051 56935 11054
rect 57094 11052 57100 11054
rect 57164 11052 57170 11116
rect 15390 10912 15706 10913
rect 15390 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15706 10912
rect 15390 10847 15706 10848
rect 29834 10912 30150 10913
rect 29834 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30150 10912
rect 29834 10847 30150 10848
rect 44278 10912 44594 10913
rect 44278 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44594 10912
rect 44278 10847 44594 10848
rect 58722 10912 59038 10913
rect 58722 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59038 10912
rect 58722 10847 59038 10848
rect 9489 10706 9555 10709
rect 18413 10706 18479 10709
rect 9489 10704 18479 10706
rect 9489 10648 9494 10704
rect 9550 10648 18418 10704
rect 18474 10648 18479 10704
rect 9489 10646 18479 10648
rect 9489 10643 9555 10646
rect 18413 10643 18479 10646
rect 17677 10570 17743 10573
rect 19057 10570 19123 10573
rect 17677 10568 19123 10570
rect 17677 10512 17682 10568
rect 17738 10512 19062 10568
rect 19118 10512 19123 10568
rect 17677 10510 19123 10512
rect 17677 10507 17743 10510
rect 19057 10507 19123 10510
rect 8168 10368 8484 10369
rect 8168 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8484 10368
rect 8168 10303 8484 10304
rect 22612 10368 22928 10369
rect 22612 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22928 10368
rect 22612 10303 22928 10304
rect 37056 10368 37372 10369
rect 37056 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37372 10368
rect 37056 10303 37372 10304
rect 51500 10368 51816 10369
rect 51500 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51816 10368
rect 51500 10303 51816 10304
rect 17033 10298 17099 10301
rect 18597 10298 18663 10301
rect 17033 10296 18663 10298
rect 17033 10240 17038 10296
rect 17094 10240 18602 10296
rect 18658 10240 18663 10296
rect 17033 10238 18663 10240
rect 17033 10235 17099 10238
rect 18597 10235 18663 10238
rect 6821 10026 6887 10029
rect 29913 10026 29979 10029
rect 6821 10024 29979 10026
rect 6821 9968 6826 10024
rect 6882 9968 29918 10024
rect 29974 9968 29979 10024
rect 6821 9966 29979 9968
rect 6821 9963 6887 9966
rect 29913 9963 29979 9966
rect 15390 9824 15706 9825
rect 15390 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15706 9824
rect 15390 9759 15706 9760
rect 29834 9824 30150 9825
rect 29834 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30150 9824
rect 29834 9759 30150 9760
rect 44278 9824 44594 9825
rect 44278 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44594 9824
rect 44278 9759 44594 9760
rect 58722 9824 59038 9825
rect 58722 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59038 9824
rect 58722 9759 59038 9760
rect 9765 9618 9831 9621
rect 16021 9618 16087 9621
rect 9765 9616 16087 9618
rect 9765 9560 9770 9616
rect 9826 9560 16026 9616
rect 16082 9560 16087 9616
rect 9765 9558 16087 9560
rect 9765 9555 9831 9558
rect 16021 9555 16087 9558
rect 8168 9280 8484 9281
rect 8168 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8484 9280
rect 8168 9215 8484 9216
rect 22612 9280 22928 9281
rect 22612 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22928 9280
rect 22612 9215 22928 9216
rect 37056 9280 37372 9281
rect 37056 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37372 9280
rect 37056 9215 37372 9216
rect 51500 9280 51816 9281
rect 51500 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51816 9280
rect 51500 9215 51816 9216
rect 23289 8802 23355 8805
rect 28901 8802 28967 8805
rect 23289 8800 28967 8802
rect 23289 8744 23294 8800
rect 23350 8744 28906 8800
rect 28962 8744 28967 8800
rect 23289 8742 28967 8744
rect 23289 8739 23355 8742
rect 28901 8739 28967 8742
rect 15390 8736 15706 8737
rect 15390 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15706 8736
rect 15390 8671 15706 8672
rect 29834 8736 30150 8737
rect 29834 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30150 8736
rect 29834 8671 30150 8672
rect 44278 8736 44594 8737
rect 44278 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44594 8736
rect 44278 8671 44594 8672
rect 58722 8736 59038 8737
rect 58722 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59038 8736
rect 58722 8671 59038 8672
rect 8168 8192 8484 8193
rect 8168 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8484 8192
rect 8168 8127 8484 8128
rect 22612 8192 22928 8193
rect 22612 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22928 8192
rect 22612 8127 22928 8128
rect 37056 8192 37372 8193
rect 37056 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37372 8192
rect 37056 8127 37372 8128
rect 51500 8192 51816 8193
rect 51500 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51816 8192
rect 51500 8127 51816 8128
rect 15390 7648 15706 7649
rect 15390 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15706 7648
rect 15390 7583 15706 7584
rect 29834 7648 30150 7649
rect 29834 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30150 7648
rect 29834 7583 30150 7584
rect 44278 7648 44594 7649
rect 44278 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44594 7648
rect 44278 7583 44594 7584
rect 58722 7648 59038 7649
rect 58722 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59038 7648
rect 58722 7583 59038 7584
rect 49509 7306 49575 7309
rect 54937 7306 55003 7309
rect 49509 7304 55003 7306
rect 49509 7248 49514 7304
rect 49570 7248 54942 7304
rect 54998 7248 55003 7304
rect 49509 7246 55003 7248
rect 49509 7243 49575 7246
rect 54937 7243 55003 7246
rect 8168 7104 8484 7105
rect 8168 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8484 7104
rect 8168 7039 8484 7040
rect 22612 7104 22928 7105
rect 22612 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22928 7104
rect 22612 7039 22928 7040
rect 37056 7104 37372 7105
rect 37056 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37372 7104
rect 37056 7039 37372 7040
rect 51500 7104 51816 7105
rect 51500 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51816 7104
rect 51500 7039 51816 7040
rect 37457 6898 37523 6901
rect 41965 6898 42031 6901
rect 37457 6896 42031 6898
rect 37457 6840 37462 6896
rect 37518 6840 41970 6896
rect 42026 6840 42031 6896
rect 37457 6838 42031 6840
rect 37457 6835 37523 6838
rect 41965 6835 42031 6838
rect 49141 6626 49207 6629
rect 57237 6626 57303 6629
rect 49141 6624 57303 6626
rect 49141 6568 49146 6624
rect 49202 6568 57242 6624
rect 57298 6568 57303 6624
rect 49141 6566 57303 6568
rect 49141 6563 49207 6566
rect 57237 6563 57303 6566
rect 15390 6560 15706 6561
rect 15390 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15706 6560
rect 15390 6495 15706 6496
rect 29834 6560 30150 6561
rect 29834 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30150 6560
rect 29834 6495 30150 6496
rect 44278 6560 44594 6561
rect 44278 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44594 6560
rect 44278 6495 44594 6496
rect 58722 6560 59038 6561
rect 58722 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59038 6560
rect 58722 6495 59038 6496
rect 8661 6354 8727 6357
rect 33409 6354 33475 6357
rect 8661 6352 33475 6354
rect 8661 6296 8666 6352
rect 8722 6296 33414 6352
rect 33470 6296 33475 6352
rect 8661 6294 33475 6296
rect 8661 6291 8727 6294
rect 33409 6291 33475 6294
rect 30465 6218 30531 6221
rect 32765 6218 32831 6221
rect 30465 6216 32831 6218
rect 30465 6160 30470 6216
rect 30526 6160 32770 6216
rect 32826 6160 32831 6216
rect 30465 6158 32831 6160
rect 30465 6155 30531 6158
rect 32765 6155 32831 6158
rect 30005 6082 30071 6085
rect 31845 6082 31911 6085
rect 30005 6080 31911 6082
rect 30005 6024 30010 6080
rect 30066 6024 31850 6080
rect 31906 6024 31911 6080
rect 30005 6022 31911 6024
rect 30005 6019 30071 6022
rect 31845 6019 31911 6022
rect 8168 6016 8484 6017
rect 8168 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8484 6016
rect 8168 5951 8484 5952
rect 22612 6016 22928 6017
rect 22612 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22928 6016
rect 22612 5951 22928 5952
rect 37056 6016 37372 6017
rect 37056 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37372 6016
rect 37056 5951 37372 5952
rect 51500 6016 51816 6017
rect 51500 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51816 6016
rect 51500 5951 51816 5952
rect 30557 5946 30623 5949
rect 32949 5946 33015 5949
rect 30557 5944 33015 5946
rect 30557 5888 30562 5944
rect 30618 5888 32954 5944
rect 33010 5888 33015 5944
rect 30557 5886 33015 5888
rect 30557 5883 30623 5886
rect 32949 5883 33015 5886
rect 8937 5810 9003 5813
rect 34697 5810 34763 5813
rect 8937 5808 34763 5810
rect 8937 5752 8942 5808
rect 8998 5752 34702 5808
rect 34758 5752 34763 5808
rect 8937 5750 34763 5752
rect 8937 5747 9003 5750
rect 34697 5747 34763 5750
rect 20253 5674 20319 5677
rect 23381 5674 23447 5677
rect 24761 5674 24827 5677
rect 20253 5672 24827 5674
rect 20253 5616 20258 5672
rect 20314 5616 23386 5672
rect 23442 5616 24766 5672
rect 24822 5616 24827 5672
rect 20253 5614 24827 5616
rect 20253 5611 20319 5614
rect 23381 5611 23447 5614
rect 24761 5611 24827 5614
rect 39021 5674 39087 5677
rect 44725 5674 44791 5677
rect 48221 5674 48287 5677
rect 39021 5672 48287 5674
rect 39021 5616 39026 5672
rect 39082 5616 44730 5672
rect 44786 5616 48226 5672
rect 48282 5616 48287 5672
rect 39021 5614 48287 5616
rect 39021 5611 39087 5614
rect 44725 5611 44791 5614
rect 48221 5611 48287 5614
rect 55121 5674 55187 5677
rect 57973 5674 58039 5677
rect 55121 5672 58039 5674
rect 55121 5616 55126 5672
rect 55182 5616 57978 5672
rect 58034 5616 58039 5672
rect 55121 5614 58039 5616
rect 55121 5611 55187 5614
rect 57973 5611 58039 5614
rect 15390 5472 15706 5473
rect 15390 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15706 5472
rect 15390 5407 15706 5408
rect 29834 5472 30150 5473
rect 29834 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30150 5472
rect 29834 5407 30150 5408
rect 44278 5472 44594 5473
rect 44278 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44594 5472
rect 44278 5407 44594 5408
rect 58722 5472 59038 5473
rect 58722 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59038 5472
rect 58722 5407 59038 5408
rect 13721 5266 13787 5269
rect 56961 5266 57027 5269
rect 13721 5264 57027 5266
rect 13721 5208 13726 5264
rect 13782 5208 56966 5264
rect 57022 5208 57027 5264
rect 13721 5206 57027 5208
rect 13721 5203 13787 5206
rect 56961 5203 57027 5206
rect 11145 5130 11211 5133
rect 56409 5130 56475 5133
rect 11145 5128 56475 5130
rect 11145 5072 11150 5128
rect 11206 5072 56414 5128
rect 56470 5072 56475 5128
rect 11145 5070 56475 5072
rect 11145 5067 11211 5070
rect 56409 5067 56475 5070
rect 8168 4928 8484 4929
rect 8168 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8484 4928
rect 8168 4863 8484 4864
rect 22612 4928 22928 4929
rect 22612 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22928 4928
rect 22612 4863 22928 4864
rect 37056 4928 37372 4929
rect 37056 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37372 4928
rect 37056 4863 37372 4864
rect 51500 4928 51816 4929
rect 51500 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51816 4928
rect 51500 4863 51816 4864
rect 34881 4858 34947 4861
rect 26926 4856 34947 4858
rect 26926 4800 34886 4856
rect 34942 4800 34947 4856
rect 26926 4798 34947 4800
rect 9121 4722 9187 4725
rect 26926 4722 26986 4798
rect 34881 4795 34947 4798
rect 9121 4720 26986 4722
rect 9121 4664 9126 4720
rect 9182 4664 26986 4720
rect 9121 4662 26986 4664
rect 31201 4722 31267 4725
rect 38009 4722 38075 4725
rect 31201 4720 38075 4722
rect 31201 4664 31206 4720
rect 31262 4664 38014 4720
rect 38070 4664 38075 4720
rect 31201 4662 38075 4664
rect 9121 4659 9187 4662
rect 31201 4659 31267 4662
rect 38009 4659 38075 4662
rect 33317 4586 33383 4589
rect 42425 4586 42491 4589
rect 33317 4584 42491 4586
rect 33317 4528 33322 4584
rect 33378 4528 42430 4584
rect 42486 4528 42491 4584
rect 33317 4526 42491 4528
rect 33317 4523 33383 4526
rect 42425 4523 42491 4526
rect 15390 4384 15706 4385
rect 15390 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15706 4384
rect 15390 4319 15706 4320
rect 29834 4384 30150 4385
rect 29834 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30150 4384
rect 29834 4319 30150 4320
rect 44278 4384 44594 4385
rect 44278 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44594 4384
rect 44278 4319 44594 4320
rect 58722 4384 59038 4385
rect 58722 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59038 4384
rect 58722 4319 59038 4320
rect 55305 4314 55371 4317
rect 57881 4314 57947 4317
rect 55305 4312 57947 4314
rect 55305 4256 55310 4312
rect 55366 4256 57886 4312
rect 57942 4256 57947 4312
rect 55305 4254 57947 4256
rect 55305 4251 55371 4254
rect 57881 4251 57947 4254
rect 5441 4178 5507 4181
rect 33409 4178 33475 4181
rect 5441 4176 33475 4178
rect 5441 4120 5446 4176
rect 5502 4120 33414 4176
rect 33470 4120 33475 4176
rect 5441 4118 33475 4120
rect 5441 4115 5507 4118
rect 33409 4115 33475 4118
rect 27337 4042 27403 4045
rect 35157 4042 35223 4045
rect 37273 4042 37339 4045
rect 27337 4040 35223 4042
rect 27337 3984 27342 4040
rect 27398 3984 35162 4040
rect 35218 3984 35223 4040
rect 27337 3982 35223 3984
rect 27337 3979 27403 3982
rect 35157 3979 35223 3982
rect 35390 4040 37339 4042
rect 35390 3984 37278 4040
rect 37334 3984 37339 4040
rect 35390 3982 37339 3984
rect 32949 3906 33015 3909
rect 35390 3906 35450 3982
rect 37273 3979 37339 3982
rect 41321 4042 41387 4045
rect 42885 4042 42951 4045
rect 41321 4040 42951 4042
rect 41321 3984 41326 4040
rect 41382 3984 42890 4040
rect 42946 3984 42951 4040
rect 41321 3982 42951 3984
rect 41321 3979 41387 3982
rect 42885 3979 42951 3982
rect 47577 4042 47643 4045
rect 51257 4042 51323 4045
rect 47577 4040 51323 4042
rect 47577 3984 47582 4040
rect 47638 3984 51262 4040
rect 51318 3984 51323 4040
rect 47577 3982 51323 3984
rect 47577 3979 47643 3982
rect 51257 3979 51323 3982
rect 53649 4042 53715 4045
rect 55397 4042 55463 4045
rect 56593 4042 56659 4045
rect 57145 4044 57211 4045
rect 53649 4040 56659 4042
rect 53649 3984 53654 4040
rect 53710 3984 55402 4040
rect 55458 3984 56598 4040
rect 56654 3984 56659 4040
rect 53649 3982 56659 3984
rect 53649 3979 53715 3982
rect 55397 3979 55463 3982
rect 56593 3979 56659 3982
rect 57094 3980 57100 4044
rect 57164 4042 57211 4044
rect 57164 4040 57256 4042
rect 57206 3984 57256 4040
rect 57164 3982 57256 3984
rect 57164 3980 57211 3982
rect 57145 3979 57211 3980
rect 32949 3904 35450 3906
rect 32949 3848 32954 3904
rect 33010 3848 35450 3904
rect 32949 3846 35450 3848
rect 49325 3906 49391 3909
rect 51073 3906 51139 3909
rect 49325 3904 51139 3906
rect 49325 3848 49330 3904
rect 49386 3848 51078 3904
rect 51134 3848 51139 3904
rect 49325 3846 51139 3848
rect 32949 3843 33015 3846
rect 49325 3843 49391 3846
rect 51073 3843 51139 3846
rect 52545 3906 52611 3909
rect 58433 3906 58499 3909
rect 52545 3904 58499 3906
rect 52545 3848 52550 3904
rect 52606 3848 58438 3904
rect 58494 3848 58499 3904
rect 52545 3846 58499 3848
rect 52545 3843 52611 3846
rect 58433 3843 58499 3846
rect 8168 3840 8484 3841
rect 8168 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8484 3840
rect 8168 3775 8484 3776
rect 22612 3840 22928 3841
rect 22612 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22928 3840
rect 22612 3775 22928 3776
rect 37056 3840 37372 3841
rect 37056 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37372 3840
rect 37056 3775 37372 3776
rect 51500 3840 51816 3841
rect 51500 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51816 3840
rect 51500 3775 51816 3776
rect 48129 3770 48195 3773
rect 50705 3770 50771 3773
rect 48129 3768 50771 3770
rect 48129 3712 48134 3768
rect 48190 3712 50710 3768
rect 50766 3712 50771 3768
rect 48129 3710 50771 3712
rect 48129 3707 48195 3710
rect 50705 3707 50771 3710
rect 5993 3634 6059 3637
rect 46749 3634 46815 3637
rect 52085 3634 52151 3637
rect 5993 3632 52151 3634
rect 5993 3576 5998 3632
rect 6054 3576 46754 3632
rect 46810 3576 52090 3632
rect 52146 3576 52151 3632
rect 5993 3574 52151 3576
rect 5993 3571 6059 3574
rect 46749 3571 46815 3574
rect 52085 3571 52151 3574
rect 933 3498 999 3501
rect 30189 3498 30255 3501
rect 933 3496 30255 3498
rect 933 3440 938 3496
rect 994 3440 30194 3496
rect 30250 3440 30255 3496
rect 933 3438 30255 3440
rect 933 3435 999 3438
rect 30189 3435 30255 3438
rect 43805 3498 43871 3501
rect 46473 3498 46539 3501
rect 43805 3496 46539 3498
rect 43805 3440 43810 3496
rect 43866 3440 46478 3496
rect 46534 3440 46539 3496
rect 43805 3438 46539 3440
rect 43805 3435 43871 3438
rect 46473 3435 46539 3438
rect 51993 3498 52059 3501
rect 58341 3498 58407 3501
rect 51993 3496 58407 3498
rect 51993 3440 51998 3496
rect 52054 3440 58346 3496
rect 58402 3440 58407 3496
rect 51993 3438 58407 3440
rect 51993 3435 52059 3438
rect 58341 3435 58407 3438
rect 15390 3296 15706 3297
rect 15390 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15706 3296
rect 15390 3231 15706 3232
rect 29834 3296 30150 3297
rect 29834 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30150 3296
rect 29834 3231 30150 3232
rect 44278 3296 44594 3297
rect 44278 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44594 3296
rect 44278 3231 44594 3232
rect 58722 3296 59038 3297
rect 58722 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59038 3296
rect 58722 3231 59038 3232
rect 31201 3226 31267 3229
rect 34053 3226 34119 3229
rect 31201 3224 34119 3226
rect 31201 3168 31206 3224
rect 31262 3168 34058 3224
rect 34114 3168 34119 3224
rect 31201 3166 34119 3168
rect 31201 3163 31267 3166
rect 34053 3163 34119 3166
rect 34881 3226 34947 3229
rect 39481 3226 39547 3229
rect 34881 3224 39547 3226
rect 34881 3168 34886 3224
rect 34942 3168 39486 3224
rect 39542 3168 39547 3224
rect 34881 3166 39547 3168
rect 34881 3163 34947 3166
rect 39481 3163 39547 3166
rect 9489 3090 9555 3093
rect 11605 3090 11671 3093
rect 12341 3090 12407 3093
rect 9489 3088 12407 3090
rect 9489 3032 9494 3088
rect 9550 3032 11610 3088
rect 11666 3032 12346 3088
rect 12402 3032 12407 3088
rect 9489 3030 12407 3032
rect 9489 3027 9555 3030
rect 11605 3027 11671 3030
rect 12341 3027 12407 3030
rect 16297 3090 16363 3093
rect 27337 3090 27403 3093
rect 16297 3088 27403 3090
rect 16297 3032 16302 3088
rect 16358 3032 27342 3088
rect 27398 3032 27403 3088
rect 16297 3030 27403 3032
rect 16297 3027 16363 3030
rect 27337 3027 27403 3030
rect 27797 3090 27863 3093
rect 42333 3090 42399 3093
rect 27797 3088 42399 3090
rect 27797 3032 27802 3088
rect 27858 3032 42338 3088
rect 42394 3032 42399 3088
rect 27797 3030 42399 3032
rect 27797 3027 27863 3030
rect 42333 3027 42399 3030
rect 42885 3090 42951 3093
rect 46381 3090 46447 3093
rect 48037 3090 48103 3093
rect 42885 3088 48103 3090
rect 42885 3032 42890 3088
rect 42946 3032 46386 3088
rect 46442 3032 48042 3088
rect 48098 3032 48103 3088
rect 42885 3030 48103 3032
rect 42885 3027 42951 3030
rect 46381 3027 46447 3030
rect 48037 3027 48103 3030
rect 15101 2954 15167 2957
rect 18965 2954 19031 2957
rect 15101 2952 19031 2954
rect 15101 2896 15106 2952
rect 15162 2896 18970 2952
rect 19026 2896 19031 2952
rect 15101 2894 19031 2896
rect 15101 2891 15167 2894
rect 18965 2891 19031 2894
rect 32305 2954 32371 2957
rect 34605 2954 34671 2957
rect 32305 2952 34671 2954
rect 32305 2896 32310 2952
rect 32366 2896 34610 2952
rect 34666 2896 34671 2952
rect 32305 2894 34671 2896
rect 32305 2891 32371 2894
rect 34605 2891 34671 2894
rect 35157 2954 35223 2957
rect 38745 2954 38811 2957
rect 35157 2952 38811 2954
rect 35157 2896 35162 2952
rect 35218 2896 38750 2952
rect 38806 2896 38811 2952
rect 35157 2894 38811 2896
rect 35157 2891 35223 2894
rect 38745 2891 38811 2894
rect 42793 2954 42859 2957
rect 55121 2954 55187 2957
rect 42793 2952 55187 2954
rect 42793 2896 42798 2952
rect 42854 2896 55126 2952
rect 55182 2896 55187 2952
rect 42793 2894 55187 2896
rect 42793 2891 42859 2894
rect 55121 2891 55187 2894
rect 53373 2818 53439 2821
rect 57881 2818 57947 2821
rect 53373 2816 57947 2818
rect 53373 2760 53378 2816
rect 53434 2760 57886 2816
rect 57942 2760 57947 2816
rect 53373 2758 57947 2760
rect 53373 2755 53439 2758
rect 57881 2755 57947 2758
rect 8168 2752 8484 2753
rect 8168 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8484 2752
rect 8168 2687 8484 2688
rect 22612 2752 22928 2753
rect 22612 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22928 2752
rect 22612 2687 22928 2688
rect 37056 2752 37372 2753
rect 37056 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37372 2752
rect 37056 2687 37372 2688
rect 51500 2752 51816 2753
rect 51500 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51816 2752
rect 51500 2687 51816 2688
rect 15390 2208 15706 2209
rect 15390 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15706 2208
rect 15390 2143 15706 2144
rect 29834 2208 30150 2209
rect 29834 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30150 2208
rect 29834 2143 30150 2144
rect 44278 2208 44594 2209
rect 44278 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44594 2208
rect 44278 2143 44594 2144
rect 58722 2208 59038 2209
rect 58722 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59038 2208
rect 58722 2143 59038 2144
<< via3 >>
rect 8174 27772 8238 27776
rect 8174 27716 8178 27772
rect 8178 27716 8234 27772
rect 8234 27716 8238 27772
rect 8174 27712 8238 27716
rect 8254 27772 8318 27776
rect 8254 27716 8258 27772
rect 8258 27716 8314 27772
rect 8314 27716 8318 27772
rect 8254 27712 8318 27716
rect 8334 27772 8398 27776
rect 8334 27716 8338 27772
rect 8338 27716 8394 27772
rect 8394 27716 8398 27772
rect 8334 27712 8398 27716
rect 8414 27772 8478 27776
rect 8414 27716 8418 27772
rect 8418 27716 8474 27772
rect 8474 27716 8478 27772
rect 8414 27712 8478 27716
rect 22618 27772 22682 27776
rect 22618 27716 22622 27772
rect 22622 27716 22678 27772
rect 22678 27716 22682 27772
rect 22618 27712 22682 27716
rect 22698 27772 22762 27776
rect 22698 27716 22702 27772
rect 22702 27716 22758 27772
rect 22758 27716 22762 27772
rect 22698 27712 22762 27716
rect 22778 27772 22842 27776
rect 22778 27716 22782 27772
rect 22782 27716 22838 27772
rect 22838 27716 22842 27772
rect 22778 27712 22842 27716
rect 22858 27772 22922 27776
rect 22858 27716 22862 27772
rect 22862 27716 22918 27772
rect 22918 27716 22922 27772
rect 22858 27712 22922 27716
rect 37062 27772 37126 27776
rect 37062 27716 37066 27772
rect 37066 27716 37122 27772
rect 37122 27716 37126 27772
rect 37062 27712 37126 27716
rect 37142 27772 37206 27776
rect 37142 27716 37146 27772
rect 37146 27716 37202 27772
rect 37202 27716 37206 27772
rect 37142 27712 37206 27716
rect 37222 27772 37286 27776
rect 37222 27716 37226 27772
rect 37226 27716 37282 27772
rect 37282 27716 37286 27772
rect 37222 27712 37286 27716
rect 37302 27772 37366 27776
rect 37302 27716 37306 27772
rect 37306 27716 37362 27772
rect 37362 27716 37366 27772
rect 37302 27712 37366 27716
rect 51506 27772 51570 27776
rect 51506 27716 51510 27772
rect 51510 27716 51566 27772
rect 51566 27716 51570 27772
rect 51506 27712 51570 27716
rect 51586 27772 51650 27776
rect 51586 27716 51590 27772
rect 51590 27716 51646 27772
rect 51646 27716 51650 27772
rect 51586 27712 51650 27716
rect 51666 27772 51730 27776
rect 51666 27716 51670 27772
rect 51670 27716 51726 27772
rect 51726 27716 51730 27772
rect 51666 27712 51730 27716
rect 51746 27772 51810 27776
rect 51746 27716 51750 27772
rect 51750 27716 51806 27772
rect 51806 27716 51810 27772
rect 51746 27712 51810 27716
rect 15396 27228 15460 27232
rect 15396 27172 15400 27228
rect 15400 27172 15456 27228
rect 15456 27172 15460 27228
rect 15396 27168 15460 27172
rect 15476 27228 15540 27232
rect 15476 27172 15480 27228
rect 15480 27172 15536 27228
rect 15536 27172 15540 27228
rect 15476 27168 15540 27172
rect 15556 27228 15620 27232
rect 15556 27172 15560 27228
rect 15560 27172 15616 27228
rect 15616 27172 15620 27228
rect 15556 27168 15620 27172
rect 15636 27228 15700 27232
rect 15636 27172 15640 27228
rect 15640 27172 15696 27228
rect 15696 27172 15700 27228
rect 15636 27168 15700 27172
rect 29840 27228 29904 27232
rect 29840 27172 29844 27228
rect 29844 27172 29900 27228
rect 29900 27172 29904 27228
rect 29840 27168 29904 27172
rect 29920 27228 29984 27232
rect 29920 27172 29924 27228
rect 29924 27172 29980 27228
rect 29980 27172 29984 27228
rect 29920 27168 29984 27172
rect 30000 27228 30064 27232
rect 30000 27172 30004 27228
rect 30004 27172 30060 27228
rect 30060 27172 30064 27228
rect 30000 27168 30064 27172
rect 30080 27228 30144 27232
rect 30080 27172 30084 27228
rect 30084 27172 30140 27228
rect 30140 27172 30144 27228
rect 30080 27168 30144 27172
rect 44284 27228 44348 27232
rect 44284 27172 44288 27228
rect 44288 27172 44344 27228
rect 44344 27172 44348 27228
rect 44284 27168 44348 27172
rect 44364 27228 44428 27232
rect 44364 27172 44368 27228
rect 44368 27172 44424 27228
rect 44424 27172 44428 27228
rect 44364 27168 44428 27172
rect 44444 27228 44508 27232
rect 44444 27172 44448 27228
rect 44448 27172 44504 27228
rect 44504 27172 44508 27228
rect 44444 27168 44508 27172
rect 44524 27228 44588 27232
rect 44524 27172 44528 27228
rect 44528 27172 44584 27228
rect 44584 27172 44588 27228
rect 44524 27168 44588 27172
rect 58728 27228 58792 27232
rect 58728 27172 58732 27228
rect 58732 27172 58788 27228
rect 58788 27172 58792 27228
rect 58728 27168 58792 27172
rect 58808 27228 58872 27232
rect 58808 27172 58812 27228
rect 58812 27172 58868 27228
rect 58868 27172 58872 27228
rect 58808 27168 58872 27172
rect 58888 27228 58952 27232
rect 58888 27172 58892 27228
rect 58892 27172 58948 27228
rect 58948 27172 58952 27228
rect 58888 27168 58952 27172
rect 58968 27228 59032 27232
rect 58968 27172 58972 27228
rect 58972 27172 59028 27228
rect 59028 27172 59032 27228
rect 58968 27168 59032 27172
rect 8174 26684 8238 26688
rect 8174 26628 8178 26684
rect 8178 26628 8234 26684
rect 8234 26628 8238 26684
rect 8174 26624 8238 26628
rect 8254 26684 8318 26688
rect 8254 26628 8258 26684
rect 8258 26628 8314 26684
rect 8314 26628 8318 26684
rect 8254 26624 8318 26628
rect 8334 26684 8398 26688
rect 8334 26628 8338 26684
rect 8338 26628 8394 26684
rect 8394 26628 8398 26684
rect 8334 26624 8398 26628
rect 8414 26684 8478 26688
rect 8414 26628 8418 26684
rect 8418 26628 8474 26684
rect 8474 26628 8478 26684
rect 8414 26624 8478 26628
rect 22618 26684 22682 26688
rect 22618 26628 22622 26684
rect 22622 26628 22678 26684
rect 22678 26628 22682 26684
rect 22618 26624 22682 26628
rect 22698 26684 22762 26688
rect 22698 26628 22702 26684
rect 22702 26628 22758 26684
rect 22758 26628 22762 26684
rect 22698 26624 22762 26628
rect 22778 26684 22842 26688
rect 22778 26628 22782 26684
rect 22782 26628 22838 26684
rect 22838 26628 22842 26684
rect 22778 26624 22842 26628
rect 22858 26684 22922 26688
rect 22858 26628 22862 26684
rect 22862 26628 22918 26684
rect 22918 26628 22922 26684
rect 22858 26624 22922 26628
rect 37062 26684 37126 26688
rect 37062 26628 37066 26684
rect 37066 26628 37122 26684
rect 37122 26628 37126 26684
rect 37062 26624 37126 26628
rect 37142 26684 37206 26688
rect 37142 26628 37146 26684
rect 37146 26628 37202 26684
rect 37202 26628 37206 26684
rect 37142 26624 37206 26628
rect 37222 26684 37286 26688
rect 37222 26628 37226 26684
rect 37226 26628 37282 26684
rect 37282 26628 37286 26684
rect 37222 26624 37286 26628
rect 37302 26684 37366 26688
rect 37302 26628 37306 26684
rect 37306 26628 37362 26684
rect 37362 26628 37366 26684
rect 37302 26624 37366 26628
rect 51506 26684 51570 26688
rect 51506 26628 51510 26684
rect 51510 26628 51566 26684
rect 51566 26628 51570 26684
rect 51506 26624 51570 26628
rect 51586 26684 51650 26688
rect 51586 26628 51590 26684
rect 51590 26628 51646 26684
rect 51646 26628 51650 26684
rect 51586 26624 51650 26628
rect 51666 26684 51730 26688
rect 51666 26628 51670 26684
rect 51670 26628 51726 26684
rect 51726 26628 51730 26684
rect 51666 26624 51730 26628
rect 51746 26684 51810 26688
rect 51746 26628 51750 26684
rect 51750 26628 51806 26684
rect 51806 26628 51810 26684
rect 51746 26624 51810 26628
rect 15396 26140 15460 26144
rect 15396 26084 15400 26140
rect 15400 26084 15456 26140
rect 15456 26084 15460 26140
rect 15396 26080 15460 26084
rect 15476 26140 15540 26144
rect 15476 26084 15480 26140
rect 15480 26084 15536 26140
rect 15536 26084 15540 26140
rect 15476 26080 15540 26084
rect 15556 26140 15620 26144
rect 15556 26084 15560 26140
rect 15560 26084 15616 26140
rect 15616 26084 15620 26140
rect 15556 26080 15620 26084
rect 15636 26140 15700 26144
rect 15636 26084 15640 26140
rect 15640 26084 15696 26140
rect 15696 26084 15700 26140
rect 15636 26080 15700 26084
rect 29840 26140 29904 26144
rect 29840 26084 29844 26140
rect 29844 26084 29900 26140
rect 29900 26084 29904 26140
rect 29840 26080 29904 26084
rect 29920 26140 29984 26144
rect 29920 26084 29924 26140
rect 29924 26084 29980 26140
rect 29980 26084 29984 26140
rect 29920 26080 29984 26084
rect 30000 26140 30064 26144
rect 30000 26084 30004 26140
rect 30004 26084 30060 26140
rect 30060 26084 30064 26140
rect 30000 26080 30064 26084
rect 30080 26140 30144 26144
rect 30080 26084 30084 26140
rect 30084 26084 30140 26140
rect 30140 26084 30144 26140
rect 30080 26080 30144 26084
rect 44284 26140 44348 26144
rect 44284 26084 44288 26140
rect 44288 26084 44344 26140
rect 44344 26084 44348 26140
rect 44284 26080 44348 26084
rect 44364 26140 44428 26144
rect 44364 26084 44368 26140
rect 44368 26084 44424 26140
rect 44424 26084 44428 26140
rect 44364 26080 44428 26084
rect 44444 26140 44508 26144
rect 44444 26084 44448 26140
rect 44448 26084 44504 26140
rect 44504 26084 44508 26140
rect 44444 26080 44508 26084
rect 44524 26140 44588 26144
rect 44524 26084 44528 26140
rect 44528 26084 44584 26140
rect 44584 26084 44588 26140
rect 44524 26080 44588 26084
rect 58728 26140 58792 26144
rect 58728 26084 58732 26140
rect 58732 26084 58788 26140
rect 58788 26084 58792 26140
rect 58728 26080 58792 26084
rect 58808 26140 58872 26144
rect 58808 26084 58812 26140
rect 58812 26084 58868 26140
rect 58868 26084 58872 26140
rect 58808 26080 58872 26084
rect 58888 26140 58952 26144
rect 58888 26084 58892 26140
rect 58892 26084 58948 26140
rect 58948 26084 58952 26140
rect 58888 26080 58952 26084
rect 58968 26140 59032 26144
rect 58968 26084 58972 26140
rect 58972 26084 59028 26140
rect 59028 26084 59032 26140
rect 58968 26080 59032 26084
rect 8174 25596 8238 25600
rect 8174 25540 8178 25596
rect 8178 25540 8234 25596
rect 8234 25540 8238 25596
rect 8174 25536 8238 25540
rect 8254 25596 8318 25600
rect 8254 25540 8258 25596
rect 8258 25540 8314 25596
rect 8314 25540 8318 25596
rect 8254 25536 8318 25540
rect 8334 25596 8398 25600
rect 8334 25540 8338 25596
rect 8338 25540 8394 25596
rect 8394 25540 8398 25596
rect 8334 25536 8398 25540
rect 8414 25596 8478 25600
rect 8414 25540 8418 25596
rect 8418 25540 8474 25596
rect 8474 25540 8478 25596
rect 8414 25536 8478 25540
rect 22618 25596 22682 25600
rect 22618 25540 22622 25596
rect 22622 25540 22678 25596
rect 22678 25540 22682 25596
rect 22618 25536 22682 25540
rect 22698 25596 22762 25600
rect 22698 25540 22702 25596
rect 22702 25540 22758 25596
rect 22758 25540 22762 25596
rect 22698 25536 22762 25540
rect 22778 25596 22842 25600
rect 22778 25540 22782 25596
rect 22782 25540 22838 25596
rect 22838 25540 22842 25596
rect 22778 25536 22842 25540
rect 22858 25596 22922 25600
rect 22858 25540 22862 25596
rect 22862 25540 22918 25596
rect 22918 25540 22922 25596
rect 22858 25536 22922 25540
rect 37062 25596 37126 25600
rect 37062 25540 37066 25596
rect 37066 25540 37122 25596
rect 37122 25540 37126 25596
rect 37062 25536 37126 25540
rect 37142 25596 37206 25600
rect 37142 25540 37146 25596
rect 37146 25540 37202 25596
rect 37202 25540 37206 25596
rect 37142 25536 37206 25540
rect 37222 25596 37286 25600
rect 37222 25540 37226 25596
rect 37226 25540 37282 25596
rect 37282 25540 37286 25596
rect 37222 25536 37286 25540
rect 37302 25596 37366 25600
rect 37302 25540 37306 25596
rect 37306 25540 37362 25596
rect 37362 25540 37366 25596
rect 37302 25536 37366 25540
rect 51506 25596 51570 25600
rect 51506 25540 51510 25596
rect 51510 25540 51566 25596
rect 51566 25540 51570 25596
rect 51506 25536 51570 25540
rect 51586 25596 51650 25600
rect 51586 25540 51590 25596
rect 51590 25540 51646 25596
rect 51646 25540 51650 25596
rect 51586 25536 51650 25540
rect 51666 25596 51730 25600
rect 51666 25540 51670 25596
rect 51670 25540 51726 25596
rect 51726 25540 51730 25596
rect 51666 25536 51730 25540
rect 51746 25596 51810 25600
rect 51746 25540 51750 25596
rect 51750 25540 51806 25596
rect 51806 25540 51810 25596
rect 51746 25536 51810 25540
rect 15396 25052 15460 25056
rect 15396 24996 15400 25052
rect 15400 24996 15456 25052
rect 15456 24996 15460 25052
rect 15396 24992 15460 24996
rect 15476 25052 15540 25056
rect 15476 24996 15480 25052
rect 15480 24996 15536 25052
rect 15536 24996 15540 25052
rect 15476 24992 15540 24996
rect 15556 25052 15620 25056
rect 15556 24996 15560 25052
rect 15560 24996 15616 25052
rect 15616 24996 15620 25052
rect 15556 24992 15620 24996
rect 15636 25052 15700 25056
rect 15636 24996 15640 25052
rect 15640 24996 15696 25052
rect 15696 24996 15700 25052
rect 15636 24992 15700 24996
rect 29840 25052 29904 25056
rect 29840 24996 29844 25052
rect 29844 24996 29900 25052
rect 29900 24996 29904 25052
rect 29840 24992 29904 24996
rect 29920 25052 29984 25056
rect 29920 24996 29924 25052
rect 29924 24996 29980 25052
rect 29980 24996 29984 25052
rect 29920 24992 29984 24996
rect 30000 25052 30064 25056
rect 30000 24996 30004 25052
rect 30004 24996 30060 25052
rect 30060 24996 30064 25052
rect 30000 24992 30064 24996
rect 30080 25052 30144 25056
rect 30080 24996 30084 25052
rect 30084 24996 30140 25052
rect 30140 24996 30144 25052
rect 30080 24992 30144 24996
rect 44284 25052 44348 25056
rect 44284 24996 44288 25052
rect 44288 24996 44344 25052
rect 44344 24996 44348 25052
rect 44284 24992 44348 24996
rect 44364 25052 44428 25056
rect 44364 24996 44368 25052
rect 44368 24996 44424 25052
rect 44424 24996 44428 25052
rect 44364 24992 44428 24996
rect 44444 25052 44508 25056
rect 44444 24996 44448 25052
rect 44448 24996 44504 25052
rect 44504 24996 44508 25052
rect 44444 24992 44508 24996
rect 44524 25052 44588 25056
rect 44524 24996 44528 25052
rect 44528 24996 44584 25052
rect 44584 24996 44588 25052
rect 44524 24992 44588 24996
rect 58728 25052 58792 25056
rect 58728 24996 58732 25052
rect 58732 24996 58788 25052
rect 58788 24996 58792 25052
rect 58728 24992 58792 24996
rect 58808 25052 58872 25056
rect 58808 24996 58812 25052
rect 58812 24996 58868 25052
rect 58868 24996 58872 25052
rect 58808 24992 58872 24996
rect 58888 25052 58952 25056
rect 58888 24996 58892 25052
rect 58892 24996 58948 25052
rect 58948 24996 58952 25052
rect 58888 24992 58952 24996
rect 58968 25052 59032 25056
rect 58968 24996 58972 25052
rect 58972 24996 59028 25052
rect 59028 24996 59032 25052
rect 58968 24992 59032 24996
rect 8174 24508 8238 24512
rect 8174 24452 8178 24508
rect 8178 24452 8234 24508
rect 8234 24452 8238 24508
rect 8174 24448 8238 24452
rect 8254 24508 8318 24512
rect 8254 24452 8258 24508
rect 8258 24452 8314 24508
rect 8314 24452 8318 24508
rect 8254 24448 8318 24452
rect 8334 24508 8398 24512
rect 8334 24452 8338 24508
rect 8338 24452 8394 24508
rect 8394 24452 8398 24508
rect 8334 24448 8398 24452
rect 8414 24508 8478 24512
rect 8414 24452 8418 24508
rect 8418 24452 8474 24508
rect 8474 24452 8478 24508
rect 8414 24448 8478 24452
rect 22618 24508 22682 24512
rect 22618 24452 22622 24508
rect 22622 24452 22678 24508
rect 22678 24452 22682 24508
rect 22618 24448 22682 24452
rect 22698 24508 22762 24512
rect 22698 24452 22702 24508
rect 22702 24452 22758 24508
rect 22758 24452 22762 24508
rect 22698 24448 22762 24452
rect 22778 24508 22842 24512
rect 22778 24452 22782 24508
rect 22782 24452 22838 24508
rect 22838 24452 22842 24508
rect 22778 24448 22842 24452
rect 22858 24508 22922 24512
rect 22858 24452 22862 24508
rect 22862 24452 22918 24508
rect 22918 24452 22922 24508
rect 22858 24448 22922 24452
rect 37062 24508 37126 24512
rect 37062 24452 37066 24508
rect 37066 24452 37122 24508
rect 37122 24452 37126 24508
rect 37062 24448 37126 24452
rect 37142 24508 37206 24512
rect 37142 24452 37146 24508
rect 37146 24452 37202 24508
rect 37202 24452 37206 24508
rect 37142 24448 37206 24452
rect 37222 24508 37286 24512
rect 37222 24452 37226 24508
rect 37226 24452 37282 24508
rect 37282 24452 37286 24508
rect 37222 24448 37286 24452
rect 37302 24508 37366 24512
rect 37302 24452 37306 24508
rect 37306 24452 37362 24508
rect 37362 24452 37366 24508
rect 37302 24448 37366 24452
rect 51506 24508 51570 24512
rect 51506 24452 51510 24508
rect 51510 24452 51566 24508
rect 51566 24452 51570 24508
rect 51506 24448 51570 24452
rect 51586 24508 51650 24512
rect 51586 24452 51590 24508
rect 51590 24452 51646 24508
rect 51646 24452 51650 24508
rect 51586 24448 51650 24452
rect 51666 24508 51730 24512
rect 51666 24452 51670 24508
rect 51670 24452 51726 24508
rect 51726 24452 51730 24508
rect 51666 24448 51730 24452
rect 51746 24508 51810 24512
rect 51746 24452 51750 24508
rect 51750 24452 51806 24508
rect 51806 24452 51810 24508
rect 51746 24448 51810 24452
rect 15396 23964 15460 23968
rect 15396 23908 15400 23964
rect 15400 23908 15456 23964
rect 15456 23908 15460 23964
rect 15396 23904 15460 23908
rect 15476 23964 15540 23968
rect 15476 23908 15480 23964
rect 15480 23908 15536 23964
rect 15536 23908 15540 23964
rect 15476 23904 15540 23908
rect 15556 23964 15620 23968
rect 15556 23908 15560 23964
rect 15560 23908 15616 23964
rect 15616 23908 15620 23964
rect 15556 23904 15620 23908
rect 15636 23964 15700 23968
rect 15636 23908 15640 23964
rect 15640 23908 15696 23964
rect 15696 23908 15700 23964
rect 15636 23904 15700 23908
rect 29840 23964 29904 23968
rect 29840 23908 29844 23964
rect 29844 23908 29900 23964
rect 29900 23908 29904 23964
rect 29840 23904 29904 23908
rect 29920 23964 29984 23968
rect 29920 23908 29924 23964
rect 29924 23908 29980 23964
rect 29980 23908 29984 23964
rect 29920 23904 29984 23908
rect 30000 23964 30064 23968
rect 30000 23908 30004 23964
rect 30004 23908 30060 23964
rect 30060 23908 30064 23964
rect 30000 23904 30064 23908
rect 30080 23964 30144 23968
rect 30080 23908 30084 23964
rect 30084 23908 30140 23964
rect 30140 23908 30144 23964
rect 30080 23904 30144 23908
rect 44284 23964 44348 23968
rect 44284 23908 44288 23964
rect 44288 23908 44344 23964
rect 44344 23908 44348 23964
rect 44284 23904 44348 23908
rect 44364 23964 44428 23968
rect 44364 23908 44368 23964
rect 44368 23908 44424 23964
rect 44424 23908 44428 23964
rect 44364 23904 44428 23908
rect 44444 23964 44508 23968
rect 44444 23908 44448 23964
rect 44448 23908 44504 23964
rect 44504 23908 44508 23964
rect 44444 23904 44508 23908
rect 44524 23964 44588 23968
rect 44524 23908 44528 23964
rect 44528 23908 44584 23964
rect 44584 23908 44588 23964
rect 44524 23904 44588 23908
rect 58728 23964 58792 23968
rect 58728 23908 58732 23964
rect 58732 23908 58788 23964
rect 58788 23908 58792 23964
rect 58728 23904 58792 23908
rect 58808 23964 58872 23968
rect 58808 23908 58812 23964
rect 58812 23908 58868 23964
rect 58868 23908 58872 23964
rect 58808 23904 58872 23908
rect 58888 23964 58952 23968
rect 58888 23908 58892 23964
rect 58892 23908 58948 23964
rect 58948 23908 58952 23964
rect 58888 23904 58952 23908
rect 58968 23964 59032 23968
rect 58968 23908 58972 23964
rect 58972 23908 59028 23964
rect 59028 23908 59032 23964
rect 58968 23904 59032 23908
rect 8174 23420 8238 23424
rect 8174 23364 8178 23420
rect 8178 23364 8234 23420
rect 8234 23364 8238 23420
rect 8174 23360 8238 23364
rect 8254 23420 8318 23424
rect 8254 23364 8258 23420
rect 8258 23364 8314 23420
rect 8314 23364 8318 23420
rect 8254 23360 8318 23364
rect 8334 23420 8398 23424
rect 8334 23364 8338 23420
rect 8338 23364 8394 23420
rect 8394 23364 8398 23420
rect 8334 23360 8398 23364
rect 8414 23420 8478 23424
rect 8414 23364 8418 23420
rect 8418 23364 8474 23420
rect 8474 23364 8478 23420
rect 8414 23360 8478 23364
rect 22618 23420 22682 23424
rect 22618 23364 22622 23420
rect 22622 23364 22678 23420
rect 22678 23364 22682 23420
rect 22618 23360 22682 23364
rect 22698 23420 22762 23424
rect 22698 23364 22702 23420
rect 22702 23364 22758 23420
rect 22758 23364 22762 23420
rect 22698 23360 22762 23364
rect 22778 23420 22842 23424
rect 22778 23364 22782 23420
rect 22782 23364 22838 23420
rect 22838 23364 22842 23420
rect 22778 23360 22842 23364
rect 22858 23420 22922 23424
rect 22858 23364 22862 23420
rect 22862 23364 22918 23420
rect 22918 23364 22922 23420
rect 22858 23360 22922 23364
rect 37062 23420 37126 23424
rect 37062 23364 37066 23420
rect 37066 23364 37122 23420
rect 37122 23364 37126 23420
rect 37062 23360 37126 23364
rect 37142 23420 37206 23424
rect 37142 23364 37146 23420
rect 37146 23364 37202 23420
rect 37202 23364 37206 23420
rect 37142 23360 37206 23364
rect 37222 23420 37286 23424
rect 37222 23364 37226 23420
rect 37226 23364 37282 23420
rect 37282 23364 37286 23420
rect 37222 23360 37286 23364
rect 37302 23420 37366 23424
rect 37302 23364 37306 23420
rect 37306 23364 37362 23420
rect 37362 23364 37366 23420
rect 37302 23360 37366 23364
rect 51506 23420 51570 23424
rect 51506 23364 51510 23420
rect 51510 23364 51566 23420
rect 51566 23364 51570 23420
rect 51506 23360 51570 23364
rect 51586 23420 51650 23424
rect 51586 23364 51590 23420
rect 51590 23364 51646 23420
rect 51646 23364 51650 23420
rect 51586 23360 51650 23364
rect 51666 23420 51730 23424
rect 51666 23364 51670 23420
rect 51670 23364 51726 23420
rect 51726 23364 51730 23420
rect 51666 23360 51730 23364
rect 51746 23420 51810 23424
rect 51746 23364 51750 23420
rect 51750 23364 51806 23420
rect 51806 23364 51810 23420
rect 51746 23360 51810 23364
rect 15396 22876 15460 22880
rect 15396 22820 15400 22876
rect 15400 22820 15456 22876
rect 15456 22820 15460 22876
rect 15396 22816 15460 22820
rect 15476 22876 15540 22880
rect 15476 22820 15480 22876
rect 15480 22820 15536 22876
rect 15536 22820 15540 22876
rect 15476 22816 15540 22820
rect 15556 22876 15620 22880
rect 15556 22820 15560 22876
rect 15560 22820 15616 22876
rect 15616 22820 15620 22876
rect 15556 22816 15620 22820
rect 15636 22876 15700 22880
rect 15636 22820 15640 22876
rect 15640 22820 15696 22876
rect 15696 22820 15700 22876
rect 15636 22816 15700 22820
rect 29840 22876 29904 22880
rect 29840 22820 29844 22876
rect 29844 22820 29900 22876
rect 29900 22820 29904 22876
rect 29840 22816 29904 22820
rect 29920 22876 29984 22880
rect 29920 22820 29924 22876
rect 29924 22820 29980 22876
rect 29980 22820 29984 22876
rect 29920 22816 29984 22820
rect 30000 22876 30064 22880
rect 30000 22820 30004 22876
rect 30004 22820 30060 22876
rect 30060 22820 30064 22876
rect 30000 22816 30064 22820
rect 30080 22876 30144 22880
rect 30080 22820 30084 22876
rect 30084 22820 30140 22876
rect 30140 22820 30144 22876
rect 30080 22816 30144 22820
rect 44284 22876 44348 22880
rect 44284 22820 44288 22876
rect 44288 22820 44344 22876
rect 44344 22820 44348 22876
rect 44284 22816 44348 22820
rect 44364 22876 44428 22880
rect 44364 22820 44368 22876
rect 44368 22820 44424 22876
rect 44424 22820 44428 22876
rect 44364 22816 44428 22820
rect 44444 22876 44508 22880
rect 44444 22820 44448 22876
rect 44448 22820 44504 22876
rect 44504 22820 44508 22876
rect 44444 22816 44508 22820
rect 44524 22876 44588 22880
rect 44524 22820 44528 22876
rect 44528 22820 44584 22876
rect 44584 22820 44588 22876
rect 44524 22816 44588 22820
rect 58728 22876 58792 22880
rect 58728 22820 58732 22876
rect 58732 22820 58788 22876
rect 58788 22820 58792 22876
rect 58728 22816 58792 22820
rect 58808 22876 58872 22880
rect 58808 22820 58812 22876
rect 58812 22820 58868 22876
rect 58868 22820 58872 22876
rect 58808 22816 58872 22820
rect 58888 22876 58952 22880
rect 58888 22820 58892 22876
rect 58892 22820 58948 22876
rect 58948 22820 58952 22876
rect 58888 22816 58952 22820
rect 58968 22876 59032 22880
rect 58968 22820 58972 22876
rect 58972 22820 59028 22876
rect 59028 22820 59032 22876
rect 58968 22816 59032 22820
rect 8174 22332 8238 22336
rect 8174 22276 8178 22332
rect 8178 22276 8234 22332
rect 8234 22276 8238 22332
rect 8174 22272 8238 22276
rect 8254 22332 8318 22336
rect 8254 22276 8258 22332
rect 8258 22276 8314 22332
rect 8314 22276 8318 22332
rect 8254 22272 8318 22276
rect 8334 22332 8398 22336
rect 8334 22276 8338 22332
rect 8338 22276 8394 22332
rect 8394 22276 8398 22332
rect 8334 22272 8398 22276
rect 8414 22332 8478 22336
rect 8414 22276 8418 22332
rect 8418 22276 8474 22332
rect 8474 22276 8478 22332
rect 8414 22272 8478 22276
rect 22618 22332 22682 22336
rect 22618 22276 22622 22332
rect 22622 22276 22678 22332
rect 22678 22276 22682 22332
rect 22618 22272 22682 22276
rect 22698 22332 22762 22336
rect 22698 22276 22702 22332
rect 22702 22276 22758 22332
rect 22758 22276 22762 22332
rect 22698 22272 22762 22276
rect 22778 22332 22842 22336
rect 22778 22276 22782 22332
rect 22782 22276 22838 22332
rect 22838 22276 22842 22332
rect 22778 22272 22842 22276
rect 22858 22332 22922 22336
rect 22858 22276 22862 22332
rect 22862 22276 22918 22332
rect 22918 22276 22922 22332
rect 22858 22272 22922 22276
rect 37062 22332 37126 22336
rect 37062 22276 37066 22332
rect 37066 22276 37122 22332
rect 37122 22276 37126 22332
rect 37062 22272 37126 22276
rect 37142 22332 37206 22336
rect 37142 22276 37146 22332
rect 37146 22276 37202 22332
rect 37202 22276 37206 22332
rect 37142 22272 37206 22276
rect 37222 22332 37286 22336
rect 37222 22276 37226 22332
rect 37226 22276 37282 22332
rect 37282 22276 37286 22332
rect 37222 22272 37286 22276
rect 37302 22332 37366 22336
rect 37302 22276 37306 22332
rect 37306 22276 37362 22332
rect 37362 22276 37366 22332
rect 37302 22272 37366 22276
rect 51506 22332 51570 22336
rect 51506 22276 51510 22332
rect 51510 22276 51566 22332
rect 51566 22276 51570 22332
rect 51506 22272 51570 22276
rect 51586 22332 51650 22336
rect 51586 22276 51590 22332
rect 51590 22276 51646 22332
rect 51646 22276 51650 22332
rect 51586 22272 51650 22276
rect 51666 22332 51730 22336
rect 51666 22276 51670 22332
rect 51670 22276 51726 22332
rect 51726 22276 51730 22332
rect 51666 22272 51730 22276
rect 51746 22332 51810 22336
rect 51746 22276 51750 22332
rect 51750 22276 51806 22332
rect 51806 22276 51810 22332
rect 51746 22272 51810 22276
rect 15396 21788 15460 21792
rect 15396 21732 15400 21788
rect 15400 21732 15456 21788
rect 15456 21732 15460 21788
rect 15396 21728 15460 21732
rect 15476 21788 15540 21792
rect 15476 21732 15480 21788
rect 15480 21732 15536 21788
rect 15536 21732 15540 21788
rect 15476 21728 15540 21732
rect 15556 21788 15620 21792
rect 15556 21732 15560 21788
rect 15560 21732 15616 21788
rect 15616 21732 15620 21788
rect 15556 21728 15620 21732
rect 15636 21788 15700 21792
rect 15636 21732 15640 21788
rect 15640 21732 15696 21788
rect 15696 21732 15700 21788
rect 15636 21728 15700 21732
rect 29840 21788 29904 21792
rect 29840 21732 29844 21788
rect 29844 21732 29900 21788
rect 29900 21732 29904 21788
rect 29840 21728 29904 21732
rect 29920 21788 29984 21792
rect 29920 21732 29924 21788
rect 29924 21732 29980 21788
rect 29980 21732 29984 21788
rect 29920 21728 29984 21732
rect 30000 21788 30064 21792
rect 30000 21732 30004 21788
rect 30004 21732 30060 21788
rect 30060 21732 30064 21788
rect 30000 21728 30064 21732
rect 30080 21788 30144 21792
rect 30080 21732 30084 21788
rect 30084 21732 30140 21788
rect 30140 21732 30144 21788
rect 30080 21728 30144 21732
rect 44284 21788 44348 21792
rect 44284 21732 44288 21788
rect 44288 21732 44344 21788
rect 44344 21732 44348 21788
rect 44284 21728 44348 21732
rect 44364 21788 44428 21792
rect 44364 21732 44368 21788
rect 44368 21732 44424 21788
rect 44424 21732 44428 21788
rect 44364 21728 44428 21732
rect 44444 21788 44508 21792
rect 44444 21732 44448 21788
rect 44448 21732 44504 21788
rect 44504 21732 44508 21788
rect 44444 21728 44508 21732
rect 44524 21788 44588 21792
rect 44524 21732 44528 21788
rect 44528 21732 44584 21788
rect 44584 21732 44588 21788
rect 44524 21728 44588 21732
rect 58728 21788 58792 21792
rect 58728 21732 58732 21788
rect 58732 21732 58788 21788
rect 58788 21732 58792 21788
rect 58728 21728 58792 21732
rect 58808 21788 58872 21792
rect 58808 21732 58812 21788
rect 58812 21732 58868 21788
rect 58868 21732 58872 21788
rect 58808 21728 58872 21732
rect 58888 21788 58952 21792
rect 58888 21732 58892 21788
rect 58892 21732 58948 21788
rect 58948 21732 58952 21788
rect 58888 21728 58952 21732
rect 58968 21788 59032 21792
rect 58968 21732 58972 21788
rect 58972 21732 59028 21788
rect 59028 21732 59032 21788
rect 58968 21728 59032 21732
rect 8174 21244 8238 21248
rect 8174 21188 8178 21244
rect 8178 21188 8234 21244
rect 8234 21188 8238 21244
rect 8174 21184 8238 21188
rect 8254 21244 8318 21248
rect 8254 21188 8258 21244
rect 8258 21188 8314 21244
rect 8314 21188 8318 21244
rect 8254 21184 8318 21188
rect 8334 21244 8398 21248
rect 8334 21188 8338 21244
rect 8338 21188 8394 21244
rect 8394 21188 8398 21244
rect 8334 21184 8398 21188
rect 8414 21244 8478 21248
rect 8414 21188 8418 21244
rect 8418 21188 8474 21244
rect 8474 21188 8478 21244
rect 8414 21184 8478 21188
rect 22618 21244 22682 21248
rect 22618 21188 22622 21244
rect 22622 21188 22678 21244
rect 22678 21188 22682 21244
rect 22618 21184 22682 21188
rect 22698 21244 22762 21248
rect 22698 21188 22702 21244
rect 22702 21188 22758 21244
rect 22758 21188 22762 21244
rect 22698 21184 22762 21188
rect 22778 21244 22842 21248
rect 22778 21188 22782 21244
rect 22782 21188 22838 21244
rect 22838 21188 22842 21244
rect 22778 21184 22842 21188
rect 22858 21244 22922 21248
rect 22858 21188 22862 21244
rect 22862 21188 22918 21244
rect 22918 21188 22922 21244
rect 22858 21184 22922 21188
rect 37062 21244 37126 21248
rect 37062 21188 37066 21244
rect 37066 21188 37122 21244
rect 37122 21188 37126 21244
rect 37062 21184 37126 21188
rect 37142 21244 37206 21248
rect 37142 21188 37146 21244
rect 37146 21188 37202 21244
rect 37202 21188 37206 21244
rect 37142 21184 37206 21188
rect 37222 21244 37286 21248
rect 37222 21188 37226 21244
rect 37226 21188 37282 21244
rect 37282 21188 37286 21244
rect 37222 21184 37286 21188
rect 37302 21244 37366 21248
rect 37302 21188 37306 21244
rect 37306 21188 37362 21244
rect 37362 21188 37366 21244
rect 37302 21184 37366 21188
rect 51506 21244 51570 21248
rect 51506 21188 51510 21244
rect 51510 21188 51566 21244
rect 51566 21188 51570 21244
rect 51506 21184 51570 21188
rect 51586 21244 51650 21248
rect 51586 21188 51590 21244
rect 51590 21188 51646 21244
rect 51646 21188 51650 21244
rect 51586 21184 51650 21188
rect 51666 21244 51730 21248
rect 51666 21188 51670 21244
rect 51670 21188 51726 21244
rect 51726 21188 51730 21244
rect 51666 21184 51730 21188
rect 51746 21244 51810 21248
rect 51746 21188 51750 21244
rect 51750 21188 51806 21244
rect 51806 21188 51810 21244
rect 51746 21184 51810 21188
rect 15396 20700 15460 20704
rect 15396 20644 15400 20700
rect 15400 20644 15456 20700
rect 15456 20644 15460 20700
rect 15396 20640 15460 20644
rect 15476 20700 15540 20704
rect 15476 20644 15480 20700
rect 15480 20644 15536 20700
rect 15536 20644 15540 20700
rect 15476 20640 15540 20644
rect 15556 20700 15620 20704
rect 15556 20644 15560 20700
rect 15560 20644 15616 20700
rect 15616 20644 15620 20700
rect 15556 20640 15620 20644
rect 15636 20700 15700 20704
rect 15636 20644 15640 20700
rect 15640 20644 15696 20700
rect 15696 20644 15700 20700
rect 15636 20640 15700 20644
rect 29840 20700 29904 20704
rect 29840 20644 29844 20700
rect 29844 20644 29900 20700
rect 29900 20644 29904 20700
rect 29840 20640 29904 20644
rect 29920 20700 29984 20704
rect 29920 20644 29924 20700
rect 29924 20644 29980 20700
rect 29980 20644 29984 20700
rect 29920 20640 29984 20644
rect 30000 20700 30064 20704
rect 30000 20644 30004 20700
rect 30004 20644 30060 20700
rect 30060 20644 30064 20700
rect 30000 20640 30064 20644
rect 30080 20700 30144 20704
rect 30080 20644 30084 20700
rect 30084 20644 30140 20700
rect 30140 20644 30144 20700
rect 30080 20640 30144 20644
rect 44284 20700 44348 20704
rect 44284 20644 44288 20700
rect 44288 20644 44344 20700
rect 44344 20644 44348 20700
rect 44284 20640 44348 20644
rect 44364 20700 44428 20704
rect 44364 20644 44368 20700
rect 44368 20644 44424 20700
rect 44424 20644 44428 20700
rect 44364 20640 44428 20644
rect 44444 20700 44508 20704
rect 44444 20644 44448 20700
rect 44448 20644 44504 20700
rect 44504 20644 44508 20700
rect 44444 20640 44508 20644
rect 44524 20700 44588 20704
rect 44524 20644 44528 20700
rect 44528 20644 44584 20700
rect 44584 20644 44588 20700
rect 44524 20640 44588 20644
rect 58728 20700 58792 20704
rect 58728 20644 58732 20700
rect 58732 20644 58788 20700
rect 58788 20644 58792 20700
rect 58728 20640 58792 20644
rect 58808 20700 58872 20704
rect 58808 20644 58812 20700
rect 58812 20644 58868 20700
rect 58868 20644 58872 20700
rect 58808 20640 58872 20644
rect 58888 20700 58952 20704
rect 58888 20644 58892 20700
rect 58892 20644 58948 20700
rect 58948 20644 58952 20700
rect 58888 20640 58952 20644
rect 58968 20700 59032 20704
rect 58968 20644 58972 20700
rect 58972 20644 59028 20700
rect 59028 20644 59032 20700
rect 58968 20640 59032 20644
rect 8174 20156 8238 20160
rect 8174 20100 8178 20156
rect 8178 20100 8234 20156
rect 8234 20100 8238 20156
rect 8174 20096 8238 20100
rect 8254 20156 8318 20160
rect 8254 20100 8258 20156
rect 8258 20100 8314 20156
rect 8314 20100 8318 20156
rect 8254 20096 8318 20100
rect 8334 20156 8398 20160
rect 8334 20100 8338 20156
rect 8338 20100 8394 20156
rect 8394 20100 8398 20156
rect 8334 20096 8398 20100
rect 8414 20156 8478 20160
rect 8414 20100 8418 20156
rect 8418 20100 8474 20156
rect 8474 20100 8478 20156
rect 8414 20096 8478 20100
rect 22618 20156 22682 20160
rect 22618 20100 22622 20156
rect 22622 20100 22678 20156
rect 22678 20100 22682 20156
rect 22618 20096 22682 20100
rect 22698 20156 22762 20160
rect 22698 20100 22702 20156
rect 22702 20100 22758 20156
rect 22758 20100 22762 20156
rect 22698 20096 22762 20100
rect 22778 20156 22842 20160
rect 22778 20100 22782 20156
rect 22782 20100 22838 20156
rect 22838 20100 22842 20156
rect 22778 20096 22842 20100
rect 22858 20156 22922 20160
rect 22858 20100 22862 20156
rect 22862 20100 22918 20156
rect 22918 20100 22922 20156
rect 22858 20096 22922 20100
rect 37062 20156 37126 20160
rect 37062 20100 37066 20156
rect 37066 20100 37122 20156
rect 37122 20100 37126 20156
rect 37062 20096 37126 20100
rect 37142 20156 37206 20160
rect 37142 20100 37146 20156
rect 37146 20100 37202 20156
rect 37202 20100 37206 20156
rect 37142 20096 37206 20100
rect 37222 20156 37286 20160
rect 37222 20100 37226 20156
rect 37226 20100 37282 20156
rect 37282 20100 37286 20156
rect 37222 20096 37286 20100
rect 37302 20156 37366 20160
rect 37302 20100 37306 20156
rect 37306 20100 37362 20156
rect 37362 20100 37366 20156
rect 37302 20096 37366 20100
rect 51506 20156 51570 20160
rect 51506 20100 51510 20156
rect 51510 20100 51566 20156
rect 51566 20100 51570 20156
rect 51506 20096 51570 20100
rect 51586 20156 51650 20160
rect 51586 20100 51590 20156
rect 51590 20100 51646 20156
rect 51646 20100 51650 20156
rect 51586 20096 51650 20100
rect 51666 20156 51730 20160
rect 51666 20100 51670 20156
rect 51670 20100 51726 20156
rect 51726 20100 51730 20156
rect 51666 20096 51730 20100
rect 51746 20156 51810 20160
rect 51746 20100 51750 20156
rect 51750 20100 51806 20156
rect 51806 20100 51810 20156
rect 51746 20096 51810 20100
rect 15396 19612 15460 19616
rect 15396 19556 15400 19612
rect 15400 19556 15456 19612
rect 15456 19556 15460 19612
rect 15396 19552 15460 19556
rect 15476 19612 15540 19616
rect 15476 19556 15480 19612
rect 15480 19556 15536 19612
rect 15536 19556 15540 19612
rect 15476 19552 15540 19556
rect 15556 19612 15620 19616
rect 15556 19556 15560 19612
rect 15560 19556 15616 19612
rect 15616 19556 15620 19612
rect 15556 19552 15620 19556
rect 15636 19612 15700 19616
rect 15636 19556 15640 19612
rect 15640 19556 15696 19612
rect 15696 19556 15700 19612
rect 15636 19552 15700 19556
rect 29840 19612 29904 19616
rect 29840 19556 29844 19612
rect 29844 19556 29900 19612
rect 29900 19556 29904 19612
rect 29840 19552 29904 19556
rect 29920 19612 29984 19616
rect 29920 19556 29924 19612
rect 29924 19556 29980 19612
rect 29980 19556 29984 19612
rect 29920 19552 29984 19556
rect 30000 19612 30064 19616
rect 30000 19556 30004 19612
rect 30004 19556 30060 19612
rect 30060 19556 30064 19612
rect 30000 19552 30064 19556
rect 30080 19612 30144 19616
rect 30080 19556 30084 19612
rect 30084 19556 30140 19612
rect 30140 19556 30144 19612
rect 30080 19552 30144 19556
rect 44284 19612 44348 19616
rect 44284 19556 44288 19612
rect 44288 19556 44344 19612
rect 44344 19556 44348 19612
rect 44284 19552 44348 19556
rect 44364 19612 44428 19616
rect 44364 19556 44368 19612
rect 44368 19556 44424 19612
rect 44424 19556 44428 19612
rect 44364 19552 44428 19556
rect 44444 19612 44508 19616
rect 44444 19556 44448 19612
rect 44448 19556 44504 19612
rect 44504 19556 44508 19612
rect 44444 19552 44508 19556
rect 44524 19612 44588 19616
rect 44524 19556 44528 19612
rect 44528 19556 44584 19612
rect 44584 19556 44588 19612
rect 44524 19552 44588 19556
rect 58728 19612 58792 19616
rect 58728 19556 58732 19612
rect 58732 19556 58788 19612
rect 58788 19556 58792 19612
rect 58728 19552 58792 19556
rect 58808 19612 58872 19616
rect 58808 19556 58812 19612
rect 58812 19556 58868 19612
rect 58868 19556 58872 19612
rect 58808 19552 58872 19556
rect 58888 19612 58952 19616
rect 58888 19556 58892 19612
rect 58892 19556 58948 19612
rect 58948 19556 58952 19612
rect 58888 19552 58952 19556
rect 58968 19612 59032 19616
rect 58968 19556 58972 19612
rect 58972 19556 59028 19612
rect 59028 19556 59032 19612
rect 58968 19552 59032 19556
rect 8174 19068 8238 19072
rect 8174 19012 8178 19068
rect 8178 19012 8234 19068
rect 8234 19012 8238 19068
rect 8174 19008 8238 19012
rect 8254 19068 8318 19072
rect 8254 19012 8258 19068
rect 8258 19012 8314 19068
rect 8314 19012 8318 19068
rect 8254 19008 8318 19012
rect 8334 19068 8398 19072
rect 8334 19012 8338 19068
rect 8338 19012 8394 19068
rect 8394 19012 8398 19068
rect 8334 19008 8398 19012
rect 8414 19068 8478 19072
rect 8414 19012 8418 19068
rect 8418 19012 8474 19068
rect 8474 19012 8478 19068
rect 8414 19008 8478 19012
rect 22618 19068 22682 19072
rect 22618 19012 22622 19068
rect 22622 19012 22678 19068
rect 22678 19012 22682 19068
rect 22618 19008 22682 19012
rect 22698 19068 22762 19072
rect 22698 19012 22702 19068
rect 22702 19012 22758 19068
rect 22758 19012 22762 19068
rect 22698 19008 22762 19012
rect 22778 19068 22842 19072
rect 22778 19012 22782 19068
rect 22782 19012 22838 19068
rect 22838 19012 22842 19068
rect 22778 19008 22842 19012
rect 22858 19068 22922 19072
rect 22858 19012 22862 19068
rect 22862 19012 22918 19068
rect 22918 19012 22922 19068
rect 22858 19008 22922 19012
rect 37062 19068 37126 19072
rect 37062 19012 37066 19068
rect 37066 19012 37122 19068
rect 37122 19012 37126 19068
rect 37062 19008 37126 19012
rect 37142 19068 37206 19072
rect 37142 19012 37146 19068
rect 37146 19012 37202 19068
rect 37202 19012 37206 19068
rect 37142 19008 37206 19012
rect 37222 19068 37286 19072
rect 37222 19012 37226 19068
rect 37226 19012 37282 19068
rect 37282 19012 37286 19068
rect 37222 19008 37286 19012
rect 37302 19068 37366 19072
rect 37302 19012 37306 19068
rect 37306 19012 37362 19068
rect 37362 19012 37366 19068
rect 37302 19008 37366 19012
rect 51506 19068 51570 19072
rect 51506 19012 51510 19068
rect 51510 19012 51566 19068
rect 51566 19012 51570 19068
rect 51506 19008 51570 19012
rect 51586 19068 51650 19072
rect 51586 19012 51590 19068
rect 51590 19012 51646 19068
rect 51646 19012 51650 19068
rect 51586 19008 51650 19012
rect 51666 19068 51730 19072
rect 51666 19012 51670 19068
rect 51670 19012 51726 19068
rect 51726 19012 51730 19068
rect 51666 19008 51730 19012
rect 51746 19068 51810 19072
rect 51746 19012 51750 19068
rect 51750 19012 51806 19068
rect 51806 19012 51810 19068
rect 51746 19008 51810 19012
rect 15396 18524 15460 18528
rect 15396 18468 15400 18524
rect 15400 18468 15456 18524
rect 15456 18468 15460 18524
rect 15396 18464 15460 18468
rect 15476 18524 15540 18528
rect 15476 18468 15480 18524
rect 15480 18468 15536 18524
rect 15536 18468 15540 18524
rect 15476 18464 15540 18468
rect 15556 18524 15620 18528
rect 15556 18468 15560 18524
rect 15560 18468 15616 18524
rect 15616 18468 15620 18524
rect 15556 18464 15620 18468
rect 15636 18524 15700 18528
rect 15636 18468 15640 18524
rect 15640 18468 15696 18524
rect 15696 18468 15700 18524
rect 15636 18464 15700 18468
rect 29840 18524 29904 18528
rect 29840 18468 29844 18524
rect 29844 18468 29900 18524
rect 29900 18468 29904 18524
rect 29840 18464 29904 18468
rect 29920 18524 29984 18528
rect 29920 18468 29924 18524
rect 29924 18468 29980 18524
rect 29980 18468 29984 18524
rect 29920 18464 29984 18468
rect 30000 18524 30064 18528
rect 30000 18468 30004 18524
rect 30004 18468 30060 18524
rect 30060 18468 30064 18524
rect 30000 18464 30064 18468
rect 30080 18524 30144 18528
rect 30080 18468 30084 18524
rect 30084 18468 30140 18524
rect 30140 18468 30144 18524
rect 30080 18464 30144 18468
rect 44284 18524 44348 18528
rect 44284 18468 44288 18524
rect 44288 18468 44344 18524
rect 44344 18468 44348 18524
rect 44284 18464 44348 18468
rect 44364 18524 44428 18528
rect 44364 18468 44368 18524
rect 44368 18468 44424 18524
rect 44424 18468 44428 18524
rect 44364 18464 44428 18468
rect 44444 18524 44508 18528
rect 44444 18468 44448 18524
rect 44448 18468 44504 18524
rect 44504 18468 44508 18524
rect 44444 18464 44508 18468
rect 44524 18524 44588 18528
rect 44524 18468 44528 18524
rect 44528 18468 44584 18524
rect 44584 18468 44588 18524
rect 44524 18464 44588 18468
rect 58728 18524 58792 18528
rect 58728 18468 58732 18524
rect 58732 18468 58788 18524
rect 58788 18468 58792 18524
rect 58728 18464 58792 18468
rect 58808 18524 58872 18528
rect 58808 18468 58812 18524
rect 58812 18468 58868 18524
rect 58868 18468 58872 18524
rect 58808 18464 58872 18468
rect 58888 18524 58952 18528
rect 58888 18468 58892 18524
rect 58892 18468 58948 18524
rect 58948 18468 58952 18524
rect 58888 18464 58952 18468
rect 58968 18524 59032 18528
rect 58968 18468 58972 18524
rect 58972 18468 59028 18524
rect 59028 18468 59032 18524
rect 58968 18464 59032 18468
rect 8174 17980 8238 17984
rect 8174 17924 8178 17980
rect 8178 17924 8234 17980
rect 8234 17924 8238 17980
rect 8174 17920 8238 17924
rect 8254 17980 8318 17984
rect 8254 17924 8258 17980
rect 8258 17924 8314 17980
rect 8314 17924 8318 17980
rect 8254 17920 8318 17924
rect 8334 17980 8398 17984
rect 8334 17924 8338 17980
rect 8338 17924 8394 17980
rect 8394 17924 8398 17980
rect 8334 17920 8398 17924
rect 8414 17980 8478 17984
rect 8414 17924 8418 17980
rect 8418 17924 8474 17980
rect 8474 17924 8478 17980
rect 8414 17920 8478 17924
rect 22618 17980 22682 17984
rect 22618 17924 22622 17980
rect 22622 17924 22678 17980
rect 22678 17924 22682 17980
rect 22618 17920 22682 17924
rect 22698 17980 22762 17984
rect 22698 17924 22702 17980
rect 22702 17924 22758 17980
rect 22758 17924 22762 17980
rect 22698 17920 22762 17924
rect 22778 17980 22842 17984
rect 22778 17924 22782 17980
rect 22782 17924 22838 17980
rect 22838 17924 22842 17980
rect 22778 17920 22842 17924
rect 22858 17980 22922 17984
rect 22858 17924 22862 17980
rect 22862 17924 22918 17980
rect 22918 17924 22922 17980
rect 22858 17920 22922 17924
rect 37062 17980 37126 17984
rect 37062 17924 37066 17980
rect 37066 17924 37122 17980
rect 37122 17924 37126 17980
rect 37062 17920 37126 17924
rect 37142 17980 37206 17984
rect 37142 17924 37146 17980
rect 37146 17924 37202 17980
rect 37202 17924 37206 17980
rect 37142 17920 37206 17924
rect 37222 17980 37286 17984
rect 37222 17924 37226 17980
rect 37226 17924 37282 17980
rect 37282 17924 37286 17980
rect 37222 17920 37286 17924
rect 37302 17980 37366 17984
rect 37302 17924 37306 17980
rect 37306 17924 37362 17980
rect 37362 17924 37366 17980
rect 37302 17920 37366 17924
rect 51506 17980 51570 17984
rect 51506 17924 51510 17980
rect 51510 17924 51566 17980
rect 51566 17924 51570 17980
rect 51506 17920 51570 17924
rect 51586 17980 51650 17984
rect 51586 17924 51590 17980
rect 51590 17924 51646 17980
rect 51646 17924 51650 17980
rect 51586 17920 51650 17924
rect 51666 17980 51730 17984
rect 51666 17924 51670 17980
rect 51670 17924 51726 17980
rect 51726 17924 51730 17980
rect 51666 17920 51730 17924
rect 51746 17980 51810 17984
rect 51746 17924 51750 17980
rect 51750 17924 51806 17980
rect 51806 17924 51810 17980
rect 51746 17920 51810 17924
rect 15396 17436 15460 17440
rect 15396 17380 15400 17436
rect 15400 17380 15456 17436
rect 15456 17380 15460 17436
rect 15396 17376 15460 17380
rect 15476 17436 15540 17440
rect 15476 17380 15480 17436
rect 15480 17380 15536 17436
rect 15536 17380 15540 17436
rect 15476 17376 15540 17380
rect 15556 17436 15620 17440
rect 15556 17380 15560 17436
rect 15560 17380 15616 17436
rect 15616 17380 15620 17436
rect 15556 17376 15620 17380
rect 15636 17436 15700 17440
rect 15636 17380 15640 17436
rect 15640 17380 15696 17436
rect 15696 17380 15700 17436
rect 15636 17376 15700 17380
rect 29840 17436 29904 17440
rect 29840 17380 29844 17436
rect 29844 17380 29900 17436
rect 29900 17380 29904 17436
rect 29840 17376 29904 17380
rect 29920 17436 29984 17440
rect 29920 17380 29924 17436
rect 29924 17380 29980 17436
rect 29980 17380 29984 17436
rect 29920 17376 29984 17380
rect 30000 17436 30064 17440
rect 30000 17380 30004 17436
rect 30004 17380 30060 17436
rect 30060 17380 30064 17436
rect 30000 17376 30064 17380
rect 30080 17436 30144 17440
rect 30080 17380 30084 17436
rect 30084 17380 30140 17436
rect 30140 17380 30144 17436
rect 30080 17376 30144 17380
rect 44284 17436 44348 17440
rect 44284 17380 44288 17436
rect 44288 17380 44344 17436
rect 44344 17380 44348 17436
rect 44284 17376 44348 17380
rect 44364 17436 44428 17440
rect 44364 17380 44368 17436
rect 44368 17380 44424 17436
rect 44424 17380 44428 17436
rect 44364 17376 44428 17380
rect 44444 17436 44508 17440
rect 44444 17380 44448 17436
rect 44448 17380 44504 17436
rect 44504 17380 44508 17436
rect 44444 17376 44508 17380
rect 44524 17436 44588 17440
rect 44524 17380 44528 17436
rect 44528 17380 44584 17436
rect 44584 17380 44588 17436
rect 44524 17376 44588 17380
rect 58728 17436 58792 17440
rect 58728 17380 58732 17436
rect 58732 17380 58788 17436
rect 58788 17380 58792 17436
rect 58728 17376 58792 17380
rect 58808 17436 58872 17440
rect 58808 17380 58812 17436
rect 58812 17380 58868 17436
rect 58868 17380 58872 17436
rect 58808 17376 58872 17380
rect 58888 17436 58952 17440
rect 58888 17380 58892 17436
rect 58892 17380 58948 17436
rect 58948 17380 58952 17436
rect 58888 17376 58952 17380
rect 58968 17436 59032 17440
rect 58968 17380 58972 17436
rect 58972 17380 59028 17436
rect 59028 17380 59032 17436
rect 58968 17376 59032 17380
rect 8174 16892 8238 16896
rect 8174 16836 8178 16892
rect 8178 16836 8234 16892
rect 8234 16836 8238 16892
rect 8174 16832 8238 16836
rect 8254 16892 8318 16896
rect 8254 16836 8258 16892
rect 8258 16836 8314 16892
rect 8314 16836 8318 16892
rect 8254 16832 8318 16836
rect 8334 16892 8398 16896
rect 8334 16836 8338 16892
rect 8338 16836 8394 16892
rect 8394 16836 8398 16892
rect 8334 16832 8398 16836
rect 8414 16892 8478 16896
rect 8414 16836 8418 16892
rect 8418 16836 8474 16892
rect 8474 16836 8478 16892
rect 8414 16832 8478 16836
rect 22618 16892 22682 16896
rect 22618 16836 22622 16892
rect 22622 16836 22678 16892
rect 22678 16836 22682 16892
rect 22618 16832 22682 16836
rect 22698 16892 22762 16896
rect 22698 16836 22702 16892
rect 22702 16836 22758 16892
rect 22758 16836 22762 16892
rect 22698 16832 22762 16836
rect 22778 16892 22842 16896
rect 22778 16836 22782 16892
rect 22782 16836 22838 16892
rect 22838 16836 22842 16892
rect 22778 16832 22842 16836
rect 22858 16892 22922 16896
rect 22858 16836 22862 16892
rect 22862 16836 22918 16892
rect 22918 16836 22922 16892
rect 22858 16832 22922 16836
rect 37062 16892 37126 16896
rect 37062 16836 37066 16892
rect 37066 16836 37122 16892
rect 37122 16836 37126 16892
rect 37062 16832 37126 16836
rect 37142 16892 37206 16896
rect 37142 16836 37146 16892
rect 37146 16836 37202 16892
rect 37202 16836 37206 16892
rect 37142 16832 37206 16836
rect 37222 16892 37286 16896
rect 37222 16836 37226 16892
rect 37226 16836 37282 16892
rect 37282 16836 37286 16892
rect 37222 16832 37286 16836
rect 37302 16892 37366 16896
rect 37302 16836 37306 16892
rect 37306 16836 37362 16892
rect 37362 16836 37366 16892
rect 37302 16832 37366 16836
rect 51506 16892 51570 16896
rect 51506 16836 51510 16892
rect 51510 16836 51566 16892
rect 51566 16836 51570 16892
rect 51506 16832 51570 16836
rect 51586 16892 51650 16896
rect 51586 16836 51590 16892
rect 51590 16836 51646 16892
rect 51646 16836 51650 16892
rect 51586 16832 51650 16836
rect 51666 16892 51730 16896
rect 51666 16836 51670 16892
rect 51670 16836 51726 16892
rect 51726 16836 51730 16892
rect 51666 16832 51730 16836
rect 51746 16892 51810 16896
rect 51746 16836 51750 16892
rect 51750 16836 51806 16892
rect 51806 16836 51810 16892
rect 51746 16832 51810 16836
rect 15396 16348 15460 16352
rect 15396 16292 15400 16348
rect 15400 16292 15456 16348
rect 15456 16292 15460 16348
rect 15396 16288 15460 16292
rect 15476 16348 15540 16352
rect 15476 16292 15480 16348
rect 15480 16292 15536 16348
rect 15536 16292 15540 16348
rect 15476 16288 15540 16292
rect 15556 16348 15620 16352
rect 15556 16292 15560 16348
rect 15560 16292 15616 16348
rect 15616 16292 15620 16348
rect 15556 16288 15620 16292
rect 15636 16348 15700 16352
rect 15636 16292 15640 16348
rect 15640 16292 15696 16348
rect 15696 16292 15700 16348
rect 15636 16288 15700 16292
rect 29840 16348 29904 16352
rect 29840 16292 29844 16348
rect 29844 16292 29900 16348
rect 29900 16292 29904 16348
rect 29840 16288 29904 16292
rect 29920 16348 29984 16352
rect 29920 16292 29924 16348
rect 29924 16292 29980 16348
rect 29980 16292 29984 16348
rect 29920 16288 29984 16292
rect 30000 16348 30064 16352
rect 30000 16292 30004 16348
rect 30004 16292 30060 16348
rect 30060 16292 30064 16348
rect 30000 16288 30064 16292
rect 30080 16348 30144 16352
rect 30080 16292 30084 16348
rect 30084 16292 30140 16348
rect 30140 16292 30144 16348
rect 30080 16288 30144 16292
rect 44284 16348 44348 16352
rect 44284 16292 44288 16348
rect 44288 16292 44344 16348
rect 44344 16292 44348 16348
rect 44284 16288 44348 16292
rect 44364 16348 44428 16352
rect 44364 16292 44368 16348
rect 44368 16292 44424 16348
rect 44424 16292 44428 16348
rect 44364 16288 44428 16292
rect 44444 16348 44508 16352
rect 44444 16292 44448 16348
rect 44448 16292 44504 16348
rect 44504 16292 44508 16348
rect 44444 16288 44508 16292
rect 44524 16348 44588 16352
rect 44524 16292 44528 16348
rect 44528 16292 44584 16348
rect 44584 16292 44588 16348
rect 44524 16288 44588 16292
rect 58728 16348 58792 16352
rect 58728 16292 58732 16348
rect 58732 16292 58788 16348
rect 58788 16292 58792 16348
rect 58728 16288 58792 16292
rect 58808 16348 58872 16352
rect 58808 16292 58812 16348
rect 58812 16292 58868 16348
rect 58868 16292 58872 16348
rect 58808 16288 58872 16292
rect 58888 16348 58952 16352
rect 58888 16292 58892 16348
rect 58892 16292 58948 16348
rect 58948 16292 58952 16348
rect 58888 16288 58952 16292
rect 58968 16348 59032 16352
rect 58968 16292 58972 16348
rect 58972 16292 59028 16348
rect 59028 16292 59032 16348
rect 58968 16288 59032 16292
rect 8174 15804 8238 15808
rect 8174 15748 8178 15804
rect 8178 15748 8234 15804
rect 8234 15748 8238 15804
rect 8174 15744 8238 15748
rect 8254 15804 8318 15808
rect 8254 15748 8258 15804
rect 8258 15748 8314 15804
rect 8314 15748 8318 15804
rect 8254 15744 8318 15748
rect 8334 15804 8398 15808
rect 8334 15748 8338 15804
rect 8338 15748 8394 15804
rect 8394 15748 8398 15804
rect 8334 15744 8398 15748
rect 8414 15804 8478 15808
rect 8414 15748 8418 15804
rect 8418 15748 8474 15804
rect 8474 15748 8478 15804
rect 8414 15744 8478 15748
rect 22618 15804 22682 15808
rect 22618 15748 22622 15804
rect 22622 15748 22678 15804
rect 22678 15748 22682 15804
rect 22618 15744 22682 15748
rect 22698 15804 22762 15808
rect 22698 15748 22702 15804
rect 22702 15748 22758 15804
rect 22758 15748 22762 15804
rect 22698 15744 22762 15748
rect 22778 15804 22842 15808
rect 22778 15748 22782 15804
rect 22782 15748 22838 15804
rect 22838 15748 22842 15804
rect 22778 15744 22842 15748
rect 22858 15804 22922 15808
rect 22858 15748 22862 15804
rect 22862 15748 22918 15804
rect 22918 15748 22922 15804
rect 22858 15744 22922 15748
rect 37062 15804 37126 15808
rect 37062 15748 37066 15804
rect 37066 15748 37122 15804
rect 37122 15748 37126 15804
rect 37062 15744 37126 15748
rect 37142 15804 37206 15808
rect 37142 15748 37146 15804
rect 37146 15748 37202 15804
rect 37202 15748 37206 15804
rect 37142 15744 37206 15748
rect 37222 15804 37286 15808
rect 37222 15748 37226 15804
rect 37226 15748 37282 15804
rect 37282 15748 37286 15804
rect 37222 15744 37286 15748
rect 37302 15804 37366 15808
rect 37302 15748 37306 15804
rect 37306 15748 37362 15804
rect 37362 15748 37366 15804
rect 37302 15744 37366 15748
rect 51506 15804 51570 15808
rect 51506 15748 51510 15804
rect 51510 15748 51566 15804
rect 51566 15748 51570 15804
rect 51506 15744 51570 15748
rect 51586 15804 51650 15808
rect 51586 15748 51590 15804
rect 51590 15748 51646 15804
rect 51646 15748 51650 15804
rect 51586 15744 51650 15748
rect 51666 15804 51730 15808
rect 51666 15748 51670 15804
rect 51670 15748 51726 15804
rect 51726 15748 51730 15804
rect 51666 15744 51730 15748
rect 51746 15804 51810 15808
rect 51746 15748 51750 15804
rect 51750 15748 51806 15804
rect 51806 15748 51810 15804
rect 51746 15744 51810 15748
rect 15396 15260 15460 15264
rect 15396 15204 15400 15260
rect 15400 15204 15456 15260
rect 15456 15204 15460 15260
rect 15396 15200 15460 15204
rect 15476 15260 15540 15264
rect 15476 15204 15480 15260
rect 15480 15204 15536 15260
rect 15536 15204 15540 15260
rect 15476 15200 15540 15204
rect 15556 15260 15620 15264
rect 15556 15204 15560 15260
rect 15560 15204 15616 15260
rect 15616 15204 15620 15260
rect 15556 15200 15620 15204
rect 15636 15260 15700 15264
rect 15636 15204 15640 15260
rect 15640 15204 15696 15260
rect 15696 15204 15700 15260
rect 15636 15200 15700 15204
rect 29840 15260 29904 15264
rect 29840 15204 29844 15260
rect 29844 15204 29900 15260
rect 29900 15204 29904 15260
rect 29840 15200 29904 15204
rect 29920 15260 29984 15264
rect 29920 15204 29924 15260
rect 29924 15204 29980 15260
rect 29980 15204 29984 15260
rect 29920 15200 29984 15204
rect 30000 15260 30064 15264
rect 30000 15204 30004 15260
rect 30004 15204 30060 15260
rect 30060 15204 30064 15260
rect 30000 15200 30064 15204
rect 30080 15260 30144 15264
rect 30080 15204 30084 15260
rect 30084 15204 30140 15260
rect 30140 15204 30144 15260
rect 30080 15200 30144 15204
rect 44284 15260 44348 15264
rect 44284 15204 44288 15260
rect 44288 15204 44344 15260
rect 44344 15204 44348 15260
rect 44284 15200 44348 15204
rect 44364 15260 44428 15264
rect 44364 15204 44368 15260
rect 44368 15204 44424 15260
rect 44424 15204 44428 15260
rect 44364 15200 44428 15204
rect 44444 15260 44508 15264
rect 44444 15204 44448 15260
rect 44448 15204 44504 15260
rect 44504 15204 44508 15260
rect 44444 15200 44508 15204
rect 44524 15260 44588 15264
rect 44524 15204 44528 15260
rect 44528 15204 44584 15260
rect 44584 15204 44588 15260
rect 44524 15200 44588 15204
rect 58728 15260 58792 15264
rect 58728 15204 58732 15260
rect 58732 15204 58788 15260
rect 58788 15204 58792 15260
rect 58728 15200 58792 15204
rect 58808 15260 58872 15264
rect 58808 15204 58812 15260
rect 58812 15204 58868 15260
rect 58868 15204 58872 15260
rect 58808 15200 58872 15204
rect 58888 15260 58952 15264
rect 58888 15204 58892 15260
rect 58892 15204 58948 15260
rect 58948 15204 58952 15260
rect 58888 15200 58952 15204
rect 58968 15260 59032 15264
rect 58968 15204 58972 15260
rect 58972 15204 59028 15260
rect 59028 15204 59032 15260
rect 58968 15200 59032 15204
rect 8174 14716 8238 14720
rect 8174 14660 8178 14716
rect 8178 14660 8234 14716
rect 8234 14660 8238 14716
rect 8174 14656 8238 14660
rect 8254 14716 8318 14720
rect 8254 14660 8258 14716
rect 8258 14660 8314 14716
rect 8314 14660 8318 14716
rect 8254 14656 8318 14660
rect 8334 14716 8398 14720
rect 8334 14660 8338 14716
rect 8338 14660 8394 14716
rect 8394 14660 8398 14716
rect 8334 14656 8398 14660
rect 8414 14716 8478 14720
rect 8414 14660 8418 14716
rect 8418 14660 8474 14716
rect 8474 14660 8478 14716
rect 8414 14656 8478 14660
rect 22618 14716 22682 14720
rect 22618 14660 22622 14716
rect 22622 14660 22678 14716
rect 22678 14660 22682 14716
rect 22618 14656 22682 14660
rect 22698 14716 22762 14720
rect 22698 14660 22702 14716
rect 22702 14660 22758 14716
rect 22758 14660 22762 14716
rect 22698 14656 22762 14660
rect 22778 14716 22842 14720
rect 22778 14660 22782 14716
rect 22782 14660 22838 14716
rect 22838 14660 22842 14716
rect 22778 14656 22842 14660
rect 22858 14716 22922 14720
rect 22858 14660 22862 14716
rect 22862 14660 22918 14716
rect 22918 14660 22922 14716
rect 22858 14656 22922 14660
rect 37062 14716 37126 14720
rect 37062 14660 37066 14716
rect 37066 14660 37122 14716
rect 37122 14660 37126 14716
rect 37062 14656 37126 14660
rect 37142 14716 37206 14720
rect 37142 14660 37146 14716
rect 37146 14660 37202 14716
rect 37202 14660 37206 14716
rect 37142 14656 37206 14660
rect 37222 14716 37286 14720
rect 37222 14660 37226 14716
rect 37226 14660 37282 14716
rect 37282 14660 37286 14716
rect 37222 14656 37286 14660
rect 37302 14716 37366 14720
rect 37302 14660 37306 14716
rect 37306 14660 37362 14716
rect 37362 14660 37366 14716
rect 37302 14656 37366 14660
rect 51506 14716 51570 14720
rect 51506 14660 51510 14716
rect 51510 14660 51566 14716
rect 51566 14660 51570 14716
rect 51506 14656 51570 14660
rect 51586 14716 51650 14720
rect 51586 14660 51590 14716
rect 51590 14660 51646 14716
rect 51646 14660 51650 14716
rect 51586 14656 51650 14660
rect 51666 14716 51730 14720
rect 51666 14660 51670 14716
rect 51670 14660 51726 14716
rect 51726 14660 51730 14716
rect 51666 14656 51730 14660
rect 51746 14716 51810 14720
rect 51746 14660 51750 14716
rect 51750 14660 51806 14716
rect 51806 14660 51810 14716
rect 51746 14656 51810 14660
rect 15396 14172 15460 14176
rect 15396 14116 15400 14172
rect 15400 14116 15456 14172
rect 15456 14116 15460 14172
rect 15396 14112 15460 14116
rect 15476 14172 15540 14176
rect 15476 14116 15480 14172
rect 15480 14116 15536 14172
rect 15536 14116 15540 14172
rect 15476 14112 15540 14116
rect 15556 14172 15620 14176
rect 15556 14116 15560 14172
rect 15560 14116 15616 14172
rect 15616 14116 15620 14172
rect 15556 14112 15620 14116
rect 15636 14172 15700 14176
rect 15636 14116 15640 14172
rect 15640 14116 15696 14172
rect 15696 14116 15700 14172
rect 15636 14112 15700 14116
rect 29840 14172 29904 14176
rect 29840 14116 29844 14172
rect 29844 14116 29900 14172
rect 29900 14116 29904 14172
rect 29840 14112 29904 14116
rect 29920 14172 29984 14176
rect 29920 14116 29924 14172
rect 29924 14116 29980 14172
rect 29980 14116 29984 14172
rect 29920 14112 29984 14116
rect 30000 14172 30064 14176
rect 30000 14116 30004 14172
rect 30004 14116 30060 14172
rect 30060 14116 30064 14172
rect 30000 14112 30064 14116
rect 30080 14172 30144 14176
rect 30080 14116 30084 14172
rect 30084 14116 30140 14172
rect 30140 14116 30144 14172
rect 30080 14112 30144 14116
rect 44284 14172 44348 14176
rect 44284 14116 44288 14172
rect 44288 14116 44344 14172
rect 44344 14116 44348 14172
rect 44284 14112 44348 14116
rect 44364 14172 44428 14176
rect 44364 14116 44368 14172
rect 44368 14116 44424 14172
rect 44424 14116 44428 14172
rect 44364 14112 44428 14116
rect 44444 14172 44508 14176
rect 44444 14116 44448 14172
rect 44448 14116 44504 14172
rect 44504 14116 44508 14172
rect 44444 14112 44508 14116
rect 44524 14172 44588 14176
rect 44524 14116 44528 14172
rect 44528 14116 44584 14172
rect 44584 14116 44588 14172
rect 44524 14112 44588 14116
rect 58728 14172 58792 14176
rect 58728 14116 58732 14172
rect 58732 14116 58788 14172
rect 58788 14116 58792 14172
rect 58728 14112 58792 14116
rect 58808 14172 58872 14176
rect 58808 14116 58812 14172
rect 58812 14116 58868 14172
rect 58868 14116 58872 14172
rect 58808 14112 58872 14116
rect 58888 14172 58952 14176
rect 58888 14116 58892 14172
rect 58892 14116 58948 14172
rect 58948 14116 58952 14172
rect 58888 14112 58952 14116
rect 58968 14172 59032 14176
rect 58968 14116 58972 14172
rect 58972 14116 59028 14172
rect 59028 14116 59032 14172
rect 58968 14112 59032 14116
rect 8174 13628 8238 13632
rect 8174 13572 8178 13628
rect 8178 13572 8234 13628
rect 8234 13572 8238 13628
rect 8174 13568 8238 13572
rect 8254 13628 8318 13632
rect 8254 13572 8258 13628
rect 8258 13572 8314 13628
rect 8314 13572 8318 13628
rect 8254 13568 8318 13572
rect 8334 13628 8398 13632
rect 8334 13572 8338 13628
rect 8338 13572 8394 13628
rect 8394 13572 8398 13628
rect 8334 13568 8398 13572
rect 8414 13628 8478 13632
rect 8414 13572 8418 13628
rect 8418 13572 8474 13628
rect 8474 13572 8478 13628
rect 8414 13568 8478 13572
rect 22618 13628 22682 13632
rect 22618 13572 22622 13628
rect 22622 13572 22678 13628
rect 22678 13572 22682 13628
rect 22618 13568 22682 13572
rect 22698 13628 22762 13632
rect 22698 13572 22702 13628
rect 22702 13572 22758 13628
rect 22758 13572 22762 13628
rect 22698 13568 22762 13572
rect 22778 13628 22842 13632
rect 22778 13572 22782 13628
rect 22782 13572 22838 13628
rect 22838 13572 22842 13628
rect 22778 13568 22842 13572
rect 22858 13628 22922 13632
rect 22858 13572 22862 13628
rect 22862 13572 22918 13628
rect 22918 13572 22922 13628
rect 22858 13568 22922 13572
rect 37062 13628 37126 13632
rect 37062 13572 37066 13628
rect 37066 13572 37122 13628
rect 37122 13572 37126 13628
rect 37062 13568 37126 13572
rect 37142 13628 37206 13632
rect 37142 13572 37146 13628
rect 37146 13572 37202 13628
rect 37202 13572 37206 13628
rect 37142 13568 37206 13572
rect 37222 13628 37286 13632
rect 37222 13572 37226 13628
rect 37226 13572 37282 13628
rect 37282 13572 37286 13628
rect 37222 13568 37286 13572
rect 37302 13628 37366 13632
rect 37302 13572 37306 13628
rect 37306 13572 37362 13628
rect 37362 13572 37366 13628
rect 37302 13568 37366 13572
rect 51506 13628 51570 13632
rect 51506 13572 51510 13628
rect 51510 13572 51566 13628
rect 51566 13572 51570 13628
rect 51506 13568 51570 13572
rect 51586 13628 51650 13632
rect 51586 13572 51590 13628
rect 51590 13572 51646 13628
rect 51646 13572 51650 13628
rect 51586 13568 51650 13572
rect 51666 13628 51730 13632
rect 51666 13572 51670 13628
rect 51670 13572 51726 13628
rect 51726 13572 51730 13628
rect 51666 13568 51730 13572
rect 51746 13628 51810 13632
rect 51746 13572 51750 13628
rect 51750 13572 51806 13628
rect 51806 13572 51810 13628
rect 51746 13568 51810 13572
rect 15396 13084 15460 13088
rect 15396 13028 15400 13084
rect 15400 13028 15456 13084
rect 15456 13028 15460 13084
rect 15396 13024 15460 13028
rect 15476 13084 15540 13088
rect 15476 13028 15480 13084
rect 15480 13028 15536 13084
rect 15536 13028 15540 13084
rect 15476 13024 15540 13028
rect 15556 13084 15620 13088
rect 15556 13028 15560 13084
rect 15560 13028 15616 13084
rect 15616 13028 15620 13084
rect 15556 13024 15620 13028
rect 15636 13084 15700 13088
rect 15636 13028 15640 13084
rect 15640 13028 15696 13084
rect 15696 13028 15700 13084
rect 15636 13024 15700 13028
rect 29840 13084 29904 13088
rect 29840 13028 29844 13084
rect 29844 13028 29900 13084
rect 29900 13028 29904 13084
rect 29840 13024 29904 13028
rect 29920 13084 29984 13088
rect 29920 13028 29924 13084
rect 29924 13028 29980 13084
rect 29980 13028 29984 13084
rect 29920 13024 29984 13028
rect 30000 13084 30064 13088
rect 30000 13028 30004 13084
rect 30004 13028 30060 13084
rect 30060 13028 30064 13084
rect 30000 13024 30064 13028
rect 30080 13084 30144 13088
rect 30080 13028 30084 13084
rect 30084 13028 30140 13084
rect 30140 13028 30144 13084
rect 30080 13024 30144 13028
rect 44284 13084 44348 13088
rect 44284 13028 44288 13084
rect 44288 13028 44344 13084
rect 44344 13028 44348 13084
rect 44284 13024 44348 13028
rect 44364 13084 44428 13088
rect 44364 13028 44368 13084
rect 44368 13028 44424 13084
rect 44424 13028 44428 13084
rect 44364 13024 44428 13028
rect 44444 13084 44508 13088
rect 44444 13028 44448 13084
rect 44448 13028 44504 13084
rect 44504 13028 44508 13084
rect 44444 13024 44508 13028
rect 44524 13084 44588 13088
rect 44524 13028 44528 13084
rect 44528 13028 44584 13084
rect 44584 13028 44588 13084
rect 44524 13024 44588 13028
rect 58728 13084 58792 13088
rect 58728 13028 58732 13084
rect 58732 13028 58788 13084
rect 58788 13028 58792 13084
rect 58728 13024 58792 13028
rect 58808 13084 58872 13088
rect 58808 13028 58812 13084
rect 58812 13028 58868 13084
rect 58868 13028 58872 13084
rect 58808 13024 58872 13028
rect 58888 13084 58952 13088
rect 58888 13028 58892 13084
rect 58892 13028 58948 13084
rect 58948 13028 58952 13084
rect 58888 13024 58952 13028
rect 58968 13084 59032 13088
rect 58968 13028 58972 13084
rect 58972 13028 59028 13084
rect 59028 13028 59032 13084
rect 58968 13024 59032 13028
rect 8174 12540 8238 12544
rect 8174 12484 8178 12540
rect 8178 12484 8234 12540
rect 8234 12484 8238 12540
rect 8174 12480 8238 12484
rect 8254 12540 8318 12544
rect 8254 12484 8258 12540
rect 8258 12484 8314 12540
rect 8314 12484 8318 12540
rect 8254 12480 8318 12484
rect 8334 12540 8398 12544
rect 8334 12484 8338 12540
rect 8338 12484 8394 12540
rect 8394 12484 8398 12540
rect 8334 12480 8398 12484
rect 8414 12540 8478 12544
rect 8414 12484 8418 12540
rect 8418 12484 8474 12540
rect 8474 12484 8478 12540
rect 8414 12480 8478 12484
rect 22618 12540 22682 12544
rect 22618 12484 22622 12540
rect 22622 12484 22678 12540
rect 22678 12484 22682 12540
rect 22618 12480 22682 12484
rect 22698 12540 22762 12544
rect 22698 12484 22702 12540
rect 22702 12484 22758 12540
rect 22758 12484 22762 12540
rect 22698 12480 22762 12484
rect 22778 12540 22842 12544
rect 22778 12484 22782 12540
rect 22782 12484 22838 12540
rect 22838 12484 22842 12540
rect 22778 12480 22842 12484
rect 22858 12540 22922 12544
rect 22858 12484 22862 12540
rect 22862 12484 22918 12540
rect 22918 12484 22922 12540
rect 22858 12480 22922 12484
rect 37062 12540 37126 12544
rect 37062 12484 37066 12540
rect 37066 12484 37122 12540
rect 37122 12484 37126 12540
rect 37062 12480 37126 12484
rect 37142 12540 37206 12544
rect 37142 12484 37146 12540
rect 37146 12484 37202 12540
rect 37202 12484 37206 12540
rect 37142 12480 37206 12484
rect 37222 12540 37286 12544
rect 37222 12484 37226 12540
rect 37226 12484 37282 12540
rect 37282 12484 37286 12540
rect 37222 12480 37286 12484
rect 37302 12540 37366 12544
rect 37302 12484 37306 12540
rect 37306 12484 37362 12540
rect 37362 12484 37366 12540
rect 37302 12480 37366 12484
rect 51506 12540 51570 12544
rect 51506 12484 51510 12540
rect 51510 12484 51566 12540
rect 51566 12484 51570 12540
rect 51506 12480 51570 12484
rect 51586 12540 51650 12544
rect 51586 12484 51590 12540
rect 51590 12484 51646 12540
rect 51646 12484 51650 12540
rect 51586 12480 51650 12484
rect 51666 12540 51730 12544
rect 51666 12484 51670 12540
rect 51670 12484 51726 12540
rect 51726 12484 51730 12540
rect 51666 12480 51730 12484
rect 51746 12540 51810 12544
rect 51746 12484 51750 12540
rect 51750 12484 51806 12540
rect 51806 12484 51810 12540
rect 51746 12480 51810 12484
rect 15396 11996 15460 12000
rect 15396 11940 15400 11996
rect 15400 11940 15456 11996
rect 15456 11940 15460 11996
rect 15396 11936 15460 11940
rect 15476 11996 15540 12000
rect 15476 11940 15480 11996
rect 15480 11940 15536 11996
rect 15536 11940 15540 11996
rect 15476 11936 15540 11940
rect 15556 11996 15620 12000
rect 15556 11940 15560 11996
rect 15560 11940 15616 11996
rect 15616 11940 15620 11996
rect 15556 11936 15620 11940
rect 15636 11996 15700 12000
rect 15636 11940 15640 11996
rect 15640 11940 15696 11996
rect 15696 11940 15700 11996
rect 15636 11936 15700 11940
rect 29840 11996 29904 12000
rect 29840 11940 29844 11996
rect 29844 11940 29900 11996
rect 29900 11940 29904 11996
rect 29840 11936 29904 11940
rect 29920 11996 29984 12000
rect 29920 11940 29924 11996
rect 29924 11940 29980 11996
rect 29980 11940 29984 11996
rect 29920 11936 29984 11940
rect 30000 11996 30064 12000
rect 30000 11940 30004 11996
rect 30004 11940 30060 11996
rect 30060 11940 30064 11996
rect 30000 11936 30064 11940
rect 30080 11996 30144 12000
rect 30080 11940 30084 11996
rect 30084 11940 30140 11996
rect 30140 11940 30144 11996
rect 30080 11936 30144 11940
rect 44284 11996 44348 12000
rect 44284 11940 44288 11996
rect 44288 11940 44344 11996
rect 44344 11940 44348 11996
rect 44284 11936 44348 11940
rect 44364 11996 44428 12000
rect 44364 11940 44368 11996
rect 44368 11940 44424 11996
rect 44424 11940 44428 11996
rect 44364 11936 44428 11940
rect 44444 11996 44508 12000
rect 44444 11940 44448 11996
rect 44448 11940 44504 11996
rect 44504 11940 44508 11996
rect 44444 11936 44508 11940
rect 44524 11996 44588 12000
rect 44524 11940 44528 11996
rect 44528 11940 44584 11996
rect 44584 11940 44588 11996
rect 44524 11936 44588 11940
rect 58728 11996 58792 12000
rect 58728 11940 58732 11996
rect 58732 11940 58788 11996
rect 58788 11940 58792 11996
rect 58728 11936 58792 11940
rect 58808 11996 58872 12000
rect 58808 11940 58812 11996
rect 58812 11940 58868 11996
rect 58868 11940 58872 11996
rect 58808 11936 58872 11940
rect 58888 11996 58952 12000
rect 58888 11940 58892 11996
rect 58892 11940 58948 11996
rect 58948 11940 58952 11996
rect 58888 11936 58952 11940
rect 58968 11996 59032 12000
rect 58968 11940 58972 11996
rect 58972 11940 59028 11996
rect 59028 11940 59032 11996
rect 58968 11936 59032 11940
rect 8174 11452 8238 11456
rect 8174 11396 8178 11452
rect 8178 11396 8234 11452
rect 8234 11396 8238 11452
rect 8174 11392 8238 11396
rect 8254 11452 8318 11456
rect 8254 11396 8258 11452
rect 8258 11396 8314 11452
rect 8314 11396 8318 11452
rect 8254 11392 8318 11396
rect 8334 11452 8398 11456
rect 8334 11396 8338 11452
rect 8338 11396 8394 11452
rect 8394 11396 8398 11452
rect 8334 11392 8398 11396
rect 8414 11452 8478 11456
rect 8414 11396 8418 11452
rect 8418 11396 8474 11452
rect 8474 11396 8478 11452
rect 8414 11392 8478 11396
rect 22618 11452 22682 11456
rect 22618 11396 22622 11452
rect 22622 11396 22678 11452
rect 22678 11396 22682 11452
rect 22618 11392 22682 11396
rect 22698 11452 22762 11456
rect 22698 11396 22702 11452
rect 22702 11396 22758 11452
rect 22758 11396 22762 11452
rect 22698 11392 22762 11396
rect 22778 11452 22842 11456
rect 22778 11396 22782 11452
rect 22782 11396 22838 11452
rect 22838 11396 22842 11452
rect 22778 11392 22842 11396
rect 22858 11452 22922 11456
rect 22858 11396 22862 11452
rect 22862 11396 22918 11452
rect 22918 11396 22922 11452
rect 22858 11392 22922 11396
rect 37062 11452 37126 11456
rect 37062 11396 37066 11452
rect 37066 11396 37122 11452
rect 37122 11396 37126 11452
rect 37062 11392 37126 11396
rect 37142 11452 37206 11456
rect 37142 11396 37146 11452
rect 37146 11396 37202 11452
rect 37202 11396 37206 11452
rect 37142 11392 37206 11396
rect 37222 11452 37286 11456
rect 37222 11396 37226 11452
rect 37226 11396 37282 11452
rect 37282 11396 37286 11452
rect 37222 11392 37286 11396
rect 37302 11452 37366 11456
rect 37302 11396 37306 11452
rect 37306 11396 37362 11452
rect 37362 11396 37366 11452
rect 37302 11392 37366 11396
rect 51506 11452 51570 11456
rect 51506 11396 51510 11452
rect 51510 11396 51566 11452
rect 51566 11396 51570 11452
rect 51506 11392 51570 11396
rect 51586 11452 51650 11456
rect 51586 11396 51590 11452
rect 51590 11396 51646 11452
rect 51646 11396 51650 11452
rect 51586 11392 51650 11396
rect 51666 11452 51730 11456
rect 51666 11396 51670 11452
rect 51670 11396 51726 11452
rect 51726 11396 51730 11452
rect 51666 11392 51730 11396
rect 51746 11452 51810 11456
rect 51746 11396 51750 11452
rect 51750 11396 51806 11452
rect 51806 11396 51810 11452
rect 51746 11392 51810 11396
rect 57100 11052 57164 11116
rect 15396 10908 15460 10912
rect 15396 10852 15400 10908
rect 15400 10852 15456 10908
rect 15456 10852 15460 10908
rect 15396 10848 15460 10852
rect 15476 10908 15540 10912
rect 15476 10852 15480 10908
rect 15480 10852 15536 10908
rect 15536 10852 15540 10908
rect 15476 10848 15540 10852
rect 15556 10908 15620 10912
rect 15556 10852 15560 10908
rect 15560 10852 15616 10908
rect 15616 10852 15620 10908
rect 15556 10848 15620 10852
rect 15636 10908 15700 10912
rect 15636 10852 15640 10908
rect 15640 10852 15696 10908
rect 15696 10852 15700 10908
rect 15636 10848 15700 10852
rect 29840 10908 29904 10912
rect 29840 10852 29844 10908
rect 29844 10852 29900 10908
rect 29900 10852 29904 10908
rect 29840 10848 29904 10852
rect 29920 10908 29984 10912
rect 29920 10852 29924 10908
rect 29924 10852 29980 10908
rect 29980 10852 29984 10908
rect 29920 10848 29984 10852
rect 30000 10908 30064 10912
rect 30000 10852 30004 10908
rect 30004 10852 30060 10908
rect 30060 10852 30064 10908
rect 30000 10848 30064 10852
rect 30080 10908 30144 10912
rect 30080 10852 30084 10908
rect 30084 10852 30140 10908
rect 30140 10852 30144 10908
rect 30080 10848 30144 10852
rect 44284 10908 44348 10912
rect 44284 10852 44288 10908
rect 44288 10852 44344 10908
rect 44344 10852 44348 10908
rect 44284 10848 44348 10852
rect 44364 10908 44428 10912
rect 44364 10852 44368 10908
rect 44368 10852 44424 10908
rect 44424 10852 44428 10908
rect 44364 10848 44428 10852
rect 44444 10908 44508 10912
rect 44444 10852 44448 10908
rect 44448 10852 44504 10908
rect 44504 10852 44508 10908
rect 44444 10848 44508 10852
rect 44524 10908 44588 10912
rect 44524 10852 44528 10908
rect 44528 10852 44584 10908
rect 44584 10852 44588 10908
rect 44524 10848 44588 10852
rect 58728 10908 58792 10912
rect 58728 10852 58732 10908
rect 58732 10852 58788 10908
rect 58788 10852 58792 10908
rect 58728 10848 58792 10852
rect 58808 10908 58872 10912
rect 58808 10852 58812 10908
rect 58812 10852 58868 10908
rect 58868 10852 58872 10908
rect 58808 10848 58872 10852
rect 58888 10908 58952 10912
rect 58888 10852 58892 10908
rect 58892 10852 58948 10908
rect 58948 10852 58952 10908
rect 58888 10848 58952 10852
rect 58968 10908 59032 10912
rect 58968 10852 58972 10908
rect 58972 10852 59028 10908
rect 59028 10852 59032 10908
rect 58968 10848 59032 10852
rect 8174 10364 8238 10368
rect 8174 10308 8178 10364
rect 8178 10308 8234 10364
rect 8234 10308 8238 10364
rect 8174 10304 8238 10308
rect 8254 10364 8318 10368
rect 8254 10308 8258 10364
rect 8258 10308 8314 10364
rect 8314 10308 8318 10364
rect 8254 10304 8318 10308
rect 8334 10364 8398 10368
rect 8334 10308 8338 10364
rect 8338 10308 8394 10364
rect 8394 10308 8398 10364
rect 8334 10304 8398 10308
rect 8414 10364 8478 10368
rect 8414 10308 8418 10364
rect 8418 10308 8474 10364
rect 8474 10308 8478 10364
rect 8414 10304 8478 10308
rect 22618 10364 22682 10368
rect 22618 10308 22622 10364
rect 22622 10308 22678 10364
rect 22678 10308 22682 10364
rect 22618 10304 22682 10308
rect 22698 10364 22762 10368
rect 22698 10308 22702 10364
rect 22702 10308 22758 10364
rect 22758 10308 22762 10364
rect 22698 10304 22762 10308
rect 22778 10364 22842 10368
rect 22778 10308 22782 10364
rect 22782 10308 22838 10364
rect 22838 10308 22842 10364
rect 22778 10304 22842 10308
rect 22858 10364 22922 10368
rect 22858 10308 22862 10364
rect 22862 10308 22918 10364
rect 22918 10308 22922 10364
rect 22858 10304 22922 10308
rect 37062 10364 37126 10368
rect 37062 10308 37066 10364
rect 37066 10308 37122 10364
rect 37122 10308 37126 10364
rect 37062 10304 37126 10308
rect 37142 10364 37206 10368
rect 37142 10308 37146 10364
rect 37146 10308 37202 10364
rect 37202 10308 37206 10364
rect 37142 10304 37206 10308
rect 37222 10364 37286 10368
rect 37222 10308 37226 10364
rect 37226 10308 37282 10364
rect 37282 10308 37286 10364
rect 37222 10304 37286 10308
rect 37302 10364 37366 10368
rect 37302 10308 37306 10364
rect 37306 10308 37362 10364
rect 37362 10308 37366 10364
rect 37302 10304 37366 10308
rect 51506 10364 51570 10368
rect 51506 10308 51510 10364
rect 51510 10308 51566 10364
rect 51566 10308 51570 10364
rect 51506 10304 51570 10308
rect 51586 10364 51650 10368
rect 51586 10308 51590 10364
rect 51590 10308 51646 10364
rect 51646 10308 51650 10364
rect 51586 10304 51650 10308
rect 51666 10364 51730 10368
rect 51666 10308 51670 10364
rect 51670 10308 51726 10364
rect 51726 10308 51730 10364
rect 51666 10304 51730 10308
rect 51746 10364 51810 10368
rect 51746 10308 51750 10364
rect 51750 10308 51806 10364
rect 51806 10308 51810 10364
rect 51746 10304 51810 10308
rect 15396 9820 15460 9824
rect 15396 9764 15400 9820
rect 15400 9764 15456 9820
rect 15456 9764 15460 9820
rect 15396 9760 15460 9764
rect 15476 9820 15540 9824
rect 15476 9764 15480 9820
rect 15480 9764 15536 9820
rect 15536 9764 15540 9820
rect 15476 9760 15540 9764
rect 15556 9820 15620 9824
rect 15556 9764 15560 9820
rect 15560 9764 15616 9820
rect 15616 9764 15620 9820
rect 15556 9760 15620 9764
rect 15636 9820 15700 9824
rect 15636 9764 15640 9820
rect 15640 9764 15696 9820
rect 15696 9764 15700 9820
rect 15636 9760 15700 9764
rect 29840 9820 29904 9824
rect 29840 9764 29844 9820
rect 29844 9764 29900 9820
rect 29900 9764 29904 9820
rect 29840 9760 29904 9764
rect 29920 9820 29984 9824
rect 29920 9764 29924 9820
rect 29924 9764 29980 9820
rect 29980 9764 29984 9820
rect 29920 9760 29984 9764
rect 30000 9820 30064 9824
rect 30000 9764 30004 9820
rect 30004 9764 30060 9820
rect 30060 9764 30064 9820
rect 30000 9760 30064 9764
rect 30080 9820 30144 9824
rect 30080 9764 30084 9820
rect 30084 9764 30140 9820
rect 30140 9764 30144 9820
rect 30080 9760 30144 9764
rect 44284 9820 44348 9824
rect 44284 9764 44288 9820
rect 44288 9764 44344 9820
rect 44344 9764 44348 9820
rect 44284 9760 44348 9764
rect 44364 9820 44428 9824
rect 44364 9764 44368 9820
rect 44368 9764 44424 9820
rect 44424 9764 44428 9820
rect 44364 9760 44428 9764
rect 44444 9820 44508 9824
rect 44444 9764 44448 9820
rect 44448 9764 44504 9820
rect 44504 9764 44508 9820
rect 44444 9760 44508 9764
rect 44524 9820 44588 9824
rect 44524 9764 44528 9820
rect 44528 9764 44584 9820
rect 44584 9764 44588 9820
rect 44524 9760 44588 9764
rect 58728 9820 58792 9824
rect 58728 9764 58732 9820
rect 58732 9764 58788 9820
rect 58788 9764 58792 9820
rect 58728 9760 58792 9764
rect 58808 9820 58872 9824
rect 58808 9764 58812 9820
rect 58812 9764 58868 9820
rect 58868 9764 58872 9820
rect 58808 9760 58872 9764
rect 58888 9820 58952 9824
rect 58888 9764 58892 9820
rect 58892 9764 58948 9820
rect 58948 9764 58952 9820
rect 58888 9760 58952 9764
rect 58968 9820 59032 9824
rect 58968 9764 58972 9820
rect 58972 9764 59028 9820
rect 59028 9764 59032 9820
rect 58968 9760 59032 9764
rect 8174 9276 8238 9280
rect 8174 9220 8178 9276
rect 8178 9220 8234 9276
rect 8234 9220 8238 9276
rect 8174 9216 8238 9220
rect 8254 9276 8318 9280
rect 8254 9220 8258 9276
rect 8258 9220 8314 9276
rect 8314 9220 8318 9276
rect 8254 9216 8318 9220
rect 8334 9276 8398 9280
rect 8334 9220 8338 9276
rect 8338 9220 8394 9276
rect 8394 9220 8398 9276
rect 8334 9216 8398 9220
rect 8414 9276 8478 9280
rect 8414 9220 8418 9276
rect 8418 9220 8474 9276
rect 8474 9220 8478 9276
rect 8414 9216 8478 9220
rect 22618 9276 22682 9280
rect 22618 9220 22622 9276
rect 22622 9220 22678 9276
rect 22678 9220 22682 9276
rect 22618 9216 22682 9220
rect 22698 9276 22762 9280
rect 22698 9220 22702 9276
rect 22702 9220 22758 9276
rect 22758 9220 22762 9276
rect 22698 9216 22762 9220
rect 22778 9276 22842 9280
rect 22778 9220 22782 9276
rect 22782 9220 22838 9276
rect 22838 9220 22842 9276
rect 22778 9216 22842 9220
rect 22858 9276 22922 9280
rect 22858 9220 22862 9276
rect 22862 9220 22918 9276
rect 22918 9220 22922 9276
rect 22858 9216 22922 9220
rect 37062 9276 37126 9280
rect 37062 9220 37066 9276
rect 37066 9220 37122 9276
rect 37122 9220 37126 9276
rect 37062 9216 37126 9220
rect 37142 9276 37206 9280
rect 37142 9220 37146 9276
rect 37146 9220 37202 9276
rect 37202 9220 37206 9276
rect 37142 9216 37206 9220
rect 37222 9276 37286 9280
rect 37222 9220 37226 9276
rect 37226 9220 37282 9276
rect 37282 9220 37286 9276
rect 37222 9216 37286 9220
rect 37302 9276 37366 9280
rect 37302 9220 37306 9276
rect 37306 9220 37362 9276
rect 37362 9220 37366 9276
rect 37302 9216 37366 9220
rect 51506 9276 51570 9280
rect 51506 9220 51510 9276
rect 51510 9220 51566 9276
rect 51566 9220 51570 9276
rect 51506 9216 51570 9220
rect 51586 9276 51650 9280
rect 51586 9220 51590 9276
rect 51590 9220 51646 9276
rect 51646 9220 51650 9276
rect 51586 9216 51650 9220
rect 51666 9276 51730 9280
rect 51666 9220 51670 9276
rect 51670 9220 51726 9276
rect 51726 9220 51730 9276
rect 51666 9216 51730 9220
rect 51746 9276 51810 9280
rect 51746 9220 51750 9276
rect 51750 9220 51806 9276
rect 51806 9220 51810 9276
rect 51746 9216 51810 9220
rect 15396 8732 15460 8736
rect 15396 8676 15400 8732
rect 15400 8676 15456 8732
rect 15456 8676 15460 8732
rect 15396 8672 15460 8676
rect 15476 8732 15540 8736
rect 15476 8676 15480 8732
rect 15480 8676 15536 8732
rect 15536 8676 15540 8732
rect 15476 8672 15540 8676
rect 15556 8732 15620 8736
rect 15556 8676 15560 8732
rect 15560 8676 15616 8732
rect 15616 8676 15620 8732
rect 15556 8672 15620 8676
rect 15636 8732 15700 8736
rect 15636 8676 15640 8732
rect 15640 8676 15696 8732
rect 15696 8676 15700 8732
rect 15636 8672 15700 8676
rect 29840 8732 29904 8736
rect 29840 8676 29844 8732
rect 29844 8676 29900 8732
rect 29900 8676 29904 8732
rect 29840 8672 29904 8676
rect 29920 8732 29984 8736
rect 29920 8676 29924 8732
rect 29924 8676 29980 8732
rect 29980 8676 29984 8732
rect 29920 8672 29984 8676
rect 30000 8732 30064 8736
rect 30000 8676 30004 8732
rect 30004 8676 30060 8732
rect 30060 8676 30064 8732
rect 30000 8672 30064 8676
rect 30080 8732 30144 8736
rect 30080 8676 30084 8732
rect 30084 8676 30140 8732
rect 30140 8676 30144 8732
rect 30080 8672 30144 8676
rect 44284 8732 44348 8736
rect 44284 8676 44288 8732
rect 44288 8676 44344 8732
rect 44344 8676 44348 8732
rect 44284 8672 44348 8676
rect 44364 8732 44428 8736
rect 44364 8676 44368 8732
rect 44368 8676 44424 8732
rect 44424 8676 44428 8732
rect 44364 8672 44428 8676
rect 44444 8732 44508 8736
rect 44444 8676 44448 8732
rect 44448 8676 44504 8732
rect 44504 8676 44508 8732
rect 44444 8672 44508 8676
rect 44524 8732 44588 8736
rect 44524 8676 44528 8732
rect 44528 8676 44584 8732
rect 44584 8676 44588 8732
rect 44524 8672 44588 8676
rect 58728 8732 58792 8736
rect 58728 8676 58732 8732
rect 58732 8676 58788 8732
rect 58788 8676 58792 8732
rect 58728 8672 58792 8676
rect 58808 8732 58872 8736
rect 58808 8676 58812 8732
rect 58812 8676 58868 8732
rect 58868 8676 58872 8732
rect 58808 8672 58872 8676
rect 58888 8732 58952 8736
rect 58888 8676 58892 8732
rect 58892 8676 58948 8732
rect 58948 8676 58952 8732
rect 58888 8672 58952 8676
rect 58968 8732 59032 8736
rect 58968 8676 58972 8732
rect 58972 8676 59028 8732
rect 59028 8676 59032 8732
rect 58968 8672 59032 8676
rect 8174 8188 8238 8192
rect 8174 8132 8178 8188
rect 8178 8132 8234 8188
rect 8234 8132 8238 8188
rect 8174 8128 8238 8132
rect 8254 8188 8318 8192
rect 8254 8132 8258 8188
rect 8258 8132 8314 8188
rect 8314 8132 8318 8188
rect 8254 8128 8318 8132
rect 8334 8188 8398 8192
rect 8334 8132 8338 8188
rect 8338 8132 8394 8188
rect 8394 8132 8398 8188
rect 8334 8128 8398 8132
rect 8414 8188 8478 8192
rect 8414 8132 8418 8188
rect 8418 8132 8474 8188
rect 8474 8132 8478 8188
rect 8414 8128 8478 8132
rect 22618 8188 22682 8192
rect 22618 8132 22622 8188
rect 22622 8132 22678 8188
rect 22678 8132 22682 8188
rect 22618 8128 22682 8132
rect 22698 8188 22762 8192
rect 22698 8132 22702 8188
rect 22702 8132 22758 8188
rect 22758 8132 22762 8188
rect 22698 8128 22762 8132
rect 22778 8188 22842 8192
rect 22778 8132 22782 8188
rect 22782 8132 22838 8188
rect 22838 8132 22842 8188
rect 22778 8128 22842 8132
rect 22858 8188 22922 8192
rect 22858 8132 22862 8188
rect 22862 8132 22918 8188
rect 22918 8132 22922 8188
rect 22858 8128 22922 8132
rect 37062 8188 37126 8192
rect 37062 8132 37066 8188
rect 37066 8132 37122 8188
rect 37122 8132 37126 8188
rect 37062 8128 37126 8132
rect 37142 8188 37206 8192
rect 37142 8132 37146 8188
rect 37146 8132 37202 8188
rect 37202 8132 37206 8188
rect 37142 8128 37206 8132
rect 37222 8188 37286 8192
rect 37222 8132 37226 8188
rect 37226 8132 37282 8188
rect 37282 8132 37286 8188
rect 37222 8128 37286 8132
rect 37302 8188 37366 8192
rect 37302 8132 37306 8188
rect 37306 8132 37362 8188
rect 37362 8132 37366 8188
rect 37302 8128 37366 8132
rect 51506 8188 51570 8192
rect 51506 8132 51510 8188
rect 51510 8132 51566 8188
rect 51566 8132 51570 8188
rect 51506 8128 51570 8132
rect 51586 8188 51650 8192
rect 51586 8132 51590 8188
rect 51590 8132 51646 8188
rect 51646 8132 51650 8188
rect 51586 8128 51650 8132
rect 51666 8188 51730 8192
rect 51666 8132 51670 8188
rect 51670 8132 51726 8188
rect 51726 8132 51730 8188
rect 51666 8128 51730 8132
rect 51746 8188 51810 8192
rect 51746 8132 51750 8188
rect 51750 8132 51806 8188
rect 51806 8132 51810 8188
rect 51746 8128 51810 8132
rect 15396 7644 15460 7648
rect 15396 7588 15400 7644
rect 15400 7588 15456 7644
rect 15456 7588 15460 7644
rect 15396 7584 15460 7588
rect 15476 7644 15540 7648
rect 15476 7588 15480 7644
rect 15480 7588 15536 7644
rect 15536 7588 15540 7644
rect 15476 7584 15540 7588
rect 15556 7644 15620 7648
rect 15556 7588 15560 7644
rect 15560 7588 15616 7644
rect 15616 7588 15620 7644
rect 15556 7584 15620 7588
rect 15636 7644 15700 7648
rect 15636 7588 15640 7644
rect 15640 7588 15696 7644
rect 15696 7588 15700 7644
rect 15636 7584 15700 7588
rect 29840 7644 29904 7648
rect 29840 7588 29844 7644
rect 29844 7588 29900 7644
rect 29900 7588 29904 7644
rect 29840 7584 29904 7588
rect 29920 7644 29984 7648
rect 29920 7588 29924 7644
rect 29924 7588 29980 7644
rect 29980 7588 29984 7644
rect 29920 7584 29984 7588
rect 30000 7644 30064 7648
rect 30000 7588 30004 7644
rect 30004 7588 30060 7644
rect 30060 7588 30064 7644
rect 30000 7584 30064 7588
rect 30080 7644 30144 7648
rect 30080 7588 30084 7644
rect 30084 7588 30140 7644
rect 30140 7588 30144 7644
rect 30080 7584 30144 7588
rect 44284 7644 44348 7648
rect 44284 7588 44288 7644
rect 44288 7588 44344 7644
rect 44344 7588 44348 7644
rect 44284 7584 44348 7588
rect 44364 7644 44428 7648
rect 44364 7588 44368 7644
rect 44368 7588 44424 7644
rect 44424 7588 44428 7644
rect 44364 7584 44428 7588
rect 44444 7644 44508 7648
rect 44444 7588 44448 7644
rect 44448 7588 44504 7644
rect 44504 7588 44508 7644
rect 44444 7584 44508 7588
rect 44524 7644 44588 7648
rect 44524 7588 44528 7644
rect 44528 7588 44584 7644
rect 44584 7588 44588 7644
rect 44524 7584 44588 7588
rect 58728 7644 58792 7648
rect 58728 7588 58732 7644
rect 58732 7588 58788 7644
rect 58788 7588 58792 7644
rect 58728 7584 58792 7588
rect 58808 7644 58872 7648
rect 58808 7588 58812 7644
rect 58812 7588 58868 7644
rect 58868 7588 58872 7644
rect 58808 7584 58872 7588
rect 58888 7644 58952 7648
rect 58888 7588 58892 7644
rect 58892 7588 58948 7644
rect 58948 7588 58952 7644
rect 58888 7584 58952 7588
rect 58968 7644 59032 7648
rect 58968 7588 58972 7644
rect 58972 7588 59028 7644
rect 59028 7588 59032 7644
rect 58968 7584 59032 7588
rect 8174 7100 8238 7104
rect 8174 7044 8178 7100
rect 8178 7044 8234 7100
rect 8234 7044 8238 7100
rect 8174 7040 8238 7044
rect 8254 7100 8318 7104
rect 8254 7044 8258 7100
rect 8258 7044 8314 7100
rect 8314 7044 8318 7100
rect 8254 7040 8318 7044
rect 8334 7100 8398 7104
rect 8334 7044 8338 7100
rect 8338 7044 8394 7100
rect 8394 7044 8398 7100
rect 8334 7040 8398 7044
rect 8414 7100 8478 7104
rect 8414 7044 8418 7100
rect 8418 7044 8474 7100
rect 8474 7044 8478 7100
rect 8414 7040 8478 7044
rect 22618 7100 22682 7104
rect 22618 7044 22622 7100
rect 22622 7044 22678 7100
rect 22678 7044 22682 7100
rect 22618 7040 22682 7044
rect 22698 7100 22762 7104
rect 22698 7044 22702 7100
rect 22702 7044 22758 7100
rect 22758 7044 22762 7100
rect 22698 7040 22762 7044
rect 22778 7100 22842 7104
rect 22778 7044 22782 7100
rect 22782 7044 22838 7100
rect 22838 7044 22842 7100
rect 22778 7040 22842 7044
rect 22858 7100 22922 7104
rect 22858 7044 22862 7100
rect 22862 7044 22918 7100
rect 22918 7044 22922 7100
rect 22858 7040 22922 7044
rect 37062 7100 37126 7104
rect 37062 7044 37066 7100
rect 37066 7044 37122 7100
rect 37122 7044 37126 7100
rect 37062 7040 37126 7044
rect 37142 7100 37206 7104
rect 37142 7044 37146 7100
rect 37146 7044 37202 7100
rect 37202 7044 37206 7100
rect 37142 7040 37206 7044
rect 37222 7100 37286 7104
rect 37222 7044 37226 7100
rect 37226 7044 37282 7100
rect 37282 7044 37286 7100
rect 37222 7040 37286 7044
rect 37302 7100 37366 7104
rect 37302 7044 37306 7100
rect 37306 7044 37362 7100
rect 37362 7044 37366 7100
rect 37302 7040 37366 7044
rect 51506 7100 51570 7104
rect 51506 7044 51510 7100
rect 51510 7044 51566 7100
rect 51566 7044 51570 7100
rect 51506 7040 51570 7044
rect 51586 7100 51650 7104
rect 51586 7044 51590 7100
rect 51590 7044 51646 7100
rect 51646 7044 51650 7100
rect 51586 7040 51650 7044
rect 51666 7100 51730 7104
rect 51666 7044 51670 7100
rect 51670 7044 51726 7100
rect 51726 7044 51730 7100
rect 51666 7040 51730 7044
rect 51746 7100 51810 7104
rect 51746 7044 51750 7100
rect 51750 7044 51806 7100
rect 51806 7044 51810 7100
rect 51746 7040 51810 7044
rect 15396 6556 15460 6560
rect 15396 6500 15400 6556
rect 15400 6500 15456 6556
rect 15456 6500 15460 6556
rect 15396 6496 15460 6500
rect 15476 6556 15540 6560
rect 15476 6500 15480 6556
rect 15480 6500 15536 6556
rect 15536 6500 15540 6556
rect 15476 6496 15540 6500
rect 15556 6556 15620 6560
rect 15556 6500 15560 6556
rect 15560 6500 15616 6556
rect 15616 6500 15620 6556
rect 15556 6496 15620 6500
rect 15636 6556 15700 6560
rect 15636 6500 15640 6556
rect 15640 6500 15696 6556
rect 15696 6500 15700 6556
rect 15636 6496 15700 6500
rect 29840 6556 29904 6560
rect 29840 6500 29844 6556
rect 29844 6500 29900 6556
rect 29900 6500 29904 6556
rect 29840 6496 29904 6500
rect 29920 6556 29984 6560
rect 29920 6500 29924 6556
rect 29924 6500 29980 6556
rect 29980 6500 29984 6556
rect 29920 6496 29984 6500
rect 30000 6556 30064 6560
rect 30000 6500 30004 6556
rect 30004 6500 30060 6556
rect 30060 6500 30064 6556
rect 30000 6496 30064 6500
rect 30080 6556 30144 6560
rect 30080 6500 30084 6556
rect 30084 6500 30140 6556
rect 30140 6500 30144 6556
rect 30080 6496 30144 6500
rect 44284 6556 44348 6560
rect 44284 6500 44288 6556
rect 44288 6500 44344 6556
rect 44344 6500 44348 6556
rect 44284 6496 44348 6500
rect 44364 6556 44428 6560
rect 44364 6500 44368 6556
rect 44368 6500 44424 6556
rect 44424 6500 44428 6556
rect 44364 6496 44428 6500
rect 44444 6556 44508 6560
rect 44444 6500 44448 6556
rect 44448 6500 44504 6556
rect 44504 6500 44508 6556
rect 44444 6496 44508 6500
rect 44524 6556 44588 6560
rect 44524 6500 44528 6556
rect 44528 6500 44584 6556
rect 44584 6500 44588 6556
rect 44524 6496 44588 6500
rect 58728 6556 58792 6560
rect 58728 6500 58732 6556
rect 58732 6500 58788 6556
rect 58788 6500 58792 6556
rect 58728 6496 58792 6500
rect 58808 6556 58872 6560
rect 58808 6500 58812 6556
rect 58812 6500 58868 6556
rect 58868 6500 58872 6556
rect 58808 6496 58872 6500
rect 58888 6556 58952 6560
rect 58888 6500 58892 6556
rect 58892 6500 58948 6556
rect 58948 6500 58952 6556
rect 58888 6496 58952 6500
rect 58968 6556 59032 6560
rect 58968 6500 58972 6556
rect 58972 6500 59028 6556
rect 59028 6500 59032 6556
rect 58968 6496 59032 6500
rect 8174 6012 8238 6016
rect 8174 5956 8178 6012
rect 8178 5956 8234 6012
rect 8234 5956 8238 6012
rect 8174 5952 8238 5956
rect 8254 6012 8318 6016
rect 8254 5956 8258 6012
rect 8258 5956 8314 6012
rect 8314 5956 8318 6012
rect 8254 5952 8318 5956
rect 8334 6012 8398 6016
rect 8334 5956 8338 6012
rect 8338 5956 8394 6012
rect 8394 5956 8398 6012
rect 8334 5952 8398 5956
rect 8414 6012 8478 6016
rect 8414 5956 8418 6012
rect 8418 5956 8474 6012
rect 8474 5956 8478 6012
rect 8414 5952 8478 5956
rect 22618 6012 22682 6016
rect 22618 5956 22622 6012
rect 22622 5956 22678 6012
rect 22678 5956 22682 6012
rect 22618 5952 22682 5956
rect 22698 6012 22762 6016
rect 22698 5956 22702 6012
rect 22702 5956 22758 6012
rect 22758 5956 22762 6012
rect 22698 5952 22762 5956
rect 22778 6012 22842 6016
rect 22778 5956 22782 6012
rect 22782 5956 22838 6012
rect 22838 5956 22842 6012
rect 22778 5952 22842 5956
rect 22858 6012 22922 6016
rect 22858 5956 22862 6012
rect 22862 5956 22918 6012
rect 22918 5956 22922 6012
rect 22858 5952 22922 5956
rect 37062 6012 37126 6016
rect 37062 5956 37066 6012
rect 37066 5956 37122 6012
rect 37122 5956 37126 6012
rect 37062 5952 37126 5956
rect 37142 6012 37206 6016
rect 37142 5956 37146 6012
rect 37146 5956 37202 6012
rect 37202 5956 37206 6012
rect 37142 5952 37206 5956
rect 37222 6012 37286 6016
rect 37222 5956 37226 6012
rect 37226 5956 37282 6012
rect 37282 5956 37286 6012
rect 37222 5952 37286 5956
rect 37302 6012 37366 6016
rect 37302 5956 37306 6012
rect 37306 5956 37362 6012
rect 37362 5956 37366 6012
rect 37302 5952 37366 5956
rect 51506 6012 51570 6016
rect 51506 5956 51510 6012
rect 51510 5956 51566 6012
rect 51566 5956 51570 6012
rect 51506 5952 51570 5956
rect 51586 6012 51650 6016
rect 51586 5956 51590 6012
rect 51590 5956 51646 6012
rect 51646 5956 51650 6012
rect 51586 5952 51650 5956
rect 51666 6012 51730 6016
rect 51666 5956 51670 6012
rect 51670 5956 51726 6012
rect 51726 5956 51730 6012
rect 51666 5952 51730 5956
rect 51746 6012 51810 6016
rect 51746 5956 51750 6012
rect 51750 5956 51806 6012
rect 51806 5956 51810 6012
rect 51746 5952 51810 5956
rect 15396 5468 15460 5472
rect 15396 5412 15400 5468
rect 15400 5412 15456 5468
rect 15456 5412 15460 5468
rect 15396 5408 15460 5412
rect 15476 5468 15540 5472
rect 15476 5412 15480 5468
rect 15480 5412 15536 5468
rect 15536 5412 15540 5468
rect 15476 5408 15540 5412
rect 15556 5468 15620 5472
rect 15556 5412 15560 5468
rect 15560 5412 15616 5468
rect 15616 5412 15620 5468
rect 15556 5408 15620 5412
rect 15636 5468 15700 5472
rect 15636 5412 15640 5468
rect 15640 5412 15696 5468
rect 15696 5412 15700 5468
rect 15636 5408 15700 5412
rect 29840 5468 29904 5472
rect 29840 5412 29844 5468
rect 29844 5412 29900 5468
rect 29900 5412 29904 5468
rect 29840 5408 29904 5412
rect 29920 5468 29984 5472
rect 29920 5412 29924 5468
rect 29924 5412 29980 5468
rect 29980 5412 29984 5468
rect 29920 5408 29984 5412
rect 30000 5468 30064 5472
rect 30000 5412 30004 5468
rect 30004 5412 30060 5468
rect 30060 5412 30064 5468
rect 30000 5408 30064 5412
rect 30080 5468 30144 5472
rect 30080 5412 30084 5468
rect 30084 5412 30140 5468
rect 30140 5412 30144 5468
rect 30080 5408 30144 5412
rect 44284 5468 44348 5472
rect 44284 5412 44288 5468
rect 44288 5412 44344 5468
rect 44344 5412 44348 5468
rect 44284 5408 44348 5412
rect 44364 5468 44428 5472
rect 44364 5412 44368 5468
rect 44368 5412 44424 5468
rect 44424 5412 44428 5468
rect 44364 5408 44428 5412
rect 44444 5468 44508 5472
rect 44444 5412 44448 5468
rect 44448 5412 44504 5468
rect 44504 5412 44508 5468
rect 44444 5408 44508 5412
rect 44524 5468 44588 5472
rect 44524 5412 44528 5468
rect 44528 5412 44584 5468
rect 44584 5412 44588 5468
rect 44524 5408 44588 5412
rect 58728 5468 58792 5472
rect 58728 5412 58732 5468
rect 58732 5412 58788 5468
rect 58788 5412 58792 5468
rect 58728 5408 58792 5412
rect 58808 5468 58872 5472
rect 58808 5412 58812 5468
rect 58812 5412 58868 5468
rect 58868 5412 58872 5468
rect 58808 5408 58872 5412
rect 58888 5468 58952 5472
rect 58888 5412 58892 5468
rect 58892 5412 58948 5468
rect 58948 5412 58952 5468
rect 58888 5408 58952 5412
rect 58968 5468 59032 5472
rect 58968 5412 58972 5468
rect 58972 5412 59028 5468
rect 59028 5412 59032 5468
rect 58968 5408 59032 5412
rect 8174 4924 8238 4928
rect 8174 4868 8178 4924
rect 8178 4868 8234 4924
rect 8234 4868 8238 4924
rect 8174 4864 8238 4868
rect 8254 4924 8318 4928
rect 8254 4868 8258 4924
rect 8258 4868 8314 4924
rect 8314 4868 8318 4924
rect 8254 4864 8318 4868
rect 8334 4924 8398 4928
rect 8334 4868 8338 4924
rect 8338 4868 8394 4924
rect 8394 4868 8398 4924
rect 8334 4864 8398 4868
rect 8414 4924 8478 4928
rect 8414 4868 8418 4924
rect 8418 4868 8474 4924
rect 8474 4868 8478 4924
rect 8414 4864 8478 4868
rect 22618 4924 22682 4928
rect 22618 4868 22622 4924
rect 22622 4868 22678 4924
rect 22678 4868 22682 4924
rect 22618 4864 22682 4868
rect 22698 4924 22762 4928
rect 22698 4868 22702 4924
rect 22702 4868 22758 4924
rect 22758 4868 22762 4924
rect 22698 4864 22762 4868
rect 22778 4924 22842 4928
rect 22778 4868 22782 4924
rect 22782 4868 22838 4924
rect 22838 4868 22842 4924
rect 22778 4864 22842 4868
rect 22858 4924 22922 4928
rect 22858 4868 22862 4924
rect 22862 4868 22918 4924
rect 22918 4868 22922 4924
rect 22858 4864 22922 4868
rect 37062 4924 37126 4928
rect 37062 4868 37066 4924
rect 37066 4868 37122 4924
rect 37122 4868 37126 4924
rect 37062 4864 37126 4868
rect 37142 4924 37206 4928
rect 37142 4868 37146 4924
rect 37146 4868 37202 4924
rect 37202 4868 37206 4924
rect 37142 4864 37206 4868
rect 37222 4924 37286 4928
rect 37222 4868 37226 4924
rect 37226 4868 37282 4924
rect 37282 4868 37286 4924
rect 37222 4864 37286 4868
rect 37302 4924 37366 4928
rect 37302 4868 37306 4924
rect 37306 4868 37362 4924
rect 37362 4868 37366 4924
rect 37302 4864 37366 4868
rect 51506 4924 51570 4928
rect 51506 4868 51510 4924
rect 51510 4868 51566 4924
rect 51566 4868 51570 4924
rect 51506 4864 51570 4868
rect 51586 4924 51650 4928
rect 51586 4868 51590 4924
rect 51590 4868 51646 4924
rect 51646 4868 51650 4924
rect 51586 4864 51650 4868
rect 51666 4924 51730 4928
rect 51666 4868 51670 4924
rect 51670 4868 51726 4924
rect 51726 4868 51730 4924
rect 51666 4864 51730 4868
rect 51746 4924 51810 4928
rect 51746 4868 51750 4924
rect 51750 4868 51806 4924
rect 51806 4868 51810 4924
rect 51746 4864 51810 4868
rect 15396 4380 15460 4384
rect 15396 4324 15400 4380
rect 15400 4324 15456 4380
rect 15456 4324 15460 4380
rect 15396 4320 15460 4324
rect 15476 4380 15540 4384
rect 15476 4324 15480 4380
rect 15480 4324 15536 4380
rect 15536 4324 15540 4380
rect 15476 4320 15540 4324
rect 15556 4380 15620 4384
rect 15556 4324 15560 4380
rect 15560 4324 15616 4380
rect 15616 4324 15620 4380
rect 15556 4320 15620 4324
rect 15636 4380 15700 4384
rect 15636 4324 15640 4380
rect 15640 4324 15696 4380
rect 15696 4324 15700 4380
rect 15636 4320 15700 4324
rect 29840 4380 29904 4384
rect 29840 4324 29844 4380
rect 29844 4324 29900 4380
rect 29900 4324 29904 4380
rect 29840 4320 29904 4324
rect 29920 4380 29984 4384
rect 29920 4324 29924 4380
rect 29924 4324 29980 4380
rect 29980 4324 29984 4380
rect 29920 4320 29984 4324
rect 30000 4380 30064 4384
rect 30000 4324 30004 4380
rect 30004 4324 30060 4380
rect 30060 4324 30064 4380
rect 30000 4320 30064 4324
rect 30080 4380 30144 4384
rect 30080 4324 30084 4380
rect 30084 4324 30140 4380
rect 30140 4324 30144 4380
rect 30080 4320 30144 4324
rect 44284 4380 44348 4384
rect 44284 4324 44288 4380
rect 44288 4324 44344 4380
rect 44344 4324 44348 4380
rect 44284 4320 44348 4324
rect 44364 4380 44428 4384
rect 44364 4324 44368 4380
rect 44368 4324 44424 4380
rect 44424 4324 44428 4380
rect 44364 4320 44428 4324
rect 44444 4380 44508 4384
rect 44444 4324 44448 4380
rect 44448 4324 44504 4380
rect 44504 4324 44508 4380
rect 44444 4320 44508 4324
rect 44524 4380 44588 4384
rect 44524 4324 44528 4380
rect 44528 4324 44584 4380
rect 44584 4324 44588 4380
rect 44524 4320 44588 4324
rect 58728 4380 58792 4384
rect 58728 4324 58732 4380
rect 58732 4324 58788 4380
rect 58788 4324 58792 4380
rect 58728 4320 58792 4324
rect 58808 4380 58872 4384
rect 58808 4324 58812 4380
rect 58812 4324 58868 4380
rect 58868 4324 58872 4380
rect 58808 4320 58872 4324
rect 58888 4380 58952 4384
rect 58888 4324 58892 4380
rect 58892 4324 58948 4380
rect 58948 4324 58952 4380
rect 58888 4320 58952 4324
rect 58968 4380 59032 4384
rect 58968 4324 58972 4380
rect 58972 4324 59028 4380
rect 59028 4324 59032 4380
rect 58968 4320 59032 4324
rect 57100 4040 57164 4044
rect 57100 3984 57150 4040
rect 57150 3984 57164 4040
rect 57100 3980 57164 3984
rect 8174 3836 8238 3840
rect 8174 3780 8178 3836
rect 8178 3780 8234 3836
rect 8234 3780 8238 3836
rect 8174 3776 8238 3780
rect 8254 3836 8318 3840
rect 8254 3780 8258 3836
rect 8258 3780 8314 3836
rect 8314 3780 8318 3836
rect 8254 3776 8318 3780
rect 8334 3836 8398 3840
rect 8334 3780 8338 3836
rect 8338 3780 8394 3836
rect 8394 3780 8398 3836
rect 8334 3776 8398 3780
rect 8414 3836 8478 3840
rect 8414 3780 8418 3836
rect 8418 3780 8474 3836
rect 8474 3780 8478 3836
rect 8414 3776 8478 3780
rect 22618 3836 22682 3840
rect 22618 3780 22622 3836
rect 22622 3780 22678 3836
rect 22678 3780 22682 3836
rect 22618 3776 22682 3780
rect 22698 3836 22762 3840
rect 22698 3780 22702 3836
rect 22702 3780 22758 3836
rect 22758 3780 22762 3836
rect 22698 3776 22762 3780
rect 22778 3836 22842 3840
rect 22778 3780 22782 3836
rect 22782 3780 22838 3836
rect 22838 3780 22842 3836
rect 22778 3776 22842 3780
rect 22858 3836 22922 3840
rect 22858 3780 22862 3836
rect 22862 3780 22918 3836
rect 22918 3780 22922 3836
rect 22858 3776 22922 3780
rect 37062 3836 37126 3840
rect 37062 3780 37066 3836
rect 37066 3780 37122 3836
rect 37122 3780 37126 3836
rect 37062 3776 37126 3780
rect 37142 3836 37206 3840
rect 37142 3780 37146 3836
rect 37146 3780 37202 3836
rect 37202 3780 37206 3836
rect 37142 3776 37206 3780
rect 37222 3836 37286 3840
rect 37222 3780 37226 3836
rect 37226 3780 37282 3836
rect 37282 3780 37286 3836
rect 37222 3776 37286 3780
rect 37302 3836 37366 3840
rect 37302 3780 37306 3836
rect 37306 3780 37362 3836
rect 37362 3780 37366 3836
rect 37302 3776 37366 3780
rect 51506 3836 51570 3840
rect 51506 3780 51510 3836
rect 51510 3780 51566 3836
rect 51566 3780 51570 3836
rect 51506 3776 51570 3780
rect 51586 3836 51650 3840
rect 51586 3780 51590 3836
rect 51590 3780 51646 3836
rect 51646 3780 51650 3836
rect 51586 3776 51650 3780
rect 51666 3836 51730 3840
rect 51666 3780 51670 3836
rect 51670 3780 51726 3836
rect 51726 3780 51730 3836
rect 51666 3776 51730 3780
rect 51746 3836 51810 3840
rect 51746 3780 51750 3836
rect 51750 3780 51806 3836
rect 51806 3780 51810 3836
rect 51746 3776 51810 3780
rect 15396 3292 15460 3296
rect 15396 3236 15400 3292
rect 15400 3236 15456 3292
rect 15456 3236 15460 3292
rect 15396 3232 15460 3236
rect 15476 3292 15540 3296
rect 15476 3236 15480 3292
rect 15480 3236 15536 3292
rect 15536 3236 15540 3292
rect 15476 3232 15540 3236
rect 15556 3292 15620 3296
rect 15556 3236 15560 3292
rect 15560 3236 15616 3292
rect 15616 3236 15620 3292
rect 15556 3232 15620 3236
rect 15636 3292 15700 3296
rect 15636 3236 15640 3292
rect 15640 3236 15696 3292
rect 15696 3236 15700 3292
rect 15636 3232 15700 3236
rect 29840 3292 29904 3296
rect 29840 3236 29844 3292
rect 29844 3236 29900 3292
rect 29900 3236 29904 3292
rect 29840 3232 29904 3236
rect 29920 3292 29984 3296
rect 29920 3236 29924 3292
rect 29924 3236 29980 3292
rect 29980 3236 29984 3292
rect 29920 3232 29984 3236
rect 30000 3292 30064 3296
rect 30000 3236 30004 3292
rect 30004 3236 30060 3292
rect 30060 3236 30064 3292
rect 30000 3232 30064 3236
rect 30080 3292 30144 3296
rect 30080 3236 30084 3292
rect 30084 3236 30140 3292
rect 30140 3236 30144 3292
rect 30080 3232 30144 3236
rect 44284 3292 44348 3296
rect 44284 3236 44288 3292
rect 44288 3236 44344 3292
rect 44344 3236 44348 3292
rect 44284 3232 44348 3236
rect 44364 3292 44428 3296
rect 44364 3236 44368 3292
rect 44368 3236 44424 3292
rect 44424 3236 44428 3292
rect 44364 3232 44428 3236
rect 44444 3292 44508 3296
rect 44444 3236 44448 3292
rect 44448 3236 44504 3292
rect 44504 3236 44508 3292
rect 44444 3232 44508 3236
rect 44524 3292 44588 3296
rect 44524 3236 44528 3292
rect 44528 3236 44584 3292
rect 44584 3236 44588 3292
rect 44524 3232 44588 3236
rect 58728 3292 58792 3296
rect 58728 3236 58732 3292
rect 58732 3236 58788 3292
rect 58788 3236 58792 3292
rect 58728 3232 58792 3236
rect 58808 3292 58872 3296
rect 58808 3236 58812 3292
rect 58812 3236 58868 3292
rect 58868 3236 58872 3292
rect 58808 3232 58872 3236
rect 58888 3292 58952 3296
rect 58888 3236 58892 3292
rect 58892 3236 58948 3292
rect 58948 3236 58952 3292
rect 58888 3232 58952 3236
rect 58968 3292 59032 3296
rect 58968 3236 58972 3292
rect 58972 3236 59028 3292
rect 59028 3236 59032 3292
rect 58968 3232 59032 3236
rect 8174 2748 8238 2752
rect 8174 2692 8178 2748
rect 8178 2692 8234 2748
rect 8234 2692 8238 2748
rect 8174 2688 8238 2692
rect 8254 2748 8318 2752
rect 8254 2692 8258 2748
rect 8258 2692 8314 2748
rect 8314 2692 8318 2748
rect 8254 2688 8318 2692
rect 8334 2748 8398 2752
rect 8334 2692 8338 2748
rect 8338 2692 8394 2748
rect 8394 2692 8398 2748
rect 8334 2688 8398 2692
rect 8414 2748 8478 2752
rect 8414 2692 8418 2748
rect 8418 2692 8474 2748
rect 8474 2692 8478 2748
rect 8414 2688 8478 2692
rect 22618 2748 22682 2752
rect 22618 2692 22622 2748
rect 22622 2692 22678 2748
rect 22678 2692 22682 2748
rect 22618 2688 22682 2692
rect 22698 2748 22762 2752
rect 22698 2692 22702 2748
rect 22702 2692 22758 2748
rect 22758 2692 22762 2748
rect 22698 2688 22762 2692
rect 22778 2748 22842 2752
rect 22778 2692 22782 2748
rect 22782 2692 22838 2748
rect 22838 2692 22842 2748
rect 22778 2688 22842 2692
rect 22858 2748 22922 2752
rect 22858 2692 22862 2748
rect 22862 2692 22918 2748
rect 22918 2692 22922 2748
rect 22858 2688 22922 2692
rect 37062 2748 37126 2752
rect 37062 2692 37066 2748
rect 37066 2692 37122 2748
rect 37122 2692 37126 2748
rect 37062 2688 37126 2692
rect 37142 2748 37206 2752
rect 37142 2692 37146 2748
rect 37146 2692 37202 2748
rect 37202 2692 37206 2748
rect 37142 2688 37206 2692
rect 37222 2748 37286 2752
rect 37222 2692 37226 2748
rect 37226 2692 37282 2748
rect 37282 2692 37286 2748
rect 37222 2688 37286 2692
rect 37302 2748 37366 2752
rect 37302 2692 37306 2748
rect 37306 2692 37362 2748
rect 37362 2692 37366 2748
rect 37302 2688 37366 2692
rect 51506 2748 51570 2752
rect 51506 2692 51510 2748
rect 51510 2692 51566 2748
rect 51566 2692 51570 2748
rect 51506 2688 51570 2692
rect 51586 2748 51650 2752
rect 51586 2692 51590 2748
rect 51590 2692 51646 2748
rect 51646 2692 51650 2748
rect 51586 2688 51650 2692
rect 51666 2748 51730 2752
rect 51666 2692 51670 2748
rect 51670 2692 51726 2748
rect 51726 2692 51730 2748
rect 51666 2688 51730 2692
rect 51746 2748 51810 2752
rect 51746 2692 51750 2748
rect 51750 2692 51806 2748
rect 51806 2692 51810 2748
rect 51746 2688 51810 2692
rect 15396 2204 15460 2208
rect 15396 2148 15400 2204
rect 15400 2148 15456 2204
rect 15456 2148 15460 2204
rect 15396 2144 15460 2148
rect 15476 2204 15540 2208
rect 15476 2148 15480 2204
rect 15480 2148 15536 2204
rect 15536 2148 15540 2204
rect 15476 2144 15540 2148
rect 15556 2204 15620 2208
rect 15556 2148 15560 2204
rect 15560 2148 15616 2204
rect 15616 2148 15620 2204
rect 15556 2144 15620 2148
rect 15636 2204 15700 2208
rect 15636 2148 15640 2204
rect 15640 2148 15696 2204
rect 15696 2148 15700 2204
rect 15636 2144 15700 2148
rect 29840 2204 29904 2208
rect 29840 2148 29844 2204
rect 29844 2148 29900 2204
rect 29900 2148 29904 2204
rect 29840 2144 29904 2148
rect 29920 2204 29984 2208
rect 29920 2148 29924 2204
rect 29924 2148 29980 2204
rect 29980 2148 29984 2204
rect 29920 2144 29984 2148
rect 30000 2204 30064 2208
rect 30000 2148 30004 2204
rect 30004 2148 30060 2204
rect 30060 2148 30064 2204
rect 30000 2144 30064 2148
rect 30080 2204 30144 2208
rect 30080 2148 30084 2204
rect 30084 2148 30140 2204
rect 30140 2148 30144 2204
rect 30080 2144 30144 2148
rect 44284 2204 44348 2208
rect 44284 2148 44288 2204
rect 44288 2148 44344 2204
rect 44344 2148 44348 2204
rect 44284 2144 44348 2148
rect 44364 2204 44428 2208
rect 44364 2148 44368 2204
rect 44368 2148 44424 2204
rect 44424 2148 44428 2204
rect 44364 2144 44428 2148
rect 44444 2204 44508 2208
rect 44444 2148 44448 2204
rect 44448 2148 44504 2204
rect 44504 2148 44508 2204
rect 44444 2144 44508 2148
rect 44524 2204 44588 2208
rect 44524 2148 44528 2204
rect 44528 2148 44584 2204
rect 44584 2148 44588 2204
rect 44524 2144 44588 2148
rect 58728 2204 58792 2208
rect 58728 2148 58732 2204
rect 58732 2148 58788 2204
rect 58788 2148 58792 2204
rect 58728 2144 58792 2148
rect 58808 2204 58872 2208
rect 58808 2148 58812 2204
rect 58812 2148 58868 2204
rect 58868 2148 58872 2204
rect 58808 2144 58872 2148
rect 58888 2204 58952 2208
rect 58888 2148 58892 2204
rect 58892 2148 58948 2204
rect 58948 2148 58952 2204
rect 58888 2144 58952 2148
rect 58968 2204 59032 2208
rect 58968 2148 58972 2204
rect 58972 2148 59028 2204
rect 59028 2148 59032 2204
rect 58968 2144 59032 2148
<< metal4 >>
rect 8166 27776 8486 27792
rect 8166 27712 8174 27776
rect 8238 27712 8254 27776
rect 8318 27712 8334 27776
rect 8398 27712 8414 27776
rect 8478 27712 8486 27776
rect 8166 26688 8486 27712
rect 8166 26624 8174 26688
rect 8238 26624 8254 26688
rect 8318 26624 8334 26688
rect 8398 26624 8414 26688
rect 8478 26624 8486 26688
rect 8166 25600 8486 26624
rect 8166 25536 8174 25600
rect 8238 25536 8254 25600
rect 8318 25536 8334 25600
rect 8398 25536 8414 25600
rect 8478 25536 8486 25600
rect 8166 24512 8486 25536
rect 8166 24448 8174 24512
rect 8238 24448 8254 24512
rect 8318 24448 8334 24512
rect 8398 24448 8414 24512
rect 8478 24448 8486 24512
rect 8166 23424 8486 24448
rect 8166 23360 8174 23424
rect 8238 23360 8254 23424
rect 8318 23360 8334 23424
rect 8398 23360 8414 23424
rect 8478 23360 8486 23424
rect 8166 22336 8486 23360
rect 8166 22272 8174 22336
rect 8238 22272 8254 22336
rect 8318 22272 8334 22336
rect 8398 22272 8414 22336
rect 8478 22272 8486 22336
rect 8166 21248 8486 22272
rect 8166 21184 8174 21248
rect 8238 21184 8254 21248
rect 8318 21184 8334 21248
rect 8398 21184 8414 21248
rect 8478 21184 8486 21248
rect 8166 20160 8486 21184
rect 8166 20096 8174 20160
rect 8238 20096 8254 20160
rect 8318 20096 8334 20160
rect 8398 20096 8414 20160
rect 8478 20096 8486 20160
rect 8166 19072 8486 20096
rect 8166 19008 8174 19072
rect 8238 19008 8254 19072
rect 8318 19008 8334 19072
rect 8398 19008 8414 19072
rect 8478 19008 8486 19072
rect 8166 17984 8486 19008
rect 8166 17920 8174 17984
rect 8238 17920 8254 17984
rect 8318 17920 8334 17984
rect 8398 17920 8414 17984
rect 8478 17920 8486 17984
rect 8166 16896 8486 17920
rect 8166 16832 8174 16896
rect 8238 16832 8254 16896
rect 8318 16832 8334 16896
rect 8398 16832 8414 16896
rect 8478 16832 8486 16896
rect 8166 15808 8486 16832
rect 8166 15744 8174 15808
rect 8238 15744 8254 15808
rect 8318 15744 8334 15808
rect 8398 15744 8414 15808
rect 8478 15744 8486 15808
rect 8166 14720 8486 15744
rect 8166 14656 8174 14720
rect 8238 14656 8254 14720
rect 8318 14656 8334 14720
rect 8398 14656 8414 14720
rect 8478 14656 8486 14720
rect 8166 13632 8486 14656
rect 8166 13568 8174 13632
rect 8238 13568 8254 13632
rect 8318 13568 8334 13632
rect 8398 13568 8414 13632
rect 8478 13568 8486 13632
rect 8166 12544 8486 13568
rect 8166 12480 8174 12544
rect 8238 12480 8254 12544
rect 8318 12480 8334 12544
rect 8398 12480 8414 12544
rect 8478 12480 8486 12544
rect 8166 11456 8486 12480
rect 8166 11392 8174 11456
rect 8238 11392 8254 11456
rect 8318 11392 8334 11456
rect 8398 11392 8414 11456
rect 8478 11392 8486 11456
rect 8166 10368 8486 11392
rect 8166 10304 8174 10368
rect 8238 10304 8254 10368
rect 8318 10304 8334 10368
rect 8398 10304 8414 10368
rect 8478 10304 8486 10368
rect 8166 9280 8486 10304
rect 8166 9216 8174 9280
rect 8238 9216 8254 9280
rect 8318 9216 8334 9280
rect 8398 9216 8414 9280
rect 8478 9216 8486 9280
rect 8166 8192 8486 9216
rect 8166 8128 8174 8192
rect 8238 8128 8254 8192
rect 8318 8128 8334 8192
rect 8398 8128 8414 8192
rect 8478 8128 8486 8192
rect 8166 7104 8486 8128
rect 8166 7040 8174 7104
rect 8238 7040 8254 7104
rect 8318 7040 8334 7104
rect 8398 7040 8414 7104
rect 8478 7040 8486 7104
rect 8166 6016 8486 7040
rect 8166 5952 8174 6016
rect 8238 5952 8254 6016
rect 8318 5952 8334 6016
rect 8398 5952 8414 6016
rect 8478 5952 8486 6016
rect 8166 4928 8486 5952
rect 8166 4864 8174 4928
rect 8238 4864 8254 4928
rect 8318 4864 8334 4928
rect 8398 4864 8414 4928
rect 8478 4864 8486 4928
rect 8166 3840 8486 4864
rect 8166 3776 8174 3840
rect 8238 3776 8254 3840
rect 8318 3776 8334 3840
rect 8398 3776 8414 3840
rect 8478 3776 8486 3840
rect 8166 2752 8486 3776
rect 8166 2688 8174 2752
rect 8238 2688 8254 2752
rect 8318 2688 8334 2752
rect 8398 2688 8414 2752
rect 8478 2688 8486 2752
rect 8166 2128 8486 2688
rect 15388 27232 15708 27792
rect 15388 27168 15396 27232
rect 15460 27168 15476 27232
rect 15540 27168 15556 27232
rect 15620 27168 15636 27232
rect 15700 27168 15708 27232
rect 15388 26144 15708 27168
rect 15388 26080 15396 26144
rect 15460 26080 15476 26144
rect 15540 26080 15556 26144
rect 15620 26080 15636 26144
rect 15700 26080 15708 26144
rect 15388 25056 15708 26080
rect 15388 24992 15396 25056
rect 15460 24992 15476 25056
rect 15540 24992 15556 25056
rect 15620 24992 15636 25056
rect 15700 24992 15708 25056
rect 15388 23968 15708 24992
rect 15388 23904 15396 23968
rect 15460 23904 15476 23968
rect 15540 23904 15556 23968
rect 15620 23904 15636 23968
rect 15700 23904 15708 23968
rect 15388 22880 15708 23904
rect 15388 22816 15396 22880
rect 15460 22816 15476 22880
rect 15540 22816 15556 22880
rect 15620 22816 15636 22880
rect 15700 22816 15708 22880
rect 15388 21792 15708 22816
rect 15388 21728 15396 21792
rect 15460 21728 15476 21792
rect 15540 21728 15556 21792
rect 15620 21728 15636 21792
rect 15700 21728 15708 21792
rect 15388 20704 15708 21728
rect 15388 20640 15396 20704
rect 15460 20640 15476 20704
rect 15540 20640 15556 20704
rect 15620 20640 15636 20704
rect 15700 20640 15708 20704
rect 15388 19616 15708 20640
rect 15388 19552 15396 19616
rect 15460 19552 15476 19616
rect 15540 19552 15556 19616
rect 15620 19552 15636 19616
rect 15700 19552 15708 19616
rect 15388 18528 15708 19552
rect 15388 18464 15396 18528
rect 15460 18464 15476 18528
rect 15540 18464 15556 18528
rect 15620 18464 15636 18528
rect 15700 18464 15708 18528
rect 15388 17440 15708 18464
rect 15388 17376 15396 17440
rect 15460 17376 15476 17440
rect 15540 17376 15556 17440
rect 15620 17376 15636 17440
rect 15700 17376 15708 17440
rect 15388 16352 15708 17376
rect 15388 16288 15396 16352
rect 15460 16288 15476 16352
rect 15540 16288 15556 16352
rect 15620 16288 15636 16352
rect 15700 16288 15708 16352
rect 15388 15264 15708 16288
rect 15388 15200 15396 15264
rect 15460 15200 15476 15264
rect 15540 15200 15556 15264
rect 15620 15200 15636 15264
rect 15700 15200 15708 15264
rect 15388 14176 15708 15200
rect 15388 14112 15396 14176
rect 15460 14112 15476 14176
rect 15540 14112 15556 14176
rect 15620 14112 15636 14176
rect 15700 14112 15708 14176
rect 15388 13088 15708 14112
rect 15388 13024 15396 13088
rect 15460 13024 15476 13088
rect 15540 13024 15556 13088
rect 15620 13024 15636 13088
rect 15700 13024 15708 13088
rect 15388 12000 15708 13024
rect 15388 11936 15396 12000
rect 15460 11936 15476 12000
rect 15540 11936 15556 12000
rect 15620 11936 15636 12000
rect 15700 11936 15708 12000
rect 15388 10912 15708 11936
rect 15388 10848 15396 10912
rect 15460 10848 15476 10912
rect 15540 10848 15556 10912
rect 15620 10848 15636 10912
rect 15700 10848 15708 10912
rect 15388 9824 15708 10848
rect 15388 9760 15396 9824
rect 15460 9760 15476 9824
rect 15540 9760 15556 9824
rect 15620 9760 15636 9824
rect 15700 9760 15708 9824
rect 15388 8736 15708 9760
rect 15388 8672 15396 8736
rect 15460 8672 15476 8736
rect 15540 8672 15556 8736
rect 15620 8672 15636 8736
rect 15700 8672 15708 8736
rect 15388 7648 15708 8672
rect 15388 7584 15396 7648
rect 15460 7584 15476 7648
rect 15540 7584 15556 7648
rect 15620 7584 15636 7648
rect 15700 7584 15708 7648
rect 15388 6560 15708 7584
rect 15388 6496 15396 6560
rect 15460 6496 15476 6560
rect 15540 6496 15556 6560
rect 15620 6496 15636 6560
rect 15700 6496 15708 6560
rect 15388 5472 15708 6496
rect 15388 5408 15396 5472
rect 15460 5408 15476 5472
rect 15540 5408 15556 5472
rect 15620 5408 15636 5472
rect 15700 5408 15708 5472
rect 15388 4384 15708 5408
rect 15388 4320 15396 4384
rect 15460 4320 15476 4384
rect 15540 4320 15556 4384
rect 15620 4320 15636 4384
rect 15700 4320 15708 4384
rect 15388 3296 15708 4320
rect 15388 3232 15396 3296
rect 15460 3232 15476 3296
rect 15540 3232 15556 3296
rect 15620 3232 15636 3296
rect 15700 3232 15708 3296
rect 15388 2208 15708 3232
rect 15388 2144 15396 2208
rect 15460 2144 15476 2208
rect 15540 2144 15556 2208
rect 15620 2144 15636 2208
rect 15700 2144 15708 2208
rect 15388 2128 15708 2144
rect 22610 27776 22930 27792
rect 22610 27712 22618 27776
rect 22682 27712 22698 27776
rect 22762 27712 22778 27776
rect 22842 27712 22858 27776
rect 22922 27712 22930 27776
rect 22610 26688 22930 27712
rect 22610 26624 22618 26688
rect 22682 26624 22698 26688
rect 22762 26624 22778 26688
rect 22842 26624 22858 26688
rect 22922 26624 22930 26688
rect 22610 25600 22930 26624
rect 22610 25536 22618 25600
rect 22682 25536 22698 25600
rect 22762 25536 22778 25600
rect 22842 25536 22858 25600
rect 22922 25536 22930 25600
rect 22610 24512 22930 25536
rect 22610 24448 22618 24512
rect 22682 24448 22698 24512
rect 22762 24448 22778 24512
rect 22842 24448 22858 24512
rect 22922 24448 22930 24512
rect 22610 23424 22930 24448
rect 22610 23360 22618 23424
rect 22682 23360 22698 23424
rect 22762 23360 22778 23424
rect 22842 23360 22858 23424
rect 22922 23360 22930 23424
rect 22610 22336 22930 23360
rect 22610 22272 22618 22336
rect 22682 22272 22698 22336
rect 22762 22272 22778 22336
rect 22842 22272 22858 22336
rect 22922 22272 22930 22336
rect 22610 21248 22930 22272
rect 22610 21184 22618 21248
rect 22682 21184 22698 21248
rect 22762 21184 22778 21248
rect 22842 21184 22858 21248
rect 22922 21184 22930 21248
rect 22610 20160 22930 21184
rect 22610 20096 22618 20160
rect 22682 20096 22698 20160
rect 22762 20096 22778 20160
rect 22842 20096 22858 20160
rect 22922 20096 22930 20160
rect 22610 19072 22930 20096
rect 22610 19008 22618 19072
rect 22682 19008 22698 19072
rect 22762 19008 22778 19072
rect 22842 19008 22858 19072
rect 22922 19008 22930 19072
rect 22610 17984 22930 19008
rect 22610 17920 22618 17984
rect 22682 17920 22698 17984
rect 22762 17920 22778 17984
rect 22842 17920 22858 17984
rect 22922 17920 22930 17984
rect 22610 16896 22930 17920
rect 22610 16832 22618 16896
rect 22682 16832 22698 16896
rect 22762 16832 22778 16896
rect 22842 16832 22858 16896
rect 22922 16832 22930 16896
rect 22610 15808 22930 16832
rect 22610 15744 22618 15808
rect 22682 15744 22698 15808
rect 22762 15744 22778 15808
rect 22842 15744 22858 15808
rect 22922 15744 22930 15808
rect 22610 14720 22930 15744
rect 22610 14656 22618 14720
rect 22682 14656 22698 14720
rect 22762 14656 22778 14720
rect 22842 14656 22858 14720
rect 22922 14656 22930 14720
rect 22610 13632 22930 14656
rect 22610 13568 22618 13632
rect 22682 13568 22698 13632
rect 22762 13568 22778 13632
rect 22842 13568 22858 13632
rect 22922 13568 22930 13632
rect 22610 12544 22930 13568
rect 22610 12480 22618 12544
rect 22682 12480 22698 12544
rect 22762 12480 22778 12544
rect 22842 12480 22858 12544
rect 22922 12480 22930 12544
rect 22610 11456 22930 12480
rect 22610 11392 22618 11456
rect 22682 11392 22698 11456
rect 22762 11392 22778 11456
rect 22842 11392 22858 11456
rect 22922 11392 22930 11456
rect 22610 10368 22930 11392
rect 22610 10304 22618 10368
rect 22682 10304 22698 10368
rect 22762 10304 22778 10368
rect 22842 10304 22858 10368
rect 22922 10304 22930 10368
rect 22610 9280 22930 10304
rect 22610 9216 22618 9280
rect 22682 9216 22698 9280
rect 22762 9216 22778 9280
rect 22842 9216 22858 9280
rect 22922 9216 22930 9280
rect 22610 8192 22930 9216
rect 22610 8128 22618 8192
rect 22682 8128 22698 8192
rect 22762 8128 22778 8192
rect 22842 8128 22858 8192
rect 22922 8128 22930 8192
rect 22610 7104 22930 8128
rect 22610 7040 22618 7104
rect 22682 7040 22698 7104
rect 22762 7040 22778 7104
rect 22842 7040 22858 7104
rect 22922 7040 22930 7104
rect 22610 6016 22930 7040
rect 22610 5952 22618 6016
rect 22682 5952 22698 6016
rect 22762 5952 22778 6016
rect 22842 5952 22858 6016
rect 22922 5952 22930 6016
rect 22610 4928 22930 5952
rect 22610 4864 22618 4928
rect 22682 4864 22698 4928
rect 22762 4864 22778 4928
rect 22842 4864 22858 4928
rect 22922 4864 22930 4928
rect 22610 3840 22930 4864
rect 22610 3776 22618 3840
rect 22682 3776 22698 3840
rect 22762 3776 22778 3840
rect 22842 3776 22858 3840
rect 22922 3776 22930 3840
rect 22610 2752 22930 3776
rect 22610 2688 22618 2752
rect 22682 2688 22698 2752
rect 22762 2688 22778 2752
rect 22842 2688 22858 2752
rect 22922 2688 22930 2752
rect 22610 2128 22930 2688
rect 29832 27232 30152 27792
rect 29832 27168 29840 27232
rect 29904 27168 29920 27232
rect 29984 27168 30000 27232
rect 30064 27168 30080 27232
rect 30144 27168 30152 27232
rect 29832 26144 30152 27168
rect 29832 26080 29840 26144
rect 29904 26080 29920 26144
rect 29984 26080 30000 26144
rect 30064 26080 30080 26144
rect 30144 26080 30152 26144
rect 29832 25056 30152 26080
rect 29832 24992 29840 25056
rect 29904 24992 29920 25056
rect 29984 24992 30000 25056
rect 30064 24992 30080 25056
rect 30144 24992 30152 25056
rect 29832 23968 30152 24992
rect 29832 23904 29840 23968
rect 29904 23904 29920 23968
rect 29984 23904 30000 23968
rect 30064 23904 30080 23968
rect 30144 23904 30152 23968
rect 29832 22880 30152 23904
rect 29832 22816 29840 22880
rect 29904 22816 29920 22880
rect 29984 22816 30000 22880
rect 30064 22816 30080 22880
rect 30144 22816 30152 22880
rect 29832 21792 30152 22816
rect 29832 21728 29840 21792
rect 29904 21728 29920 21792
rect 29984 21728 30000 21792
rect 30064 21728 30080 21792
rect 30144 21728 30152 21792
rect 29832 20704 30152 21728
rect 29832 20640 29840 20704
rect 29904 20640 29920 20704
rect 29984 20640 30000 20704
rect 30064 20640 30080 20704
rect 30144 20640 30152 20704
rect 29832 19616 30152 20640
rect 29832 19552 29840 19616
rect 29904 19552 29920 19616
rect 29984 19552 30000 19616
rect 30064 19552 30080 19616
rect 30144 19552 30152 19616
rect 29832 18528 30152 19552
rect 29832 18464 29840 18528
rect 29904 18464 29920 18528
rect 29984 18464 30000 18528
rect 30064 18464 30080 18528
rect 30144 18464 30152 18528
rect 29832 17440 30152 18464
rect 29832 17376 29840 17440
rect 29904 17376 29920 17440
rect 29984 17376 30000 17440
rect 30064 17376 30080 17440
rect 30144 17376 30152 17440
rect 29832 16352 30152 17376
rect 29832 16288 29840 16352
rect 29904 16288 29920 16352
rect 29984 16288 30000 16352
rect 30064 16288 30080 16352
rect 30144 16288 30152 16352
rect 29832 15264 30152 16288
rect 29832 15200 29840 15264
rect 29904 15200 29920 15264
rect 29984 15200 30000 15264
rect 30064 15200 30080 15264
rect 30144 15200 30152 15264
rect 29832 14176 30152 15200
rect 29832 14112 29840 14176
rect 29904 14112 29920 14176
rect 29984 14112 30000 14176
rect 30064 14112 30080 14176
rect 30144 14112 30152 14176
rect 29832 13088 30152 14112
rect 29832 13024 29840 13088
rect 29904 13024 29920 13088
rect 29984 13024 30000 13088
rect 30064 13024 30080 13088
rect 30144 13024 30152 13088
rect 29832 12000 30152 13024
rect 29832 11936 29840 12000
rect 29904 11936 29920 12000
rect 29984 11936 30000 12000
rect 30064 11936 30080 12000
rect 30144 11936 30152 12000
rect 29832 10912 30152 11936
rect 29832 10848 29840 10912
rect 29904 10848 29920 10912
rect 29984 10848 30000 10912
rect 30064 10848 30080 10912
rect 30144 10848 30152 10912
rect 29832 9824 30152 10848
rect 29832 9760 29840 9824
rect 29904 9760 29920 9824
rect 29984 9760 30000 9824
rect 30064 9760 30080 9824
rect 30144 9760 30152 9824
rect 29832 8736 30152 9760
rect 29832 8672 29840 8736
rect 29904 8672 29920 8736
rect 29984 8672 30000 8736
rect 30064 8672 30080 8736
rect 30144 8672 30152 8736
rect 29832 7648 30152 8672
rect 29832 7584 29840 7648
rect 29904 7584 29920 7648
rect 29984 7584 30000 7648
rect 30064 7584 30080 7648
rect 30144 7584 30152 7648
rect 29832 6560 30152 7584
rect 29832 6496 29840 6560
rect 29904 6496 29920 6560
rect 29984 6496 30000 6560
rect 30064 6496 30080 6560
rect 30144 6496 30152 6560
rect 29832 5472 30152 6496
rect 29832 5408 29840 5472
rect 29904 5408 29920 5472
rect 29984 5408 30000 5472
rect 30064 5408 30080 5472
rect 30144 5408 30152 5472
rect 29832 4384 30152 5408
rect 29832 4320 29840 4384
rect 29904 4320 29920 4384
rect 29984 4320 30000 4384
rect 30064 4320 30080 4384
rect 30144 4320 30152 4384
rect 29832 3296 30152 4320
rect 29832 3232 29840 3296
rect 29904 3232 29920 3296
rect 29984 3232 30000 3296
rect 30064 3232 30080 3296
rect 30144 3232 30152 3296
rect 29832 2208 30152 3232
rect 29832 2144 29840 2208
rect 29904 2144 29920 2208
rect 29984 2144 30000 2208
rect 30064 2144 30080 2208
rect 30144 2144 30152 2208
rect 29832 2128 30152 2144
rect 37054 27776 37374 27792
rect 37054 27712 37062 27776
rect 37126 27712 37142 27776
rect 37206 27712 37222 27776
rect 37286 27712 37302 27776
rect 37366 27712 37374 27776
rect 37054 26688 37374 27712
rect 37054 26624 37062 26688
rect 37126 26624 37142 26688
rect 37206 26624 37222 26688
rect 37286 26624 37302 26688
rect 37366 26624 37374 26688
rect 37054 25600 37374 26624
rect 37054 25536 37062 25600
rect 37126 25536 37142 25600
rect 37206 25536 37222 25600
rect 37286 25536 37302 25600
rect 37366 25536 37374 25600
rect 37054 24512 37374 25536
rect 37054 24448 37062 24512
rect 37126 24448 37142 24512
rect 37206 24448 37222 24512
rect 37286 24448 37302 24512
rect 37366 24448 37374 24512
rect 37054 23424 37374 24448
rect 37054 23360 37062 23424
rect 37126 23360 37142 23424
rect 37206 23360 37222 23424
rect 37286 23360 37302 23424
rect 37366 23360 37374 23424
rect 37054 22336 37374 23360
rect 37054 22272 37062 22336
rect 37126 22272 37142 22336
rect 37206 22272 37222 22336
rect 37286 22272 37302 22336
rect 37366 22272 37374 22336
rect 37054 21248 37374 22272
rect 37054 21184 37062 21248
rect 37126 21184 37142 21248
rect 37206 21184 37222 21248
rect 37286 21184 37302 21248
rect 37366 21184 37374 21248
rect 37054 20160 37374 21184
rect 37054 20096 37062 20160
rect 37126 20096 37142 20160
rect 37206 20096 37222 20160
rect 37286 20096 37302 20160
rect 37366 20096 37374 20160
rect 37054 19072 37374 20096
rect 37054 19008 37062 19072
rect 37126 19008 37142 19072
rect 37206 19008 37222 19072
rect 37286 19008 37302 19072
rect 37366 19008 37374 19072
rect 37054 17984 37374 19008
rect 37054 17920 37062 17984
rect 37126 17920 37142 17984
rect 37206 17920 37222 17984
rect 37286 17920 37302 17984
rect 37366 17920 37374 17984
rect 37054 16896 37374 17920
rect 37054 16832 37062 16896
rect 37126 16832 37142 16896
rect 37206 16832 37222 16896
rect 37286 16832 37302 16896
rect 37366 16832 37374 16896
rect 37054 15808 37374 16832
rect 37054 15744 37062 15808
rect 37126 15744 37142 15808
rect 37206 15744 37222 15808
rect 37286 15744 37302 15808
rect 37366 15744 37374 15808
rect 37054 14720 37374 15744
rect 37054 14656 37062 14720
rect 37126 14656 37142 14720
rect 37206 14656 37222 14720
rect 37286 14656 37302 14720
rect 37366 14656 37374 14720
rect 37054 13632 37374 14656
rect 37054 13568 37062 13632
rect 37126 13568 37142 13632
rect 37206 13568 37222 13632
rect 37286 13568 37302 13632
rect 37366 13568 37374 13632
rect 37054 12544 37374 13568
rect 37054 12480 37062 12544
rect 37126 12480 37142 12544
rect 37206 12480 37222 12544
rect 37286 12480 37302 12544
rect 37366 12480 37374 12544
rect 37054 11456 37374 12480
rect 37054 11392 37062 11456
rect 37126 11392 37142 11456
rect 37206 11392 37222 11456
rect 37286 11392 37302 11456
rect 37366 11392 37374 11456
rect 37054 10368 37374 11392
rect 37054 10304 37062 10368
rect 37126 10304 37142 10368
rect 37206 10304 37222 10368
rect 37286 10304 37302 10368
rect 37366 10304 37374 10368
rect 37054 9280 37374 10304
rect 37054 9216 37062 9280
rect 37126 9216 37142 9280
rect 37206 9216 37222 9280
rect 37286 9216 37302 9280
rect 37366 9216 37374 9280
rect 37054 8192 37374 9216
rect 37054 8128 37062 8192
rect 37126 8128 37142 8192
rect 37206 8128 37222 8192
rect 37286 8128 37302 8192
rect 37366 8128 37374 8192
rect 37054 7104 37374 8128
rect 37054 7040 37062 7104
rect 37126 7040 37142 7104
rect 37206 7040 37222 7104
rect 37286 7040 37302 7104
rect 37366 7040 37374 7104
rect 37054 6016 37374 7040
rect 37054 5952 37062 6016
rect 37126 5952 37142 6016
rect 37206 5952 37222 6016
rect 37286 5952 37302 6016
rect 37366 5952 37374 6016
rect 37054 4928 37374 5952
rect 37054 4864 37062 4928
rect 37126 4864 37142 4928
rect 37206 4864 37222 4928
rect 37286 4864 37302 4928
rect 37366 4864 37374 4928
rect 37054 3840 37374 4864
rect 37054 3776 37062 3840
rect 37126 3776 37142 3840
rect 37206 3776 37222 3840
rect 37286 3776 37302 3840
rect 37366 3776 37374 3840
rect 37054 2752 37374 3776
rect 37054 2688 37062 2752
rect 37126 2688 37142 2752
rect 37206 2688 37222 2752
rect 37286 2688 37302 2752
rect 37366 2688 37374 2752
rect 37054 2128 37374 2688
rect 44276 27232 44596 27792
rect 44276 27168 44284 27232
rect 44348 27168 44364 27232
rect 44428 27168 44444 27232
rect 44508 27168 44524 27232
rect 44588 27168 44596 27232
rect 44276 26144 44596 27168
rect 44276 26080 44284 26144
rect 44348 26080 44364 26144
rect 44428 26080 44444 26144
rect 44508 26080 44524 26144
rect 44588 26080 44596 26144
rect 44276 25056 44596 26080
rect 44276 24992 44284 25056
rect 44348 24992 44364 25056
rect 44428 24992 44444 25056
rect 44508 24992 44524 25056
rect 44588 24992 44596 25056
rect 44276 23968 44596 24992
rect 44276 23904 44284 23968
rect 44348 23904 44364 23968
rect 44428 23904 44444 23968
rect 44508 23904 44524 23968
rect 44588 23904 44596 23968
rect 44276 22880 44596 23904
rect 44276 22816 44284 22880
rect 44348 22816 44364 22880
rect 44428 22816 44444 22880
rect 44508 22816 44524 22880
rect 44588 22816 44596 22880
rect 44276 21792 44596 22816
rect 44276 21728 44284 21792
rect 44348 21728 44364 21792
rect 44428 21728 44444 21792
rect 44508 21728 44524 21792
rect 44588 21728 44596 21792
rect 44276 20704 44596 21728
rect 44276 20640 44284 20704
rect 44348 20640 44364 20704
rect 44428 20640 44444 20704
rect 44508 20640 44524 20704
rect 44588 20640 44596 20704
rect 44276 19616 44596 20640
rect 44276 19552 44284 19616
rect 44348 19552 44364 19616
rect 44428 19552 44444 19616
rect 44508 19552 44524 19616
rect 44588 19552 44596 19616
rect 44276 18528 44596 19552
rect 44276 18464 44284 18528
rect 44348 18464 44364 18528
rect 44428 18464 44444 18528
rect 44508 18464 44524 18528
rect 44588 18464 44596 18528
rect 44276 17440 44596 18464
rect 44276 17376 44284 17440
rect 44348 17376 44364 17440
rect 44428 17376 44444 17440
rect 44508 17376 44524 17440
rect 44588 17376 44596 17440
rect 44276 16352 44596 17376
rect 44276 16288 44284 16352
rect 44348 16288 44364 16352
rect 44428 16288 44444 16352
rect 44508 16288 44524 16352
rect 44588 16288 44596 16352
rect 44276 15264 44596 16288
rect 44276 15200 44284 15264
rect 44348 15200 44364 15264
rect 44428 15200 44444 15264
rect 44508 15200 44524 15264
rect 44588 15200 44596 15264
rect 44276 14176 44596 15200
rect 44276 14112 44284 14176
rect 44348 14112 44364 14176
rect 44428 14112 44444 14176
rect 44508 14112 44524 14176
rect 44588 14112 44596 14176
rect 44276 13088 44596 14112
rect 44276 13024 44284 13088
rect 44348 13024 44364 13088
rect 44428 13024 44444 13088
rect 44508 13024 44524 13088
rect 44588 13024 44596 13088
rect 44276 12000 44596 13024
rect 44276 11936 44284 12000
rect 44348 11936 44364 12000
rect 44428 11936 44444 12000
rect 44508 11936 44524 12000
rect 44588 11936 44596 12000
rect 44276 10912 44596 11936
rect 44276 10848 44284 10912
rect 44348 10848 44364 10912
rect 44428 10848 44444 10912
rect 44508 10848 44524 10912
rect 44588 10848 44596 10912
rect 44276 9824 44596 10848
rect 44276 9760 44284 9824
rect 44348 9760 44364 9824
rect 44428 9760 44444 9824
rect 44508 9760 44524 9824
rect 44588 9760 44596 9824
rect 44276 8736 44596 9760
rect 44276 8672 44284 8736
rect 44348 8672 44364 8736
rect 44428 8672 44444 8736
rect 44508 8672 44524 8736
rect 44588 8672 44596 8736
rect 44276 7648 44596 8672
rect 44276 7584 44284 7648
rect 44348 7584 44364 7648
rect 44428 7584 44444 7648
rect 44508 7584 44524 7648
rect 44588 7584 44596 7648
rect 44276 6560 44596 7584
rect 44276 6496 44284 6560
rect 44348 6496 44364 6560
rect 44428 6496 44444 6560
rect 44508 6496 44524 6560
rect 44588 6496 44596 6560
rect 44276 5472 44596 6496
rect 44276 5408 44284 5472
rect 44348 5408 44364 5472
rect 44428 5408 44444 5472
rect 44508 5408 44524 5472
rect 44588 5408 44596 5472
rect 44276 4384 44596 5408
rect 44276 4320 44284 4384
rect 44348 4320 44364 4384
rect 44428 4320 44444 4384
rect 44508 4320 44524 4384
rect 44588 4320 44596 4384
rect 44276 3296 44596 4320
rect 44276 3232 44284 3296
rect 44348 3232 44364 3296
rect 44428 3232 44444 3296
rect 44508 3232 44524 3296
rect 44588 3232 44596 3296
rect 44276 2208 44596 3232
rect 44276 2144 44284 2208
rect 44348 2144 44364 2208
rect 44428 2144 44444 2208
rect 44508 2144 44524 2208
rect 44588 2144 44596 2208
rect 44276 2128 44596 2144
rect 51498 27776 51818 27792
rect 51498 27712 51506 27776
rect 51570 27712 51586 27776
rect 51650 27712 51666 27776
rect 51730 27712 51746 27776
rect 51810 27712 51818 27776
rect 51498 26688 51818 27712
rect 51498 26624 51506 26688
rect 51570 26624 51586 26688
rect 51650 26624 51666 26688
rect 51730 26624 51746 26688
rect 51810 26624 51818 26688
rect 51498 25600 51818 26624
rect 51498 25536 51506 25600
rect 51570 25536 51586 25600
rect 51650 25536 51666 25600
rect 51730 25536 51746 25600
rect 51810 25536 51818 25600
rect 51498 24512 51818 25536
rect 51498 24448 51506 24512
rect 51570 24448 51586 24512
rect 51650 24448 51666 24512
rect 51730 24448 51746 24512
rect 51810 24448 51818 24512
rect 51498 23424 51818 24448
rect 51498 23360 51506 23424
rect 51570 23360 51586 23424
rect 51650 23360 51666 23424
rect 51730 23360 51746 23424
rect 51810 23360 51818 23424
rect 51498 22336 51818 23360
rect 51498 22272 51506 22336
rect 51570 22272 51586 22336
rect 51650 22272 51666 22336
rect 51730 22272 51746 22336
rect 51810 22272 51818 22336
rect 51498 21248 51818 22272
rect 51498 21184 51506 21248
rect 51570 21184 51586 21248
rect 51650 21184 51666 21248
rect 51730 21184 51746 21248
rect 51810 21184 51818 21248
rect 51498 20160 51818 21184
rect 51498 20096 51506 20160
rect 51570 20096 51586 20160
rect 51650 20096 51666 20160
rect 51730 20096 51746 20160
rect 51810 20096 51818 20160
rect 51498 19072 51818 20096
rect 51498 19008 51506 19072
rect 51570 19008 51586 19072
rect 51650 19008 51666 19072
rect 51730 19008 51746 19072
rect 51810 19008 51818 19072
rect 51498 17984 51818 19008
rect 51498 17920 51506 17984
rect 51570 17920 51586 17984
rect 51650 17920 51666 17984
rect 51730 17920 51746 17984
rect 51810 17920 51818 17984
rect 51498 16896 51818 17920
rect 51498 16832 51506 16896
rect 51570 16832 51586 16896
rect 51650 16832 51666 16896
rect 51730 16832 51746 16896
rect 51810 16832 51818 16896
rect 51498 15808 51818 16832
rect 51498 15744 51506 15808
rect 51570 15744 51586 15808
rect 51650 15744 51666 15808
rect 51730 15744 51746 15808
rect 51810 15744 51818 15808
rect 51498 14720 51818 15744
rect 51498 14656 51506 14720
rect 51570 14656 51586 14720
rect 51650 14656 51666 14720
rect 51730 14656 51746 14720
rect 51810 14656 51818 14720
rect 51498 13632 51818 14656
rect 51498 13568 51506 13632
rect 51570 13568 51586 13632
rect 51650 13568 51666 13632
rect 51730 13568 51746 13632
rect 51810 13568 51818 13632
rect 51498 12544 51818 13568
rect 51498 12480 51506 12544
rect 51570 12480 51586 12544
rect 51650 12480 51666 12544
rect 51730 12480 51746 12544
rect 51810 12480 51818 12544
rect 51498 11456 51818 12480
rect 51498 11392 51506 11456
rect 51570 11392 51586 11456
rect 51650 11392 51666 11456
rect 51730 11392 51746 11456
rect 51810 11392 51818 11456
rect 51498 10368 51818 11392
rect 58720 27232 59040 27792
rect 58720 27168 58728 27232
rect 58792 27168 58808 27232
rect 58872 27168 58888 27232
rect 58952 27168 58968 27232
rect 59032 27168 59040 27232
rect 58720 26144 59040 27168
rect 58720 26080 58728 26144
rect 58792 26080 58808 26144
rect 58872 26080 58888 26144
rect 58952 26080 58968 26144
rect 59032 26080 59040 26144
rect 58720 25056 59040 26080
rect 58720 24992 58728 25056
rect 58792 24992 58808 25056
rect 58872 24992 58888 25056
rect 58952 24992 58968 25056
rect 59032 24992 59040 25056
rect 58720 23968 59040 24992
rect 58720 23904 58728 23968
rect 58792 23904 58808 23968
rect 58872 23904 58888 23968
rect 58952 23904 58968 23968
rect 59032 23904 59040 23968
rect 58720 22880 59040 23904
rect 58720 22816 58728 22880
rect 58792 22816 58808 22880
rect 58872 22816 58888 22880
rect 58952 22816 58968 22880
rect 59032 22816 59040 22880
rect 58720 21792 59040 22816
rect 58720 21728 58728 21792
rect 58792 21728 58808 21792
rect 58872 21728 58888 21792
rect 58952 21728 58968 21792
rect 59032 21728 59040 21792
rect 58720 20704 59040 21728
rect 58720 20640 58728 20704
rect 58792 20640 58808 20704
rect 58872 20640 58888 20704
rect 58952 20640 58968 20704
rect 59032 20640 59040 20704
rect 58720 19616 59040 20640
rect 58720 19552 58728 19616
rect 58792 19552 58808 19616
rect 58872 19552 58888 19616
rect 58952 19552 58968 19616
rect 59032 19552 59040 19616
rect 58720 18528 59040 19552
rect 58720 18464 58728 18528
rect 58792 18464 58808 18528
rect 58872 18464 58888 18528
rect 58952 18464 58968 18528
rect 59032 18464 59040 18528
rect 58720 17440 59040 18464
rect 58720 17376 58728 17440
rect 58792 17376 58808 17440
rect 58872 17376 58888 17440
rect 58952 17376 58968 17440
rect 59032 17376 59040 17440
rect 58720 16352 59040 17376
rect 58720 16288 58728 16352
rect 58792 16288 58808 16352
rect 58872 16288 58888 16352
rect 58952 16288 58968 16352
rect 59032 16288 59040 16352
rect 58720 15264 59040 16288
rect 58720 15200 58728 15264
rect 58792 15200 58808 15264
rect 58872 15200 58888 15264
rect 58952 15200 58968 15264
rect 59032 15200 59040 15264
rect 58720 14176 59040 15200
rect 58720 14112 58728 14176
rect 58792 14112 58808 14176
rect 58872 14112 58888 14176
rect 58952 14112 58968 14176
rect 59032 14112 59040 14176
rect 58720 13088 59040 14112
rect 58720 13024 58728 13088
rect 58792 13024 58808 13088
rect 58872 13024 58888 13088
rect 58952 13024 58968 13088
rect 59032 13024 59040 13088
rect 58720 12000 59040 13024
rect 58720 11936 58728 12000
rect 58792 11936 58808 12000
rect 58872 11936 58888 12000
rect 58952 11936 58968 12000
rect 59032 11936 59040 12000
rect 57099 11116 57165 11117
rect 57099 11052 57100 11116
rect 57164 11052 57165 11116
rect 57099 11051 57165 11052
rect 51498 10304 51506 10368
rect 51570 10304 51586 10368
rect 51650 10304 51666 10368
rect 51730 10304 51746 10368
rect 51810 10304 51818 10368
rect 51498 9280 51818 10304
rect 51498 9216 51506 9280
rect 51570 9216 51586 9280
rect 51650 9216 51666 9280
rect 51730 9216 51746 9280
rect 51810 9216 51818 9280
rect 51498 8192 51818 9216
rect 51498 8128 51506 8192
rect 51570 8128 51586 8192
rect 51650 8128 51666 8192
rect 51730 8128 51746 8192
rect 51810 8128 51818 8192
rect 51498 7104 51818 8128
rect 51498 7040 51506 7104
rect 51570 7040 51586 7104
rect 51650 7040 51666 7104
rect 51730 7040 51746 7104
rect 51810 7040 51818 7104
rect 51498 6016 51818 7040
rect 51498 5952 51506 6016
rect 51570 5952 51586 6016
rect 51650 5952 51666 6016
rect 51730 5952 51746 6016
rect 51810 5952 51818 6016
rect 51498 4928 51818 5952
rect 51498 4864 51506 4928
rect 51570 4864 51586 4928
rect 51650 4864 51666 4928
rect 51730 4864 51746 4928
rect 51810 4864 51818 4928
rect 51498 3840 51818 4864
rect 57102 4045 57162 11051
rect 58720 10912 59040 11936
rect 58720 10848 58728 10912
rect 58792 10848 58808 10912
rect 58872 10848 58888 10912
rect 58952 10848 58968 10912
rect 59032 10848 59040 10912
rect 58720 9824 59040 10848
rect 58720 9760 58728 9824
rect 58792 9760 58808 9824
rect 58872 9760 58888 9824
rect 58952 9760 58968 9824
rect 59032 9760 59040 9824
rect 58720 8736 59040 9760
rect 58720 8672 58728 8736
rect 58792 8672 58808 8736
rect 58872 8672 58888 8736
rect 58952 8672 58968 8736
rect 59032 8672 59040 8736
rect 58720 7648 59040 8672
rect 58720 7584 58728 7648
rect 58792 7584 58808 7648
rect 58872 7584 58888 7648
rect 58952 7584 58968 7648
rect 59032 7584 59040 7648
rect 58720 6560 59040 7584
rect 58720 6496 58728 6560
rect 58792 6496 58808 6560
rect 58872 6496 58888 6560
rect 58952 6496 58968 6560
rect 59032 6496 59040 6560
rect 58720 5472 59040 6496
rect 58720 5408 58728 5472
rect 58792 5408 58808 5472
rect 58872 5408 58888 5472
rect 58952 5408 58968 5472
rect 59032 5408 59040 5472
rect 58720 4384 59040 5408
rect 58720 4320 58728 4384
rect 58792 4320 58808 4384
rect 58872 4320 58888 4384
rect 58952 4320 58968 4384
rect 59032 4320 59040 4384
rect 57099 4044 57165 4045
rect 57099 3980 57100 4044
rect 57164 3980 57165 4044
rect 57099 3979 57165 3980
rect 51498 3776 51506 3840
rect 51570 3776 51586 3840
rect 51650 3776 51666 3840
rect 51730 3776 51746 3840
rect 51810 3776 51818 3840
rect 51498 2752 51818 3776
rect 51498 2688 51506 2752
rect 51570 2688 51586 2752
rect 51650 2688 51666 2752
rect 51730 2688 51746 2752
rect 51810 2688 51818 2752
rect 51498 2128 51818 2688
rect 58720 3296 59040 4320
rect 58720 3232 58728 3296
rect 58792 3232 58808 3296
rect 58872 3232 58888 3296
rect 58952 3232 58968 3296
rect 59032 3232 59040 3296
rect 58720 2208 59040 3232
rect 58720 2144 58728 2208
rect 58792 2144 58808 2208
rect 58872 2144 58888 2208
rect 58952 2144 58968 2208
rect 59032 2144 59040 2208
rect 58720 2128 59040 2144
use sky130_fd_sc_hd__or4bb_1  _0414_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 54372 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0415_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0416_
timestamp 1688980957
transform 1 0 41768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0417_
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0418_
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0419_
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0420_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0421_
timestamp 1688980957
transform 1 0 27324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _0422_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _0423_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0424_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0425_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _0426_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _0427_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0428_
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0429_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0430_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0431_
timestamp 1688980957
transform 1 0 9016 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0432_
timestamp 1688980957
transform 1 0 9476 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0433_
timestamp 1688980957
transform 1 0 9844 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0434_
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0435_
timestamp 1688980957
transform 1 0 8004 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0436_
timestamp 1688980957
transform 1 0 6716 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0437_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0438_
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0439_
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0440_
timestamp 1688980957
transform 1 0 9476 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0441_
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0442_
timestamp 1688980957
transform 1 0 11592 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0443_
timestamp 1688980957
transform 1 0 12788 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0444_
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0445_
timestamp 1688980957
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0446_
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0447_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0448_
timestamp 1688980957
transform 1 0 14260 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0449_
timestamp 1688980957
transform 1 0 16008 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0450_
timestamp 1688980957
transform 1 0 14996 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0451_
timestamp 1688980957
transform 1 0 15456 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0452_
timestamp 1688980957
transform 1 0 14996 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0453_
timestamp 1688980957
transform 1 0 17480 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0454_
timestamp 1688980957
transform 1 0 17848 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0455_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0456_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0457_
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0458_
timestamp 1688980957
transform 1 0 20516 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0459_
timestamp 1688980957
transform 1 0 17848 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0460_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0461_
timestamp 1688980957
transform 1 0 19872 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0462_
timestamp 1688980957
transform 1 0 17848 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0463_
timestamp 1688980957
transform 1 0 20240 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0464_
timestamp 1688980957
transform 1 0 19780 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0465_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0466_
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0467_
timestamp 1688980957
transform 1 0 23276 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0468_
timestamp 1688980957
transform 1 0 23460 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0469_
timestamp 1688980957
transform 1 0 24380 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0470_
timestamp 1688980957
transform 1 0 22816 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0471_
timestamp 1688980957
transform 1 0 24380 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0472_
timestamp 1688980957
transform 1 0 24748 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0473_
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0474_
timestamp 1688980957
transform 1 0 24196 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0475_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0476_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0477_
timestamp 1688980957
transform 1 0 25760 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0478_
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0479_
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0480_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0481_
timestamp 1688980957
transform 1 0 30360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0482_
timestamp 1688980957
transform 1 0 29532 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0483_
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0484_
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0485_
timestamp 1688980957
transform 1 0 31464 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0486_
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0487_
timestamp 1688980957
transform 1 0 30084 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0488_
timestamp 1688980957
transform 1 0 29900 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0489_
timestamp 1688980957
transform 1 0 31188 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0490_
timestamp 1688980957
transform 1 0 37812 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0491_
timestamp 1688980957
transform 1 0 35052 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0492_
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1688980957
transform 1 0 36156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0494_
timestamp 1688980957
transform 1 0 35236 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0495_
timestamp 1688980957
transform 1 0 33396 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0496_
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0497_
timestamp 1688980957
transform 1 0 35328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0498_
timestamp 1688980957
transform 1 0 34592 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0499_
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0500_
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0501_
timestamp 1688980957
transform 1 0 36616 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0502_
timestamp 1688980957
transform 1 0 37444 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0503_
timestamp 1688980957
transform 1 0 37904 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0504_
timestamp 1688980957
transform 1 0 38364 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0505_
timestamp 1688980957
transform 1 0 39192 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0506_
timestamp 1688980957
transform 1 0 40756 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0507_
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0508_
timestamp 1688980957
transform 1 0 39376 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0509_
timestamp 1688980957
transform 1 0 41308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0510_
timestamp 1688980957
transform 1 0 41216 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0511_
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0512_
timestamp 1688980957
transform 1 0 40388 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0513_
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0514_
timestamp 1688980957
transform 1 0 42872 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0515_
timestamp 1688980957
transform 1 0 42688 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0516_
timestamp 1688980957
transform 1 0 42688 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1688980957
transform 1 0 43884 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0518_
timestamp 1688980957
transform 1 0 46276 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0519_
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0520_
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1688980957
transform 1 0 45724 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0522_
timestamp 1688980957
transform 1 0 46736 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0523_
timestamp 1688980957
transform 1 0 46552 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0524_
timestamp 1688980957
transform 1 0 46460 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1688980957
transform 1 0 47564 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0526_
timestamp 1688980957
transform 1 0 47932 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0527_
timestamp 1688980957
transform 1 0 48484 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0528_
timestamp 1688980957
transform 1 0 48852 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0529_
timestamp 1688980957
transform 1 0 50140 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0530_
timestamp 1688980957
transform 1 0 48300 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0531_
timestamp 1688980957
transform 1 0 48116 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0532_
timestamp 1688980957
transform 1 0 47564 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0533_
timestamp 1688980957
transform 1 0 50140 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0534_
timestamp 1688980957
transform 1 0 50876 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0535_
timestamp 1688980957
transform 1 0 51336 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0536_
timestamp 1688980957
transform 1 0 51428 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0537_
timestamp 1688980957
transform 1 0 53268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0538_
timestamp 1688980957
transform 1 0 51428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0539_
timestamp 1688980957
transform 1 0 54004 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0540_
timestamp 1688980957
transform 1 0 51612 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0541_
timestamp 1688980957
transform 1 0 54280 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0542_
timestamp 1688980957
transform 1 0 53544 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0543_
timestamp 1688980957
transform 1 0 54464 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0544_
timestamp 1688980957
transform 1 0 54740 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0545_
timestamp 1688980957
transform 1 0 56396 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0546_
timestamp 1688980957
transform 1 0 57132 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0547_
timestamp 1688980957
transform 1 0 55752 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0548_
timestamp 1688980957
transform 1 0 55660 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0549_
timestamp 1688980957
transform 1 0 56856 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0550_
timestamp 1688980957
transform 1 0 57224 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0551_
timestamp 1688980957
transform 1 0 55476 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _0552_
timestamp 1688980957
transform 1 0 55660 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _0553_
timestamp 1688980957
transform 1 0 56948 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0554_
timestamp 1688980957
transform 1 0 55476 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0555_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _0556_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0557_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1688980957
transform 1 0 29256 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0559_
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1688980957
transform 1 0 30912 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0561_
timestamp 1688980957
transform 1 0 36984 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0562_
timestamp 1688980957
transform 1 0 33764 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0564_
timestamp 1688980957
transform 1 0 38916 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0565_
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0566_
timestamp 1688980957
transform 1 0 42136 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0567_
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0568_
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0569_
timestamp 1688980957
transform 1 0 48484 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1688980957
transform 1 0 50140 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0571_
timestamp 1688980957
transform 1 0 48944 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0572_
timestamp 1688980957
transform 1 0 52716 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0573_
timestamp 1688980957
transform 1 0 56028 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0574_
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0575_
timestamp 1688980957
transform 1 0 56580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0576_
timestamp 1688980957
transform 1 0 56396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0577_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_4  _0578_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0579_
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0580_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0581_
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0582_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0583_
timestamp 1688980957
transform 1 0 14720 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0584_
timestamp 1688980957
transform 1 0 15088 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0585_
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0586_
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0587_
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0588_
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0589_
timestamp 1688980957
transform 1 0 24748 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1688980957
transform 1 0 25852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0591_
timestamp 1688980957
transform 1 0 26312 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0592_
timestamp 1688980957
transform 1 0 30176 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0593_
timestamp 1688980957
transform 1 0 30360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0594_
timestamp 1688980957
transform 1 0 32292 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0595_
timestamp 1688980957
transform 1 0 36156 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0596_
timestamp 1688980957
transform 1 0 34776 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0597_
timestamp 1688980957
transform 1 0 36616 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0598_
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0599_
timestamp 1688980957
transform 1 0 41124 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0600_
timestamp 1688980957
transform 1 0 42228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0601_
timestamp 1688980957
transform 1 0 43884 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0602_
timestamp 1688980957
transform 1 0 45724 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0603_
timestamp 1688980957
transform 1 0 48392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1688980957
transform 1 0 48944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0605_
timestamp 1688980957
transform 1 0 50140 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0606_
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1688980957
transform 1 0 56856 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0608_
timestamp 1688980957
transform 1 0 56304 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0609_
timestamp 1688980957
transform 1 0 56856 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0610_
timestamp 1688980957
transform 1 0 57500 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0611_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0612_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0613_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0615_
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 1688980957
transform 1 0 5520 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0617_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0618_
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0619_
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0620_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0621_
timestamp 1688980957
transform 1 0 18032 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1688980957
transform 1 0 17940 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0623_
timestamp 1688980957
transform 1 0 19320 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0624_
timestamp 1688980957
transform 1 0 23184 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0625_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0626_
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0627_
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0628_
timestamp 1688980957
transform 1 0 28152 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0629_
timestamp 1688980957
transform 1 0 28704 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 1688980957
transform 1 0 33120 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0631_
timestamp 1688980957
transform 1 0 32936 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0632_
timestamp 1688980957
transform 1 0 33856 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0633_
timestamp 1688980957
transform 1 0 38916 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0634_
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0635_
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0637_
timestamp 1688980957
transform 1 0 43332 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0638_
timestamp 1688980957
transform 1 0 45080 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 1688980957
transform 1 0 48024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0640_
timestamp 1688980957
transform 1 0 46736 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0641_
timestamp 1688980957
transform 1 0 50692 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1688980957
transform 1 0 51704 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 1688980957
transform 1 0 53636 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0644_
timestamp 1688980957
transform 1 0 55292 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0645_
timestamp 1688980957
transform 1 0 55292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0646_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0647_
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0648_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0649_
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0650_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0651_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0652_
timestamp 1688980957
transform 1 0 5152 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0653_
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0654_
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0655_
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0656_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0657_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0658_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0659_
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0660_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0661_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0662_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0663_
timestamp 1688980957
transform 1 0 2760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0664_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0665_
timestamp 1688980957
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0666_
timestamp 1688980957
transform 1 0 2668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0667_
timestamp 1688980957
transform 1 0 3404 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _0668_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1688980957
transform 1 0 2944 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0670_
timestamp 1688980957
transform 1 0 8004 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0671_
timestamp 1688980957
transform 1 0 6992 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0672_
timestamp 1688980957
transform 1 0 8372 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0673_
timestamp 1688980957
transform 1 0 12604 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0674_
timestamp 1688980957
transform 1 0 12972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0675_
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0676_
timestamp 1688980957
transform 1 0 17664 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0677_
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0678_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0679_
timestamp 1688980957
transform 1 0 22356 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0680_
timestamp 1688980957
transform 1 0 23460 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0681_
timestamp 1688980957
transform 1 0 23644 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0682_
timestamp 1688980957
transform 1 0 27600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0683_
timestamp 1688980957
transform 1 0 28704 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0684_
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0685_
timestamp 1688980957
transform 1 0 34500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1688980957
transform 1 0 32384 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0687_
timestamp 1688980957
transform 1 0 33948 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0688_
timestamp 1688980957
transform 1 0 38456 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0689_
timestamp 1688980957
transform 1 0 39284 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0691_
timestamp 1688980957
transform 1 0 41492 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 43332 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0693_
timestamp 1688980957
transform 1 0 46000 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1688980957
transform 1 0 48392 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0695_
timestamp 1688980957
transform 1 0 47012 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 1688980957
transform 1 0 51612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0697_
timestamp 1688980957
transform 1 0 53912 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 1688980957
transform 1 0 52532 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1688980957
transform 1 0 55292 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 1688980957
transform 1 0 54188 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0701_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1688980957
transform 1 0 5428 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0705_
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0706_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0708_
timestamp 1688980957
transform 1 0 13156 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 1688980957
transform 1 0 18676 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0710_
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 1688980957
transform 1 0 23460 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1688980957
transform 1 0 23736 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 1688980957
transform 1 0 28704 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1688980957
transform 1 0 28704 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0717_
timestamp 1688980957
transform 1 0 28428 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1688980957
transform 1 0 32660 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1688980957
transform 1 0 33028 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform 1 0 37536 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0722_
timestamp 1688980957
transform 1 0 38732 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0724_
timestamp 1688980957
transform 1 0 41492 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1688980957
transform 1 0 43884 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0726_
timestamp 1688980957
transform 1 0 45816 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1688980957
transform 1 0 47932 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 1688980957
transform 1 0 47380 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1688980957
transform 1 0 51428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 1688980957
transform 1 0 50968 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1688980957
transform 1 0 52808 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1688980957
transform 1 0 55292 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0733_
timestamp 1688980957
transform 1 0 54648 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0734_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0735_
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0737_
timestamp 1688980957
transform 1 0 7268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1688980957
transform 1 0 10488 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0739_
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform 1 0 14996 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1688980957
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0745_
timestamp 1688980957
transform 1 0 26036 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1688980957
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform 1 0 30176 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0749_
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1688980957
transform 1 0 30820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1688980957
transform 1 0 36616 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1688980957
transform 1 0 35972 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1688980957
transform 1 0 38824 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1688980957
transform 1 0 41860 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0757_
timestamp 1688980957
transform 1 0 44988 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1688980957
transform 1 0 46092 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0759_
timestamp 1688980957
transform 1 0 49220 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1688980957
transform 1 0 49220 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1688980957
transform 1 0 47748 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1688980957
transform 1 0 51612 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1688980957
transform 1 0 51060 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1688980957
transform 1 0 56672 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1688980957
transform 1 0 56488 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1688980957
transform 1 0 56488 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_4  _0767_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1688980957
transform 1 0 13800 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1688980957
transform 1 0 16376 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 1688980957
transform 1 0 21160 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1688980957
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1688980957
transform 1 0 22080 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1688980957
transform 1 0 25392 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1688980957
transform 1 0 25300 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1688980957
transform 1 0 26312 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1688980957
transform 1 0 30176 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1688980957
transform 1 0 31464 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1688980957
transform 1 0 32016 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1688980957
transform 1 0 36064 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1688980957
transform 1 0 35788 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1688980957
transform 1 0 38916 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1688980957
transform 1 0 41124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1688980957
transform 1 0 42688 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1688980957
transform 1 0 44620 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1688980957
transform 1 0 45448 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1688980957
transform 1 0 48392 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1688980957
transform 1 0 50784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1688980957
transform 1 0 49496 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1688980957
transform 1 0 52716 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1688980957
transform 1 0 52716 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1688980957
transform 1 0 57408 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1688980957
transform 1 0 57592 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1688980957
transform 1 0 57592 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0800_
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0801_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1688980957
transform 1 0 2668 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0803_
timestamp 1688980957
transform 1 0 2300 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0804_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0805_
timestamp 1688980957
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0806_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0807_
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0809_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0810_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0811_
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0812_
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0813_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0814_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0815_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1688980957
transform 1 0 7728 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1688980957
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp 1688980957
transform 1 0 13524 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp 1688980957
transform 1 0 18400 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 1688980957
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp 1688980957
transform 1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp 1688980957
transform 1 0 23184 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 1688980957
transform 1 0 22816 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform 1 0 28152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1688980957
transform 1 0 27784 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp 1688980957
transform 1 0 28520 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp 1688980957
transform 1 0 33580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0833_
timestamp 1688980957
transform 1 0 32200 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0834_
timestamp 1688980957
transform 1 0 33120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp 1688980957
transform 1 0 38088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp 1688980957
transform 1 0 38456 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp 1688980957
transform 1 0 39192 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 1688980957
transform 1 0 41492 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp 1688980957
transform 1 0 43792 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 1688980957
transform 1 0 45172 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp 1688980957
transform 1 0 47656 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1688980957
transform 1 0 47564 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0843_
timestamp 1688980957
transform 1 0 50692 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 1688980957
transform 1 0 52992 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1688980957
transform 1 0 52808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1688980957
transform 1 0 54372 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0847_
timestamp 1688980957
transform 1 0 54096 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1688980957
transform 1 0 4416 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1688980957
transform 1 0 10488 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1688980957
transform 1 0 9016 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1688980957
transform 1 0 14076 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1688980957
transform 1 0 14720 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1688980957
transform 1 0 20056 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1688980957
transform 1 0 25024 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1688980957
transform 1 0 24564 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1688980957
transform 1 0 25024 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _0861_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0862_
timestamp 1688980957
transform 1 0 28612 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0863_
timestamp 1688980957
transform 1 0 30360 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0864_
timestamp 1688980957
transform 1 0 35880 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0865_
timestamp 1688980957
transform 1 0 33120 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0866_
timestamp 1688980957
transform 1 0 35236 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0867_
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0868_
timestamp 1688980957
transform 1 0 39284 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0869_
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0870_
timestamp 1688980957
transform 1 0 43516 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0871_
timestamp 1688980957
transform 1 0 44252 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0872_
timestamp 1688980957
transform 1 0 47564 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0873_
timestamp 1688980957
transform 1 0 50416 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0874_
timestamp 1688980957
transform 1 0 48392 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0875_
timestamp 1688980957
transform 1 0 51704 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0876_
timestamp 1688980957
transform 1 0 55936 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0877_
timestamp 1688980957
transform 1 0 55292 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0878_
timestamp 1688980957
transform 1 0 56396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0879_
timestamp 1688980957
transform 1 0 56028 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0880_
timestamp 1688980957
transform 1 0 5704 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0881_
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0882_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0883_
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0884_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0885_
timestamp 1688980957
transform 1 0 14720 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0886_
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0887_
timestamp 1688980957
transform 1 0 19596 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0888_
timestamp 1688980957
transform 1 0 19320 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0889_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0890_
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0891_
timestamp 1688980957
transform 1 0 25392 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0892_
timestamp 1688980957
transform 1 0 25208 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0893_
timestamp 1688980957
transform 1 0 29900 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0894_
timestamp 1688980957
transform 1 0 30084 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0895_
timestamp 1688980957
transform 1 0 32200 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0896_
timestamp 1688980957
transform 1 0 35880 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0897_
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0898_
timestamp 1688980957
transform 1 0 35880 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0899_
timestamp 1688980957
transform 1 0 39836 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0900_
timestamp 1688980957
transform 1 0 40848 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0901_
timestamp 1688980957
transform 1 0 42872 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0902_
timestamp 1688980957
transform 1 0 43516 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0903_
timestamp 1688980957
transform 1 0 45080 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0904_
timestamp 1688980957
transform 1 0 47564 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0905_
timestamp 1688980957
transform 1 0 48392 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0906_
timestamp 1688980957
transform 1 0 49588 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0907_
timestamp 1688980957
transform 1 0 51704 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0908_
timestamp 1688980957
transform 1 0 56396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0909_
timestamp 1688980957
transform 1 0 56856 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0910_
timestamp 1688980957
transform 1 0 56304 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0911_
timestamp 1688980957
transform 1 0 56488 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0912_
timestamp 1688980957
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0913_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0914_
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0915_
timestamp 1688980957
transform 1 0 7360 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0916_
timestamp 1688980957
transform 1 0 10488 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0917_
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0918_
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0919_
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0920_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0921_
timestamp 1688980957
transform 1 0 18308 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0922_
timestamp 1688980957
transform 1 0 21988 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0923_
timestamp 1688980957
transform 1 0 23276 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0924_
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0925_
timestamp 1688980957
transform 1 0 27416 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0926_
timestamp 1688980957
transform 1 0 27416 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0927_
timestamp 1688980957
transform 1 0 27968 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0928_
timestamp 1688980957
transform 1 0 32384 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0929_
timestamp 1688980957
transform 1 0 32292 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0930_
timestamp 1688980957
transform 1 0 32476 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0931_
timestamp 1688980957
transform 1 0 37444 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0932_
timestamp 1688980957
transform 1 0 38272 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0933_
timestamp 1688980957
transform 1 0 38456 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0934_
timestamp 1688980957
transform 1 0 40848 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0935_
timestamp 1688980957
transform 1 0 42688 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0936_
timestamp 1688980957
transform 1 0 44988 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0937_
timestamp 1688980957
transform 1 0 47472 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0938_
timestamp 1688980957
transform 1 0 46000 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0939_
timestamp 1688980957
transform 1 0 50140 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0940_
timestamp 1688980957
transform 1 0 50140 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0941_
timestamp 1688980957
transform 1 0 52624 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0942_
timestamp 1688980957
transform 1 0 53728 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0943_
timestamp 1688980957
transform 1 0 54280 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0944_
timestamp 1688980957
transform 1 0 1840 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0945_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0946_
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0947_
timestamp 1688980957
transform 1 0 1840 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0948_
timestamp 1688980957
transform 1 0 7544 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0949_
timestamp 1688980957
transform 1 0 6440 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0950_
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0951_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0952_
timestamp 1688980957
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0953_
timestamp 1688980957
transform 1 0 13248 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0954_
timestamp 1688980957
transform 1 0 16928 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0955_
timestamp 1688980957
transform 1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0956_
timestamp 1688980957
transform 1 0 18400 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0957_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0958_
timestamp 1688980957
transform 1 0 22724 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0959_
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0960_
timestamp 1688980957
transform 1 0 27324 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0961_
timestamp 1688980957
transform 1 0 27416 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 1688980957
transform 1 0 32568 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 1688980957
transform 1 0 36984 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 1688980957
transform 1 0 38272 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 1688980957
transform 1 0 40848 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0970_
timestamp 1688980957
transform 1 0 42688 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0971_
timestamp 1688980957
transform 1 0 44804 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1688980957
transform 1 0 47196 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1688980957
transform 1 0 46460 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1688980957
transform 1 0 50232 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1688980957
transform 1 0 52808 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1688980957
transform 1 0 52716 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0977_
timestamp 1688980957
transform 1 0 54280 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1688980957
transform 1 0 53636 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1688980957
transform 1 0 2024 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1688980957
transform 1 0 4692 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1688980957
transform 1 0 7636 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1688980957
transform 1 0 9936 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1688980957
transform 1 0 17204 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1688980957
transform 1 0 16468 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1688980957
transform 1 0 22264 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1688980957
transform 1 0 27232 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1688980957
transform 1 0 27232 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1688980957
transform 1 0 27784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1688980957
transform 1 0 32016 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1688980957
transform 1 0 32384 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1688980957
transform 1 0 36984 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1688980957
transform 1 0 37904 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1688980957
transform 1 0 38272 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1688980957
transform 1 0 40756 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1688980957
transform 1 0 42412 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1688980957
transform 1 0 44344 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1688980957
transform 1 0 47564 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1688980957
transform 1 0 45908 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1688980957
transform 1 0 50876 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1688980957
transform 1 0 50232 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1688980957
transform 1 0 53912 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1688980957
transform 1 0 53728 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1688980957
transform 1 0 4784 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1688980957
transform 1 0 12420 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1688980957
transform 1 0 19504 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1688980957
transform 1 0 18584 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1688980957
transform 1 0 24288 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1688980957
transform 1 0 24932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1688980957
transform 1 0 29808 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1688980957
transform 1 0 29532 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1688980957
transform 1 0 35604 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1688980957
transform 1 0 38272 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1688980957
transform 1 0 38272 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1688980957
transform 1 0 40664 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1688980957
transform 1 0 43148 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1688980957
transform 1 0 44528 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1688980957
transform 1 0 49312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1688980957
transform 1 0 47564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1688980957
transform 1 0 51612 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1688980957
transform 1 0 50416 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1688980957
transform 1 0 55936 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1688980957
transform 1 0 56120 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1688980957
transform 1 0 56120 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1688980957
transform 1 0 5244 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1688980957
transform 1 0 8648 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1688980957
transform 1 0 10488 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1688980957
transform 1 0 15088 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1688980957
transform 1 0 19780 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1688980957
transform 1 0 19596 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1688980957
transform 1 0 20884 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1688980957
transform 1 0 24564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1688980957
transform 1 0 26128 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1688980957
transform 1 0 25300 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1688980957
transform 1 0 29808 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1688980957
transform 1 0 29992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1688980957
transform 1 0 30544 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1688980957
transform 1 0 35328 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1688980957
transform 1 0 34500 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1688980957
transform 1 0 35880 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1688980957
transform 1 0 43332 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1688980957
transform 1 0 45080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1688980957
transform 1 0 47564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1688980957
transform 1 0 50140 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1688980957
transform 1 0 48300 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1688980957
transform 1 0 52716 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1688980957
transform 1 0 52256 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1688980957
transform 1 0 56764 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1688980957
transform 1 0 56764 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1688980957
transform 1 0 56856 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1688980957
transform 1 0 1748 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1076_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1077_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1688980957
transform 1 0 6900 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1080_
timestamp 1688980957
transform 1 0 8096 0 -1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1688980957
transform 1 0 7268 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1688980957
transform 1 0 6256 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1688980957
transform 1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1688980957
transform 1 0 12052 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1688980957
transform 1 0 13248 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1688980957
transform 1 0 16928 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1688980957
transform 1 0 15640 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1688980957
transform 1 0 21712 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1688980957
transform 1 0 22816 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1688980957
transform 1 0 26680 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1688980957
transform 1 0 27232 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1688980957
transform 1 0 27048 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1688980957
transform 1 0 33028 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1688980957
transform 1 0 31464 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1688980957
transform 1 0 32476 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1688980957
transform 1 0 36616 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1688980957
transform 1 0 37720 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1688980957
transform 1 0 38272 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1688980957
transform 1 0 40756 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1688980957
transform 1 0 42320 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1688980957
transform 1 0 44988 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1688980957
transform 1 0 46920 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1688980957
transform 1 0 46000 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1688980957
transform 1 0 50140 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1688980957
transform 1 0 52440 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1688980957
transform 1 0 51336 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1688980957
transform 1 0 53912 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1688980957
transform 1 0 53452 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1688980957
transform 1 0 3496 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1688980957
transform 1 0 14168 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1688980957
transform 1 0 19504 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1688980957
transform 1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1688980957
transform 1 0 20792 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1688980957
transform 1 0 25208 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1688980957
transform 1 0 24472 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 51520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0424__C
timestamp 1688980957
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0426__B
timestamp 1688980957
transform 1 0 5336 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__S0
timestamp 1688980957
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0427__S1
timestamp 1688980957
transform 1 0 5704 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__S0
timestamp 1688980957
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0428__S1
timestamp 1688980957
transform 1 0 5060 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0429__S
timestamp 1688980957
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0430__A
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0431__S0
timestamp 1688980957
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0431__S1
timestamp 1688980957
transform 1 0 9476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__S0
timestamp 1688980957
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0432__S1
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0433__S
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0434__A
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0435__S0
timestamp 1688980957
transform 1 0 6808 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0435__S1
timestamp 1688980957
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__S0
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0436__S1
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0437__S
timestamp 1688980957
transform 1 0 8740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0438__A
timestamp 1688980957
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0439__S0
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0439__S1
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__S0
timestamp 1688980957
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0440__S1
timestamp 1688980957
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0441__S
timestamp 1688980957
transform 1 0 12512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0442__A
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__S0
timestamp 1688980957
transform 1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0443__S1
timestamp 1688980957
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__S0
timestamp 1688980957
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0444__S1
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0445__S
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0446__A
timestamp 1688980957
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__S0
timestamp 1688980957
transform 1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0447__S1
timestamp 1688980957
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__S0
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0448__S1
timestamp 1688980957
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0449__S
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0450__A
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__S0
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0451__S1
timestamp 1688980957
transform 1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__S0
timestamp 1688980957
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0452__S1
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0453__S
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0454__A
timestamp 1688980957
transform 1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__S0
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0455__S1
timestamp 1688980957
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__S0
timestamp 1688980957
transform 1 0 19412 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0456__S1
timestamp 1688980957
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0457__S
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0458__A
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__S0
timestamp 1688980957
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0459__S1
timestamp 1688980957
transform 1 0 17664 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__S0
timestamp 1688980957
transform 1 0 18400 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0460__S1
timestamp 1688980957
transform 1 0 19044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0461__S
timestamp 1688980957
transform 1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0462__A
timestamp 1688980957
transform 1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__S0
timestamp 1688980957
transform 1 0 20148 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0463__S1
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__S0
timestamp 1688980957
transform 1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0464__S1
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0465__S
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0466__A
timestamp 1688980957
transform 1 0 17296 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__S0
timestamp 1688980957
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0467__S1
timestamp 1688980957
transform 1 0 22172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__S0
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0468__S1
timestamp 1688980957
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0469__S
timestamp 1688980957
transform 1 0 24196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0470__A
timestamp 1688980957
transform 1 0 22816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__S0
timestamp 1688980957
transform 1 0 23368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0471__S1
timestamp 1688980957
transform 1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__S0
timestamp 1688980957
transform 1 0 23920 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0472__S1
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0473__S
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0474__A
timestamp 1688980957
transform 1 0 24564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__S0
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0475__S1
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0476__S0
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0476__S1
timestamp 1688980957
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0477__S
timestamp 1688980957
transform 1 0 25576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0478__A
timestamp 1688980957
transform 1 0 22540 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__S0
timestamp 1688980957
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0479__S1
timestamp 1688980957
transform 1 0 27416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__S0
timestamp 1688980957
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0480__S1
timestamp 1688980957
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0481__S
timestamp 1688980957
transform 1 0 30176 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0482__A
timestamp 1688980957
transform 1 0 27876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__S0
timestamp 1688980957
transform 1 0 29716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0483__S1
timestamp 1688980957
transform 1 0 31740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__S0
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0484__S1
timestamp 1688980957
transform 1 0 32292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__S
timestamp 1688980957
transform 1 0 31464 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1688980957
transform 1 0 31648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__S0
timestamp 1688980957
transform 1 0 33304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__S1
timestamp 1688980957
transform 1 0 32936 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__S0
timestamp 1688980957
transform 1 0 33028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__S1
timestamp 1688980957
transform 1 0 32200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__S
timestamp 1688980957
transform 1 0 32660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__S0
timestamp 1688980957
transform 1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__S1
timestamp 1688980957
transform 1 0 38548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__S0
timestamp 1688980957
transform 1 0 34408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__S1
timestamp 1688980957
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__S
timestamp 1688980957
transform 1 0 39744 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1688980957
transform 1 0 40112 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__S0
timestamp 1688980957
transform 1 0 33856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__S1
timestamp 1688980957
transform 1 0 33396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__S0
timestamp 1688980957
transform 1 0 34868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__S1
timestamp 1688980957
transform 1 0 35236 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__S
timestamp 1688980957
transform 1 0 35236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__S0
timestamp 1688980957
transform 1 0 34960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__S1
timestamp 1688980957
transform 1 0 34960 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__S0
timestamp 1688980957
transform 1 0 34316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__S1
timestamp 1688980957
transform 1 0 34868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__S
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1688980957
transform 1 0 40480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__S0
timestamp 1688980957
transform 1 0 37536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__S1
timestamp 1688980957
transform 1 0 37720 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__S0
timestamp 1688980957
transform 1 0 37996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__S1
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__S
timestamp 1688980957
transform 1 0 40204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1688980957
transform 1 0 43700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__S0
timestamp 1688980957
transform 1 0 40020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__S1
timestamp 1688980957
transform 1 0 41032 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__S0
timestamp 1688980957
transform 1 0 42872 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__S1
timestamp 1688980957
transform 1 0 42596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__S
timestamp 1688980957
transform 1 0 42504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A
timestamp 1688980957
transform 1 0 42596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__S0
timestamp 1688980957
transform 1 0 41032 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__S1
timestamp 1688980957
transform 1 0 41400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__S0
timestamp 1688980957
transform 1 0 40020 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__S1
timestamp 1688980957
transform 1 0 40388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__S
timestamp 1688980957
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1688980957
transform 1 0 44436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__S0
timestamp 1688980957
transform 1 0 45908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__S1
timestamp 1688980957
transform 1 0 46000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__S0
timestamp 1688980957
transform 1 0 45172 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__S1
timestamp 1688980957
transform 1 0 44620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__S
timestamp 1688980957
transform 1 0 43700 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1688980957
transform 1 0 51704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__S0
timestamp 1688980957
transform 1 0 48852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__S1
timestamp 1688980957
transform 1 0 49588 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__S0
timestamp 1688980957
transform 1 0 47748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__S1
timestamp 1688980957
transform 1 0 47104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__S
timestamp 1688980957
transform 1 0 47104 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1688980957
transform 1 0 52072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__S0
timestamp 1688980957
transform 1 0 46368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__S1
timestamp 1688980957
transform 1 0 49220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__S0
timestamp 1688980957
transform 1 0 46276 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__S1
timestamp 1688980957
transform 1 0 48576 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__S
timestamp 1688980957
transform 1 0 47748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1688980957
transform 1 0 52440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__S0
timestamp 1688980957
transform 1 0 49220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__S1
timestamp 1688980957
transform 1 0 49588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__S0
timestamp 1688980957
transform 1 0 48484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__S1
timestamp 1688980957
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__S
timestamp 1688980957
transform 1 0 52900 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1688980957
transform 1 0 52072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__S0
timestamp 1688980957
transform 1 0 48484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__S1
timestamp 1688980957
transform 1 0 47288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__S0
timestamp 1688980957
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__S1
timestamp 1688980957
transform 1 0 48484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__S
timestamp 1688980957
transform 1 0 51152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1688980957
transform 1 0 51060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__S0
timestamp 1688980957
transform 1 0 50968 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__S1
timestamp 1688980957
transform 1 0 51336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__S0
timestamp 1688980957
transform 1 0 51060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__S1
timestamp 1688980957
transform 1 0 50692 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__S
timestamp 1688980957
transform 1 0 53084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1688980957
transform 1 0 51428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__S0
timestamp 1688980957
transform 1 0 54924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__S1
timestamp 1688980957
transform 1 0 55476 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__S0
timestamp 1688980957
transform 1 0 50508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__S1
timestamp 1688980957
transform 1 0 52072 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__S
timestamp 1688980957
transform 1 0 55476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1688980957
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__S0
timestamp 1688980957
transform 1 0 56580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__S1
timestamp 1688980957
transform 1 0 56028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__S0
timestamp 1688980957
transform 1 0 55844 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__S1
timestamp 1688980957
transform 1 0 56212 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__S
timestamp 1688980957
transform 1 0 56212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1688980957
transform 1 0 58052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__S0
timestamp 1688980957
transform 1 0 55568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__S1
timestamp 1688980957
transform 1 0 56212 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__S0
timestamp 1688980957
transform 1 0 56304 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__S1
timestamp 1688980957
transform 1 0 53728 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__S
timestamp 1688980957
transform 1 0 57868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1688980957
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S0
timestamp 1688980957
transform 1 0 55108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__S1
timestamp 1688980957
transform 1 0 55476 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__S0
timestamp 1688980957
transform 1 0 55476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__S1
timestamp 1688980957
transform 1 0 55936 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__S
timestamp 1688980957
transform 1 0 56764 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1688980957
transform 1 0 55660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__S
timestamp 1688980957
transform 1 0 29072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__S
timestamp 1688980957
transform 1 0 28520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__S
timestamp 1688980957
transform 1 0 28520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__S
timestamp 1688980957
transform 1 0 41308 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__S
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__S
timestamp 1688980957
transform 1 0 38272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__S
timestamp 1688980957
transform 1 0 38916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__S
timestamp 1688980957
transform 1 0 40848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__S
timestamp 1688980957
transform 1 0 41584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__S
timestamp 1688980957
transform 1 0 46276 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__S
timestamp 1688980957
transform 1 0 46368 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__S
timestamp 1688980957
transform 1 0 48300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__S
timestamp 1688980957
transform 1 0 50324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__S
timestamp 1688980957
transform 1 0 48760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__S
timestamp 1688980957
transform 1 0 52440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__S
timestamp 1688980957
transform 1 0 55844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__S
timestamp 1688980957
transform 1 0 55844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__S
timestamp 1688980957
transform 1 0 55660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__S
timestamp 1688980957
transform 1 0 56212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__S
timestamp 1688980957
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__S
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__S
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__S
timestamp 1688980957
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__S
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__S
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__S
timestamp 1688980957
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__S
timestamp 1688980957
transform 1 0 19780 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__S
timestamp 1688980957
transform 1 0 19596 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__S
timestamp 1688980957
transform 1 0 20608 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__S
timestamp 1688980957
transform 1 0 24564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__S
timestamp 1688980957
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__S
timestamp 1688980957
transform 1 0 26128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__S
timestamp 1688980957
transform 1 0 29992 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__S
timestamp 1688980957
transform 1 0 30176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__S
timestamp 1688980957
transform 1 0 30360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__S
timestamp 1688980957
transform 1 0 41124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__S
timestamp 1688980957
transform 1 0 34868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__S
timestamp 1688980957
transform 1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__S
timestamp 1688980957
transform 1 0 40020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__S
timestamp 1688980957
transform 1 0 40940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__S
timestamp 1688980957
transform 1 0 42044 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__S
timestamp 1688980957
transform 1 0 43700 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__S
timestamp 1688980957
transform 1 0 53268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__S
timestamp 1688980957
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__S
timestamp 1688980957
transform 1 0 52072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__S
timestamp 1688980957
transform 1 0 49864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__S
timestamp 1688980957
transform 1 0 52440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__S
timestamp 1688980957
transform 1 0 57040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__S
timestamp 1688980957
transform 1 0 56396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__S
timestamp 1688980957
transform 1 0 56672 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__S
timestamp 1688980957
transform 1 0 57408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__S
timestamp 1688980957
transform 1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__S
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__S
timestamp 1688980957
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__S
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__S
timestamp 1688980957
transform 1 0 10580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__S
timestamp 1688980957
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__S
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__S
timestamp 1688980957
transform 1 0 17848 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__S
timestamp 1688980957
transform 1 0 16928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__S
timestamp 1688980957
transform 1 0 19596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__S
timestamp 1688980957
transform 1 0 22264 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__S
timestamp 1688980957
transform 1 0 24564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__S
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__S
timestamp 1688980957
transform 1 0 27876 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__S
timestamp 1688980957
transform 1 0 27232 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__S
timestamp 1688980957
transform 1 0 28520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__S
timestamp 1688980957
transform 1 0 35236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__S
timestamp 1688980957
transform 1 0 32752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__S
timestamp 1688980957
transform 1 0 35052 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__S
timestamp 1688980957
transform 1 0 38088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__S
timestamp 1688980957
transform 1 0 42136 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__S
timestamp 1688980957
transform 1 0 39100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__S
timestamp 1688980957
transform 1 0 40664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__S
timestamp 1688980957
transform 1 0 43148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__S
timestamp 1688980957
transform 1 0 44896 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__S
timestamp 1688980957
transform 1 0 47840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__S
timestamp 1688980957
transform 1 0 46368 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__S
timestamp 1688980957
transform 1 0 50508 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__S
timestamp 1688980957
transform 1 0 51704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__S
timestamp 1688980957
transform 1 0 55476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__S
timestamp 1688980957
transform 1 0 55108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__S
timestamp 1688980957
transform 1 0 56304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A_N
timestamp 1688980957
transform 1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A_N
timestamp 1688980957
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A_N
timestamp 1688980957
transform 1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B
timestamp 1688980957
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__S
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__S
timestamp 1688980957
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__S
timestamp 1688980957
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__S
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__S
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__S
timestamp 1688980957
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__S
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__S
timestamp 1688980957
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__S
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__S
timestamp 1688980957
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__S
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__S
timestamp 1688980957
transform 1 0 23276 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__S
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__S
timestamp 1688980957
transform 1 0 27416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__S
timestamp 1688980957
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__S
timestamp 1688980957
transform 1 0 26496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__S
timestamp 1688980957
transform 1 0 39376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__S
timestamp 1688980957
transform 1 0 34132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__S
timestamp 1688980957
transform 1 0 35696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__S
timestamp 1688980957
transform 1 0 38272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__S
timestamp 1688980957
transform 1 0 40388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__S
timestamp 1688980957
transform 1 0 38824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__S
timestamp 1688980957
transform 1 0 41308 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__S
timestamp 1688980957
transform 1 0 44068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__S
timestamp 1688980957
transform 1 0 47012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__S
timestamp 1688980957
transform 1 0 49956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__S
timestamp 1688980957
transform 1 0 46828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__S
timestamp 1688980957
transform 1 0 51428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__S
timestamp 1688980957
transform 1 0 55292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__S
timestamp 1688980957
transform 1 0 51520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__S
timestamp 1688980957
transform 1 0 55936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__S
timestamp 1688980957
transform 1 0 54464 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__S
timestamp 1688980957
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__S
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__S
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__S
timestamp 1688980957
transform 1 0 9752 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__S
timestamp 1688980957
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__S
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__S
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__S
timestamp 1688980957
transform 1 0 18216 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__S
timestamp 1688980957
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__S
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__S
timestamp 1688980957
transform 1 0 22080 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__S
timestamp 1688980957
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__S
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__S
timestamp 1688980957
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__S
timestamp 1688980957
transform 1 0 28520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__S
timestamp 1688980957
transform 1 0 28244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__S
timestamp 1688980957
transform 1 0 35144 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__S
timestamp 1688980957
transform 1 0 36800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__S
timestamp 1688980957
transform 1 0 35604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__S
timestamp 1688980957
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__S
timestamp 1688980957
transform 1 0 40756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__S
timestamp 1688980957
transform 1 0 39652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__S
timestamp 1688980957
transform 1 0 42504 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__S
timestamp 1688980957
transform 1 0 43700 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__S
timestamp 1688980957
transform 1 0 46184 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__S
timestamp 1688980957
transform 1 0 47748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__S
timestamp 1688980957
transform 1 0 47196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__S
timestamp 1688980957
transform 1 0 50324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__S
timestamp 1688980957
transform 1 0 50784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__S
timestamp 1688980957
transform 1 0 51888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__S
timestamp 1688980957
transform 1 0 54556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__S
timestamp 1688980957
transform 1 0 54188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__S
timestamp 1688980957
transform 1 0 7360 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__S
timestamp 1688980957
transform 1 0 12788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__S
timestamp 1688980957
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__S
timestamp 1688980957
transform 1 0 11316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__S
timestamp 1688980957
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__S
timestamp 1688980957
transform 1 0 14812 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__S
timestamp 1688980957
transform 1 0 15364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__S
timestamp 1688980957
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__S
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__S
timestamp 1688980957
transform 1 0 20516 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__S
timestamp 1688980957
transform 1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__S
timestamp 1688980957
transform 1 0 27968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__S
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__S
timestamp 1688980957
transform 1 0 29992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__S
timestamp 1688980957
transform 1 0 29808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__S
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__S
timestamp 1688980957
transform 1 0 36984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__S
timestamp 1688980957
transform 1 0 35512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__S
timestamp 1688980957
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__S
timestamp 1688980957
transform 1 0 39100 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__S
timestamp 1688980957
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__S
timestamp 1688980957
transform 1 0 41676 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__S
timestamp 1688980957
transform 1 0 45724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S
timestamp 1688980957
transform 1 0 46368 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__S
timestamp 1688980957
transform 1 0 49036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__S
timestamp 1688980957
transform 1 0 49036 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__S
timestamp 1688980957
transform 1 0 47564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S
timestamp 1688980957
transform 1 0 50140 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__S
timestamp 1688980957
transform 1 0 50876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__S
timestamp 1688980957
transform 1 0 58052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S
timestamp 1688980957
transform 1 0 56304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S
timestamp 1688980957
transform 1 0 56672 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__S
timestamp 1688980957
transform 1 0 7268 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S
timestamp 1688980957
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__S
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S
timestamp 1688980957
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S
timestamp 1688980957
transform 1 0 16192 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__S
timestamp 1688980957
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__S
timestamp 1688980957
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__S
timestamp 1688980957
transform 1 0 22448 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__S
timestamp 1688980957
transform 1 0 26036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S
timestamp 1688980957
transform 1 0 25668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__S
timestamp 1688980957
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__S
timestamp 1688980957
transform 1 0 29992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S
timestamp 1688980957
transform 1 0 31372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S
timestamp 1688980957
transform 1 0 31832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__S
timestamp 1688980957
transform 1 0 37352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__S
timestamp 1688980957
transform 1 0 37444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S
timestamp 1688980957
transform 1 0 38272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S
timestamp 1688980957
transform 1 0 39008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp 1688980957
transform 1 0 41768 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__S
timestamp 1688980957
transform 1 0 42596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S
timestamp 1688980957
transform 1 0 44436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S
timestamp 1688980957
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp 1688980957
transform 1 0 48208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__S
timestamp 1688980957
transform 1 0 50600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S
timestamp 1688980957
transform 1 0 48852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S
timestamp 1688980957
transform 1 0 52440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__S
timestamp 1688980957
transform 1 0 53728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__S
timestamp 1688980957
transform 1 0 58420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__S
timestamp 1688980957
transform 1 0 57500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__S
timestamp 1688980957
transform 1 0 56856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1688980957
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__S
timestamp 1688980957
transform 1 0 3680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__S
timestamp 1688980957
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S
timestamp 1688980957
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__S
timestamp 1688980957
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__S
timestamp 1688980957
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__S
timestamp 1688980957
transform 1 0 18216 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__S
timestamp 1688980957
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__S
timestamp 1688980957
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__S
timestamp 1688980957
transform 1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__S
timestamp 1688980957
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__S
timestamp 1688980957
transform 1 0 22632 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__S
timestamp 1688980957
transform 1 0 29716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__S
timestamp 1688980957
transform 1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__S
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__S
timestamp 1688980957
transform 1 0 38180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__S
timestamp 1688980957
transform 1 0 33028 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__S
timestamp 1688980957
transform 1 0 35328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__S
timestamp 1688980957
transform 1 0 38088 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__S
timestamp 1688980957
transform 1 0 38088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__S
timestamp 1688980957
transform 1 0 39008 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__S
timestamp 1688980957
transform 1 0 41308 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S
timestamp 1688980957
transform 1 0 50692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__S
timestamp 1688980957
transform 1 0 44988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__S
timestamp 1688980957
transform 1 0 48116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__S
timestamp 1688980957
transform 1 0 48576 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__S
timestamp 1688980957
transform 1 0 50416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__S
timestamp 1688980957
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__S
timestamp 1688980957
transform 1 0 52072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__S
timestamp 1688980957
transform 1 0 54188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__S
timestamp 1688980957
transform 1 0 53912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__S
timestamp 1688980957
transform 1 0 5244 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__S
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__S
timestamp 1688980957
transform 1 0 9844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__S
timestamp 1688980957
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__S
timestamp 1688980957
transform 1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__S
timestamp 1688980957
transform 1 0 16192 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__S
timestamp 1688980957
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__S
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__S
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__S
timestamp 1688980957
transform 1 0 19688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__S
timestamp 1688980957
transform 1 0 24840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__S
timestamp 1688980957
transform 1 0 23276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__S
timestamp 1688980957
transform 1 0 24840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__CLK
timestamp 1688980957
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__CLK
timestamp 1688980957
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__CLK
timestamp 1688980957
transform 1 0 33396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__CLK
timestamp 1688980957
transform 1 0 37720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__CLK
timestamp 1688980957
transform 1 0 32936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__CLK
timestamp 1688980957
transform 1 0 36892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__CLK
timestamp 1688980957
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__CLK
timestamp 1688980957
transform 1 0 39376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__CLK
timestamp 1688980957
transform 1 0 43976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__CLK
timestamp 1688980957
transform 1 0 43332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__CLK
timestamp 1688980957
transform 1 0 47196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__CLK
timestamp 1688980957
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__CLK
timestamp 1688980957
transform 1 0 50692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__CLK
timestamp 1688980957
transform 1 0 56764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__CLK
timestamp 1688980957
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__CLK
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__CLK
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__CLK
timestamp 1688980957
transform 1 0 23276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__CLK
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__CLK
timestamp 1688980957
transform 1 0 27324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__CLK
timestamp 1688980957
transform 1 0 31556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__CLK
timestamp 1688980957
transform 1 0 29992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__CLK
timestamp 1688980957
transform 1 0 42044 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__CLK
timestamp 1688980957
transform 1 0 34868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__CLK
timestamp 1688980957
transform 1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__CLK
timestamp 1688980957
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__CLK
timestamp 1688980957
transform 1 0 41400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__CLK
timestamp 1688980957
transform 1 0 43332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__CLK
timestamp 1688980957
transform 1 0 48116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__CLK
timestamp 1688980957
transform 1 0 53636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__CLK
timestamp 1688980957
transform 1 0 57408 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__CLK
timestamp 1688980957
transform 1 0 3680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__CLK
timestamp 1688980957
transform 1 0 8096 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__CLK
timestamp 1688980957
transform 1 0 11960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__CLK
timestamp 1688980957
transform 1 0 12880 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__CLK
timestamp 1688980957
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__CLK
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__CLK
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__CLK
timestamp 1688980957
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__CLK
timestamp 1688980957
transform 1 0 22264 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__CLK
timestamp 1688980957
transform 1 0 27232 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__CLK
timestamp 1688980957
transform 1 0 27232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__CLK
timestamp 1688980957
transform 1 0 34868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__CLK
timestamp 1688980957
transform 1 0 33948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__CLK
timestamp 1688980957
transform 1 0 35420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__CLK
timestamp 1688980957
transform 1 0 39468 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__CLK
timestamp 1688980957
transform 1 0 43332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__CLK
timestamp 1688980957
transform 1 0 40112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__CLK
timestamp 1688980957
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__CLK
timestamp 1688980957
transform 1 0 44344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__CLK
timestamp 1688980957
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__CLK
timestamp 1688980957
transform 1 0 45816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__CLK
timestamp 1688980957
transform 1 0 49864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__CLK
timestamp 1688980957
transform 1 0 54740 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__CLK
timestamp 1688980957
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__CLK
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__CLK
timestamp 1688980957
transform 1 0 17572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__CLK
timestamp 1688980957
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__CLK
timestamp 1688980957
transform 1 0 24012 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__CLK
timestamp 1688980957
transform 1 0 29716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__CLK
timestamp 1688980957
transform 1 0 27232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__CLK
timestamp 1688980957
transform 1 0 40756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__CLK
timestamp 1688980957
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__CLK
timestamp 1688980957
transform 1 0 32384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__CLK
timestamp 1688980957
transform 1 0 38640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__CLK
timestamp 1688980957
transform 1 0 37628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__CLK
timestamp 1688980957
transform 1 0 40388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__CLK
timestamp 1688980957
transform 1 0 42412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__CLK
timestamp 1688980957
transform 1 0 46736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__CLK
timestamp 1688980957
transform 1 0 44620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__CLK
timestamp 1688980957
transform 1 0 47748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__CLK
timestamp 1688980957
transform 1 0 46644 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__CLK
timestamp 1688980957
transform 1 0 54372 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__CLK
timestamp 1688980957
transform 1 0 3956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__CLK
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__CLK
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__CLK
timestamp 1688980957
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__CLK
timestamp 1688980957
transform 1 0 17940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__CLK
timestamp 1688980957
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__CLK
timestamp 1688980957
transform 1 0 22080 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__CLK
timestamp 1688980957
transform 1 0 27968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__CLK
timestamp 1688980957
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__CLK
timestamp 1688980957
transform 1 0 34132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__CLK
timestamp 1688980957
transform 1 0 33488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__CLK
timestamp 1688980957
transform 1 0 34132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__CLK
timestamp 1688980957
transform 1 0 38640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__CLK
timestamp 1688980957
transform 1 0 42964 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__CLK
timestamp 1688980957
transform 1 0 40020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__CLK
timestamp 1688980957
transform 1 0 42228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__CLK
timestamp 1688980957
transform 1 0 42228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__CLK
timestamp 1688980957
transform 1 0 44160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__CLK
timestamp 1688980957
transform 1 0 46368 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__CLK
timestamp 1688980957
transform 1 0 50048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__CLK
timestamp 1688980957
transform 1 0 6256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__CLK
timestamp 1688980957
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__CLK
timestamp 1688980957
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__CLK
timestamp 1688980957
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__CLK
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__CLK
timestamp 1688980957
transform 1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__CLK
timestamp 1688980957
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__CLK
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__CLK
timestamp 1688980957
transform 1 0 24196 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__CLK
timestamp 1688980957
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__CLK
timestamp 1688980957
transform 1 0 31004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__CLK
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__CLK
timestamp 1688980957
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__CLK
timestamp 1688980957
transform 1 0 36800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__CLK
timestamp 1688980957
transform 1 0 35420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__CLK
timestamp 1688980957
transform 1 0 40020 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__CLK
timestamp 1688980957
transform 1 0 42872 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__CLK
timestamp 1688980957
transform 1 0 41216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__CLK
timestamp 1688980957
transform 1 0 42964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__CLK
timestamp 1688980957
transform 1 0 44344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__CLK
timestamp 1688980957
transform 1 0 47380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__CLK
timestamp 1688980957
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__CLK
timestamp 1688980957
transform 1 0 52256 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__CLK
timestamp 1688980957
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__CLK
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__CLK
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__CLK
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__CLK
timestamp 1688980957
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__CLK
timestamp 1688980957
transform 1 0 19412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__CLK
timestamp 1688980957
transform 1 0 24564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__CLK
timestamp 1688980957
transform 1 0 27140 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__CLK
timestamp 1688980957
transform 1 0 31648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__CLK
timestamp 1688980957
transform 1 0 31464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__CLK
timestamp 1688980957
transform 1 0 32108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__CLK
timestamp 1688980957
transform 1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__CLK
timestamp 1688980957
transform 1 0 36892 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__CLK
timestamp 1688980957
transform 1 0 35696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__CLK
timestamp 1688980957
transform 1 0 41308 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__CLK
timestamp 1688980957
transform 1 0 43240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__CLK
timestamp 1688980957
transform 1 0 44068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__CLK
timestamp 1688980957
transform 1 0 43516 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__CLK
timestamp 1688980957
transform 1 0 45172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__CLK
timestamp 1688980957
transform 1 0 47380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__CLK
timestamp 1688980957
transform 1 0 48300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__CLK
timestamp 1688980957
transform 1 0 53544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1688980957
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1688980957
transform 1 0 21528 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__CLK
timestamp 1688980957
transform 1 0 21988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1688980957
transform 1 0 29164 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__CLK
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1688980957
transform 1 0 37444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1688980957
transform 1 0 31280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__CLK
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1688980957
transform 1 0 36432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__CLK
timestamp 1688980957
transform 1 0 38180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1688980957
transform 1 0 40204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__CLK
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1688980957
transform 1 0 46736 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1688980957
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1688980957
transform 1 0 48484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__CLK
timestamp 1688980957
transform 1 0 54372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__CLK
timestamp 1688980957
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1688980957
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1688980957
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__CLK
timestamp 1688980957
transform 1 0 22724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__CLK
timestamp 1688980957
transform 1 0 27140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1688980957
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1688980957
transform 1 0 14996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1688980957
transform 1 0 29532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1688980957
transform 1 0 41768 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1688980957
transform 1 0 52440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1688980957
transform 1 0 41952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1688980957
transform 1 0 52440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1688980957
transform 1 0 34868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1688980957
transform 1 0 22080 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout1_A
timestamp 1688980957
transform 1 0 27140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout2_A
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1688980957
transform 1 0 34776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1688980957
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 1688980957
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 1688980957
transform 1 0 35236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 1688980957
transform 1 0 34868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 1688980957
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1688980957
transform 1 0 36156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 1688980957
transform 1 0 27508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp 1688980957
transform 1 0 12420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 1688980957
transform 1 0 32568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 1688980957
transform 1 0 32292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 1688980957
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 1688980957
transform 1 0 6808 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout123_A
timestamp 1688980957
transform 1 0 30084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 1688980957
transform 1 0 47196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp 1688980957
transform 1 0 44896 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout129_A
timestamp 1688980957
transform 1 0 29532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold558_A
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1688980957
transform 1 0 19780 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 39008 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1688980957
transform 1 0 9016 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1688980957
transform 1 0 13156 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1688980957
transform 1 0 29716 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1688980957
transform 1 0 42412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1688980957
transform 1 0 53176 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1688980957
transform 1 0 42136 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1688980957
transform 1 0 52716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1688980957
transform 1 0 43884 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1688980957
transform 1 0 32476 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1688980957
transform 1 0 20240 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout2
timestamp 1688980957
transform 1 0 5888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout102 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout103
timestamp 1688980957
transform 1 0 33488 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout104
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout105
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout106
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout107
timestamp 1688980957
transform 1 0 36524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout108
timestamp 1688980957
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout109
timestamp 1688980957
transform 1 0 35420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout110
timestamp 1688980957
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout111
timestamp 1688980957
transform 1 0 33580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout112
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout113
timestamp 1688980957
transform 1 0 34868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout114
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout115
timestamp 1688980957
transform 1 0 12052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout116
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout117
timestamp 1688980957
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout119 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout120
timestamp 1688980957
transform 1 0 32016 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout121 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6440 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout122
timestamp 1688980957
transform 1 0 6624 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout123
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout124
timestamp 1688980957
transform 1 0 46000 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout125 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout126
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout127
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout128
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout129
timestamp 1688980957
transform 1 0 29716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout130
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_36
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_465
timestamp 1688980957
transform 1 0 43884 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_474
timestamp 1688980957
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_533
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_537
timestamp 1688980957
transform 1 0 50508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_555
timestamp 1688980957
transform 1 0 52164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_559
timestamp 1688980957
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_577
timestamp 1688980957
transform 1 0 54188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_581
timestamp 1688980957
transform 1 0 54556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_586
timestamp 1688980957
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_614
timestamp 1688980957
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_122
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_172
timestamp 1688980957
transform 1 0 16928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_185
timestamp 1688980957
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_229 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_380
timestamp 1688980957
transform 1 0 36064 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1688980957
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_430
timestamp 1688980957
transform 1 0 40664 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_466
timestamp 1688980957
transform 1 0 43976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_545
timestamp 1688980957
transform 1 0 51244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_569
timestamp 1688980957
transform 1 0 53452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_599
timestamp 1688980957
transform 1 0 56212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_23
timestamp 1688980957
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_58
timestamp 1688980957
transform 1 0 6440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_100 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_131
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_193
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_274
timestamp 1688980957
transform 1 0 26312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_281
timestamp 1688980957
transform 1 0 26956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_337
timestamp 1688980957
transform 1 0 32108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_354
timestamp 1688980957
transform 1 0 33672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_376
timestamp 1688980957
transform 1 0 35696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_402
timestamp 1688980957
transform 1 0 38088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_446
timestamp 1688980957
transform 1 0 42136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_502
timestamp 1688980957
transform 1 0 47288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_530
timestamp 1688980957
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_537
timestamp 1688980957
transform 1 0 50508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_605
timestamp 1688980957
transform 1 0 56764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_11
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_24
timestamp 1688980957
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_28
timestamp 1688980957
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_44
timestamp 1688980957
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_48
timestamp 1688980957
transform 1 0 5520 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_52
timestamp 1688980957
transform 1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_62
timestamp 1688980957
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_67
timestamp 1688980957
transform 1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_195
timestamp 1688980957
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_233
timestamp 1688980957
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_267
timestamp 1688980957
transform 1 0 25668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_276
timestamp 1688980957
transform 1 0 26496 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_284
timestamp 1688980957
transform 1 0 27232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_291
timestamp 1688980957
transform 1 0 27876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_314
timestamp 1688980957
transform 1 0 29992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_388
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_413
timestamp 1688980957
transform 1 0 39100 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_422
timestamp 1688980957
transform 1 0 39928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_502
timestamp 1688980957
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_505
timestamp 1688980957
transform 1 0 47564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_509
timestamp 1688980957
transform 1 0 47932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_545
timestamp 1688980957
transform 1 0 51244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_550
timestamp 1688980957
transform 1 0 51704 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1688980957
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_34
timestamp 1688980957
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_40
timestamp 1688980957
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_64
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_68
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_71
timestamp 1688980957
transform 1 0 7636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_131
timestamp 1688980957
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_158
timestamp 1688980957
transform 1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_185
timestamp 1688980957
transform 1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_213
timestamp 1688980957
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_239
timestamp 1688980957
transform 1 0 23092 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_280
timestamp 1688980957
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_285
timestamp 1688980957
transform 1 0 27324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_296
timestamp 1688980957
transform 1 0 28336 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_348
timestamp 1688980957
transform 1 0 33120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_362
timestamp 1688980957
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_471
timestamp 1688980957
transform 1 0 44436 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1688980957
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_542
timestamp 1688980957
transform 1 0 50968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_548
timestamp 1688980957
transform 1 0 51520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_552
timestamp 1688980957
transform 1 0 51888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_556
timestamp 1688980957
transform 1 0 52256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_584
timestamp 1688980957
transform 1 0 54832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_598
timestamp 1688980957
transform 1 0 56120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_38
timestamp 1688980957
transform 1 0 4600 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_67
timestamp 1688980957
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_71
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_82
timestamp 1688980957
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_91
timestamp 1688980957
transform 1 0 9476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_96
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_100
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_131
timestamp 1688980957
transform 1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_135
timestamp 1688980957
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_139
timestamp 1688980957
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_156
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_160
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_174
timestamp 1688980957
transform 1 0 17112 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_178
timestamp 1688980957
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_234
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_251
timestamp 1688980957
transform 1 0 24196 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_274
timestamp 1688980957
transform 1 0 26312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_290
timestamp 1688980957
transform 1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_306
timestamp 1688980957
transform 1 0 29256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_322
timestamp 1688980957
transform 1 0 30728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_330
timestamp 1688980957
transform 1 0 31464 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_334
timestamp 1688980957
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_341
timestamp 1688980957
transform 1 0 32476 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_345
timestamp 1688980957
transform 1 0 32844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_363
timestamp 1688980957
transform 1 0 34500 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 1688980957
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_446
timestamp 1688980957
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_468
timestamp 1688980957
transform 1 0 44160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_494
timestamp 1688980957
transform 1 0 46552 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_505
timestamp 1688980957
transform 1 0 47564 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_552
timestamp 1688980957
transform 1 0 51888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_556
timestamp 1688980957
transform 1 0 52256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_561
timestamp 1688980957
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_565
timestamp 1688980957
transform 1 0 53084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_569
timestamp 1688980957
transform 1 0 53452 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_36
timestamp 1688980957
transform 1 0 4416 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_42
timestamp 1688980957
transform 1 0 4968 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_64
timestamp 1688980957
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_78
timestamp 1688980957
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_89
timestamp 1688980957
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_105
timestamp 1688980957
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_113
timestamp 1688980957
transform 1 0 11500 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_123
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_127
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_131
timestamp 1688980957
transform 1 0 13156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_149
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_157
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_161
timestamp 1688980957
transform 1 0 15916 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_175
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_179
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_187
timestamp 1688980957
transform 1 0 18308 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_207
timestamp 1688980957
transform 1 0 20148 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_237
timestamp 1688980957
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_241
timestamp 1688980957
transform 1 0 23276 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_286
timestamp 1688980957
transform 1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_294
timestamp 1688980957
transform 1 0 28152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 1688980957
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_332
timestamp 1688980957
transform 1 0 31648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_336
timestamp 1688980957
transform 1 0 32016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_340
timestamp 1688980957
transform 1 0 32384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_344
timestamp 1688980957
transform 1 0 32752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_348
timestamp 1688980957
transform 1 0 33120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_360
timestamp 1688980957
transform 1 0 34224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_405
timestamp 1688980957
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_418
timestamp 1688980957
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_429
timestamp 1688980957
transform 1 0 40572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_452
timestamp 1688980957
transform 1 0 42688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_456
timestamp 1688980957
transform 1 0 43056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_465
timestamp 1688980957
transform 1 0 43884 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_474
timestamp 1688980957
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_494
timestamp 1688980957
transform 1 0 46552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_498
timestamp 1688980957
transform 1 0 46920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_525
timestamp 1688980957
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_529
timestamp 1688980957
transform 1 0 49772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_558
timestamp 1688980957
transform 1 0 52440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_584
timestamp 1688980957
transform 1 0 54832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_589
timestamp 1688980957
transform 1 0 55292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_624
timestamp 1688980957
transform 1 0 58512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_25
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_32
timestamp 1688980957
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_44
timestamp 1688980957
transform 1 0 5152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_92
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_100
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_122
timestamp 1688980957
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_155
timestamp 1688980957
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_173
timestamp 1688980957
transform 1 0 17020 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_179
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_182
timestamp 1688980957
transform 1 0 17848 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_188
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_191
timestamp 1688980957
transform 1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_199
timestamp 1688980957
transform 1 0 19412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_216
timestamp 1688980957
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_230
timestamp 1688980957
transform 1 0 22264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_234
timestamp 1688980957
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_238
timestamp 1688980957
transform 1 0 23000 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_243
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_257
timestamp 1688980957
transform 1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_272
timestamp 1688980957
transform 1 0 26128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_276
timestamp 1688980957
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_289
timestamp 1688980957
transform 1 0 27692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_306
timestamp 1688980957
transform 1 0 29256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_311
timestamp 1688980957
transform 1 0 29716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_334
timestamp 1688980957
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_345
timestamp 1688980957
transform 1 0 32844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_353
timestamp 1688980957
transform 1 0 33580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_360
timestamp 1688980957
transform 1 0 34224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_364
timestamp 1688980957
transform 1 0 34592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_379
timestamp 1688980957
transform 1 0 35972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_383
timestamp 1688980957
transform 1 0 36340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_387
timestamp 1688980957
transform 1 0 36708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_397
timestamp 1688980957
transform 1 0 37628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_401
timestamp 1688980957
transform 1 0 37996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_414
timestamp 1688980957
transform 1 0 39192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_418
timestamp 1688980957
transform 1 0 39560 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_422
timestamp 1688980957
transform 1 0 39928 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_426
timestamp 1688980957
transform 1 0 40296 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_430
timestamp 1688980957
transform 1 0 40664 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_435
timestamp 1688980957
transform 1 0 41124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_439
timestamp 1688980957
transform 1 0 41492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_443
timestamp 1688980957
transform 1 0 41860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_453
timestamp 1688980957
transform 1 0 42780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_457
timestamp 1688980957
transform 1 0 43148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_465
timestamp 1688980957
transform 1 0 43884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_469
timestamp 1688980957
transform 1 0 44252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_483
timestamp 1688980957
transform 1 0 45540 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_490
timestamp 1688980957
transform 1 0 46184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_494
timestamp 1688980957
transform 1 0 46552 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_498
timestamp 1688980957
transform 1 0 46920 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_502
timestamp 1688980957
transform 1 0 47288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_505
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_509
timestamp 1688980957
transform 1 0 47932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_513
timestamp 1688980957
transform 1 0 48300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_517
timestamp 1688980957
transform 1 0 48668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_521
timestamp 1688980957
transform 1 0 49036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_525
timestamp 1688980957
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_529
timestamp 1688980957
transform 1 0 49772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_533
timestamp 1688980957
transform 1 0 50140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_537
timestamp 1688980957
transform 1 0 50508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_541
timestamp 1688980957
transform 1 0 50876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_545
timestamp 1688980957
transform 1 0 51244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_549
timestamp 1688980957
transform 1 0 51612 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_553
timestamp 1688980957
transform 1 0 51980 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_577
timestamp 1688980957
transform 1 0 54188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_581
timestamp 1688980957
transform 1 0 54556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_37
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_49
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_57
timestamp 1688980957
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_90
timestamp 1688980957
transform 1 0 9384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_128
timestamp 1688980957
transform 1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_172
timestamp 1688980957
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_184
timestamp 1688980957
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_187
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_205
timestamp 1688980957
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_213
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_225
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_237
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1688980957
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_261
timestamp 1688980957
transform 1 0 25116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_273
timestamp 1688980957
transform 1 0 26220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_285
timestamp 1688980957
transform 1 0 27324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_291
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_313
timestamp 1688980957
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_316
timestamp 1688980957
transform 1 0 30176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_353
timestamp 1688980957
transform 1 0 33580 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_362
timestamp 1688980957
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_369
timestamp 1688980957
transform 1 0 35052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_373
timestamp 1688980957
transform 1 0 35420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_388
timestamp 1688980957
transform 1 0 36800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_392
timestamp 1688980957
transform 1 0 37168 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_396
timestamp 1688980957
transform 1 0 37536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_400
timestamp 1688980957
transform 1 0 37904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_425
timestamp 1688980957
transform 1 0 40204 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_429
timestamp 1688980957
transform 1 0 40572 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_437
timestamp 1688980957
transform 1 0 41308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_444
timestamp 1688980957
transform 1 0 41952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_448
timestamp 1688980957
transform 1 0 42320 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_452
timestamp 1688980957
transform 1 0 42688 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_456
timestamp 1688980957
transform 1 0 43056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_460
timestamp 1688980957
transform 1 0 43424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_465
timestamp 1688980957
transform 1 0 43884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_472
timestamp 1688980957
transform 1 0 44528 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_481
timestamp 1688980957
transform 1 0 45356 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_499
timestamp 1688980957
transform 1 0 47012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_503
timestamp 1688980957
transform 1 0 47380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_509
timestamp 1688980957
transform 1 0 47932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_513
timestamp 1688980957
transform 1 0 48300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_517
timestamp 1688980957
transform 1 0 48668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_523
timestamp 1688980957
transform 1 0 49220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_527
timestamp 1688980957
transform 1 0 49588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 1688980957
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_537
timestamp 1688980957
transform 1 0 50508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_540
timestamp 1688980957
transform 1 0 50784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_550
timestamp 1688980957
transform 1 0 51704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_589
timestamp 1688980957
transform 1 0 55292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_593
timestamp 1688980957
transform 1 0 55660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_597
timestamp 1688980957
transform 1 0 56028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_601
timestamp 1688980957
transform 1 0 56396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_624
timestamp 1688980957
transform 1 0 58512 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_24
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1688980957
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 1688980957
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_64
timestamp 1688980957
transform 1 0 6992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_129
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_146
timestamp 1688980957
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_185
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_212
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_216
timestamp 1688980957
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_265
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_269
timestamp 1688980957
transform 1 0 25852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_289
timestamp 1688980957
transform 1 0 27692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_297
timestamp 1688980957
transform 1 0 28428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_333
timestamp 1688980957
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_345
timestamp 1688980957
transform 1 0 32844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_357
timestamp 1688980957
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_389
timestamp 1688980957
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_401
timestamp 1688980957
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_432
timestamp 1688980957
transform 1 0 40848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_436
timestamp 1688980957
transform 1 0 41216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_440
timestamp 1688980957
transform 1 0 41584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_444
timestamp 1688980957
transform 1 0 41952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_453
timestamp 1688980957
transform 1 0 42780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_475
timestamp 1688980957
transform 1 0 44804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_502
timestamp 1688980957
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_505
timestamp 1688980957
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_518
timestamp 1688980957
transform 1 0 48760 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_549
timestamp 1688980957
transform 1 0 51612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_553
timestamp 1688980957
transform 1 0 51980 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_556
timestamp 1688980957
transform 1 0 52256 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_561
timestamp 1688980957
transform 1 0 52716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_587
timestamp 1688980957
transform 1 0 55108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_591
timestamp 1688980957
transform 1 0 55476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_595
timestamp 1688980957
transform 1 0 55844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_599
timestamp 1688980957
transform 1 0 56212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_603
timestamp 1688980957
transform 1 0 56580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_607
timestamp 1688980957
transform 1 0 56948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_617
timestamp 1688980957
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1688980957
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 1688980957
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_36
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_40
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_68
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_72
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_75
timestamp 1688980957
transform 1 0 8004 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_79
timestamp 1688980957
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_101
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_106
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_130
timestamp 1688980957
transform 1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_175
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_186
timestamp 1688980957
transform 1 0 18216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_206
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_235
timestamp 1688980957
transform 1 0 22724 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_262
timestamp 1688980957
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_288
timestamp 1688980957
transform 1 0 27600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_296
timestamp 1688980957
transform 1 0 28336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_306
timestamp 1688980957
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_313
timestamp 1688980957
transform 1 0 29900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_318
timestamp 1688980957
transform 1 0 30360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_322
timestamp 1688980957
transform 1 0 30728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_331
timestamp 1688980957
transform 1 0 31556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_335
timestamp 1688980957
transform 1 0 31924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_339
timestamp 1688980957
transform 1 0 32292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_395
timestamp 1688980957
transform 1 0 37444 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_414
timestamp 1688980957
transform 1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_418
timestamp 1688980957
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_442
timestamp 1688980957
transform 1 0 41768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_446
timestamp 1688980957
transform 1 0 42136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_474
timestamp 1688980957
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_498
timestamp 1688980957
transform 1 0 46920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_502
timestamp 1688980957
transform 1 0 47288 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_520
timestamp 1688980957
transform 1 0 48944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_557
timestamp 1688980957
transform 1 0 52348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_583
timestamp 1688980957
transform 1 0 54740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1688980957
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_589
timestamp 1688980957
transform 1 0 55292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_593
timestamp 1688980957
transform 1 0 55660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_597
timestamp 1688980957
transform 1 0 56028 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 1688980957
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_78
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_122
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_136
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_152
timestamp 1688980957
transform 1 0 15088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_178
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_290
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_294
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_302
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_307
timestamp 1688980957
transform 1 0 29348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_326
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_365
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_369
timestamp 1688980957
transform 1 0 35052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_388
timestamp 1688980957
transform 1 0 36800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_397
timestamp 1688980957
transform 1 0 37628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_431
timestamp 1688980957
transform 1 0 40756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_468
timestamp 1688980957
transform 1 0 44160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_499
timestamp 1688980957
transform 1 0 47012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 1688980957
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_521
timestamp 1688980957
transform 1 0 49036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_556
timestamp 1688980957
transform 1 0 52256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_561
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_573
timestamp 1688980957
transform 1 0 53820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_612
timestamp 1688980957
transform 1 0 57408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_11
timestamp 1688980957
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_34
timestamp 1688980957
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_38
timestamp 1688980957
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_79
timestamp 1688980957
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_101
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_117
timestamp 1688980957
transform 1 0 11868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_126
timestamp 1688980957
transform 1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_149
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_161
timestamp 1688980957
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_166
timestamp 1688980957
transform 1 0 16376 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_174
timestamp 1688980957
transform 1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_187
timestamp 1688980957
transform 1 0 18308 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_208
timestamp 1688980957
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_230
timestamp 1688980957
transform 1 0 22264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_239
timestamp 1688980957
transform 1 0 23092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_275
timestamp 1688980957
transform 1 0 26404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_279
timestamp 1688980957
transform 1 0 26772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_288
timestamp 1688980957
transform 1 0 27600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_296
timestamp 1688980957
transform 1 0 28336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_335
timestamp 1688980957
transform 1 0 31924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_361
timestamp 1688980957
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_369
timestamp 1688980957
transform 1 0 35052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_405
timestamp 1688980957
transform 1 0 38364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_417
timestamp 1688980957
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_430
timestamp 1688980957
transform 1 0 40664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_434
timestamp 1688980957
transform 1 0 41032 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_452
timestamp 1688980957
transform 1 0 42688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_456
timestamp 1688980957
transform 1 0 43056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_506
timestamp 1688980957
transform 1 0 47656 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_527
timestamp 1688980957
transform 1 0 49588 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1688980957
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_541
timestamp 1688980957
transform 1 0 50876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_553
timestamp 1688980957
transform 1 0 51980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_561
timestamp 1688980957
transform 1 0 52716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1688980957
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_589
timestamp 1688980957
transform 1 0 55292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_593
timestamp 1688980957
transform 1 0 55660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_623
timestamp 1688980957
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_30
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_42
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_122
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_148
timestamp 1688980957
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_152
timestamp 1688980957
transform 1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_159
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_163
timestamp 1688980957
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_198
timestamp 1688980957
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_202
timestamp 1688980957
transform 1 0 19688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_211
timestamp 1688980957
transform 1 0 20516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_233
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_243
timestamp 1688980957
transform 1 0 23460 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_247
timestamp 1688980957
transform 1 0 23828 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_258
timestamp 1688980957
transform 1 0 24840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_262
timestamp 1688980957
transform 1 0 25208 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_270
timestamp 1688980957
transform 1 0 25944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_331
timestamp 1688980957
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_341
timestamp 1688980957
transform 1 0 32476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_364
timestamp 1688980957
transform 1 0 34592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_368
timestamp 1688980957
transform 1 0 34960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_372
timestamp 1688980957
transform 1 0 35328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_386
timestamp 1688980957
transform 1 0 36616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_390
timestamp 1688980957
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_399
timestamp 1688980957
transform 1 0 37812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_411
timestamp 1688980957
transform 1 0 38916 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_423
timestamp 1688980957
transform 1 0 40020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_443
timestamp 1688980957
transform 1 0 41860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_457
timestamp 1688980957
transform 1 0 43148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_465
timestamp 1688980957
transform 1 0 43884 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_474
timestamp 1688980957
transform 1 0 44712 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_478
timestamp 1688980957
transform 1 0 45080 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_490
timestamp 1688980957
transform 1 0 46184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_494
timestamp 1688980957
transform 1 0 46552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_499
timestamp 1688980957
transform 1 0 47012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1688980957
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_505
timestamp 1688980957
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_533
timestamp 1688980957
transform 1 0 50140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_539
timestamp 1688980957
transform 1 0 50692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_548
timestamp 1688980957
transform 1 0 51520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_552
timestamp 1688980957
transform 1 0 51888 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_589
timestamp 1688980957
transform 1 0 55292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_597
timestamp 1688980957
transform 1 0 56028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_606
timestamp 1688980957
transform 1 0 56856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_610
timestamp 1688980957
transform 1 0 57224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_614
timestamp 1688980957
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_617
timestamp 1688980957
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_621
timestamp 1688980957
transform 1 0 58236 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_34
timestamp 1688980957
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_46
timestamp 1688980957
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_51
timestamp 1688980957
transform 1 0 5796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_118
timestamp 1688980957
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_190
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1688980957
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_220
timestamp 1688980957
transform 1 0 21344 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_230
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_240
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_257
timestamp 1688980957
transform 1 0 24748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_269
timestamp 1688980957
transform 1 0 25852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_281
timestamp 1688980957
transform 1 0 26956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_302
timestamp 1688980957
transform 1 0 28888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_339
timestamp 1688980957
transform 1 0 32292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_358
timestamp 1688980957
transform 1 0 34040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_369
timestamp 1688980957
transform 1 0 35052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_375
timestamp 1688980957
transform 1 0 35604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_402
timestamp 1688980957
transform 1 0 38088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_429
timestamp 1688980957
transform 1 0 40572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_435
timestamp 1688980957
transform 1 0 41124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_443
timestamp 1688980957
transform 1 0 41860 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_464
timestamp 1688980957
transform 1 0 43792 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_468
timestamp 1688980957
transform 1 0 44160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_472
timestamp 1688980957
transform 1 0 44528 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 1688980957
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 1688980957
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_489
timestamp 1688980957
transform 1 0 46092 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_494
timestamp 1688980957
transform 1 0 46552 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_506
timestamp 1688980957
transform 1 0 47656 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_512
timestamp 1688980957
transform 1 0 48208 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_515
timestamp 1688980957
transform 1 0 48484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_523
timestamp 1688980957
transform 1 0 49220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_528
timestamp 1688980957
transform 1 0 49680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_533
timestamp 1688980957
transform 1 0 50140 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_539
timestamp 1688980957
transform 1 0 50692 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_559
timestamp 1688980957
transform 1 0 52532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_571
timestamp 1688980957
transform 1 0 53636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_583
timestamp 1688980957
transform 1 0 54740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 1688980957
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_589
timestamp 1688980957
transform 1 0 55292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_593
timestamp 1688980957
transform 1 0 55660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_602
timestamp 1688980957
transform 1 0 56488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_623
timestamp 1688980957
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_28
timestamp 1688980957
transform 1 0 3680 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_34
timestamp 1688980957
transform 1 0 4232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_42
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_61
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_82
timestamp 1688980957
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_103
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_130
timestamp 1688980957
transform 1 0 13064 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_147
timestamp 1688980957
transform 1 0 14628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_178
timestamp 1688980957
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_233
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_250
timestamp 1688980957
transform 1 0 24104 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_254
timestamp 1688980957
transform 1 0 24472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_274
timestamp 1688980957
transform 1 0 26312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_328
timestamp 1688980957
transform 1 0 31280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_332
timestamp 1688980957
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_357
timestamp 1688980957
transform 1 0 33948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_367
timestamp 1688980957
transform 1 0 34868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_371
timestamp 1688980957
transform 1 0 35236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1688980957
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_402
timestamp 1688980957
transform 1 0 38088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_406
timestamp 1688980957
transform 1 0 38456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_432
timestamp 1688980957
transform 1 0 40848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_436
timestamp 1688980957
transform 1 0 41216 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_440
timestamp 1688980957
transform 1 0 41584 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_473
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_491
timestamp 1688980957
transform 1 0 46276 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_500
timestamp 1688980957
transform 1 0 47104 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_529
timestamp 1688980957
transform 1 0 49772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 1688980957
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_569
timestamp 1688980957
transform 1 0 53452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_577
timestamp 1688980957
transform 1 0 54188 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_594
timestamp 1688980957
transform 1 0 55752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_598
timestamp 1688980957
transform 1 0 56120 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_113
timestamp 1688980957
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_120
timestamp 1688980957
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_124
timestamp 1688980957
transform 1 0 12512 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_158
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_185
timestamp 1688980957
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_193
timestamp 1688980957
transform 1 0 18860 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_214
timestamp 1688980957
transform 1 0 20792 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_249
timestamp 1688980957
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 1688980957
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_313
timestamp 1688980957
transform 1 0 29900 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_317
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_329
timestamp 1688980957
transform 1 0 31372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_337
timestamp 1688980957
transform 1 0 32108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_403
timestamp 1688980957
transform 1 0 38180 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_430
timestamp 1688980957
transform 1 0 40664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_470
timestamp 1688980957
transform 1 0 44344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_493
timestamp 1688980957
transform 1 0 46460 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_570
timestamp 1688980957
transform 1 0 53544 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_576
timestamp 1688980957
transform 1 0 54096 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_615
timestamp 1688980957
transform 1 0 57684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_619
timestamp 1688980957
transform 1 0 58052 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_26
timestamp 1688980957
transform 1 0 3496 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_74
timestamp 1688980957
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_96
timestamp 1688980957
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_100
timestamp 1688980957
transform 1 0 10304 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_103
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_145
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_154
timestamp 1688980957
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_159
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_213
timestamp 1688980957
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_220
timestamp 1688980957
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1688980957
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_303
timestamp 1688980957
transform 1 0 28980 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_307
timestamp 1688980957
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_311
timestamp 1688980957
transform 1 0 29716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_323
timestamp 1688980957
transform 1 0 30820 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_332
timestamp 1688980957
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_377
timestamp 1688980957
transform 1 0 35788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_388
timestamp 1688980957
transform 1 0 36800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_401
timestamp 1688980957
transform 1 0 37996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_439
timestamp 1688980957
transform 1 0 41492 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_445
timestamp 1688980957
transform 1 0 42044 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_474
timestamp 1688980957
transform 1 0 44712 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_497
timestamp 1688980957
transform 1 0 46828 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_501
timestamp 1688980957
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_521
timestamp 1688980957
transform 1 0 49036 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_525
timestamp 1688980957
transform 1 0 49404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_539
timestamp 1688980957
transform 1 0 50692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_570
timestamp 1688980957
transform 1 0 53544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_590
timestamp 1688980957
transform 1 0 55384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 1688980957
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_617
timestamp 1688980957
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_45
timestamp 1688980957
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_49
timestamp 1688980957
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_61
timestamp 1688980957
transform 1 0 6716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1688980957
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_94
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_106
timestamp 1688980957
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_130
timestamp 1688980957
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_134
timestamp 1688980957
transform 1 0 13432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_157
timestamp 1688980957
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_161
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_169
timestamp 1688980957
transform 1 0 16652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_180
timestamp 1688980957
transform 1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_185
timestamp 1688980957
transform 1 0 18124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_203
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_206
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_210
timestamp 1688980957
transform 1 0 20424 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_222
timestamp 1688980957
transform 1 0 21528 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_227
timestamp 1688980957
transform 1 0 21988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_248
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_257
timestamp 1688980957
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_269
timestamp 1688980957
transform 1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_280
timestamp 1688980957
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_292
timestamp 1688980957
transform 1 0 27968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_313
timestamp 1688980957
transform 1 0 29900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_338
timestamp 1688980957
transform 1 0 32200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_354
timestamp 1688980957
transform 1 0 33672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_373
timestamp 1688980957
transform 1 0 35420 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_387
timestamp 1688980957
transform 1 0 36708 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_391
timestamp 1688980957
transform 1 0 37076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_403
timestamp 1688980957
transform 1 0 38180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_411
timestamp 1688980957
transform 1 0 38916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_414
timestamp 1688980957
transform 1 0 39192 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_425
timestamp 1688980957
transform 1 0 40204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_429
timestamp 1688980957
transform 1 0 40572 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_437
timestamp 1688980957
transform 1 0 41308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_442
timestamp 1688980957
transform 1 0 41768 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_455
timestamp 1688980957
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_467
timestamp 1688980957
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 1688980957
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_477
timestamp 1688980957
transform 1 0 44988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_504
timestamp 1688980957
transform 1 0 47472 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 1688980957
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_533
timestamp 1688980957
transform 1 0 50140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_552
timestamp 1688980957
transform 1 0 51888 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_597
timestamp 1688980957
transform 1 0 56028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_617
timestamp 1688980957
transform 1 0 57868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_32
timestamp 1688980957
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_44
timestamp 1688980957
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_71
timestamp 1688980957
transform 1 0 7636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_75
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_79
timestamp 1688980957
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_85
timestamp 1688980957
transform 1 0 8924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_97
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_124
timestamp 1688980957
transform 1 0 12512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_191
timestamp 1688980957
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_197
timestamp 1688980957
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_229
timestamp 1688980957
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_238
timestamp 1688980957
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_242
timestamp 1688980957
transform 1 0 23368 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_250
timestamp 1688980957
transform 1 0 24104 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_262
timestamp 1688980957
transform 1 0 25208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_271
timestamp 1688980957
transform 1 0 26036 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_277
timestamp 1688980957
transform 1 0 26588 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_309
timestamp 1688980957
transform 1 0 29532 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_315
timestamp 1688980957
transform 1 0 30084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_345
timestamp 1688980957
transform 1 0 32844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_366
timestamp 1688980957
transform 1 0 34776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_370
timestamp 1688980957
transform 1 0 35144 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_374
timestamp 1688980957
transform 1 0 35512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_378
timestamp 1688980957
transform 1 0 35880 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_423
timestamp 1688980957
transform 1 0 40020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_432
timestamp 1688980957
transform 1 0 40848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_446
timestamp 1688980957
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_457
timestamp 1688980957
transform 1 0 43148 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_469
timestamp 1688980957
transform 1 0 44252 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_481
timestamp 1688980957
transform 1 0 45356 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_493
timestamp 1688980957
transform 1 0 46460 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_501
timestamp 1688980957
transform 1 0 47196 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_505
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_509
timestamp 1688980957
transform 1 0 47932 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_520
timestamp 1688980957
transform 1 0 48944 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_532
timestamp 1688980957
transform 1 0 50048 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_540
timestamp 1688980957
transform 1 0 50784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_549
timestamp 1688980957
transform 1 0 51612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_558
timestamp 1688980957
transform 1 0 52440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_561
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_577
timestamp 1688980957
transform 1 0 54188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_589
timestamp 1688980957
transform 1 0 55292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_612
timestamp 1688980957
transform 1 0 57408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_58
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_70
timestamp 1688980957
transform 1 0 7544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_134
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_157
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_192
timestamp 1688980957
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_218
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_226
timestamp 1688980957
transform 1 0 21896 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_246
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_257
timestamp 1688980957
transform 1 0 24748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_269
timestamp 1688980957
transform 1 0 25852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_273
timestamp 1688980957
transform 1 0 26220 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_281
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_302
timestamp 1688980957
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_339
timestamp 1688980957
transform 1 0 32292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_361
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_403
timestamp 1688980957
transform 1 0 38180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_466
timestamp 1688980957
transform 1 0 43976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_470
timestamp 1688980957
transform 1 0 44344 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_488
timestamp 1688980957
transform 1 0 46000 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_492
timestamp 1688980957
transform 1 0 46368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_500
timestamp 1688980957
transform 1 0 47104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_505
timestamp 1688980957
transform 1 0 47564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_519
timestamp 1688980957
transform 1 0 48852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_523
timestamp 1688980957
transform 1 0 49220 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_531
timestamp 1688980957
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_533
timestamp 1688980957
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_545
timestamp 1688980957
transform 1 0 51244 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_549
timestamp 1688980957
transform 1 0 51612 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_561
timestamp 1688980957
transform 1 0 52716 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_573
timestamp 1688980957
transform 1 0 53820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_585
timestamp 1688980957
transform 1 0 54924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_589
timestamp 1688980957
transform 1 0 55292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_597
timestamp 1688980957
transform 1 0 56028 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_610
timestamp 1688980957
transform 1 0 57224 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_622
timestamp 1688980957
transform 1 0 58328 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_7
timestamp 1688980957
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_32
timestamp 1688980957
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_44
timestamp 1688980957
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_65
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_74
timestamp 1688980957
transform 1 0 7912 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_86
timestamp 1688980957
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_150
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_160
timestamp 1688980957
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_185
timestamp 1688980957
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_229
timestamp 1688980957
transform 1 0 22172 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_241
timestamp 1688980957
transform 1 0 23276 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1688980957
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_303
timestamp 1688980957
transform 1 0 28980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_333
timestamp 1688980957
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_341
timestamp 1688980957
transform 1 0 32476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_366
timestamp 1688980957
transform 1 0 34776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_370
timestamp 1688980957
transform 1 0 35144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_387
timestamp 1688980957
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_402
timestamp 1688980957
transform 1 0 38088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_422
timestamp 1688980957
transform 1 0 39928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_426
timestamp 1688980957
transform 1 0 40296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_465
timestamp 1688980957
transform 1 0 43884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_469
timestamp 1688980957
transform 1 0 44252 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 1688980957
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_529
timestamp 1688980957
transform 1 0 49772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_533
timestamp 1688980957
transform 1 0 50140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_558
timestamp 1688980957
transform 1 0 52440 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_561
timestamp 1688980957
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_573
timestamp 1688980957
transform 1 0 53820 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_599
timestamp 1688980957
transform 1 0 56212 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_611
timestamp 1688980957
transform 1 0 57316 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 1688980957
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_11
timestamp 1688980957
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_20
timestamp 1688980957
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_37
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_55
timestamp 1688980957
transform 1 0 6164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_102
timestamp 1688980957
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_114
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_120
timestamp 1688980957
transform 1 0 12144 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_129
timestamp 1688980957
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_151
timestamp 1688980957
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_163
timestamp 1688980957
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_175
timestamp 1688980957
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_222
timestamp 1688980957
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_288
timestamp 1688980957
transform 1 0 27600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_327
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_331
timestamp 1688980957
transform 1 0 31556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_335
timestamp 1688980957
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_339
timestamp 1688980957
transform 1 0 32292 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_342
timestamp 1688980957
transform 1 0 32568 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_354
timestamp 1688980957
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_362
timestamp 1688980957
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_373
timestamp 1688980957
transform 1 0 35420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_402
timestamp 1688980957
transform 1 0 38088 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_410
timestamp 1688980957
transform 1 0 38824 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_438
timestamp 1688980957
transform 1 0 41400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_469
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_473
timestamp 1688980957
transform 1 0 44620 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_566
timestamp 1688980957
transform 1 0 53176 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_623
timestamp 1688980957
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_98
timestamp 1688980957
transform 1 0 10120 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_108
timestamp 1688980957
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_135
timestamp 1688980957
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_185
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_188
timestamp 1688980957
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_192
timestamp 1688980957
transform 1 0 18768 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_203
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_207
timestamp 1688980957
transform 1 0 20148 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_211
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_220
timestamp 1688980957
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_243
timestamp 1688980957
transform 1 0 23460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_276
timestamp 1688980957
transform 1 0 26496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_285
timestamp 1688980957
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_304
timestamp 1688980957
transform 1 0 29072 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_316
timestamp 1688980957
transform 1 0 30176 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_328
timestamp 1688980957
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_353
timestamp 1688980957
transform 1 0 33580 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_365
timestamp 1688980957
transform 1 0 34684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_377
timestamp 1688980957
transform 1 0 35788 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_383
timestamp 1688980957
transform 1 0 36340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_397
timestamp 1688980957
transform 1 0 37628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_409
timestamp 1688980957
transform 1 0 38732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_417
timestamp 1688980957
transform 1 0 39468 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_421
timestamp 1688980957
transform 1 0 39836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_425
timestamp 1688980957
transform 1 0 40204 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 1688980957
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 1688980957
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 1688980957
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_453
timestamp 1688980957
transform 1 0 42780 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_469
timestamp 1688980957
transform 1 0 44252 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_475
timestamp 1688980957
transform 1 0 44804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 1688980957
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_537
timestamp 1688980957
transform 1 0 50508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_556
timestamp 1688980957
transform 1 0 52256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_561
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_567
timestamp 1688980957
transform 1 0 53268 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_571
timestamp 1688980957
transform 1 0 53636 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_590
timestamp 1688980957
transform 1 0 55384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_614
timestamp 1688980957
transform 1 0 57592 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_47
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_93
timestamp 1688980957
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_126
timestamp 1688980957
transform 1 0 12696 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_145
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_172
timestamp 1688980957
transform 1 0 16928 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_180
timestamp 1688980957
transform 1 0 17664 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_190
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_201
timestamp 1688980957
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_243
timestamp 1688980957
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_261
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_272
timestamp 1688980957
transform 1 0 26128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_303
timestamp 1688980957
transform 1 0 28980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_313
timestamp 1688980957
transform 1 0 29900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_318
timestamp 1688980957
transform 1 0 30360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_326
timestamp 1688980957
transform 1 0 31096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_354
timestamp 1688980957
transform 1 0 33672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_358
timestamp 1688980957
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_369
timestamp 1688980957
transform 1 0 35052 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_373
timestamp 1688980957
transform 1 0 35420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_385
timestamp 1688980957
transform 1 0 36524 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_393
timestamp 1688980957
transform 1 0 37260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_425
timestamp 1688980957
transform 1 0 40204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_456
timestamp 1688980957
transform 1 0 43056 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_462
timestamp 1688980957
transform 1 0 43608 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_474
timestamp 1688980957
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_485
timestamp 1688980957
transform 1 0 45724 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_493
timestamp 1688980957
transform 1 0 46460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_501
timestamp 1688980957
transform 1 0 47196 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_505
timestamp 1688980957
transform 1 0 47564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_511
timestamp 1688980957
transform 1 0 48116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_514
timestamp 1688980957
transform 1 0 48392 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_518
timestamp 1688980957
transform 1 0 48760 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_530
timestamp 1688980957
transform 1 0 49864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_576
timestamp 1688980957
transform 1 0 54096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_598
timestamp 1688980957
transform 1 0 56120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_602
timestamp 1688980957
transform 1 0 56488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_621
timestamp 1688980957
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_30
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_42
timestamp 1688980957
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_75
timestamp 1688980957
transform 1 0 8004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_106
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1688980957
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_160
timestamp 1688980957
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_197
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_245
timestamp 1688980957
transform 1 0 23644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_257
timestamp 1688980957
transform 1 0 24748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_267
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_275
timestamp 1688980957
transform 1 0 26404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_285
timestamp 1688980957
transform 1 0 27324 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_327
timestamp 1688980957
transform 1 0 31188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_347
timestamp 1688980957
transform 1 0 33028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_381
timestamp 1688980957
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_389
timestamp 1688980957
transform 1 0 36892 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_409
timestamp 1688980957
transform 1 0 38732 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_413
timestamp 1688980957
transform 1 0 39100 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_423
timestamp 1688980957
transform 1 0 40020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_427
timestamp 1688980957
transform 1 0 40388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_431
timestamp 1688980957
transform 1 0 40756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_457
timestamp 1688980957
transform 1 0 43148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_485
timestamp 1688980957
transform 1 0 45724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_489
timestamp 1688980957
transform 1 0 46092 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_493
timestamp 1688980957
transform 1 0 46460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_497
timestamp 1688980957
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_503
timestamp 1688980957
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_505
timestamp 1688980957
transform 1 0 47564 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_514
timestamp 1688980957
transform 1 0 48392 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_520
timestamp 1688980957
transform 1 0 48944 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_532
timestamp 1688980957
transform 1 0 50048 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_540
timestamp 1688980957
transform 1 0 50784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_544
timestamp 1688980957
transform 1 0 51152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_548
timestamp 1688980957
transform 1 0 51520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_556
timestamp 1688980957
transform 1 0 52256 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_578
timestamp 1688980957
transform 1 0 54280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_582
timestamp 1688980957
transform 1 0 54648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_586
timestamp 1688980957
transform 1 0 55016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_589
timestamp 1688980957
transform 1 0 55292 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_600
timestamp 1688980957
transform 1 0 56304 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_612
timestamp 1688980957
transform 1 0 57408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_37
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_49
timestamp 1688980957
transform 1 0 5612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_52
timestamp 1688980957
transform 1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_64
timestamp 1688980957
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_91
timestamp 1688980957
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_95
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_107
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_118
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_171
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_227
timestamp 1688980957
transform 1 0 21988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_231
timestamp 1688980957
transform 1 0 22356 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_247
timestamp 1688980957
transform 1 0 23828 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_257
timestamp 1688980957
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_269
timestamp 1688980957
transform 1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_274
timestamp 1688980957
transform 1 0 26312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_305
timestamp 1688980957
transform 1 0 29164 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_329
timestamp 1688980957
transform 1 0 31372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_344
timestamp 1688980957
transform 1 0 32752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_381
timestamp 1688980957
transform 1 0 36156 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_430
timestamp 1688980957
transform 1 0 40664 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_447
timestamp 1688980957
transform 1 0 42228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_451
timestamp 1688980957
transform 1 0 42596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_473
timestamp 1688980957
transform 1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_486
timestamp 1688980957
transform 1 0 45816 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_490
timestamp 1688980957
transform 1 0 46184 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_509
timestamp 1688980957
transform 1 0 47932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_513
timestamp 1688980957
transform 1 0 48300 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_530
timestamp 1688980957
transform 1 0 49864 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 1688980957
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_545
timestamp 1688980957
transform 1 0 51244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_549
timestamp 1688980957
transform 1 0 51612 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_574
timestamp 1688980957
transform 1 0 53912 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_586
timestamp 1688980957
transform 1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_597
timestamp 1688980957
transform 1 0 56028 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_609
timestamp 1688980957
transform 1 0 57132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_621
timestamp 1688980957
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_66
timestamp 1688980957
transform 1 0 7176 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_70
timestamp 1688980957
transform 1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_88
timestamp 1688980957
transform 1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_122
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_126
timestamp 1688980957
transform 1 0 12696 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_157
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_162
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_177
timestamp 1688980957
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_197
timestamp 1688980957
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1688980957
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_285
timestamp 1688980957
transform 1 0 27324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_289
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_306
timestamp 1688980957
transform 1 0 29256 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_331
timestamp 1688980957
transform 1 0 31556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_353
timestamp 1688980957
transform 1 0 33580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_364
timestamp 1688980957
transform 1 0 34592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_398
timestamp 1688980957
transform 1 0 37720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_437
timestamp 1688980957
transform 1 0 41308 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_457
timestamp 1688980957
transform 1 0 43148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_485
timestamp 1688980957
transform 1 0 45724 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_514
timestamp 1688980957
transform 1 0 48392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_518
timestamp 1688980957
transform 1 0 48760 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_545
timestamp 1688980957
transform 1 0 51244 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_557
timestamp 1688980957
transform 1 0 52348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_570
timestamp 1688980957
transform 1 0 53544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_595
timestamp 1688980957
transform 1 0 55844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_610
timestamp 1688980957
transform 1 0 57224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_614
timestamp 1688980957
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_7
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_24
timestamp 1688980957
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_66
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_135
timestamp 1688980957
transform 1 0 13524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_166
timestamp 1688980957
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_186
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1688980957
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_222
timestamp 1688980957
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_226
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_283
timestamp 1688980957
transform 1 0 27140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_287
timestamp 1688980957
transform 1 0 27508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_296
timestamp 1688980957
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_313
timestamp 1688980957
transform 1 0 29900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_339
timestamp 1688980957
transform 1 0 32292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_361
timestamp 1688980957
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_373
timestamp 1688980957
transform 1 0 35420 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_385
timestamp 1688980957
transform 1 0 36524 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_397
timestamp 1688980957
transform 1 0 37628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_400
timestamp 1688980957
transform 1 0 37904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_412
timestamp 1688980957
transform 1 0 39008 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_447
timestamp 1688980957
transform 1 0 42228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_459
timestamp 1688980957
transform 1 0 43332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_474
timestamp 1688980957
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_477
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_487
timestamp 1688980957
transform 1 0 45908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_508
timestamp 1688980957
transform 1 0 47840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_542
timestamp 1688980957
transform 1 0 50968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_546
timestamp 1688980957
transform 1 0 51336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_586
timestamp 1688980957
transform 1 0 55016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_589
timestamp 1688980957
transform 1 0 55292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_593
timestamp 1688980957
transform 1 0 55660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_622
timestamp 1688980957
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_11
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_29
timestamp 1688980957
transform 1 0 3772 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_33
timestamp 1688980957
transform 1 0 4140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_68
timestamp 1688980957
transform 1 0 7360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_96
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_100
timestamp 1688980957
transform 1 0 10304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_122
timestamp 1688980957
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_126
timestamp 1688980957
transform 1 0 12696 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_138
timestamp 1688980957
transform 1 0 13800 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_141
timestamp 1688980957
transform 1 0 14076 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_155
timestamp 1688980957
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_203
timestamp 1688980957
transform 1 0 19780 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_214
timestamp 1688980957
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 1688980957
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_233
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_245
timestamp 1688980957
transform 1 0 23644 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_255
timestamp 1688980957
transform 1 0 24564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_259
timestamp 1688980957
transform 1 0 24932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_289
timestamp 1688980957
transform 1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_297
timestamp 1688980957
transform 1 0 28428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_315
timestamp 1688980957
transform 1 0 30084 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_324
timestamp 1688980957
transform 1 0 30912 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_365
timestamp 1688980957
transform 1 0 34684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_369
timestamp 1688980957
transform 1 0 35052 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_376
timestamp 1688980957
transform 1 0 35696 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_388
timestamp 1688980957
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_399
timestamp 1688980957
transform 1 0 37812 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_416
timestamp 1688980957
transform 1 0 39376 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_428
timestamp 1688980957
transform 1 0 40480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_436
timestamp 1688980957
transform 1 0 41216 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_439
timestamp 1688980957
transform 1 0 41492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 1688980957
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_473
timestamp 1688980957
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_485
timestamp 1688980957
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_499
timestamp 1688980957
transform 1 0 47012 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_513
timestamp 1688980957
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_517
timestamp 1688980957
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_525
timestamp 1688980957
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_543
timestamp 1688980957
transform 1 0 51060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_555
timestamp 1688980957
transform 1 0 52164 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_585
timestamp 1688980957
transform 1 0 54924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_589
timestamp 1688980957
transform 1 0 55292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_612
timestamp 1688980957
transform 1 0 57408 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_19
timestamp 1688980957
transform 1 0 2852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_47
timestamp 1688980957
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_51
timestamp 1688980957
transform 1 0 5796 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_54
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_66
timestamp 1688980957
transform 1 0 7176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_78
timestamp 1688980957
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_117
timestamp 1688980957
transform 1 0 11868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_120
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_124
timestamp 1688980957
transform 1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_145
timestamp 1688980957
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_151
timestamp 1688980957
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_163
timestamp 1688980957
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_173
timestamp 1688980957
transform 1 0 17020 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_185
timestamp 1688980957
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1688980957
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 1688980957
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_225
timestamp 1688980957
transform 1 0 21804 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_242
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_285
timestamp 1688980957
transform 1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_290
timestamp 1688980957
transform 1 0 27784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_302
timestamp 1688980957
transform 1 0 28888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_313
timestamp 1688980957
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_351
timestamp 1688980957
transform 1 0 33396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_362
timestamp 1688980957
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_415
timestamp 1688980957
transform 1 0 39284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1688980957
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_435
timestamp 1688980957
transform 1 0 41124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_445
timestamp 1688980957
transform 1 0 42044 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_449
timestamp 1688980957
transform 1 0 42412 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 1688980957
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_469
timestamp 1688980957
transform 1 0 44252 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_473
timestamp 1688980957
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_477
timestamp 1688980957
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_481
timestamp 1688980957
transform 1 0 45356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_493
timestamp 1688980957
transform 1 0 46460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_501
timestamp 1688980957
transform 1 0 47196 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_511
timestamp 1688980957
transform 1 0 48116 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_515
timestamp 1688980957
transform 1 0 48484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_527
timestamp 1688980957
transform 1 0 49588 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_550
timestamp 1688980957
transform 1 0 51704 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_570
timestamp 1688980957
transform 1 0 53544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_585
timestamp 1688980957
transform 1 0 54924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_597
timestamp 1688980957
transform 1 0 56028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_601
timestamp 1688980957
transform 1 0 56396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_618
timestamp 1688980957
transform 1 0 57960 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_624
timestamp 1688980957
transform 1 0 58512 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_37
timestamp 1688980957
transform 1 0 4508 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_40
timestamp 1688980957
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_52
timestamp 1688980957
transform 1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_89
timestamp 1688980957
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_96
timestamp 1688980957
transform 1 0 9936 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_130
timestamp 1688980957
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_148
timestamp 1688980957
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_200
timestamp 1688980957
transform 1 0 19504 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_219
timestamp 1688980957
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_309
timestamp 1688980957
transform 1 0 29532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_355
timestamp 1688980957
transform 1 0 33764 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_359
timestamp 1688980957
transform 1 0 34132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_386
timestamp 1688980957
transform 1 0 36616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_390
timestamp 1688980957
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_397
timestamp 1688980957
transform 1 0 37628 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_403
timestamp 1688980957
transform 1 0 38180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_406
timestamp 1688980957
transform 1 0 38456 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_410
timestamp 1688980957
transform 1 0 38824 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_414
timestamp 1688980957
transform 1 0 39192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_426
timestamp 1688980957
transform 1 0 40296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_430
timestamp 1688980957
transform 1 0 40664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 1688980957
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_490
timestamp 1688980957
transform 1 0 46184 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_494
timestamp 1688980957
transform 1 0 46552 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_500
timestamp 1688980957
transform 1 0 47104 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 1688980957
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_521
timestamp 1688980957
transform 1 0 49036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_533
timestamp 1688980957
transform 1 0 50140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_545
timestamp 1688980957
transform 1 0 51244 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_556
timestamp 1688980957
transform 1 0 52256 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_573
timestamp 1688980957
transform 1 0 53820 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_582
timestamp 1688980957
transform 1 0 54648 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_594
timestamp 1688980957
transform 1 0 55752 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_602
timestamp 1688980957
transform 1 0 56488 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_9
timestamp 1688980957
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_38
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_42
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_69
timestamp 1688980957
transform 1 0 7452 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_73
timestamp 1688980957
transform 1 0 7820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_118
timestamp 1688980957
transform 1 0 11960 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_173
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_235
timestamp 1688980957
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_239
timestamp 1688980957
transform 1 0 23092 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_248
timestamp 1688980957
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_283
timestamp 1688980957
transform 1 0 27140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_302
timestamp 1688980957
transform 1 0 28888 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_330
timestamp 1688980957
transform 1 0 31464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_334
timestamp 1688980957
transform 1 0 31832 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_361
timestamp 1688980957
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_386
timestamp 1688980957
transform 1 0 36616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_406
timestamp 1688980957
transform 1 0 38456 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_410
timestamp 1688980957
transform 1 0 38824 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_437
timestamp 1688980957
transform 1 0 41308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_448
timestamp 1688980957
transform 1 0 42320 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_473
timestamp 1688980957
transform 1 0 44620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_486
timestamp 1688980957
transform 1 0 45816 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_512
timestamp 1688980957
transform 1 0 48208 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_529
timestamp 1688980957
transform 1 0 49772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_533
timestamp 1688980957
transform 1 0 50140 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_565
timestamp 1688980957
transform 1 0 53084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 1688980957
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_589
timestamp 1688980957
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_601
timestamp 1688980957
transform 1 0 56396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_605
timestamp 1688980957
transform 1 0 56764 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_622
timestamp 1688980957
transform 1 0 58328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_9
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_26
timestamp 1688980957
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_30
timestamp 1688980957
transform 1 0 3864 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1688980957
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_66
timestamp 1688980957
transform 1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_87
timestamp 1688980957
transform 1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_173
timestamp 1688980957
transform 1 0 17020 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_197
timestamp 1688980957
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_255
timestamp 1688980957
transform 1 0 24564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_259
timestamp 1688980957
transform 1 0 24932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_285
timestamp 1688980957
transform 1 0 27324 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_310
timestamp 1688980957
transform 1 0 29624 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_328
timestamp 1688980957
transform 1 0 31280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_332
timestamp 1688980957
transform 1 0 31648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_343
timestamp 1688980957
transform 1 0 32660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_387
timestamp 1688980957
transform 1 0 36708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_426
timestamp 1688980957
transform 1 0 40296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_458
timestamp 1688980957
transform 1 0 43240 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_483
timestamp 1688980957
transform 1 0 45540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_487
timestamp 1688980957
transform 1 0 45908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_543
timestamp 1688980957
transform 1 0 51060 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_554
timestamp 1688980957
transform 1 0 52072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_570
timestamp 1688980957
transform 1 0 53544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_579
timestamp 1688980957
transform 1 0 54372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_599
timestamp 1688980957
transform 1 0 56212 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_605
timestamp 1688980957
transform 1 0 56764 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_38
timestamp 1688980957
transform 1 0 4600 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_94
timestamp 1688980957
transform 1 0 9752 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_113
timestamp 1688980957
transform 1 0 11500 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_117
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_125
timestamp 1688980957
transform 1 0 12604 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_150
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_160
timestamp 1688980957
transform 1 0 15824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_181
timestamp 1688980957
transform 1 0 17756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_184
timestamp 1688980957
transform 1 0 18032 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1688980957
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_201
timestamp 1688980957
transform 1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_220
timestamp 1688980957
transform 1 0 21344 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_228
timestamp 1688980957
transform 1 0 22080 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_248
timestamp 1688980957
transform 1 0 23920 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_299
timestamp 1688980957
transform 1 0 28612 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_313
timestamp 1688980957
transform 1 0 29900 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_341
timestamp 1688980957
transform 1 0 32476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_352
timestamp 1688980957
transform 1 0 33488 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_361
timestamp 1688980957
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_369
timestamp 1688980957
transform 1 0 35052 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_373
timestamp 1688980957
transform 1 0 35420 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_379
timestamp 1688980957
transform 1 0 35972 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_388
timestamp 1688980957
transform 1 0 36800 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_392
timestamp 1688980957
transform 1 0 37168 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_411
timestamp 1688980957
transform 1 0 38916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_415
timestamp 1688980957
transform 1 0 39284 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1688980957
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_433
timestamp 1688980957
transform 1 0 40940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_439
timestamp 1688980957
transform 1 0 41492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_469
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 1688980957
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_493
timestamp 1688980957
transform 1 0 46460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_513
timestamp 1688980957
transform 1 0 48300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_517
timestamp 1688980957
transform 1 0 48668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_529
timestamp 1688980957
transform 1 0 49772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_533
timestamp 1688980957
transform 1 0 50140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_541
timestamp 1688980957
transform 1 0 50876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_545
timestamp 1688980957
transform 1 0 51244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_568
timestamp 1688980957
transform 1 0 53360 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_589
timestamp 1688980957
transform 1 0 55292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_623
timestamp 1688980957
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_29
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_33
timestamp 1688980957
transform 1 0 4140 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_37
timestamp 1688980957
transform 1 0 4508 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_45
timestamp 1688980957
transform 1 0 5244 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_66
timestamp 1688980957
transform 1 0 7176 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_70
timestamp 1688980957
transform 1 0 7544 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_86
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_95
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_99
timestamp 1688980957
transform 1 0 10212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_133
timestamp 1688980957
transform 1 0 13340 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_146
timestamp 1688980957
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_150
timestamp 1688980957
transform 1 0 14904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_189
timestamp 1688980957
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_199
timestamp 1688980957
transform 1 0 19412 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_203
timestamp 1688980957
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_215
timestamp 1688980957
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_256
timestamp 1688980957
transform 1 0 24656 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_266
timestamp 1688980957
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1688980957
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_313
timestamp 1688980957
transform 1 0 29900 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_324
timestamp 1688980957
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_403
timestamp 1688980957
transform 1 0 38180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_407
timestamp 1688980957
transform 1 0 38548 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_427
timestamp 1688980957
transform 1 0 40388 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_439
timestamp 1688980957
transform 1 0 41492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_444
timestamp 1688980957
transform 1 0 41952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_459
timestamp 1688980957
transform 1 0 43332 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_463
timestamp 1688980957
transform 1 0 43700 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_475
timestamp 1688980957
transform 1 0 44804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_483
timestamp 1688980957
transform 1 0 45540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_488
timestamp 1688980957
transform 1 0 46000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_502
timestamp 1688980957
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_505
timestamp 1688980957
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_509
timestamp 1688980957
transform 1 0 47932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_521
timestamp 1688980957
transform 1 0 49036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_535
timestamp 1688980957
transform 1 0 50324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_548
timestamp 1688980957
transform 1 0 51520 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_558
timestamp 1688980957
transform 1 0 52440 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_577
timestamp 1688980957
transform 1 0 54188 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_594
timestamp 1688980957
transform 1 0 55752 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_614
timestamp 1688980957
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_58
timestamp 1688980957
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_70
timestamp 1688980957
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_82
timestamp 1688980957
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_113
timestamp 1688980957
transform 1 0 11500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_125
timestamp 1688980957
transform 1 0 12604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1688980957
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_151
timestamp 1688980957
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_163
timestamp 1688980957
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_175
timestamp 1688980957
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_187
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_239
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_243
timestamp 1688980957
transform 1 0 23460 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1688980957
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_429
timestamp 1688980957
transform 1 0 40572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_441
timestamp 1688980957
transform 1 0 41676 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_453
timestamp 1688980957
transform 1 0 42780 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_465
timestamp 1688980957
transform 1 0 43884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_473
timestamp 1688980957
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_477
timestamp 1688980957
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_489
timestamp 1688980957
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_501
timestamp 1688980957
transform 1 0 47196 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_516
timestamp 1688980957
transform 1 0 48576 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_528
timestamp 1688980957
transform 1 0 49680 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_581
timestamp 1688980957
transform 1 0 54556 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_585
timestamp 1688980957
transform 1 0 54924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_598
timestamp 1688980957
transform 1 0 56120 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_619
timestamp 1688980957
transform 1 0 58052 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_253
timestamp 1688980957
transform 1 0 24380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_265
timestamp 1688980957
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1688980957
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1688980957
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_401
timestamp 1688980957
transform 1 0 37996 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_428
timestamp 1688980957
transform 1 0 40480 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_440
timestamp 1688980957
transform 1 0 41584 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 1688980957
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_461
timestamp 1688980957
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_473
timestamp 1688980957
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_485
timestamp 1688980957
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_497
timestamp 1688980957
transform 1 0 46828 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_501
timestamp 1688980957
transform 1 0 47196 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_529
timestamp 1688980957
transform 1 0 49772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_537
timestamp 1688980957
transform 1 0 50508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_554
timestamp 1688980957
transform 1 0 52072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_558
timestamp 1688980957
transform 1 0 52440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_561
timestamp 1688980957
transform 1 0 52716 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_571
timestamp 1688980957
transform 1 0 53636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_583
timestamp 1688980957
transform 1 0 54740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_593
timestamp 1688980957
transform 1 0 55660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_602
timestamp 1688980957
transform 1 0 56488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_606
timestamp 1688980957
transform 1 0 56856 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_614
timestamp 1688980957
transform 1 0 57592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_617
timestamp 1688980957
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1688980957
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1688980957
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_401
timestamp 1688980957
transform 1 0 37996 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_417
timestamp 1688980957
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_421
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_425
timestamp 1688980957
transform 1 0 40204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_437
timestamp 1688980957
transform 1 0 41308 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_449
timestamp 1688980957
transform 1 0 42412 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_461
timestamp 1688980957
transform 1 0 43516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_473
timestamp 1688980957
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_477
timestamp 1688980957
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_489
timestamp 1688980957
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_501
timestamp 1688980957
transform 1 0 47196 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_507
timestamp 1688980957
transform 1 0 47748 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_516
timestamp 1688980957
transform 1 0 48576 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_528
timestamp 1688980957
transform 1 0 49680 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_533
timestamp 1688980957
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_545
timestamp 1688980957
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_557
timestamp 1688980957
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_569
timestamp 1688980957
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_581
timestamp 1688980957
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 1688980957
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_589
timestamp 1688980957
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_601
timestamp 1688980957
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_613
timestamp 1688980957
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 1688980957
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 1688980957
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 1688980957
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 1688980957
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 1688980957
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 1688980957
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 1688980957
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 1688980957
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_485
timestamp 1688980957
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_497
timestamp 1688980957
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 1688980957
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_505
timestamp 1688980957
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_517
timestamp 1688980957
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_529
timestamp 1688980957
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_541
timestamp 1688980957
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_553
timestamp 1688980957
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_559
timestamp 1688980957
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 1688980957
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_573
timestamp 1688980957
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 1688980957
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 1688980957
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 1688980957
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 1688980957
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_617
timestamp 1688980957
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 1688980957
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 1688980957
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 1688980957
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 1688980957
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 1688980957
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 1688980957
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 1688980957
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 1688980957
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 1688980957
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 1688980957
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 1688980957
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 1688980957
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 1688980957
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 1688980957
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 1688980957
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 1688980957
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 1688980957
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 1688980957
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 1688980957
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 1688980957
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 1688980957
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_613
timestamp 1688980957
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 1688980957
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 1688980957
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_441
timestamp 1688980957
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 1688980957
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 1688980957
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 1688980957
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 1688980957
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 1688980957
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 1688980957
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 1688980957
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 1688980957
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 1688980957
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 1688980957
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 1688980957
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 1688980957
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 1688980957
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 1688980957
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 1688980957
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 1688980957
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 1688980957
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_617
timestamp 1688980957
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 1688980957
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 1688980957
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 1688980957
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 1688980957
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 1688980957
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 1688980957
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 1688980957
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 1688980957
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 1688980957
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 1688980957
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 1688980957
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 1688980957
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 1688980957
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 1688980957
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1688980957
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 1688980957
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 1688980957
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 1688980957
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 1688980957
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 1688980957
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 1688980957
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 1688980957
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 1688980957
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 1688980957
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 1688980957
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 1688980957
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 1688980957
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 1688980957
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 1688980957
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 1688980957
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 1688980957
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 1688980957
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 1688980957
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 1688980957
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 1688980957
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 1688980957
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 1688980957
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 1688980957
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 1688980957
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 1688980957
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 1688980957
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_617
timestamp 1688980957
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 1688980957
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 1688980957
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 1688980957
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 1688980957
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 1688980957
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 1688980957
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 1688980957
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 1688980957
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 1688980957
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 1688980957
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 1688980957
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 1688980957
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 1688980957
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 1688980957
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 1688980957
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 1688980957
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 1688980957
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 1688980957
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 1688980957
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1688980957
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1688980957
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 1688980957
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 1688980957
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 1688980957
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 1688980957
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 1688980957
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 1688980957
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 1688980957
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 1688980957
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 1688980957
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 1688980957
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 1688980957
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 1688980957
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 1688980957
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 1688980957
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 1688980957
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 1688980957
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 1688980957
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 1688980957
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 1688980957
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 1688980957
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 1688980957
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 1688980957
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_617
timestamp 1688980957
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_57
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 1688980957
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1688980957
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_281
timestamp 1688980957
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_293
timestamp 1688980957
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_337
timestamp 1688980957
transform 1 0 32108 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_349
timestamp 1688980957
transform 1 0 33212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_393
timestamp 1688980957
transform 1 0 37260 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_405
timestamp 1688980957
transform 1 0 38364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_417
timestamp 1688980957
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 1688980957
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_445
timestamp 1688980957
transform 1 0 42044 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_449
timestamp 1688980957
transform 1 0 42412 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_461
timestamp 1688980957
transform 1 0 43516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_473
timestamp 1688980957
transform 1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1688980957
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 1688980957
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_501
timestamp 1688980957
transform 1 0 47196 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_505
timestamp 1688980957
transform 1 0 47564 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_517
timestamp 1688980957
transform 1 0 48668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_529
timestamp 1688980957
transform 1 0 49772 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 1688980957
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 1688980957
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_557
timestamp 1688980957
transform 1 0 52348 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_561
timestamp 1688980957
transform 1 0 52716 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_573
timestamp 1688980957
transform 1 0 53820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_585
timestamp 1688980957
transform 1 0 54924 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1688980957
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1688980957
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_613
timestamp 1688980957
transform 1 0 57500 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_617
timestamp 1688980957
transform 1 0 57868 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 40388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 45540 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold5
timestamp 1688980957
transform 1 0 45816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 46920 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 41952 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 43976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 44160 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold12
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold15
timestamp 1688980957
transform 1 0 16744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 16468 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 39008 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 38272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold26
timestamp 1688980957
transform 1 0 25944 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 23276 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 14904 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 14168 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 35328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold33
timestamp 1688980957
transform 1 0 31096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 28520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 25392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 24656 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 40112 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 38732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 19320 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 17572 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 41400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 39192 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 40020 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 39192 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 29532 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 28244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 22356 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 29716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 16744 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 18216 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 27692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 26680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 25760 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 25208 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 23460 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold74
timestamp 1688980957
transform 1 0 54648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 53360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 38456 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 21528 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 22356 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 42412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 41952 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 26864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 44068 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 43332 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 30820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 30452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 33856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 57040 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 55476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 45816 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 44804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold101
timestamp 1688980957
transform 1 0 50140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 51704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 50784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform 1 0 50140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 54464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform 1 0 52072 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform 1 0 55568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform 1 0 56304 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 36156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold110
timestamp 1688980957
transform 1 0 33856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 53636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 52716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform 1 0 46276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 46552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform 1 0 46552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 46552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 47932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 50508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 49772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 54096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 54096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold125
timestamp 1688980957
transform 1 0 52256 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 50784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 48208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform 1 0 46736 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 22724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold130
timestamp 1688980957
transform 1 0 24748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 51520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 51612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform 1 0 49220 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 48668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 12512 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold137
timestamp 1688980957
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 43240 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 39928 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold142
timestamp 1688980957
transform 1 0 35696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 32936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 57040 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 33120 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 34592 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 26128 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 37352 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform 1 0 36432 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 33488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform 1 0 49404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 48852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform 1 0 47564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold157
timestamp 1688980957
transform 1 0 46644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform 1 0 45908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold160
timestamp 1688980957
transform 1 0 41584 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform 1 0 40020 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform 1 0 37352 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform 1 0 37352 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform 1 0 43516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 43516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold167
timestamp 1688980957
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform 1 0 9844 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform 1 0 35972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform 1 0 25852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 25576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform 1 0 29808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold176
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform 1 0 27968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform 1 0 36064 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform 1 0 35328 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform 1 0 6900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform 1 0 37444 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 25392 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform 1 0 25760 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform 1 0 23552 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 36064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform 1 0 49036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform 1 0 49312 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold193
timestamp 1688980957
transform 1 0 19044 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform 1 0 33304 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform 1 0 32568 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold198
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 12420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform 1 0 49036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 49772 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform 1 0 20056 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform 1 0 34040 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform 1 0 40112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform 1 0 39284 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform 1 0 23000 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform 1 0 37628 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform 1 0 35880 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 37352 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 26864 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform 1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 46736 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform 1 0 45264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform 1 0 12420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform 1 0 38088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform 1 0 37352 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform 1 0 57684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform 1 0 56120 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform 1 0 41400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform 1 0 14536 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform 1 0 34684 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform 1 0 32292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform 1 0 23368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform 1 0 22632 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform 1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform 1 0 43240 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform 1 0 43976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform 1 0 51704 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform 1 0 50876 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform 1 0 14168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform 1 0 14904 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform 1 0 14996 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform 1 0 54832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold245
timestamp 1688980957
transform 1 0 58236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform 1 0 55844 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform 1 0 49036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform 1 0 48116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform 1 0 27416 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform 1 0 46368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform 1 0 46000 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform 1 0 17480 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform 1 0 17940 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform 1 0 46644 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 45264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform 1 0 29624 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform 1 0 12972 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform 1 0 6348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform 1 0 53728 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform 1 0 53452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform 1 0 31464 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform 1 0 12328 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform 1 0 11592 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform 1 0 31188 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform 1 0 20792 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform 1 0 55752 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform 1 0 56120 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform 1 0 28244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform 1 0 54372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform 1 0 52900 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform 1 0 29900 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform 1 0 38456 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform 1 0 52716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform 1 0 51888 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform 1 0 7176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform 1 0 40664 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform 1 0 39008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform 1 0 9752 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform 1 0 54556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform 1 0 53636 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform 1 0 54464 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 56488 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform 1 0 57684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform 1 0 57868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform 1 0 5244 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold316
timestamp 1688980957
transform 1 0 34500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform 1 0 33212 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform 1 0 40664 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold319
timestamp 1688980957
transform 1 0 39652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform 1 0 40020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold322
timestamp 1688980957
transform 1 0 28980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform 1 0 27600 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform 1 0 31004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform 1 0 30176 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform 1 0 39008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform 1 0 38272 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform 1 0 33948 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold331
timestamp 1688980957
transform 1 0 19872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform 1 0 38272 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform 1 0 37536 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform 1 0 27876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform 1 0 48208 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform 1 0 49220 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform 1 0 35604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform 1 0 31004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform 1 0 7912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform 1 0 32936 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform 1 0 32016 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform 1 0 55476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform 1 0 54464 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1688980957
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform 1 0 55568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1688980957
transform 1 0 54740 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1688980957
transform 1 0 43056 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1688980957
transform 1 0 43884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 1688980957
transform 1 0 31004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1688980957
transform 1 0 30176 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold359
timestamp 1688980957
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1688980957
transform 1 0 17480 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold362
timestamp 1688980957
transform 1 0 43516 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1688980957
transform 1 0 42412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1688980957
transform 1 0 28336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold365
timestamp 1688980957
transform 1 0 27600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1688980957
transform 1 0 28888 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1688980957
transform 1 0 28152 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold369
timestamp 1688980957
transform 1 0 10764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1688980957
transform 1 0 11224 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1688980957
transform 1 0 28520 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1688980957
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold375
timestamp 1688980957
transform 1 0 20056 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold376
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold377
timestamp 1688980957
transform 1 0 38640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 1688980957
transform 1 0 37904 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 1688980957
transform 1 0 39652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 1688980957
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold382
timestamp 1688980957
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold383
timestamp 1688980957
transform 1 0 44988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 1688980957
transform 1 0 44988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 1688980957
transform 1 0 50508 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold386
timestamp 1688980957
transform 1 0 49312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 1688980957
transform 1 0 46276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold388
timestamp 1688980957
transform 1 0 8648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold389
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 1688980957
transform 1 0 39744 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold391
timestamp 1688980957
transform 1 0 38732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold392
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold393
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold394
timestamp 1688980957
transform 1 0 15640 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold395
timestamp 1688980957
transform 1 0 36248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold396
timestamp 1688980957
transform 1 0 35512 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold397
timestamp 1688980957
transform 1 0 45172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold398
timestamp 1688980957
transform 1 0 44988 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold399
timestamp 1688980957
transform 1 0 38180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold400
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold401
timestamp 1688980957
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold402
timestamp 1688980957
transform 1 0 17848 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold403
timestamp 1688980957
transform 1 0 51888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold404
timestamp 1688980957
transform 1 0 53084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold405
timestamp 1688980957
transform 1 0 53084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold406
timestamp 1688980957
transform 1 0 51336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold407
timestamp 1688980957
transform 1 0 50600 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold408
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold409
timestamp 1688980957
transform 1 0 41492 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold410
timestamp 1688980957
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold411
timestamp 1688980957
transform 1 0 27324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold412
timestamp 1688980957
transform 1 0 24932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold413
timestamp 1688980957
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold414
timestamp 1688980957
transform 1 0 11592 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold415
timestamp 1688980957
transform 1 0 13800 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold416
timestamp 1688980957
transform 1 0 12788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold417
timestamp 1688980957
transform 1 0 9200 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold418
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold419
timestamp 1688980957
transform 1 0 23828 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold420
timestamp 1688980957
transform 1 0 23092 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold421
timestamp 1688980957
transform 1 0 12328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold422
timestamp 1688980957
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold423
timestamp 1688980957
transform 1 0 39560 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold424
timestamp 1688980957
transform 1 0 40388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold425
timestamp 1688980957
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold426
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold427
timestamp 1688980957
transform 1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold428
timestamp 1688980957
transform 1 0 32752 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold429
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold430
timestamp 1688980957
transform 1 0 7636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold431
timestamp 1688980957
transform 1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold432
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold433
timestamp 1688980957
transform 1 0 2208 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold434
timestamp 1688980957
transform 1 0 52716 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold435
timestamp 1688980957
transform 1 0 52808 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold436
timestamp 1688980957
transform 1 0 23460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold437
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold438
timestamp 1688980957
transform 1 0 33672 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold439
timestamp 1688980957
transform 1 0 33764 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold440
timestamp 1688980957
transform 1 0 6256 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold441
timestamp 1688980957
transform 1 0 6624 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold442
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold443
timestamp 1688980957
transform 1 0 4140 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold444
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold445
timestamp 1688980957
transform 1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold446
timestamp 1688980957
transform 1 0 27140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold447
timestamp 1688980957
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold448
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold449
timestamp 1688980957
transform 1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold450
timestamp 1688980957
transform 1 0 49036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold451
timestamp 1688980957
transform 1 0 47840 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold452
timestamp 1688980957
transform 1 0 53636 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold453
timestamp 1688980957
transform 1 0 52900 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold454
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold455
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold456
timestamp 1688980957
transform 1 0 18676 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold457
timestamp 1688980957
transform 1 0 17296 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold458
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold459
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold460
timestamp 1688980957
transform 1 0 47564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold461
timestamp 1688980957
transform 1 0 46552 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold462
timestamp 1688980957
transform 1 0 52440 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold463
timestamp 1688980957
transform 1 0 51704 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold464
timestamp 1688980957
transform 1 0 52348 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold465
timestamp 1688980957
transform 1 0 51336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold466
timestamp 1688980957
transform 1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold467
timestamp 1688980957
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold468
timestamp 1688980957
transform 1 0 51520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold469
timestamp 1688980957
transform 1 0 50600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold470
timestamp 1688980957
transform 1 0 42596 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold471
timestamp 1688980957
transform 1 0 41676 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold472
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold473
timestamp 1688980957
transform 1 0 21988 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold474
timestamp 1688980957
transform 1 0 36064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold475
timestamp 1688980957
transform 1 0 35972 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold476
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold477
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold478
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold479
timestamp 1688980957
transform 1 0 19872 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold480
timestamp 1688980957
transform 1 0 53544 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold481
timestamp 1688980957
transform 1 0 53176 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold482
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold483
timestamp 1688980957
transform 1 0 41308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold484
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold485
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold486
timestamp 1688980957
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold487
timestamp 1688980957
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold488
timestamp 1688980957
transform 1 0 9108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold489
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold490
timestamp 1688980957
transform 1 0 50508 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold491
timestamp 1688980957
transform 1 0 49772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold492
timestamp 1688980957
transform 1 0 45448 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold493
timestamp 1688980957
transform 1 0 44804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold494
timestamp 1688980957
transform 1 0 48300 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold495
timestamp 1688980957
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold496
timestamp 1688980957
transform 1 0 25852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold497
timestamp 1688980957
transform 1 0 24748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold498
timestamp 1688980957
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold499
timestamp 1688980957
transform 1 0 47380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold500
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold501
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold502
timestamp 1688980957
transform 1 0 50324 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold503
timestamp 1688980957
transform 1 0 49036 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold504
timestamp 1688980957
transform 1 0 6440 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold505
timestamp 1688980957
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold506
timestamp 1688980957
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold507
timestamp 1688980957
transform 1 0 22356 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold508
timestamp 1688980957
transform 1 0 12328 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold509
timestamp 1688980957
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold510
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold511
timestamp 1688980957
transform 1 0 6716 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold512
timestamp 1688980957
transform 1 0 51888 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold513
timestamp 1688980957
transform 1 0 58236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold514
timestamp 1688980957
transform 1 0 54924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold515
timestamp 1688980957
transform 1 0 13984 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold516
timestamp 1688980957
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold517
timestamp 1688980957
transform 1 0 45724 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold518
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold519
timestamp 1688980957
transform 1 0 50968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold520
timestamp 1688980957
transform 1 0 50508 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold521
timestamp 1688980957
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold522
timestamp 1688980957
transform 1 0 2116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold523
timestamp 1688980957
transform 1 0 9752 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold524
timestamp 1688980957
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold525
timestamp 1688980957
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold526
timestamp 1688980957
transform 1 0 56396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold527
timestamp 1688980957
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold528
timestamp 1688980957
transform 1 0 57316 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold529
timestamp 1688980957
transform 1 0 55292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold530
timestamp 1688980957
transform 1 0 55108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold531
timestamp 1688980957
transform 1 0 13800 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold532
timestamp 1688980957
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold533
timestamp 1688980957
transform 1 0 23920 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold534
timestamp 1688980957
transform 1 0 23184 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold535
timestamp 1688980957
transform 1 0 3864 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold536
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold537
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold538
timestamp 1688980957
transform 1 0 53912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold539
timestamp 1688980957
transform 1 0 55476 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold540
timestamp 1688980957
transform 1 0 54372 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold541
timestamp 1688980957
transform 1 0 57040 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold542
timestamp 1688980957
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold543
timestamp 1688980957
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold544
timestamp 1688980957
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold545
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold546
timestamp 1688980957
transform 1 0 2208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold547
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold548
timestamp 1688980957
transform 1 0 2668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold549
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold550
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold551
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold552
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold553
timestamp 1688980957
transform 1 0 2668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold554 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold555
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold556
timestamp 1688980957
transform 1 0 2116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold557
timestamp 1688980957
transform 1 0 3864 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold558
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold559
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold560
timestamp 1688980957
transform 1 0 50968 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold561
timestamp 1688980957
transform 1 0 40756 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold562
timestamp 1688980957
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold563
timestamp 1688980957
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold564
timestamp 1688980957
transform 1 0 53820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold565
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold566
timestamp 1688980957
transform 1 0 51796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold567
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold568
timestamp 1688980957
transform 1 0 41124 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold569
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold570
timestamp 1688980957
transform 1 0 55752 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold571
timestamp 1688980957
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold572
timestamp 1688980957
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold573
timestamp 1688980957
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold574
timestamp 1688980957
transform 1 0 23184 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold575
timestamp 1688980957
transform 1 0 21528 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold576
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold577
timestamp 1688980957
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold578
timestamp 1688980957
transform 1 0 54096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold579
timestamp 1688980957
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold580
timestamp 1688980957
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold581
timestamp 1688980957
transform 1 0 45448 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold582
timestamp 1688980957
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold583
timestamp 1688980957
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold584
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold585
timestamp 1688980957
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold586
timestamp 1688980957
transform 1 0 29532 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold587
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold588
timestamp 1688980957
transform 1 0 42320 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold589
timestamp 1688980957
transform 1 0 40756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold590
timestamp 1688980957
transform 1 0 47656 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 28060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 38916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 40664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 43608 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 48760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 51244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 54188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 53820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 57500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 18952 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 26680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 28980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 29072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 32200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 38088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 43332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 44160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 44528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 47656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 50232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 52256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 55384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 54924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 54924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 58236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 58236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output69 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform 1 0 4784 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform 1 0 24196 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform 1 0 30544 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform 1 0 32476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform 1 0 40756 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform 1 0 44068 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform 1 0 45724 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform 1 0 47564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform 1 0 49036 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform 1 0 50692 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1688980957
transform 1 0 52716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1688980957
transform 1 0 54004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1688980957
transform 1 0 55660 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1688980957
transform 1 0 56304 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1688980957
transform 1 0 57132 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1688980957
transform 1 0 14720 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform 1 0 19228 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 32016 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 37168 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 42320 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 47472 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 52624 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 57776 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire118
timestamp 1688980957
transform 1 0 33212 0 1 4352
box -38 -48 406 592
<< labels >>
flabel metal4 s 8166 2128 8486 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 22610 2128 22930 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 37054 2128 37374 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 51498 2128 51818 27792 0 FreeSans 1920 90 0 0 vccd1
port 0 nsew power bidirectional
flabel metal4 s 15388 2128 15708 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 29832 2128 30152 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 44276 2128 44596 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal4 s 58720 2128 59040 27792 0 FreeSans 1920 90 0 0 vssd1
port 1 nsew ground bidirectional
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 5 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 6 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 7 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 8 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 9 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 10 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 11 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 12 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 13 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 14 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 15 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 16 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 17 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 18 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 19 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 20 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 21 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 22 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 23 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 24 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 25 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 26 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 27 nsew signal input
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 28 nsew signal input
flabel metal2 s 57794 0 57850 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 29 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 30 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 31 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 32 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 33 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 34 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 35 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 36 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 37 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 38 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 40 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 41 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 42 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 43 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 44 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 45 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 46 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 47 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 48 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 49 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 50 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 51 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 52 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 53 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 54 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 55 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 56 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 57 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 58 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 59 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 60 nsew signal input
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 61 nsew signal input
flabel metal2 s 58346 0 58402 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 62 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 63 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 64 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 65 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 66 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 67 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 68 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 69 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 70 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 71 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 72 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 73 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 74 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 75 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 76 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 77 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 78 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 79 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 80 nsew signal tristate
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 81 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 82 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 83 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 84 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 85 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 86 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 87 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 88 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 89 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 90 nsew signal tristate
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 91 nsew signal tristate
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 92 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 93 nsew signal tristate
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 94 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 95 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 96 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 97 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 98 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 99 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 100 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 101 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 102 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 103 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 104 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 105 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 106 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 wbs_we_i
port 107 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 30000
<< end >>
