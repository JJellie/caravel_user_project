magic
tech sky130A
magscale 1 2
timestamp 1728393570
<< viali >>
rect 38117 34969 38151 35003
rect 38209 34901 38243 34935
rect 38117 25177 38151 25211
rect 38209 25109 38243 25143
rect 14197 15997 14231 16031
rect 14749 15861 14783 15895
rect 11805 15453 11839 15487
rect 14565 15453 14599 15487
rect 38209 15453 38243 15487
rect 12449 15317 12483 15351
rect 15117 15317 15151 15351
rect 38393 15317 38427 15351
rect 14565 15113 14599 15147
rect 14933 15113 14967 15147
rect 15025 15113 15059 15147
rect 15577 15113 15611 15147
rect 11529 14977 11563 15011
rect 11796 14977 11830 15011
rect 13093 14977 13127 15011
rect 13360 14977 13394 15011
rect 8125 14909 8159 14943
rect 8861 14909 8895 14943
rect 10333 14909 10367 14943
rect 15117 14909 15151 14943
rect 16681 14909 16715 14943
rect 8677 14773 8711 14807
rect 9413 14773 9447 14807
rect 10885 14773 10919 14807
rect 12909 14773 12943 14807
rect 14473 14773 14507 14807
rect 17325 14773 17359 14807
rect 17601 14773 17635 14807
rect 8769 14569 8803 14603
rect 11805 14569 11839 14603
rect 16773 14501 16807 14535
rect 11345 14433 11379 14467
rect 12357 14433 12391 14467
rect 12725 14433 12759 14467
rect 14749 14433 14783 14467
rect 17417 14433 17451 14467
rect 7389 14365 7423 14399
rect 9229 14365 9263 14399
rect 11069 14365 11103 14399
rect 17141 14365 17175 14399
rect 17693 14365 17727 14399
rect 18521 14365 18555 14399
rect 19349 14365 19383 14399
rect 7656 14297 7690 14331
rect 9496 14297 9530 14331
rect 12173 14297 12207 14331
rect 13277 14297 13311 14331
rect 15016 14297 15050 14331
rect 10609 14229 10643 14263
rect 10701 14229 10735 14263
rect 11161 14229 11195 14263
rect 12265 14229 12299 14263
rect 13553 14229 13587 14263
rect 16129 14229 16163 14263
rect 16497 14229 16531 14263
rect 17233 14229 17267 14263
rect 18245 14229 18279 14263
rect 19073 14229 19107 14263
rect 19993 14229 20027 14263
rect 8309 14025 8343 14059
rect 8677 14025 8711 14059
rect 11253 14025 11287 14059
rect 17325 14025 17359 14059
rect 17693 14025 17727 14059
rect 18061 14025 18095 14059
rect 19340 13957 19374 13991
rect 8769 13889 8803 13923
rect 10701 13889 10735 13923
rect 16773 13889 16807 13923
rect 18153 13889 18187 13923
rect 19073 13889 19107 13923
rect 8953 13821 8987 13855
rect 9413 13821 9447 13855
rect 11713 13821 11747 13855
rect 12173 13821 12207 13855
rect 14197 13821 14231 13855
rect 14565 13821 14599 13855
rect 14933 13821 14967 13855
rect 15301 13821 15335 13855
rect 15669 13821 15703 13855
rect 16037 13821 16071 13855
rect 16405 13821 16439 13855
rect 18245 13821 18279 13855
rect 18797 13821 18831 13855
rect 20545 13821 20579 13855
rect 12725 13685 12759 13719
rect 13093 13685 13127 13719
rect 13461 13685 13495 13719
rect 13829 13685 13863 13719
rect 20453 13685 20487 13719
rect 21189 13685 21223 13719
rect 8769 13481 8803 13515
rect 16773 13481 16807 13515
rect 18613 13481 18647 13515
rect 19349 13481 19383 13515
rect 20453 13481 20487 13515
rect 11989 13413 12023 13447
rect 15669 13413 15703 13447
rect 10609 13345 10643 13379
rect 12081 13345 12115 13379
rect 12725 13345 12759 13379
rect 13118 13345 13152 13379
rect 14289 13345 14323 13379
rect 16405 13345 16439 13379
rect 19901 13345 19935 13379
rect 9229 13277 9263 13311
rect 12265 13277 12299 13311
rect 13001 13277 13035 13311
rect 13277 13277 13311 13311
rect 17233 13277 17267 13311
rect 19717 13277 19751 13311
rect 10876 13209 10910 13243
rect 14556 13209 14590 13243
rect 17500 13209 17534 13243
rect 19809 13209 19843 13243
rect 9781 13141 9815 13175
rect 13921 13141 13955 13175
rect 15761 13141 15795 13175
rect 16129 13141 16163 13175
rect 16221 13141 16255 13175
rect 8769 12937 8803 12971
rect 12081 12937 12115 12971
rect 13737 12937 13771 12971
rect 15853 12937 15887 12971
rect 17325 12937 17359 12971
rect 7389 12801 7423 12835
rect 7656 12801 7690 12835
rect 9965 12801 9999 12835
rect 10082 12801 10116 12835
rect 10241 12801 10275 12835
rect 11989 12801 12023 12835
rect 13645 12801 13679 12835
rect 15301 12801 15335 12835
rect 18429 12801 18463 12835
rect 9045 12733 9079 12767
rect 9229 12733 9263 12767
rect 12173 12733 12207 12767
rect 13829 12733 13863 12767
rect 16681 12733 16715 12767
rect 18613 12733 18647 12767
rect 19349 12733 19383 12767
rect 19466 12733 19500 12767
rect 19625 12733 19659 12767
rect 9689 12665 9723 12699
rect 11345 12665 11379 12699
rect 19073 12665 19107 12699
rect 10885 12597 10919 12631
rect 11621 12597 11655 12631
rect 12725 12597 12759 12631
rect 13093 12597 13127 12631
rect 13277 12597 13311 12631
rect 18245 12597 18279 12631
rect 20269 12597 20303 12631
rect 8769 12393 8803 12427
rect 11161 12393 11195 12427
rect 11897 12393 11931 12427
rect 17049 12393 17083 12427
rect 8953 12325 8987 12359
rect 12725 12325 12759 12359
rect 13093 12325 13127 12359
rect 13461 12325 13495 12359
rect 15117 12325 15151 12359
rect 15853 12325 15887 12359
rect 8217 12257 8251 12291
rect 9505 12257 9539 12291
rect 10609 12257 10643 12291
rect 11345 12257 11379 12291
rect 15209 12257 15243 12291
rect 16129 12257 16163 12291
rect 16405 12257 16439 12291
rect 20729 12257 20763 12291
rect 9413 12189 9447 12223
rect 10425 12189 10459 12223
rect 10517 12189 10551 12223
rect 15393 12189 15427 12223
rect 16246 12189 16280 12223
rect 19993 12189 20027 12223
rect 9321 12121 9355 12155
rect 10057 12053 10091 12087
rect 20637 12053 20671 12087
rect 21373 12053 21407 12087
rect 4629 11849 4663 11883
rect 3801 11781 3835 11815
rect 19892 11781 19926 11815
rect 4077 11713 4111 11747
rect 4261 11713 4295 11747
rect 4445 11713 4479 11747
rect 4721 11713 4755 11747
rect 4353 11645 4387 11679
rect 9137 11645 9171 11679
rect 10149 11645 10183 11679
rect 11897 11645 11931 11679
rect 12909 11645 12943 11679
rect 14841 11645 14875 11679
rect 15669 11645 15703 11679
rect 17509 11645 17543 11679
rect 19625 11645 19659 11679
rect 4445 11577 4479 11611
rect 3893 11509 3927 11543
rect 5089 11509 5123 11543
rect 9689 11509 9723 11543
rect 10701 11509 10735 11543
rect 12541 11509 12575 11543
rect 13553 11509 13587 11543
rect 15485 11509 15519 11543
rect 16221 11509 16255 11543
rect 18153 11509 18187 11543
rect 21005 11509 21039 11543
rect 5273 11305 5307 11339
rect 6929 11305 6963 11339
rect 12357 11305 12391 11339
rect 13921 11305 13955 11339
rect 14473 11305 14507 11339
rect 16681 11305 16715 11339
rect 18613 11305 18647 11339
rect 19993 11305 20027 11339
rect 10057 11237 10091 11271
rect 14289 11237 14323 11271
rect 4169 11169 4203 11203
rect 9413 11169 9447 11203
rect 9505 11169 9539 11203
rect 15117 11169 15151 11203
rect 20453 11169 20487 11203
rect 20637 11169 20671 11203
rect 4905 11101 4939 11135
rect 4997 11101 5031 11135
rect 5365 11101 5399 11135
rect 5549 11101 5583 11135
rect 7297 11101 7331 11135
rect 9321 11101 9355 11135
rect 10241 11101 10275 11135
rect 10977 11101 11011 11135
rect 12541 11101 12575 11135
rect 15301 11101 15335 11135
rect 17233 11101 17267 11135
rect 20361 11101 20395 11135
rect 21005 11101 21039 11135
rect 5816 11033 5850 11067
rect 7564 11033 7598 11067
rect 11244 11033 11278 11067
rect 12808 11033 12842 11067
rect 14841 11033 14875 11067
rect 15568 11033 15602 11067
rect 16957 11033 16991 11067
rect 17500 11033 17534 11067
rect 4813 10965 4847 10999
rect 5089 10965 5123 10999
rect 5365 10965 5399 10999
rect 8677 10965 8711 10999
rect 8953 10965 8987 10999
rect 10885 10965 10919 10999
rect 14933 10965 14967 10999
rect 6193 10761 6227 10795
rect 8953 10761 8987 10795
rect 10609 10761 10643 10795
rect 10977 10761 11011 10795
rect 11529 10761 11563 10795
rect 16221 10761 16255 10795
rect 17509 10761 17543 10795
rect 9404 10693 9438 10727
rect 12541 10693 12575 10727
rect 15108 10693 15142 10727
rect 17877 10693 17911 10727
rect 17969 10693 18003 10727
rect 18981 10693 19015 10727
rect 2881 10625 2915 10659
rect 5181 10625 5215 10659
rect 5365 10625 5399 10659
rect 5457 10625 5491 10659
rect 5641 10625 5675 10659
rect 6653 10625 6687 10659
rect 8401 10625 8435 10659
rect 11897 10625 11931 10659
rect 13001 10625 13035 10659
rect 14749 10625 14783 10659
rect 14841 10625 14875 10659
rect 16681 10625 16715 10659
rect 18429 10625 18463 10659
rect 3157 10557 3191 10591
rect 6377 10557 6411 10591
rect 9137 10557 9171 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 11989 10557 12023 10591
rect 12173 10557 12207 10591
rect 18061 10557 18095 10591
rect 20545 10557 20579 10591
rect 4445 10489 4479 10523
rect 4905 10489 4939 10523
rect 5181 10421 5215 10455
rect 10517 10421 10551 10455
rect 17325 10421 17359 10455
rect 21189 10421 21223 10455
rect 21557 10421 21591 10455
rect 4445 10217 4479 10251
rect 4905 10217 4939 10251
rect 6561 10217 6595 10251
rect 9321 10217 9355 10251
rect 12173 10217 12207 10251
rect 12909 10217 12943 10251
rect 18521 10217 18555 10251
rect 20545 10217 20579 10251
rect 12817 10149 12851 10183
rect 11621 10081 11655 10115
rect 13553 10081 13587 10115
rect 14105 10081 14139 10115
rect 16221 10081 16255 10115
rect 16313 10081 16347 10115
rect 19901 10081 19935 10115
rect 21097 10081 21131 10115
rect 4537 10013 4571 10047
rect 7205 10013 7239 10047
rect 9505 10013 9539 10047
rect 13277 10013 13311 10047
rect 14841 10013 14875 10047
rect 16129 10013 16163 10047
rect 16773 10013 16807 10047
rect 17693 10013 17727 10047
rect 19717 10013 19751 10047
rect 20361 10013 20395 10047
rect 20913 10013 20947 10047
rect 21373 10013 21407 10047
rect 4905 9945 4939 9979
rect 5273 9945 5307 9979
rect 19625 9945 19659 9979
rect 5089 9877 5123 9911
rect 7757 9877 7791 9911
rect 10057 9877 10091 9911
rect 11345 9877 11379 9911
rect 13369 9877 13403 9911
rect 14749 9877 14783 9911
rect 15485 9877 15519 9911
rect 15761 9877 15795 9911
rect 17417 9877 17451 9911
rect 18245 9877 18279 9911
rect 19257 9877 19291 9911
rect 21005 9877 21039 9911
rect 22017 9877 22051 9911
rect 5457 9673 5491 9707
rect 7757 9673 7791 9707
rect 16773 9673 16807 9707
rect 20177 9673 20211 9707
rect 21649 9673 21683 9707
rect 13277 9605 13311 9639
rect 16313 9605 16347 9639
rect 20536 9605 20570 9639
rect 5549 9537 5583 9571
rect 6377 9537 6411 9571
rect 6633 9537 6667 9571
rect 7941 9537 7975 9571
rect 8208 9537 8242 9571
rect 9413 9537 9447 9571
rect 10333 9537 10367 9571
rect 11529 9537 11563 9571
rect 13369 9537 13403 9571
rect 13636 9537 13670 9571
rect 15761 9537 15795 9571
rect 17141 9537 17175 9571
rect 20269 9537 20303 9571
rect 3709 9469 3743 9503
rect 4905 9469 4939 9503
rect 6193 9469 6227 9503
rect 9597 9469 9631 9503
rect 10450 9469 10484 9503
rect 10609 9469 10643 9503
rect 15025 9469 15059 9503
rect 17233 9469 17267 9503
rect 17417 9469 17451 9503
rect 17601 9469 17635 9503
rect 17785 9469 17819 9503
rect 18521 9469 18555 9503
rect 18638 9469 18672 9503
rect 18797 9469 18831 9503
rect 19533 9469 19567 9503
rect 9321 9401 9355 9435
rect 10057 9401 10091 9435
rect 18245 9401 18279 9435
rect 4261 9333 4295 9367
rect 11253 9333 11287 9367
rect 14749 9333 14783 9367
rect 15577 9333 15611 9367
rect 19441 9333 19475 9367
rect 5641 9129 5675 9163
rect 8769 9129 8803 9163
rect 12817 9129 12851 9163
rect 16129 9129 16163 9163
rect 17877 9129 17911 9163
rect 20637 9129 20671 9163
rect 8953 9061 8987 9095
rect 6101 8993 6135 9027
rect 8217 8993 8251 9027
rect 9505 8993 9539 9027
rect 11989 8993 12023 9027
rect 12081 8993 12115 9027
rect 13369 8993 13403 9027
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 4905 8925 4939 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 9413 8925 9447 8959
rect 14749 8925 14783 8959
rect 16497 8925 16531 8959
rect 16764 8925 16798 8959
rect 19257 8925 19291 8959
rect 3985 8857 4019 8891
rect 9321 8857 9355 8891
rect 10057 8857 10091 8891
rect 13185 8857 13219 8891
rect 15016 8857 15050 8891
rect 19524 8857 19558 8891
rect 3899 8789 3933 8823
rect 4813 8789 4847 8823
rect 5549 8789 5583 8823
rect 6561 8789 6595 8823
rect 11529 8789 11563 8823
rect 11897 8789 11931 8823
rect 13277 8789 13311 8823
rect 13921 8789 13955 8823
rect 18245 8789 18279 8823
rect 4169 8585 4203 8619
rect 4997 8585 5031 8619
rect 5181 8585 5215 8619
rect 5733 8585 5767 8619
rect 13921 8585 13955 8619
rect 15117 8585 15151 8619
rect 15485 8585 15519 8619
rect 16221 8585 16255 8619
rect 17693 8585 17727 8619
rect 20085 8585 20119 8619
rect 3056 8517 3090 8551
rect 4261 8517 4295 8551
rect 4445 8449 4479 8483
rect 4813 8449 4847 8483
rect 4905 8449 4939 8483
rect 5365 8449 5399 8483
rect 5641 8449 5675 8483
rect 13369 8449 13403 8483
rect 15577 8449 15611 8483
rect 17325 8449 17359 8483
rect 19441 8449 19475 8483
rect 2789 8381 2823 8415
rect 4721 8381 4755 8415
rect 5181 8381 5215 8415
rect 8125 8381 8159 8415
rect 8861 8381 8895 8415
rect 11621 8381 11655 8415
rect 12265 8381 12299 8415
rect 15669 8381 15703 8415
rect 16773 8381 16807 8415
rect 20269 8381 20303 8415
rect 4629 8313 4663 8347
rect 5549 8313 5583 8347
rect 8677 8245 8711 8279
rect 9413 8245 9447 8279
rect 12173 8245 12207 8279
rect 12909 8245 12943 8279
rect 20913 8245 20947 8279
rect 5089 8041 5123 8075
rect 5641 8041 5675 8075
rect 12541 8041 12575 8075
rect 15209 8041 15243 8075
rect 18797 8041 18831 8075
rect 4721 7973 4755 8007
rect 8769 7973 8803 8007
rect 13093 7973 13127 8007
rect 4997 7905 5031 7939
rect 9413 7905 9447 7939
rect 9873 7905 9907 7939
rect 10266 7905 10300 7939
rect 10425 7905 10459 7939
rect 16037 7905 16071 7939
rect 2697 7837 2731 7871
rect 4813 7837 4847 7871
rect 5089 7837 5123 7871
rect 7389 7837 7423 7871
rect 7656 7837 7690 7871
rect 9229 7837 9263 7871
rect 10149 7837 10183 7871
rect 11161 7837 11195 7871
rect 11428 7837 11462 7871
rect 13001 7837 13035 7871
rect 13185 7837 13219 7871
rect 13461 7837 13495 7871
rect 14933 7837 14967 7871
rect 15025 7837 15059 7871
rect 15301 7837 15335 7871
rect 15669 7837 15703 7871
rect 15853 7837 15887 7871
rect 17141 7837 17175 7871
rect 17969 7837 18003 7871
rect 19901 7837 19935 7871
rect 20168 7837 20202 7871
rect 21373 7837 21407 7871
rect 3893 7769 3927 7803
rect 3249 7701 3283 7735
rect 3985 7701 4019 7735
rect 5273 7701 5307 7735
rect 11069 7701 11103 7735
rect 17693 7701 17727 7735
rect 18521 7701 18555 7735
rect 21281 7701 21315 7735
rect 22017 7701 22051 7735
rect 3255 7497 3289 7531
rect 3341 7497 3375 7531
rect 4997 7497 5031 7531
rect 8309 7497 8343 7531
rect 8769 7497 8803 7531
rect 10701 7497 10735 7531
rect 11529 7497 11563 7531
rect 11989 7497 12023 7531
rect 18061 7497 18095 7531
rect 20269 7497 20303 7531
rect 20729 7497 20763 7531
rect 8217 7429 8251 7463
rect 10609 7429 10643 7463
rect 16948 7429 16982 7463
rect 1952 7361 1986 7395
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 4629 7361 4663 7395
rect 4783 7361 4817 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 6644 7361 6678 7395
rect 8677 7361 8711 7395
rect 9321 7361 9355 7395
rect 11897 7361 11931 7395
rect 12449 7361 12483 7395
rect 12725 7361 12759 7395
rect 13093 7361 13127 7395
rect 15025 7361 15059 7395
rect 15209 7361 15243 7395
rect 18337 7361 18371 7395
rect 19190 7361 19224 7395
rect 19349 7361 19383 7395
rect 20637 7361 20671 7395
rect 21281 7361 21315 7395
rect 1685 7293 1719 7327
rect 8953 7293 8987 7327
rect 10793 7293 10827 7327
rect 12173 7293 12207 7327
rect 16681 7293 16715 7327
rect 18153 7293 18187 7327
rect 19073 7293 19107 7327
rect 20821 7293 20855 7327
rect 3065 7225 3099 7259
rect 18797 7225 18831 7259
rect 6193 7157 6227 7191
rect 7757 7157 7791 7191
rect 9873 7157 9907 7191
rect 10241 7157 10275 7191
rect 11253 7157 11287 7191
rect 12541 7157 12575 7191
rect 15025 7157 15059 7191
rect 19993 7157 20027 7191
rect 2881 6953 2915 6987
rect 7297 6953 7331 6987
rect 17141 6953 17175 6987
rect 2605 6885 2639 6919
rect 5365 6817 5399 6851
rect 5641 6817 5675 6851
rect 9689 6817 9723 6851
rect 9781 6817 9815 6851
rect 10057 6817 10091 6851
rect 17693 6817 17727 6851
rect 18245 6817 18279 6851
rect 18521 6817 18555 6851
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 5273 6749 5307 6783
rect 5457 6749 5491 6783
rect 6653 6749 6687 6783
rect 8217 6749 8251 6783
rect 9597 6749 9631 6783
rect 10793 6749 10827 6783
rect 14381 6749 14415 6783
rect 14657 6749 14691 6783
rect 15117 6749 15151 6783
rect 15669 6749 15703 6783
rect 15853 6749 15887 6783
rect 16129 6749 16163 6783
rect 16681 6749 16715 6783
rect 17601 6749 17635 6783
rect 18061 6749 18095 6783
rect 19441 6749 19475 6783
rect 16405 6681 16439 6715
rect 6285 6613 6319 6647
rect 8769 6613 8803 6647
rect 9229 6613 9263 6647
rect 10701 6613 10735 6647
rect 11437 6613 11471 6647
rect 12449 6613 12483 6647
rect 14197 6613 14231 6647
rect 17049 6613 17083 6647
rect 17509 6613 17543 6647
rect 19073 6613 19107 6647
rect 20085 6613 20119 6647
rect 9137 6409 9171 6443
rect 10057 6409 10091 6443
rect 10425 6409 10459 6443
rect 12081 6409 12115 6443
rect 17693 6409 17727 6443
rect 18061 6409 18095 6443
rect 20453 6409 20487 6443
rect 5733 6341 5767 6375
rect 8024 6341 8058 6375
rect 9781 6341 9815 6375
rect 10517 6341 10551 6375
rect 11161 6341 11195 6375
rect 11805 6341 11839 6375
rect 18153 6341 18187 6375
rect 19340 6341 19374 6375
rect 5641 6273 5675 6307
rect 5917 6273 5951 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7757 6273 7791 6307
rect 11989 6273 12023 6307
rect 12265 6273 12299 6307
rect 12731 6273 12765 6307
rect 12909 6273 12943 6307
rect 14933 6273 14967 6307
rect 17049 6273 17083 6307
rect 18797 6273 18831 6307
rect 20545 6273 20579 6307
rect 6009 6205 6043 6239
rect 6101 6205 6135 6239
rect 10701 6205 10735 6239
rect 12449 6205 12483 6239
rect 15117 6205 15151 6239
rect 15209 6205 15243 6239
rect 15301 6205 15335 6239
rect 15393 6205 15427 6239
rect 18245 6205 18279 6239
rect 19073 6205 19107 6239
rect 6377 6069 6411 6103
rect 12817 6069 12851 6103
rect 17601 6069 17635 6103
rect 21189 6069 21223 6103
rect 5181 5865 5215 5899
rect 6745 5865 6779 5899
rect 10885 5865 10919 5899
rect 15577 5865 15611 5899
rect 18889 5865 18923 5899
rect 19441 5865 19475 5899
rect 13645 5797 13679 5831
rect 20453 5797 20487 5831
rect 2605 5729 2639 5763
rect 7113 5729 7147 5763
rect 19901 5729 19935 5763
rect 20085 5729 20119 5763
rect 2697 5661 2731 5695
rect 3801 5661 3835 5695
rect 4629 5661 4663 5695
rect 5273 5661 5307 5695
rect 7297 5661 7331 5695
rect 9505 5661 9539 5695
rect 11713 5661 11747 5695
rect 11897 5661 11931 5695
rect 12449 5661 12483 5695
rect 12725 5661 12759 5695
rect 13093 5661 13127 5695
rect 13461 5661 13495 5695
rect 14197 5661 14231 5695
rect 15669 5661 15703 5695
rect 17509 5661 17543 5695
rect 17765 5661 17799 5695
rect 19809 5661 19843 5695
rect 38209 5661 38243 5695
rect 9772 5593 9806 5627
rect 14464 5593 14498 5627
rect 3065 5525 3099 5559
rect 4445 5525 4479 5559
rect 7481 5525 7515 5559
rect 11805 5525 11839 5559
rect 16957 5525 16991 5559
rect 38393 5525 38427 5559
rect 2789 5321 2823 5355
rect 3341 5321 3375 5355
rect 4261 5321 4295 5355
rect 14565 5321 14599 5355
rect 15393 5321 15427 5355
rect 3249 5253 3283 5287
rect 6561 5253 6595 5287
rect 16497 5253 16531 5287
rect 1409 5185 1443 5219
rect 1676 5185 1710 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 4445 5185 4479 5219
rect 4629 5185 4663 5219
rect 5365 5185 5399 5219
rect 6377 5185 6411 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 14381 5185 14415 5219
rect 15577 5185 15611 5219
rect 15761 5185 15795 5219
rect 16681 5185 16715 5219
rect 3525 5117 3559 5151
rect 3893 5117 3927 5151
rect 5273 5117 5307 5151
rect 6745 5117 6779 5151
rect 13093 5117 13127 5151
rect 14749 5117 14783 5151
rect 15853 5117 15887 5151
rect 16957 5117 16991 5151
rect 5733 5049 5767 5083
rect 2881 4981 2915 5015
rect 4445 4981 4479 5015
rect 4813 4981 4847 5015
rect 11897 4981 11931 5015
rect 12633 4981 12667 5015
rect 13737 4981 13771 5015
rect 15577 4981 15611 5015
rect 18061 4981 18095 5015
rect 2145 4777 2179 4811
rect 3985 4777 4019 4811
rect 4261 4777 4295 4811
rect 4905 4777 4939 4811
rect 13369 4777 13403 4811
rect 15853 4777 15887 4811
rect 17693 4777 17727 4811
rect 2053 4709 2087 4743
rect 9781 4709 9815 4743
rect 13553 4709 13587 4743
rect 1685 4641 1719 4675
rect 6745 4641 6779 4675
rect 12265 4641 12299 4675
rect 13001 4641 13035 4675
rect 15393 4641 15427 4675
rect 17049 4641 17083 4675
rect 3801 4573 3835 4607
rect 3955 4573 3989 4607
rect 4445 4573 4479 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 4813 4573 4847 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 6929 4573 6963 4607
rect 9413 4573 9447 4607
rect 10425 4573 10459 4607
rect 11253 4573 11287 4607
rect 14105 4573 14139 4607
rect 15485 4573 15519 4607
rect 8125 4505 8159 4539
rect 7113 4437 7147 4471
rect 8217 4437 8251 4471
rect 9873 4437 9907 4471
rect 10609 4437 10643 4471
rect 11805 4437 11839 4471
rect 12909 4437 12943 4471
rect 13369 4437 13403 4471
rect 14289 4437 14323 4471
rect 7665 4233 7699 4267
rect 9229 4233 9263 4267
rect 12173 4233 12207 4267
rect 14749 4233 14783 4267
rect 11989 4165 12023 4199
rect 12909 4165 12943 4199
rect 13553 4165 13587 4199
rect 4813 4097 4847 4131
rect 5181 4097 5215 4131
rect 6561 4097 6595 4131
rect 6745 4097 6779 4131
rect 6837 4097 6871 4131
rect 7849 4097 7883 4131
rect 8116 4097 8150 4131
rect 9873 4097 9907 4131
rect 10140 4097 10174 4131
rect 11621 4097 11655 4131
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 13185 4097 13219 4131
rect 13461 4097 13495 4131
rect 14381 4097 14415 4131
rect 14657 4097 14691 4131
rect 15025 4097 15059 4131
rect 15209 4097 15243 4131
rect 15393 4097 15427 4131
rect 4997 4029 5031 4063
rect 7113 4029 7147 4063
rect 12633 4029 12667 4063
rect 12725 4029 12759 4063
rect 13001 4029 13035 4063
rect 14934 4029 14968 4063
rect 15117 4029 15151 4063
rect 3065 3961 3099 3995
rect 6653 3961 6687 3995
rect 11253 3961 11287 3995
rect 13369 3961 13403 3995
rect 5089 3893 5123 3927
rect 6377 3893 6411 3927
rect 11989 3893 12023 3927
rect 12265 3893 12299 3927
rect 12909 3893 12943 3927
rect 14197 3893 14231 3927
rect 14565 3893 14599 3927
rect 15485 3893 15519 3927
rect 8769 3689 8803 3723
rect 12541 3689 12575 3723
rect 13001 3689 13035 3723
rect 15025 3689 15059 3723
rect 16037 3689 16071 3723
rect 16773 3689 16807 3723
rect 4445 3621 4479 3655
rect 5549 3621 5583 3655
rect 7481 3621 7515 3655
rect 1685 3553 1719 3587
rect 6101 3553 6135 3587
rect 7113 3553 7147 3587
rect 7573 3553 7607 3587
rect 7757 3553 7791 3587
rect 12633 3553 12667 3587
rect 13093 3553 13127 3587
rect 14289 3553 14323 3587
rect 16129 3553 16163 3587
rect 1409 3485 1443 3519
rect 2145 3485 2179 3519
rect 2421 3485 2455 3519
rect 2697 3485 2731 3519
rect 2790 3485 2824 3519
rect 3617 3485 3651 3519
rect 4629 3485 4663 3519
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 5457 3485 5491 3519
rect 6009 3485 6043 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 7021 3485 7055 3519
rect 7298 3485 7332 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 7849 3485 7883 3519
rect 8125 3485 8159 3519
rect 12817 3485 12851 3519
rect 13369 3485 13403 3519
rect 15301 3485 15335 3519
rect 15485 3485 15519 3519
rect 19349 3485 19383 3519
rect 28089 3485 28123 3519
rect 3065 3417 3099 3451
rect 7205 3417 7239 3451
rect 12541 3417 12575 3451
rect 15025 3417 15059 3451
rect 1961 3349 1995 3383
rect 2237 3349 2271 3383
rect 3433 3349 3467 3383
rect 14933 3349 14967 3383
rect 15209 3349 15243 3383
rect 17049 3349 17083 3383
rect 19901 3349 19935 3383
rect 28641 3349 28675 3383
rect 5273 3145 5307 3179
rect 5733 3145 5767 3179
rect 6653 3145 6687 3179
rect 7113 3145 7147 3179
rect 9413 3145 9447 3179
rect 10793 3145 10827 3179
rect 12265 3145 12299 3179
rect 15393 3145 15427 3179
rect 17877 3145 17911 3179
rect 20085 3145 20119 3179
rect 26801 3145 26835 3179
rect 27445 3145 27479 3179
rect 28917 3145 28951 3179
rect 29653 3145 29687 3179
rect 33885 3145 33919 3179
rect 37013 3145 37047 3179
rect 5181 3077 5215 3111
rect 5549 3077 5583 3111
rect 7481 3077 7515 3111
rect 11805 3077 11839 3111
rect 14280 3077 14314 3111
rect 26985 3077 27019 3111
rect 33241 3077 33275 3111
rect 35725 3077 35759 3111
rect 3801 3009 3835 3043
rect 5641 3009 5675 3043
rect 7021 3009 7055 3043
rect 7757 3009 7791 3043
rect 8217 3009 8251 3043
rect 8401 3009 8435 3043
rect 8953 3009 8987 3043
rect 9505 3009 9539 3043
rect 10425 3009 10459 3043
rect 10517 3009 10551 3043
rect 12081 3009 12115 3043
rect 14013 3009 14047 3043
rect 16313 3009 16347 3043
rect 17417 3009 17451 3043
rect 17693 3009 17727 3043
rect 19625 3009 19659 3043
rect 19901 3009 19935 3043
rect 25053 3009 25087 3043
rect 25329 3009 25363 3043
rect 26341 3009 26375 3043
rect 26525 3009 26559 3043
rect 26617 3009 26651 3043
rect 27261 3009 27295 3043
rect 28457 3009 28491 3043
rect 28733 3009 28767 3043
rect 33701 3009 33735 3043
rect 36001 3009 36035 3043
rect 36185 3009 36219 3043
rect 36461 3009 36495 3043
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 1869 2941 1903 2975
rect 2881 2941 2915 2975
rect 4169 2941 4203 2975
rect 5365 2941 5399 2975
rect 7297 2941 7331 2975
rect 7573 2941 7607 2975
rect 11897 2941 11931 2975
rect 15669 2941 15703 2975
rect 16773 2941 16807 2975
rect 17325 2941 17359 2975
rect 17509 2941 17543 2975
rect 19809 2941 19843 2975
rect 20177 2941 20211 2975
rect 25145 2941 25179 2975
rect 27169 2941 27203 2975
rect 28641 2941 28675 2975
rect 29101 2941 29135 2975
rect 33517 2941 33551 2975
rect 36737 2941 36771 2975
rect 8033 2873 8067 2907
rect 8769 2873 8803 2907
rect 9321 2873 9355 2907
rect 9873 2873 9907 2907
rect 20821 2873 20855 2907
rect 36369 2873 36403 2907
rect 5457 2805 5491 2839
rect 7757 2805 7791 2839
rect 7941 2805 7975 2839
rect 8861 2805 8895 2839
rect 9965 2805 9999 2839
rect 10425 2805 10459 2839
rect 12081 2805 12115 2839
rect 17417 2805 17451 2839
rect 19901 2805 19935 2839
rect 25329 2805 25363 2839
rect 25513 2805 25547 2839
rect 26341 2805 26375 2839
rect 26985 2805 27019 2839
rect 28733 2805 28767 2839
rect 33701 2805 33735 2839
rect 36185 2805 36219 2839
rect 36829 2805 36863 2839
rect 38485 2805 38519 2839
rect 1777 2601 1811 2635
rect 2605 2601 2639 2635
rect 3617 2601 3651 2635
rect 4445 2601 4479 2635
rect 6377 2601 6411 2635
rect 8309 2601 8343 2635
rect 10425 2601 10459 2635
rect 11069 2601 11103 2635
rect 12173 2601 12207 2635
rect 16681 2601 16715 2635
rect 17141 2601 17175 2635
rect 17693 2601 17727 2635
rect 19625 2601 19659 2635
rect 21005 2601 21039 2635
rect 22109 2601 22143 2635
rect 24409 2601 24443 2635
rect 25421 2601 25455 2635
rect 27629 2601 27663 2635
rect 29561 2601 29595 2635
rect 30113 2601 30147 2635
rect 30941 2601 30975 2635
rect 33149 2601 33183 2635
rect 34253 2601 34287 2635
rect 35357 2601 35391 2635
rect 36461 2601 36495 2635
rect 37565 2601 37599 2635
rect 38025 2601 38059 2635
rect 2789 2533 2823 2567
rect 4537 2533 4571 2567
rect 8769 2533 8803 2567
rect 14381 2533 14415 2567
rect 15209 2533 15243 2567
rect 17969 2533 18003 2567
rect 23213 2533 23247 2567
rect 26525 2533 26559 2567
rect 30021 2533 30055 2567
rect 32137 2533 32171 2567
rect 3801 2465 3835 2499
rect 5273 2465 5307 2499
rect 7113 2465 7147 2499
rect 9413 2465 9447 2499
rect 16129 2465 16163 2499
rect 16773 2465 16807 2499
rect 1593 2397 1627 2431
rect 1961 2397 1995 2431
rect 2053 2397 2087 2431
rect 2145 2397 2179 2431
rect 2329 2397 2363 2431
rect 2421 2397 2455 2431
rect 2605 2397 2639 2431
rect 2973 2397 3007 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 6561 2397 6595 2431
rect 6745 2397 6779 2431
rect 8493 2397 8527 2431
rect 8953 2397 8987 2431
rect 10609 2397 10643 2431
rect 10885 2397 10919 2431
rect 11253 2397 11287 2431
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 13093 2397 13127 2431
rect 13461 2397 13495 2431
rect 14289 2397 14323 2431
rect 14565 2397 14599 2431
rect 15393 2397 15427 2431
rect 15485 2397 15519 2431
rect 16497 2397 16531 2431
rect 16957 2397 16991 2431
rect 17509 2397 17543 2431
rect 17877 2397 17911 2431
rect 18153 2397 18187 2431
rect 18613 2397 18647 2431
rect 18981 2397 19015 2431
rect 19533 2397 19567 2431
rect 19809 2397 19843 2431
rect 19901 2397 19935 2431
rect 20821 2397 20855 2431
rect 21189 2397 21223 2431
rect 22017 2397 22051 2431
rect 22293 2397 22327 2431
rect 23029 2397 23063 2431
rect 23397 2397 23431 2431
rect 24133 2397 24167 2431
rect 24593 2397 24627 2431
rect 25237 2397 25271 2431
rect 25605 2397 25639 2431
rect 26341 2397 26375 2431
rect 26709 2397 26743 2431
rect 27445 2397 27479 2431
rect 27813 2397 27847 2431
rect 28549 2397 28583 2431
rect 28733 2397 28767 2431
rect 29377 2397 29411 2431
rect 29745 2397 29779 2431
rect 30297 2397 30331 2431
rect 30757 2397 30791 2431
rect 31125 2397 31159 2431
rect 31861 2397 31895 2431
rect 32321 2397 32355 2431
rect 32965 2397 32999 2431
rect 33333 2397 33367 2431
rect 34069 2397 34103 2431
rect 34437 2397 34471 2431
rect 35173 2397 35207 2431
rect 35541 2397 35575 2431
rect 36277 2397 36311 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 37749 2397 37783 2431
rect 38209 2397 38243 2431
rect 38485 2397 38519 2431
rect 16681 2329 16715 2363
rect 20545 2329 20579 2363
rect 13277 2261 13311 2295
rect 14933 2261 14967 2295
rect 18797 2261 18831 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 38102 34960 38108 35012
rect 38160 34960 38166 35012
rect 38194 34892 38200 34944
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 38105 25211 38163 25217
rect 38105 25177 38117 25211
rect 38151 25208 38163 25211
rect 38151 25180 39068 25208
rect 38151 25177 38163 25180
rect 38105 25171 38163 25177
rect 38010 25100 38016 25152
rect 38068 25140 38074 25152
rect 38197 25143 38255 25149
rect 38197 25140 38209 25143
rect 38068 25112 38209 25140
rect 38068 25100 38074 25112
rect 38197 25109 38209 25112
rect 38243 25109 38255 25143
rect 38197 25103 38255 25109
rect 39040 25084 39068 25180
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 39022 25032 39028 25084
rect 39080 25032 39086 25084
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 14458 16028 14464 16040
rect 14231 16000 14464 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14458 15988 14464 16000
rect 14516 15988 14522 16040
rect 14734 15852 14740 15904
rect 14792 15852 14798 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 11790 15444 11796 15496
rect 11848 15444 11854 15496
rect 14550 15444 14556 15496
rect 14608 15444 14614 15496
rect 38197 15487 38255 15493
rect 38197 15453 38209 15487
rect 38243 15484 38255 15487
rect 38243 15456 38976 15484
rect 38243 15453 38255 15456
rect 38197 15447 38255 15453
rect 12437 15351 12495 15357
rect 12437 15317 12449 15351
rect 12483 15348 12495 15351
rect 12526 15348 12532 15360
rect 12483 15320 12532 15348
rect 12483 15317 12495 15320
rect 12437 15311 12495 15317
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 15102 15308 15108 15360
rect 15160 15308 15166 15360
rect 38378 15308 38384 15360
rect 38436 15308 38442 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 38948 15224 38976 15456
rect 1104 15184 38824 15206
rect 38930 15172 38936 15224
rect 38988 15172 38994 15224
rect 14550 15104 14556 15156
rect 14608 15104 14614 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14792 15116 14933 15144
rect 14792 15104 14798 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15059 15116 15577 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 14090 15076 14096 15088
rect 11532 15048 14096 15076
rect 11532 15017 11560 15048
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 11784 15011 11842 15017
rect 11784 14977 11796 15011
rect 11830 15008 11842 15011
rect 12526 15008 12532 15020
rect 11830 14980 12532 15008
rect 11830 14977 11842 14980
rect 11784 14971 11842 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 13096 15017 13124 15048
rect 14090 15036 14096 15048
rect 14148 15036 14154 15088
rect 15102 15036 15108 15088
rect 15160 15036 15166 15088
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13348 15011 13406 15017
rect 13348 14977 13360 15011
rect 13394 15008 13406 15011
rect 15120 15008 15148 15036
rect 13394 14980 15148 15008
rect 13394 14977 13406 14980
rect 13348 14971 13406 14977
rect 8110 14900 8116 14952
rect 8168 14900 8174 14952
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 10594 14940 10600 14952
rect 10367 14912 10600 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 8864 14816 8892 14903
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 15120 14872 15148 14903
rect 12452 14844 13032 14872
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 8846 14764 8852 14816
rect 8904 14764 8910 14816
rect 9398 14764 9404 14816
rect 9456 14764 9462 14816
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 12452 14804 12480 14844
rect 11388 14776 12480 14804
rect 11388 14764 11394 14776
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13004 14804 13032 14844
rect 14016 14844 15148 14872
rect 15580 14872 15608 15107
rect 16114 14900 16120 14952
rect 16172 14940 16178 14952
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16172 14912 16681 14940
rect 16172 14900 16178 14912
rect 16669 14909 16681 14912
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 15580 14844 17632 14872
rect 14016 14804 14044 14844
rect 17604 14816 17632 14844
rect 13004 14776 14044 14804
rect 14458 14764 14464 14816
rect 14516 14764 14522 14816
rect 17310 14764 17316 14816
rect 17368 14764 17374 14816
rect 17586 14764 17592 14816
rect 17644 14764 17650 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 8757 14603 8815 14609
rect 8757 14569 8769 14603
rect 8803 14600 8815 14603
rect 8846 14600 8852 14612
rect 8803 14572 8852 14600
rect 8803 14569 8815 14572
rect 8757 14563 8815 14569
rect 8846 14560 8852 14572
rect 8904 14600 8910 14612
rect 9950 14600 9956 14612
rect 8904 14572 9956 14600
rect 8904 14560 8910 14572
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10870 14560 10876 14612
rect 10928 14560 10934 14612
rect 11790 14560 11796 14612
rect 11848 14560 11854 14612
rect 17310 14600 17316 14612
rect 17144 14572 17316 14600
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 7432 14368 9229 14396
rect 7432 14356 7438 14368
rect 9217 14365 9229 14368
rect 9263 14396 9275 14399
rect 10888 14396 10916 14560
rect 16758 14492 16764 14544
rect 16816 14492 16822 14544
rect 11330 14424 11336 14476
rect 11388 14424 11394 14476
rect 12342 14424 12348 14476
rect 12400 14424 12406 14476
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 12894 14464 12900 14476
rect 12759 14436 12900 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 14090 14424 14096 14476
rect 14148 14464 14154 14476
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14148 14436 14749 14464
rect 14148 14424 14154 14436
rect 14737 14433 14749 14436
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 17144 14405 17172 14572
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17405 14467 17463 14473
rect 17405 14433 17417 14467
rect 17451 14464 17463 14467
rect 19426 14464 19432 14476
rect 17451 14436 19432 14464
rect 17451 14433 17463 14436
rect 17405 14427 17463 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 20530 14424 20536 14476
rect 20588 14464 20594 14476
rect 38010 14464 38016 14476
rect 20588 14436 38016 14464
rect 20588 14424 20594 14436
rect 38010 14424 38016 14436
rect 38068 14424 38074 14476
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 9263 14368 9352 14396
rect 10888 14368 11069 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 7644 14331 7702 14337
rect 7644 14297 7656 14331
rect 7690 14328 7702 14331
rect 8662 14328 8668 14340
rect 7690 14300 8668 14328
rect 7690 14297 7702 14300
rect 7644 14291 7702 14297
rect 8662 14288 8668 14300
rect 8720 14288 8726 14340
rect 9324 14272 9352 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 17129 14359 17187 14365
rect 17678 14356 17684 14408
rect 17736 14356 17742 14408
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 19334 14356 19340 14408
rect 19392 14356 19398 14408
rect 9484 14331 9542 14337
rect 9484 14297 9496 14331
rect 9530 14328 9542 14331
rect 11238 14328 11244 14340
rect 9530 14300 11244 14328
rect 9530 14297 9542 14300
rect 9484 14291 9542 14297
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 13265 14331 13323 14337
rect 13265 14328 13277 14331
rect 12207 14300 13277 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 13265 14297 13277 14300
rect 13311 14297 13323 14331
rect 13265 14291 13323 14297
rect 15004 14331 15062 14337
rect 15004 14297 15016 14331
rect 15050 14328 15062 14331
rect 17310 14328 17316 14340
rect 15050 14300 17316 14328
rect 15050 14297 15062 14300
rect 15004 14291 15062 14297
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 17788 14300 26234 14328
rect 9306 14220 9312 14272
rect 9364 14220 9370 14272
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 10686 14220 10692 14272
rect 10744 14220 10750 14272
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11422 14260 11428 14272
rect 11195 14232 11428 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 13078 14260 13084 14272
rect 12299 14232 13084 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 13078 14220 13084 14232
rect 13136 14260 13142 14272
rect 13541 14263 13599 14269
rect 13541 14260 13553 14263
rect 13136 14232 13553 14260
rect 13136 14220 13142 14232
rect 13541 14229 13553 14232
rect 13587 14229 13599 14263
rect 13541 14223 13599 14229
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 16114 14260 16120 14272
rect 15252 14232 16120 14260
rect 15252 14220 15258 14232
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 16574 14260 16580 14272
rect 16531 14232 16580 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 16574 14220 16580 14232
rect 16632 14260 16638 14272
rect 17221 14263 17279 14269
rect 17221 14260 17233 14263
rect 16632 14232 17233 14260
rect 16632 14220 16638 14232
rect 17221 14229 17233 14232
rect 17267 14260 17279 14263
rect 17586 14260 17592 14272
rect 17267 14232 17592 14260
rect 17267 14229 17279 14232
rect 17221 14223 17279 14229
rect 17586 14220 17592 14232
rect 17644 14260 17650 14272
rect 17788 14260 17816 14300
rect 17644 14232 17816 14260
rect 17644 14220 17650 14232
rect 18230 14220 18236 14272
rect 18288 14220 18294 14272
rect 19058 14220 19064 14272
rect 19116 14220 19122 14272
rect 19978 14220 19984 14272
rect 20036 14220 20042 14272
rect 26206 14260 26234 14300
rect 38194 14260 38200 14272
rect 26206 14232 38200 14260
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 8168 14028 8309 14056
rect 8168 14016 8174 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 8297 14019 8355 14025
rect 8665 14059 8723 14065
rect 8665 14025 8677 14059
rect 8711 14056 8723 14059
rect 9398 14056 9404 14068
rect 8711 14028 9404 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 11238 14016 11244 14068
rect 11296 14016 11302 14068
rect 16574 14056 16580 14068
rect 16408 14028 16580 14056
rect 10704 13929 10732 14016
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 10689 13923 10747 13929
rect 8803 13892 9444 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 9416 13861 9444 13892
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 8941 13855 8999 13861
rect 8941 13821 8953 13855
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9490 13852 9496 13864
rect 9447 13824 9496 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 8956 13784 8984 13815
rect 9490 13812 9496 13824
rect 9548 13852 9554 13864
rect 11422 13852 11428 13864
rect 9548 13824 11428 13852
rect 9548 13812 9554 13824
rect 11422 13812 11428 13824
rect 11480 13852 11486 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11480 13824 11713 13852
rect 11480 13812 11486 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 12158 13812 12164 13864
rect 12216 13812 12222 13864
rect 16408 13861 16436 14028
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 16758 14016 16764 14068
rect 16816 14016 16822 14068
rect 17310 14016 17316 14068
rect 17368 14016 17374 14068
rect 17678 14016 17684 14068
rect 17736 14016 17742 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 19058 14056 19064 14068
rect 18095 14028 19064 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19978 14016 19984 14068
rect 20036 14016 20042 14068
rect 16776 13929 16804 14016
rect 17770 13948 17776 14000
rect 17828 13988 17834 14000
rect 19328 13991 19386 13997
rect 17828 13960 19104 13988
rect 17828 13948 17834 13960
rect 19076 13929 19104 13960
rect 19328 13957 19340 13991
rect 19374 13988 19386 13991
rect 19996 13988 20024 14016
rect 19374 13960 20024 13988
rect 19374 13957 19386 13960
rect 19328 13951 19386 13957
rect 20530 13948 20536 14000
rect 20588 13948 20594 14000
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13920 18199 13923
rect 19061 13923 19119 13929
rect 18187 13892 18828 13920
rect 18187 13889 18199 13892
rect 18141 13883 18199 13889
rect 18800 13861 18828 13892
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 20548 13920 20576 13948
rect 19061 13883 19119 13889
rect 19168 13892 20576 13920
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13832 13824 14197 13852
rect 12342 13784 12348 13796
rect 8956 13756 12348 13784
rect 9600 13728 9628 13756
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 9582 13676 9588 13728
rect 9640 13676 9646 13728
rect 12710 13676 12716 13728
rect 12768 13676 12774 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13832 13725 13860 13824
rect 14185 13821 14197 13824
rect 14231 13852 14243 13855
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 14231 13824 14565 13852
rect 14231 13821 14243 13824
rect 14185 13815 14243 13821
rect 14553 13821 14565 13824
rect 14599 13852 14611 13855
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14599 13824 14933 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14921 13821 14933 13824
rect 14967 13852 14979 13855
rect 15289 13855 15347 13861
rect 15289 13852 15301 13855
rect 14967 13824 15301 13852
rect 14967 13821 14979 13824
rect 14921 13815 14979 13821
rect 15289 13821 15301 13824
rect 15335 13852 15347 13855
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 15335 13824 15669 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15657 13821 15669 13824
rect 15703 13852 15715 13855
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15703 13824 16037 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 16025 13821 16037 13824
rect 16071 13852 16083 13855
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 16071 13824 16405 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16393 13815 16451 13821
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18233 13815 18291 13821
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13852 18843 13855
rect 19168 13852 19196 13892
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 18831 13824 19196 13852
rect 20456 13824 20545 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 18248 13784 18276 13815
rect 18156 13756 18276 13784
rect 18156 13728 18184 13756
rect 20456 13728 20484 13824
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 13136 13688 13461 13716
rect 13136 13676 13142 13688
rect 13449 13685 13461 13688
rect 13495 13716 13507 13719
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 13495 13688 13829 13716
rect 13495 13685 13507 13688
rect 13449 13679 13507 13685
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 13817 13679 13875 13685
rect 18138 13676 18144 13728
rect 18196 13676 18202 13728
rect 20438 13676 20444 13728
rect 20496 13676 20502 13728
rect 21174 13676 21180 13728
rect 21232 13676 21238 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9398 13512 9404 13524
rect 8803 13484 9404 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9398 13472 9404 13484
rect 9456 13512 9462 13524
rect 14458 13512 14464 13524
rect 9456 13484 11652 13512
rect 9456 13472 9462 13484
rect 9306 13336 9312 13388
rect 9364 13376 9370 13388
rect 10597 13379 10655 13385
rect 10597 13376 10609 13379
rect 9364 13348 10609 13376
rect 9364 13336 9370 13348
rect 10597 13345 10609 13348
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 11624 13308 11652 13484
rect 11900 13484 14464 13512
rect 11900 13376 11928 13484
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16761 13515 16819 13521
rect 16761 13512 16773 13515
rect 16632 13484 16773 13512
rect 16632 13472 16638 13484
rect 16761 13481 16773 13484
rect 16807 13481 16819 13515
rect 16761 13475 16819 13481
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 18564 13484 18613 13512
rect 18564 13472 18570 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 18601 13475 18659 13481
rect 19334 13472 19340 13524
rect 19392 13472 19398 13524
rect 20441 13515 20499 13521
rect 20441 13481 20453 13515
rect 20487 13512 20499 13515
rect 20530 13512 20536 13524
rect 20487 13484 20536 13512
rect 20487 13481 20499 13484
rect 20441 13475 20499 13481
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 11977 13447 12035 13453
rect 11977 13413 11989 13447
rect 12023 13444 12035 13447
rect 12158 13444 12164 13456
rect 12023 13416 12164 13444
rect 12023 13413 12035 13416
rect 11977 13407 12035 13413
rect 12158 13404 12164 13416
rect 12216 13444 12222 13456
rect 15657 13447 15715 13453
rect 12216 13416 12848 13444
rect 12216 13404 12222 13416
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11900 13348 12081 13376
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12618 13376 12624 13388
rect 12069 13339 12127 13345
rect 12176 13348 12624 13376
rect 12176 13308 12204 13348
rect 12618 13336 12624 13348
rect 12676 13376 12682 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12676 13348 12725 13376
rect 12676 13336 12682 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12820 13376 12848 13416
rect 15657 13413 15669 13447
rect 15703 13444 15715 13447
rect 15930 13444 15936 13456
rect 15703 13416 15936 13444
rect 15703 13413 15715 13416
rect 15657 13407 15715 13413
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 16316 13416 16574 13444
rect 13106 13379 13164 13385
rect 13106 13376 13118 13379
rect 12820 13348 13118 13376
rect 12713 13339 12771 13345
rect 13106 13345 13118 13348
rect 13152 13345 13164 13379
rect 13106 13339 13164 13345
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 14148 13348 14289 13376
rect 14148 13336 14154 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 9263 13280 10088 13308
rect 11624 13280 12204 13308
rect 12253 13311 12311 13317
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 10060 13184 10088 13280
rect 12253 13277 12265 13311
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 10864 13243 10922 13249
rect 10864 13209 10876 13243
rect 10910 13240 10922 13243
rect 11882 13240 11888 13252
rect 10910 13212 11888 13240
rect 10910 13209 10922 13212
rect 10864 13203 10922 13209
rect 11882 13200 11888 13212
rect 11940 13200 11946 13252
rect 9766 13132 9772 13184
rect 9824 13132 9830 13184
rect 10042 13132 10048 13184
rect 10100 13132 10106 13184
rect 12268 13172 12296 13271
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 14292 13308 14320 13339
rect 16316 13308 16344 13416
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 14292 13280 16344 13308
rect 14544 13243 14602 13249
rect 14544 13209 14556 13243
rect 14590 13240 14602 13243
rect 15838 13240 15844 13252
rect 14590 13212 15844 13240
rect 14590 13209 14602 13212
rect 14544 13203 14602 13209
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 16408 13240 16436 13339
rect 16546 13308 16574 13416
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19484 13348 19901 13376
rect 19484 13336 19490 13348
rect 19889 13345 19901 13348
rect 19935 13376 19947 13379
rect 20162 13376 20168 13388
rect 19935 13348 20168 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16546 13280 17233 13308
rect 17221 13277 17233 13280
rect 17267 13308 17279 13311
rect 17770 13308 17776 13320
rect 17267 13280 17776 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18230 13268 18236 13320
rect 18288 13268 18294 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 21174 13308 21180 13320
rect 19751 13280 21180 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 17488 13243 17546 13249
rect 16408 13212 17448 13240
rect 13814 13172 13820 13184
rect 12268 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 13906 13132 13912 13184
rect 13964 13132 13970 13184
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 16209 13175 16267 13181
rect 16209 13141 16221 13175
rect 16255 13172 16267 13175
rect 16574 13172 16580 13184
rect 16255 13144 16580 13172
rect 16255 13141 16267 13144
rect 16209 13135 16267 13141
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 17420 13172 17448 13212
rect 17488 13209 17500 13243
rect 17534 13240 17546 13243
rect 18248 13240 18276 13268
rect 17534 13212 18276 13240
rect 19797 13243 19855 13249
rect 17534 13209 17546 13212
rect 17488 13203 17546 13209
rect 19797 13209 19809 13243
rect 19843 13240 19855 13243
rect 20530 13240 20536 13252
rect 19843 13212 20536 13240
rect 19843 13209 19855 13212
rect 19797 13203 19855 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 18138 13172 18144 13184
rect 17420 13144 18144 13172
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 8757 12971 8815 12977
rect 8757 12937 8769 12971
rect 8803 12968 8815 12971
rect 10042 12968 10048 12980
rect 8803 12940 10048 12968
rect 8803 12937 8815 12940
rect 8757 12931 8815 12937
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 12069 12971 12127 12977
rect 10284 12940 12020 12968
rect 10284 12928 10290 12940
rect 11992 12900 12020 12940
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 12710 12968 12716 12980
rect 12115 12940 12716 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 13906 12968 13912 12980
rect 13771 12940 13912 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 15746 12928 15752 12980
rect 15804 12928 15810 12980
rect 15838 12928 15844 12980
rect 15896 12928 15902 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 16172 12940 17325 12968
rect 16172 12928 16178 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 20438 12968 20444 12980
rect 17313 12931 17371 12937
rect 18432 12940 20444 12968
rect 13262 12900 13268 12912
rect 11992 12872 13268 12900
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 7374 12792 7380 12844
rect 7432 12792 7438 12844
rect 7644 12835 7702 12841
rect 7644 12801 7656 12835
rect 7690 12832 7702 12835
rect 8754 12832 8760 12844
rect 7690 12804 8760 12832
rect 7690 12801 7702 12804
rect 7644 12795 7702 12801
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9950 12792 9956 12844
rect 10008 12792 10014 12844
rect 10042 12792 10048 12844
rect 10100 12841 10106 12844
rect 10100 12835 10128 12841
rect 10116 12801 10128 12835
rect 10100 12795 10128 12801
rect 10100 12792 10106 12795
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 13633 12835 13691 12841
rect 12023 12804 12756 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 11146 12764 11152 12776
rect 9263 12736 11152 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 9048 12628 9076 12727
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 12161 12767 12219 12773
rect 12161 12764 12173 12767
rect 11296 12736 12173 12764
rect 11296 12724 11302 12736
rect 12161 12733 12173 12736
rect 12207 12733 12219 12767
rect 12161 12727 12219 12733
rect 12618 12724 12624 12776
rect 12676 12724 12682 12776
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 9456 12668 9689 12696
rect 9456 12656 9462 12668
rect 9677 12665 9689 12668
rect 9723 12665 9735 12699
rect 9677 12659 9735 12665
rect 11333 12699 11391 12705
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 12636 12696 12664 12724
rect 11379 12668 12664 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 12728 12640 12756 12804
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15764 12832 15792 12928
rect 18432 12841 18460 12940
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 15335 12804 15792 12832
rect 18417 12835 18475 12841
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 13648 12696 13676 12795
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 18564 12804 18828 12832
rect 18564 12792 18570 12804
rect 13722 12724 13728 12776
rect 13780 12764 13786 12776
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13780 12736 13829 12764
rect 13780 12724 13786 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 16669 12767 16727 12773
rect 16669 12764 16681 12767
rect 15988 12736 16681 12764
rect 15988 12724 15994 12736
rect 16669 12733 16681 12736
rect 16715 12733 16727 12767
rect 16669 12727 16727 12733
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12733 18659 12767
rect 18800 12764 18828 12804
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 18800 12736 19349 12764
rect 18601 12727 18659 12733
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19337 12727 19395 12733
rect 17034 12696 17040 12708
rect 12860 12668 13400 12696
rect 13648 12668 17040 12696
rect 12860 12656 12866 12668
rect 10594 12628 10600 12640
rect 9048 12600 10600 12628
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 10744 12600 10885 12628
rect 10744 12588 10750 12600
rect 10873 12597 10885 12600
rect 10919 12597 10931 12631
rect 10873 12591 10931 12597
rect 11606 12588 11612 12640
rect 11664 12588 11670 12640
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 13078 12628 13084 12640
rect 12768 12600 13084 12628
rect 12768 12588 12774 12600
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13262 12588 13268 12640
rect 13320 12588 13326 12640
rect 13372 12628 13400 12668
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 15838 12628 15844 12640
rect 13372 12600 15844 12628
rect 15838 12588 15844 12600
rect 15896 12628 15902 12640
rect 18230 12628 18236 12640
rect 15896 12600 18236 12628
rect 15896 12588 15902 12600
rect 18230 12588 18236 12600
rect 18288 12628 18294 12640
rect 18506 12628 18512 12640
rect 18288 12600 18512 12628
rect 18288 12588 18294 12600
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 18616 12628 18644 12727
rect 19426 12724 19432 12776
rect 19484 12773 19490 12776
rect 19484 12767 19512 12773
rect 19500 12733 19512 12767
rect 19484 12727 19512 12733
rect 19484 12724 19490 12727
rect 19610 12724 19616 12776
rect 19668 12724 19674 12776
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 19061 12699 19119 12705
rect 19061 12696 19073 12699
rect 18748 12668 19073 12696
rect 18748 12656 18754 12668
rect 19061 12665 19073 12668
rect 19107 12665 19119 12699
rect 19061 12659 19119 12665
rect 20070 12628 20076 12640
rect 18616 12600 20076 12628
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 8754 12384 8760 12436
rect 8812 12384 8818 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11422 12424 11428 12436
rect 11195 12396 11428 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11882 12384 11888 12436
rect 11940 12384 11946 12436
rect 12406 12396 16804 12424
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 8220 12328 8953 12356
rect 8220 12297 8248 12328
rect 8941 12325 8953 12328
rect 8987 12325 8999 12359
rect 12406 12356 12434 12396
rect 8941 12319 8999 12325
rect 9508 12328 10364 12356
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12257 8263 12291
rect 8205 12251 8263 12257
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 9508 12297 9536 12328
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9272 12260 9505 12288
rect 9272 12248 9278 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9784 12220 9812 12248
rect 9447 12192 9812 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 9309 12155 9367 12161
rect 9309 12121 9321 12155
rect 9355 12152 9367 12155
rect 9490 12152 9496 12164
rect 9355 12124 9496 12152
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 10336 12152 10364 12328
rect 10428 12328 12434 12356
rect 10428 12229 10456 12328
rect 12710 12316 12716 12368
rect 12768 12356 12774 12368
rect 13081 12359 13139 12365
rect 13081 12356 13093 12359
rect 12768 12328 13093 12356
rect 12768 12316 12774 12328
rect 13081 12325 13093 12328
rect 13127 12356 13139 12359
rect 13446 12356 13452 12368
rect 13127 12328 13452 12356
rect 13127 12325 13139 12328
rect 13081 12319 13139 12325
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 15105 12359 15163 12365
rect 15105 12325 15117 12359
rect 15151 12356 15163 12359
rect 15838 12356 15844 12368
rect 15151 12328 15844 12356
rect 15151 12325 15163 12328
rect 15105 12319 15163 12325
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 16776 12356 16804 12396
rect 17034 12384 17040 12436
rect 17092 12384 17098 12436
rect 20254 12356 20260 12368
rect 16776 12328 20260 12356
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 10594 12248 10600 12300
rect 10652 12248 10658 12300
rect 10686 12248 10692 12300
rect 10744 12248 10750 12300
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 11606 12288 11612 12300
rect 11379 12260 11612 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 15194 12248 15200 12300
rect 15252 12248 15258 12300
rect 16114 12248 16120 12300
rect 16172 12248 16178 12300
rect 16393 12291 16451 12297
rect 16393 12257 16405 12291
rect 16439 12288 16451 12291
rect 19610 12288 19616 12300
rect 16439 12260 19616 12288
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10704 12220 10732 12248
rect 18800 12232 18828 12260
rect 19610 12248 19616 12260
rect 19668 12248 19674 12300
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 20530 12288 20536 12300
rect 20128 12260 20536 12288
rect 20128 12248 20134 12260
rect 20530 12248 20536 12260
rect 20588 12288 20594 12300
rect 20717 12291 20775 12297
rect 20717 12288 20729 12291
rect 20588 12260 20729 12288
rect 20588 12248 20594 12260
rect 20717 12257 20729 12260
rect 20763 12257 20775 12291
rect 20717 12251 20775 12257
rect 10551 12192 10732 12220
rect 15381 12223 15439 12229
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 15381 12189 15393 12223
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 11238 12152 11244 12164
rect 10336 12124 11244 12152
rect 11238 12112 11244 12124
rect 11296 12112 11302 12164
rect 13722 12152 13728 12164
rect 12406 12124 13728 12152
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 9916 12056 10057 12084
rect 9916 12044 9922 12056
rect 10045 12053 10057 12056
rect 10091 12053 10103 12087
rect 10045 12047 10103 12053
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 12406 12084 12434 12124
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 10652 12056 12434 12084
rect 15396 12084 15424 12183
rect 16206 12180 16212 12232
rect 16264 12229 16270 12232
rect 16264 12223 16292 12229
rect 16280 12189 16292 12223
rect 16264 12183 16292 12189
rect 16264 12180 16270 12183
rect 18782 12180 18788 12232
rect 18840 12180 18846 12232
rect 19978 12180 19984 12232
rect 20036 12180 20042 12232
rect 16666 12084 16672 12096
rect 15396 12056 16672 12084
rect 10652 12044 10658 12056
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 20622 12044 20628 12096
rect 20680 12044 20686 12096
rect 21358 12044 21364 12096
rect 21416 12044 21422 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 4172 11852 4629 11880
rect 3789 11815 3847 11821
rect 3789 11781 3801 11815
rect 3835 11812 3847 11815
rect 4172 11812 4200 11852
rect 4617 11849 4629 11852
rect 4663 11880 4675 11883
rect 4663 11852 5120 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 3835 11784 4200 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4080 11608 4108 11707
rect 4172 11676 4200 11784
rect 4264 11784 4752 11812
rect 4264 11753 4292 11784
rect 4724 11756 4752 11784
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4172 11648 4353 11676
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4448 11676 4476 11707
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 4448 11648 4660 11676
rect 4341 11639 4399 11645
rect 4433 11611 4491 11617
rect 4433 11608 4445 11611
rect 4080 11580 4445 11608
rect 4433 11577 4445 11580
rect 4479 11577 4491 11611
rect 4433 11571 4491 11577
rect 4632 11552 4660 11648
rect 3878 11500 3884 11552
rect 3936 11500 3942 11552
rect 4614 11500 4620 11552
rect 4672 11500 4678 11552
rect 5092 11549 5120 11852
rect 20622 11840 20628 11892
rect 20680 11840 20686 11892
rect 6914 11772 6920 11824
rect 6972 11812 6978 11824
rect 10226 11812 10232 11824
rect 6972 11784 10232 11812
rect 6972 11772 6978 11784
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 19880 11815 19938 11821
rect 19880 11781 19892 11815
rect 19926 11812 19938 11815
rect 20640 11812 20668 11840
rect 19926 11784 20668 11812
rect 19926 11781 19938 11784
rect 19880 11775 19938 11781
rect 9125 11679 9183 11685
rect 9125 11645 9137 11679
rect 9171 11676 9183 11679
rect 9766 11676 9772 11688
rect 9171 11648 9772 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 10134 11636 10140 11688
rect 10192 11636 10198 11688
rect 11882 11636 11888 11688
rect 11940 11636 11946 11688
rect 12894 11636 12900 11688
rect 12952 11636 12958 11688
rect 14826 11636 14832 11688
rect 14884 11636 14890 11688
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 16206 11676 16212 11688
rect 15703 11648 16212 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 17494 11636 17500 11688
rect 17552 11636 17558 11688
rect 17770 11636 17776 11688
rect 17828 11676 17834 11688
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 17828 11648 19625 11676
rect 17828 11636 17834 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5258 11540 5264 11552
rect 5123 11512 5264 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 9674 11500 9680 11552
rect 9732 11500 9738 11552
rect 10686 11500 10692 11552
rect 10744 11500 10750 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12529 11543 12587 11549
rect 12529 11540 12541 11543
rect 11848 11512 12541 11540
rect 11848 11500 11854 11512
rect 12529 11509 12541 11512
rect 12575 11509 12587 11543
rect 12529 11503 12587 11509
rect 13538 11500 13544 11552
rect 13596 11500 13602 11552
rect 15470 11500 15476 11552
rect 15528 11500 15534 11552
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 16209 11543 16267 11549
rect 16209 11540 16221 11543
rect 15712 11512 16221 11540
rect 15712 11500 15718 11512
rect 16209 11509 16221 11512
rect 16255 11509 16267 11543
rect 16209 11503 16267 11509
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 18141 11543 18199 11549
rect 18141 11540 18153 11543
rect 17920 11512 18153 11540
rect 17920 11500 17926 11512
rect 18141 11509 18153 11512
rect 18187 11509 18199 11543
rect 18141 11503 18199 11509
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 20993 11543 21051 11549
rect 20993 11540 21005 11543
rect 20588 11512 21005 11540
rect 20588 11500 20594 11512
rect 20993 11509 21005 11512
rect 21039 11509 21051 11543
rect 20993 11503 21051 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 3936 11308 4200 11336
rect 3936 11296 3942 11308
rect 4172 11209 4200 11308
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4672 11308 5273 11336
rect 4672 11296 4678 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 5261 11299 5319 11305
rect 6914 11296 6920 11348
rect 6972 11296 6978 11348
rect 9674 11336 9680 11348
rect 9324 11308 9680 11336
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11169 4215 11203
rect 4157 11163 4215 11169
rect 4706 11160 4712 11212
rect 4764 11160 4770 11212
rect 4724 11132 4752 11160
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4724 11104 4905 11132
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 5258 11132 5264 11144
rect 5031 11104 5264 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 4908 11064 4936 11095
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 7282 11132 7288 11144
rect 5592 11104 7288 11132
rect 5592 11092 5598 11104
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 9324 11141 9352 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 10778 11336 10784 11348
rect 10284 11308 10784 11336
rect 10284 11296 10290 11308
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 11606 11336 11612 11348
rect 11204 11308 11612 11336
rect 11204 11296 11210 11308
rect 11606 11296 11612 11308
rect 11664 11336 11670 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 11664 11308 12357 11336
rect 11664 11296 11670 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12345 11299 12403 11305
rect 13446 11296 13452 11348
rect 13504 11296 13510 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 13872 11308 13921 11336
rect 13872 11296 13878 11308
rect 13909 11305 13921 11308
rect 13955 11305 13967 11339
rect 13909 11299 13967 11305
rect 14461 11339 14519 11345
rect 14461 11305 14473 11339
rect 14507 11336 14519 11339
rect 14826 11336 14832 11348
rect 14507 11308 14832 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 16666 11296 16672 11348
rect 16724 11296 16730 11348
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 19242 11336 19248 11348
rect 18656 11308 19248 11336
rect 18656 11296 18662 11308
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19978 11296 19984 11348
rect 20036 11296 20042 11348
rect 21358 11336 21364 11348
rect 20456 11308 21364 11336
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 9416 11240 10057 11268
rect 9416 11209 9444 11240
rect 10045 11237 10057 11240
rect 10091 11268 10103 11271
rect 10962 11268 10968 11280
rect 10091 11240 10968 11268
rect 10091 11237 10103 11240
rect 10045 11231 10103 11237
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 13464 11268 13492 11296
rect 14277 11271 14335 11277
rect 14277 11268 14289 11271
rect 13464 11240 14289 11268
rect 14277 11237 14289 11240
rect 14323 11237 14335 11271
rect 14277 11231 14335 11237
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9490 11160 9496 11212
rect 9548 11160 9554 11212
rect 14090 11160 14096 11212
rect 14148 11160 14154 11212
rect 14292 11200 14320 11231
rect 15105 11203 15163 11209
rect 14292 11172 14412 11200
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 10965 11135 11023 11141
rect 10965 11101 10977 11135
rect 11011 11132 11023 11135
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 11011 11104 12541 11132
rect 11011 11101 11023 11104
rect 10965 11095 11023 11101
rect 12529 11101 12541 11104
rect 12575 11132 12587 11135
rect 14108 11132 14136 11160
rect 12575 11104 14136 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 5442 11064 5448 11076
rect 4908 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5804 11067 5862 11073
rect 5804 11033 5816 11067
rect 5850 11064 5862 11067
rect 6178 11064 6184 11076
rect 5850 11036 6184 11064
rect 5850 11033 5862 11036
rect 5804 11027 5862 11033
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 7552 11067 7610 11073
rect 7552 11033 7564 11067
rect 7598 11064 7610 11067
rect 8294 11064 8300 11076
rect 7598 11036 8300 11064
rect 7598 11033 7610 11036
rect 7552 11027 7610 11033
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 9766 11064 9772 11076
rect 8680 11036 9772 11064
rect 4798 10956 4804 11008
rect 4856 10956 4862 11008
rect 5077 10999 5135 11005
rect 5077 10965 5089 10999
rect 5123 10996 5135 10999
rect 5166 10996 5172 11008
rect 5123 10968 5172 10996
rect 5123 10965 5135 10968
rect 5077 10959 5135 10965
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5353 10999 5411 11005
rect 5353 10965 5365 10999
rect 5399 10996 5411 10999
rect 5626 10996 5632 11008
rect 5399 10968 5632 10996
rect 5399 10965 5411 10968
rect 5353 10959 5411 10965
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 8680 11005 8708 11036
rect 9766 11024 9772 11036
rect 9824 11064 9830 11076
rect 10318 11064 10324 11076
rect 9824 11036 10324 11064
rect 9824 11024 9830 11036
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 11232 11067 11290 11073
rect 11232 11033 11244 11067
rect 11278 11064 11290 11067
rect 11790 11064 11796 11076
rect 11278 11036 11796 11064
rect 11278 11033 11290 11036
rect 11232 11027 11290 11033
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 12796 11067 12854 11073
rect 12796 11033 12808 11067
rect 12842 11064 12854 11067
rect 13538 11064 13544 11076
rect 12842 11036 13544 11064
rect 12842 11033 12854 11036
rect 12796 11027 12854 11033
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14384 11064 14412 11172
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15194 11200 15200 11212
rect 15151 11172 15200 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 20456 11209 20484 11308
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11169 20499 11203
rect 20441 11163 20499 11169
rect 20622 11160 20628 11212
rect 20680 11160 20686 11212
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 14976 11104 15301 11132
rect 14976 11092 14982 11104
rect 15289 11101 15301 11104
rect 15335 11132 15347 11135
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 15335 11104 17233 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 17221 11101 17233 11104
rect 17267 11132 17279 11135
rect 17770 11132 17776 11144
rect 17267 11104 17776 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 17862 11092 17868 11144
rect 17920 11092 17926 11144
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20404 11104 21005 11132
rect 20404 11092 20410 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 15562 11073 15568 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 14384 11036 14841 11064
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 14936 11036 15516 11064
rect 8665 10999 8723 11005
rect 8665 10965 8677 10999
rect 8711 10965 8723 10999
rect 8665 10959 8723 10965
rect 8938 10956 8944 11008
rect 8996 10956 9002 11008
rect 10870 10956 10876 11008
rect 10928 10956 10934 11008
rect 14936 11005 14964 11036
rect 14921 10999 14979 11005
rect 14921 10965 14933 10999
rect 14967 10965 14979 10999
rect 15488 10996 15516 11036
rect 15556 11027 15568 11073
rect 15562 11024 15568 11027
rect 15620 11024 15626 11076
rect 15654 11024 15660 11076
rect 15712 11024 15718 11076
rect 16574 11064 16580 11076
rect 16546 11024 16580 11064
rect 16632 11064 16638 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16632 11036 16957 11064
rect 16632 11024 16638 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 16945 11027 17003 11033
rect 17488 11067 17546 11073
rect 17488 11033 17500 11067
rect 17534 11064 17546 11067
rect 17880 11064 17908 11092
rect 17534 11036 17908 11064
rect 17534 11033 17546 11036
rect 17488 11027 17546 11033
rect 15672 10996 15700 11024
rect 15488 10968 15700 10996
rect 14921 10959 14979 10965
rect 16114 10956 16120 11008
rect 16172 10996 16178 11008
rect 16546 10996 16574 11024
rect 16172 10968 16574 10996
rect 16172 10956 16178 10968
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 6178 10752 6184 10804
rect 6236 10752 6242 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8352 10764 8953 10792
rect 8352 10752 8358 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10192 10764 10609 10792
rect 10192 10752 10198 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10928 10764 10977 10792
rect 10928 10752 10934 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11422 10752 11428 10804
rect 11480 10752 11486 10804
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10792 11575 10795
rect 11882 10792 11888 10804
rect 11563 10764 11888 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12544 10764 16160 10792
rect 5534 10724 5540 10736
rect 5092 10696 5540 10724
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 5092 10656 5120 10696
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 9392 10727 9450 10733
rect 9392 10693 9404 10727
rect 9438 10724 9450 10727
rect 10686 10724 10692 10736
rect 9438 10696 10692 10724
rect 9438 10693 9450 10696
rect 9392 10687 9450 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 2915 10628 5120 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 5166 10616 5172 10668
rect 5224 10616 5230 10668
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5316 10628 5365 10656
rect 5316 10616 5322 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5442 10616 5448 10668
rect 5500 10616 5506 10668
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 5994 10656 6000 10668
rect 5736 10628 6000 10656
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10588 3203 10591
rect 4798 10588 4804 10600
rect 3191 10560 4804 10588
rect 3191 10557 3203 10560
rect 3145 10551 3203 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5184 10588 5212 10616
rect 5736 10588 5764 10628
rect 5994 10616 6000 10628
rect 6052 10656 6058 10668
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 6052 10628 6653 10656
rect 6052 10616 6058 10628
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8938 10656 8944 10668
rect 8435 10628 8944 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 11440 10656 11468 10752
rect 12544 10733 12572 10764
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 12406 10696 12541 10724
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11440 10628 11897 10656
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 12406 10656 12434 10696
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 12529 10687 12587 10693
rect 15096 10727 15154 10733
rect 15096 10693 15108 10727
rect 15142 10724 15154 10727
rect 15470 10724 15476 10736
rect 15142 10696 15476 10724
rect 15142 10693 15154 10696
rect 15096 10687 15154 10693
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 16132 10724 16160 10764
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 17494 10752 17500 10804
rect 17552 10752 17558 10804
rect 17862 10724 17868 10736
rect 16132 10696 17868 10724
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 17957 10727 18015 10733
rect 17957 10693 17969 10727
rect 18003 10724 18015 10727
rect 18969 10727 19027 10733
rect 18969 10724 18981 10727
rect 18003 10696 18981 10724
rect 18003 10693 18015 10696
rect 17957 10687 18015 10693
rect 18969 10693 18981 10696
rect 19015 10693 19027 10727
rect 18969 10687 19027 10693
rect 11931 10628 12434 10656
rect 12989 10659 13047 10665
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13170 10656 13176 10668
rect 13035 10628 13176 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14737 10659 14795 10665
rect 14737 10656 14749 10659
rect 14148 10628 14749 10656
rect 14148 10616 14154 10628
rect 14737 10625 14749 10628
rect 14783 10656 14795 10659
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14783 10628 14841 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 14829 10625 14841 10628
rect 14875 10656 14887 10659
rect 14918 10656 14924 10668
rect 14875 10628 14924 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 16666 10616 16672 10668
rect 16724 10616 16730 10668
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 18598 10656 18604 10668
rect 18463 10628 18604 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 5184 10560 5764 10588
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10588 6423 10591
rect 6932 10588 6960 10616
rect 6411 10560 6960 10588
rect 9125 10591 9183 10597
rect 6411 10557 6423 10560
rect 6365 10551 6423 10557
rect 9125 10557 9137 10591
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 4433 10523 4491 10529
rect 4433 10489 4445 10523
rect 4479 10520 4491 10523
rect 4706 10520 4712 10532
rect 4479 10492 4712 10520
rect 4479 10489 4491 10492
rect 4433 10483 4491 10489
rect 4706 10480 4712 10492
rect 4764 10520 4770 10532
rect 4893 10523 4951 10529
rect 4893 10520 4905 10523
rect 4764 10492 4905 10520
rect 4764 10480 4770 10492
rect 4893 10489 4905 10492
rect 4939 10520 4951 10523
rect 5258 10520 5264 10532
rect 4939 10492 5264 10520
rect 4939 10489 4951 10492
rect 4893 10483 4951 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5350 10480 5356 10532
rect 5408 10480 5414 10532
rect 9140 10520 9168 10551
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 11020 10560 11069 10588
rect 11020 10548 11026 10560
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11330 10588 11336 10600
rect 11287 10560 11336 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 6380 10492 9168 10520
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 5368 10452 5396 10480
rect 6380 10464 6408 10492
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 11256 10520 11284 10551
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 11974 10548 11980 10600
rect 12032 10548 12038 10600
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 13538 10588 13544 10600
rect 12207 10560 13544 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 13538 10548 13544 10560
rect 13596 10548 13602 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 16408 10560 18061 10588
rect 10928 10492 11284 10520
rect 10928 10480 10934 10492
rect 5215 10424 5396 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10226 10452 10232 10464
rect 9824 10424 10232 10452
rect 9824 10412 9830 10424
rect 10226 10412 10232 10424
rect 10284 10452 10290 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10284 10424 10517 10452
rect 10284 10412 10290 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 16408 10452 16436 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 20530 10548 20536 10600
rect 20588 10548 20594 10600
rect 15252 10424 16436 10452
rect 15252 10412 15258 10424
rect 17310 10412 17316 10464
rect 17368 10412 17374 10464
rect 21174 10412 21180 10464
rect 21232 10412 21238 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 38378 10452 38384 10464
rect 21600 10424 38384 10452
rect 21600 10412 21606 10424
rect 38378 10412 38384 10424
rect 38436 10412 38442 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 4433 10251 4491 10257
rect 4433 10217 4445 10251
rect 4479 10248 4491 10251
rect 4706 10248 4712 10260
rect 4479 10220 4712 10248
rect 4479 10217 4491 10220
rect 4433 10211 4491 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 4890 10208 4896 10260
rect 4948 10208 4954 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6362 10248 6368 10260
rect 5592 10220 6368 10248
rect 5592 10208 5598 10220
rect 6362 10208 6368 10220
rect 6420 10248 6426 10260
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 6420 10220 6561 10248
rect 6420 10208 6426 10220
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9950 10248 9956 10260
rect 9364 10220 9956 10248
rect 9364 10208 9370 10220
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 12032 10220 12173 10248
rect 12032 10208 12038 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 12894 10208 12900 10260
rect 12952 10208 12958 10260
rect 13446 10208 13452 10260
rect 13504 10208 13510 10260
rect 17310 10248 17316 10260
rect 16224 10220 17316 10248
rect 12805 10183 12863 10189
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 13464 10180 13492 10208
rect 12851 10152 13492 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 11606 10072 11612 10124
rect 11664 10072 11670 10124
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4614 10044 4620 10056
rect 4571 10016 4620 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 9490 10004 9496 10056
rect 9548 10004 9554 10056
rect 13280 10053 13308 10152
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 16224 10121 16252 10220
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17862 10208 17868 10260
rect 17920 10248 17926 10260
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 17920 10220 18521 10248
rect 17920 10208 17926 10220
rect 18509 10217 18521 10220
rect 18555 10248 18567 10251
rect 20346 10248 20352 10260
rect 18555 10220 20352 10248
rect 18555 10217 18567 10220
rect 18509 10211 18567 10217
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20530 10208 20536 10260
rect 20588 10208 20594 10260
rect 21542 10248 21548 10260
rect 21192 10220 21548 10248
rect 20622 10180 20628 10192
rect 16316 10152 20628 10180
rect 16316 10124 16344 10152
rect 20622 10140 20628 10152
rect 20680 10180 20686 10192
rect 20680 10152 21128 10180
rect 20680 10140 20686 10152
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13872 10084 14105 10112
rect 13872 10072 13878 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 16298 10072 16304 10124
rect 16356 10072 16362 10124
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 20162 10112 20168 10124
rect 19935 10084 20168 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 20162 10072 20168 10084
rect 20220 10072 20226 10124
rect 21100 10121 21128 10152
rect 21085 10115 21143 10121
rect 21085 10081 21097 10115
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14829 10047 14887 10053
rect 14829 10044 14841 10047
rect 13964 10016 14841 10044
rect 13964 10004 13970 10016
rect 14829 10013 14841 10016
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 16758 10004 16764 10056
rect 16816 10004 16822 10056
rect 17678 10004 17684 10056
rect 17736 10004 17742 10056
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 19978 10044 19984 10056
rect 19751 10016 19984 10044
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 19978 10004 19984 10016
rect 20036 10044 20042 10056
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 20036 10016 20361 10044
rect 20036 10004 20042 10016
rect 20349 10013 20361 10016
rect 20395 10044 20407 10047
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20395 10016 20913 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20901 10013 20913 10016
rect 20947 10044 20959 10047
rect 21192 10044 21220 10220
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 20947 10016 21220 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 21358 10004 21364 10056
rect 21416 10004 21422 10056
rect 4893 9979 4951 9985
rect 4893 9945 4905 9979
rect 4939 9976 4951 9979
rect 5166 9976 5172 9988
rect 4939 9948 5172 9976
rect 4939 9945 4951 9948
rect 4893 9939 4951 9945
rect 5166 9936 5172 9948
rect 5224 9936 5230 9988
rect 5258 9936 5264 9988
rect 5316 9976 5322 9988
rect 13170 9976 13176 9988
rect 5316 9948 13176 9976
rect 5316 9936 5322 9948
rect 13170 9936 13176 9948
rect 13228 9936 13234 9988
rect 19613 9979 19671 9985
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 20162 9976 20168 9988
rect 19659 9948 20168 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 5077 9911 5135 9917
rect 5077 9877 5089 9911
rect 5123 9908 5135 9911
rect 5534 9908 5540 9920
rect 5123 9880 5540 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 10042 9868 10048 9920
rect 10100 9868 10106 9920
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 11020 9880 11345 9908
rect 11020 9868 11026 9880
rect 11333 9877 11345 9880
rect 11379 9877 11391 9911
rect 11333 9871 11391 9877
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 14737 9911 14795 9917
rect 14737 9908 14749 9911
rect 13403 9880 14749 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 14737 9877 14749 9880
rect 14783 9877 14795 9911
rect 14737 9871 14795 9877
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 14884 9880 15485 9908
rect 14884 9868 14890 9880
rect 15473 9877 15485 9880
rect 15519 9877 15531 9911
rect 15473 9871 15531 9877
rect 15746 9868 15752 9920
rect 15804 9868 15810 9920
rect 17034 9868 17040 9920
rect 17092 9908 17098 9920
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17092 9880 17417 9908
rect 17092 9868 17098 9880
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 18012 9880 18245 9908
rect 18012 9868 18018 9880
rect 18233 9877 18245 9880
rect 18279 9877 18291 9911
rect 18233 9871 18291 9877
rect 19245 9911 19303 9917
rect 19245 9877 19257 9911
rect 19291 9908 19303 9911
rect 19426 9908 19432 9920
rect 19291 9880 19432 9908
rect 19291 9877 19303 9880
rect 19245 9871 19303 9877
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 20993 9911 21051 9917
rect 20993 9877 21005 9911
rect 21039 9908 21051 9911
rect 22005 9911 22063 9917
rect 22005 9908 22017 9911
rect 21039 9880 22017 9908
rect 21039 9877 21051 9880
rect 20993 9871 21051 9877
rect 22005 9877 22017 9880
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5445 9707 5503 9713
rect 5445 9704 5457 9707
rect 4948 9676 5457 9704
rect 4948 9664 4954 9676
rect 5445 9673 5457 9676
rect 5491 9673 5503 9707
rect 5445 9667 5503 9673
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7248 9676 7757 9704
rect 7248 9664 7254 9676
rect 7745 9673 7757 9676
rect 7791 9704 7803 9707
rect 10594 9704 10600 9716
rect 7791 9676 10600 9704
rect 7791 9673 7803 9676
rect 7745 9667 7803 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 16758 9664 16764 9716
rect 16816 9664 16822 9716
rect 17788 9676 19288 9704
rect 17788 9648 17816 9676
rect 5350 9596 5356 9648
rect 5408 9636 5414 9648
rect 5902 9636 5908 9648
rect 5408 9608 5908 9636
rect 5408 9596 5414 9608
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 6380 9608 7972 9636
rect 6380 9580 6408 9608
rect 5534 9528 5540 9580
rect 5592 9528 5598 9580
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 7944 9577 7972 9608
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 13265 9639 13323 9645
rect 13265 9636 13277 9639
rect 13228 9608 13277 9636
rect 13228 9596 13234 9608
rect 13265 9605 13277 9608
rect 13311 9636 13323 9639
rect 13311 9608 15240 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 15212 9580 15240 9608
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 15620 9608 16313 9636
rect 15620 9596 15626 9608
rect 16301 9605 16313 9608
rect 16347 9605 16359 9639
rect 16301 9599 16359 9605
rect 17770 9596 17776 9648
rect 17828 9596 17834 9648
rect 19260 9636 19288 9676
rect 20162 9664 20168 9716
rect 20220 9664 20226 9716
rect 21358 9704 21364 9716
rect 20456 9676 21364 9704
rect 20456 9636 20484 9676
rect 21358 9664 21364 9676
rect 21416 9704 21422 9716
rect 21637 9707 21695 9713
rect 21637 9704 21649 9707
rect 21416 9676 21649 9704
rect 21416 9664 21422 9676
rect 21637 9673 21649 9676
rect 21683 9673 21695 9707
rect 21637 9667 21695 9673
rect 19260 9608 20484 9636
rect 20524 9639 20582 9645
rect 20524 9605 20536 9639
rect 20570 9636 20582 9639
rect 21174 9636 21180 9648
rect 20570 9608 21180 9636
rect 20570 9605 20582 9608
rect 20524 9599 20582 9605
rect 21174 9596 21180 9608
rect 21232 9596 21238 9648
rect 6621 9571 6679 9577
rect 6621 9568 6633 9571
rect 6472 9540 6633 9568
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 3970 9500 3976 9512
rect 3743 9472 3976 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4890 9460 4896 9512
rect 4948 9460 4954 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6472 9500 6500 9540
rect 6621 9537 6633 9540
rect 6667 9537 6679 9571
rect 6621 9531 6679 9537
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 8196 9571 8254 9577
rect 8196 9537 8208 9571
rect 8242 9568 8254 9571
rect 8754 9568 8760 9580
rect 8242 9540 8760 9568
rect 8242 9537 8254 9540
rect 8196 9531 8254 9537
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9568 9459 9571
rect 9766 9568 9772 9580
rect 9447 9540 9772 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9568 13415 9571
rect 13446 9568 13452 9580
rect 13403 9540 13452 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13624 9571 13682 9577
rect 13624 9537 13636 9571
rect 13670 9568 13682 9571
rect 14826 9568 14832 9580
rect 13670 9540 14832 9568
rect 13670 9537 13682 9540
rect 13624 9531 13682 9537
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 15746 9528 15752 9580
rect 15804 9528 15810 9580
rect 17129 9571 17187 9577
rect 17129 9537 17141 9571
rect 17175 9568 17187 9571
rect 17954 9568 17960 9580
rect 17175 9540 17960 9568
rect 17175 9537 17187 9540
rect 17129 9531 17187 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19852 9540 20269 9568
rect 19852 9528 19858 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 6227 9472 6500 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 9582 9460 9588 9512
rect 9640 9460 9646 9512
rect 10438 9503 10496 9509
rect 10438 9500 10450 9503
rect 9692 9472 10450 9500
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9490 9432 9496 9444
rect 9355 9404 9496 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9490 9392 9496 9404
rect 9548 9432 9554 9444
rect 9692 9432 9720 9472
rect 10438 9469 10450 9472
rect 10484 9469 10496 9503
rect 10438 9463 10496 9469
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 10778 9500 10784 9512
rect 10643 9472 10784 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 15010 9460 15016 9512
rect 15068 9460 15074 9512
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17405 9503 17463 9509
rect 17405 9469 17417 9503
rect 17451 9500 17463 9503
rect 17494 9500 17500 9512
rect 17451 9472 17500 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 9548 9404 9720 9432
rect 9548 9392 9554 9404
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 9950 9432 9956 9444
rect 9824 9404 9956 9432
rect 9824 9392 9830 9404
rect 9950 9392 9956 9404
rect 10008 9432 10014 9444
rect 10045 9435 10103 9441
rect 10045 9432 10057 9435
rect 10008 9404 10057 9432
rect 10008 9392 10014 9404
rect 10045 9401 10057 9404
rect 10091 9401 10103 9435
rect 10045 9395 10103 9401
rect 17236 9376 17264 9463
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 17589 9463 17647 9469
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 4249 9367 4307 9373
rect 4249 9364 4261 9367
rect 3660 9336 4261 9364
rect 3660 9324 3666 9336
rect 4249 9333 4261 9336
rect 4295 9333 4307 9367
rect 4249 9327 4307 9333
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5442 9364 5448 9376
rect 4764 9336 5448 9364
rect 4764 9324 4770 9336
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 11238 9324 11244 9376
rect 11296 9324 11302 9376
rect 14734 9324 14740 9376
rect 14792 9324 14798 9376
rect 15562 9324 15568 9376
rect 15620 9324 15626 9376
rect 17218 9324 17224 9376
rect 17276 9324 17282 9376
rect 17604 9364 17632 9463
rect 17678 9460 17684 9512
rect 17736 9460 17742 9512
rect 17770 9460 17776 9512
rect 17828 9460 17834 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 17972 9472 18521 9500
rect 17696 9432 17724 9460
rect 17972 9432 18000 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 18598 9460 18604 9512
rect 18656 9509 18662 9512
rect 18656 9503 18684 9509
rect 18672 9469 18684 9503
rect 18656 9463 18684 9469
rect 18656 9460 18662 9463
rect 18782 9460 18788 9512
rect 18840 9460 18846 9512
rect 19518 9500 19524 9512
rect 19260 9472 19524 9500
rect 17696 9404 18000 9432
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9432 18291 9435
rect 18322 9432 18328 9444
rect 18279 9404 18328 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 18322 9392 18328 9404
rect 18380 9392 18386 9444
rect 19260 9364 19288 9472
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 17604 9336 19288 9364
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 19392 9336 19441 9364
rect 19392 9324 19398 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 4948 9132 5641 9160
rect 4948 9120 4954 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 8754 9120 8760 9172
rect 8812 9120 8818 9172
rect 11238 9120 11244 9172
rect 11296 9120 11302 9172
rect 12805 9163 12863 9169
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 13906 9160 13912 9172
rect 12851 9132 13912 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 16117 9163 16175 9169
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16758 9160 16764 9172
rect 16163 9132 16764 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16758 9120 16764 9132
rect 16816 9160 16822 9172
rect 16816 9132 17448 9160
rect 16816 9120 16822 9132
rect 4614 9092 4620 9104
rect 3804 9064 4620 9092
rect 3804 8965 3832 9064
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5994 9092 6000 9104
rect 5040 9064 6000 9092
rect 5040 9052 5046 9064
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 8941 9095 8999 9101
rect 8941 9061 8953 9095
rect 8987 9061 8999 9095
rect 8941 9055 8999 9061
rect 4080 8996 5212 9024
rect 4080 8965 4108 8996
rect 5184 8968 5212 8996
rect 5350 8984 5356 9036
rect 5408 8984 5414 9036
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 6089 9027 6147 9033
rect 6089 9024 6101 9027
rect 5500 8996 6101 9024
rect 5500 8984 5506 8996
rect 6089 8993 6101 8996
rect 6135 9024 6147 9027
rect 7742 9024 7748 9036
rect 6135 8996 7748 9024
rect 6135 8993 6147 8996
rect 6089 8987 6147 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8956 9024 8984 9055
rect 8251 8996 8984 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 9214 8984 9220 9036
rect 9272 9024 9278 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 9272 8996 9505 9024
rect 9272 8984 9278 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10594 8984 10600 9036
rect 10652 8984 10658 9036
rect 11256 9024 11284 9120
rect 17420 9092 17448 9132
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 17865 9163 17923 9169
rect 17865 9160 17877 9163
rect 17736 9132 17877 9160
rect 17736 9120 17742 9132
rect 17865 9129 17877 9132
rect 17911 9129 17923 9163
rect 17865 9123 17923 9129
rect 18598 9120 18604 9172
rect 18656 9120 18662 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 20625 9163 20683 9169
rect 20625 9160 20637 9163
rect 19576 9132 20637 9160
rect 19576 9120 19582 9132
rect 20625 9129 20637 9132
rect 20671 9129 20683 9163
rect 20625 9123 20683 9129
rect 18616 9092 18644 9120
rect 17420 9064 18644 9092
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11256 8996 11989 9024
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 3973 8891 4031 8897
rect 3973 8857 3985 8891
rect 4019 8888 4031 8891
rect 4908 8888 4936 8919
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 5368 8956 5396 8984
rect 5626 8956 5632 8968
rect 5368 8928 5632 8956
rect 5626 8916 5632 8928
rect 5684 8956 5690 8968
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5684 8928 5825 8956
rect 5684 8916 5690 8928
rect 5813 8925 5825 8928
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 5902 8916 5908 8968
rect 5960 8916 5966 8968
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 10060 8956 10088 8984
rect 9447 8928 10088 8956
rect 10612 8956 10640 8984
rect 12084 8956 12112 8987
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13136 8996 13369 9024
rect 13136 8984 13142 8996
rect 13357 8993 13369 8996
rect 13403 9024 13415 9027
rect 13538 9024 13544 9036
rect 13403 8996 13544 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 10612 8928 12112 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 14737 8959 14795 8965
rect 14737 8956 14749 8959
rect 13504 8928 14749 8956
rect 13504 8916 13510 8928
rect 14737 8925 14749 8928
rect 14783 8956 14795 8959
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 14783 8928 16497 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 16485 8925 16497 8928
rect 16531 8956 16543 8959
rect 16574 8956 16580 8968
rect 16531 8928 16580 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16752 8959 16810 8965
rect 16752 8925 16764 8959
rect 16798 8956 16810 8959
rect 17034 8956 17040 8968
rect 16798 8928 17040 8956
rect 16798 8925 16810 8928
rect 16752 8919 16810 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 19116 8928 19257 8956
rect 19116 8916 19122 8928
rect 19245 8925 19257 8928
rect 19291 8956 19303 8959
rect 19794 8956 19800 8968
rect 19291 8928 19800 8956
rect 19291 8925 19303 8928
rect 19245 8919 19303 8925
rect 19794 8916 19800 8928
rect 19852 8916 19858 8968
rect 5350 8888 5356 8900
rect 4019 8860 5356 8888
rect 4019 8857 4031 8860
rect 3973 8851 4031 8857
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 5920 8888 5948 8916
rect 9309 8891 9367 8897
rect 5920 8860 6592 8888
rect 6564 8832 6592 8860
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 10045 8891 10103 8897
rect 10045 8888 10057 8891
rect 9355 8860 10057 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 10045 8857 10057 8860
rect 10091 8888 10103 8891
rect 10962 8888 10968 8900
rect 10091 8860 10968 8888
rect 10091 8857 10103 8860
rect 10045 8851 10103 8857
rect 10962 8848 10968 8860
rect 11020 8888 11026 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 11020 8860 13185 8888
rect 11020 8848 11026 8860
rect 13173 8857 13185 8860
rect 13219 8888 13231 8891
rect 15004 8891 15062 8897
rect 13219 8860 13952 8888
rect 13219 8857 13231 8860
rect 13173 8851 13231 8857
rect 3878 8780 3884 8832
rect 3936 8829 3942 8832
rect 3936 8783 3945 8829
rect 3936 8780 3942 8783
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 5132 8792 5549 8820
rect 5132 8780 5138 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 5537 8783 5595 8789
rect 6546 8780 6552 8832
rect 6604 8780 6610 8832
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 11388 8792 11529 8820
rect 11388 8780 11394 8792
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 11882 8780 11888 8832
rect 11940 8780 11946 8832
rect 13262 8780 13268 8832
rect 13320 8780 13326 8832
rect 13924 8829 13952 8860
rect 15004 8857 15016 8891
rect 15050 8888 15062 8891
rect 15562 8888 15568 8900
rect 15050 8860 15568 8888
rect 15050 8857 15062 8860
rect 15004 8851 15062 8857
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 19512 8891 19570 8897
rect 19512 8857 19524 8891
rect 19558 8888 19570 8891
rect 20070 8888 20076 8900
rect 19558 8860 20076 8888
rect 19558 8857 19570 8860
rect 19512 8851 19570 8857
rect 20070 8848 20076 8860
rect 20128 8848 20134 8900
rect 13909 8823 13967 8829
rect 13909 8789 13921 8823
rect 13955 8820 13967 8823
rect 17218 8820 17224 8832
rect 13955 8792 17224 8820
rect 13955 8789 13967 8792
rect 13909 8783 13967 8789
rect 17218 8780 17224 8792
rect 17276 8820 17282 8832
rect 18233 8823 18291 8829
rect 18233 8820 18245 8823
rect 17276 8792 18245 8820
rect 17276 8780 17282 8792
rect 18233 8789 18245 8792
rect 18279 8820 18291 8823
rect 19978 8820 19984 8832
rect 18279 8792 19984 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 3602 8576 3608 8628
rect 3660 8576 3666 8628
rect 3878 8576 3884 8628
rect 3936 8576 3942 8628
rect 3970 8576 3976 8628
rect 4028 8576 4034 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 4706 8576 4712 8628
rect 4764 8576 4770 8628
rect 4798 8576 4804 8628
rect 4856 8576 4862 8628
rect 4982 8576 4988 8628
rect 5040 8576 5046 8628
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5408 8588 5733 8616
rect 5408 8576 5414 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 9582 8576 9588 8628
rect 9640 8576 9646 8628
rect 11882 8576 11888 8628
rect 11940 8616 11946 8628
rect 11940 8588 12434 8616
rect 11940 8576 11946 8588
rect 3044 8551 3102 8557
rect 3044 8517 3056 8551
rect 3090 8548 3102 8551
rect 3620 8548 3648 8576
rect 3090 8520 3648 8548
rect 3090 8517 3102 8520
rect 3044 8511 3102 8517
rect 3896 8480 3924 8576
rect 3988 8548 4016 8576
rect 4249 8551 4307 8557
rect 4249 8548 4261 8551
rect 3988 8520 4261 8548
rect 4249 8517 4261 8520
rect 4295 8517 4307 8551
rect 4249 8511 4307 8517
rect 4433 8483 4491 8489
rect 4433 8480 4445 8483
rect 3896 8452 4445 8480
rect 4433 8449 4445 8452
rect 4479 8449 4491 8483
rect 4724 8480 4752 8576
rect 4816 8548 4844 8576
rect 4816 8520 5672 8548
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4724 8452 4813 8480
rect 4433 8443 4491 8449
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5644 8489 5672 8520
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 9600 8480 9628 8576
rect 12406 8548 12434 8588
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13909 8619 13967 8625
rect 13909 8616 13921 8619
rect 13320 8588 13921 8616
rect 13320 8576 13326 8588
rect 13909 8585 13921 8588
rect 13955 8585 13967 8619
rect 13909 8579 13967 8585
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 15068 8588 15117 8616
rect 15068 8576 15074 8588
rect 15105 8585 15117 8588
rect 15151 8585 15163 8619
rect 15105 8579 15163 8585
rect 15473 8619 15531 8625
rect 15473 8585 15485 8619
rect 15519 8616 15531 8619
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 15519 8588 16221 8616
rect 15519 8585 15531 8588
rect 15473 8579 15531 8585
rect 16209 8585 16221 8588
rect 16255 8616 16267 8619
rect 17218 8616 17224 8628
rect 16255 8588 17224 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 18322 8616 18328 8628
rect 17727 8588 18328 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 19334 8576 19340 8628
rect 19392 8576 19398 8628
rect 20070 8576 20076 8628
rect 20128 8576 20134 8628
rect 19352 8548 19380 8576
rect 12406 8520 19380 8548
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 9600 8452 13369 8480
rect 5629 8443 5687 8449
rect 13357 8449 13369 8452
rect 13403 8480 13415 8483
rect 14734 8480 14740 8492
rect 13403 8452 14740 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 17313 8483 17371 8489
rect 17313 8480 17325 8483
rect 15611 8452 17325 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 17313 8449 17325 8452
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 19426 8440 19432 8492
rect 19484 8440 19490 8492
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8381 2835 8415
rect 2777 8375 2835 8381
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 5092 8412 5120 8440
rect 4755 8384 5120 8412
rect 5169 8415 5227 8421
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5169 8381 5181 8415
rect 5215 8412 5227 8415
rect 5552 8412 5580 8440
rect 5215 8384 5580 8412
rect 8113 8415 8171 8421
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 8113 8381 8125 8415
rect 8159 8412 8171 8415
rect 8294 8412 8300 8424
rect 8159 8384 8300 8412
rect 8159 8381 8171 8384
rect 8113 8375 8171 8381
rect 1394 8236 1400 8288
rect 1452 8276 1458 8288
rect 2792 8276 2820 8375
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 5074 8344 5080 8356
rect 4663 8316 5080 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 5184 8288 5212 8375
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8846 8372 8852 8424
rect 8904 8372 8910 8424
rect 11606 8372 11612 8424
rect 11664 8372 11670 8424
rect 12250 8372 12256 8424
rect 12308 8372 12314 8424
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15657 8415 15715 8421
rect 15657 8412 15669 8415
rect 15344 8384 15669 8412
rect 15344 8372 15350 8384
rect 15657 8381 15669 8384
rect 15703 8381 15715 8415
rect 15657 8375 15715 8381
rect 16758 8372 16764 8424
rect 16816 8372 16822 8424
rect 20254 8372 20260 8424
rect 20312 8372 20318 8424
rect 5537 8347 5595 8353
rect 5537 8313 5549 8347
rect 5583 8344 5595 8347
rect 5626 8344 5632 8356
rect 5583 8316 5632 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 10778 8304 10784 8356
rect 10836 8344 10842 8356
rect 18782 8344 18788 8356
rect 10836 8316 18788 8344
rect 10836 8304 10842 8316
rect 18782 8304 18788 8316
rect 18840 8344 18846 8356
rect 19334 8344 19340 8356
rect 18840 8316 19340 8344
rect 18840 8304 18846 8316
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 1452 8248 2820 8276
rect 1452 8236 1458 8248
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 8662 8236 8668 8288
rect 8720 8236 8726 8288
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 12158 8236 12164 8288
rect 12216 8236 12222 8288
rect 12894 8236 12900 8288
rect 12952 8236 12958 8288
rect 20898 8236 20904 8288
rect 20956 8236 20962 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5166 8072 5172 8084
rect 5123 8044 5172 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5629 8075 5687 8081
rect 5629 8041 5641 8075
rect 5675 8072 5687 8075
rect 6546 8072 6552 8084
rect 5675 8044 6552 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 4890 8004 4896 8016
rect 4755 7976 4896 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 2682 7828 2688 7880
rect 2740 7828 2746 7880
rect 4816 7877 4844 7976
rect 4890 7964 4896 7976
rect 4948 8004 4954 8016
rect 5644 8004 5672 8035
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 12250 8072 12256 8084
rect 9416 8044 12256 8072
rect 4948 7976 5672 8004
rect 8757 8007 8815 8013
rect 4948 7964 4954 7976
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 8846 8004 8852 8016
rect 8803 7976 8852 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 8846 7964 8852 7976
rect 8904 8004 8910 8016
rect 8904 7976 9352 8004
rect 8904 7964 8910 7976
rect 4982 7896 4988 7948
rect 5040 7896 5046 7948
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5442 7868 5448 7880
rect 5123 7840 5448 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 7374 7868 7380 7880
rect 6512 7840 7380 7868
rect 6512 7828 6518 7840
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7644 7871 7702 7877
rect 7644 7837 7656 7871
rect 7690 7868 7702 7871
rect 8662 7868 8668 7880
rect 7690 7840 8668 7868
rect 7690 7837 7702 7840
rect 7644 7831 7702 7837
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9324 7868 9352 7976
rect 9416 7945 9444 8044
rect 12250 8032 12256 8044
rect 12308 8072 12314 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12308 8044 12541 8072
rect 12308 8032 12314 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 12529 8035 12587 8041
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 15286 8072 15292 8084
rect 15243 8044 15292 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18782 8072 18788 8084
rect 18380 8044 18788 8072
rect 18380 8032 18386 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 9508 7976 9996 8004
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 9508 7868 9536 7976
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9824 7908 9873 7936
rect 9824 7896 9830 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9968 7936 9996 7976
rect 13078 7964 13084 8016
rect 13136 7964 13142 8016
rect 10254 7939 10312 7945
rect 10254 7936 10266 7939
rect 9968 7908 10266 7936
rect 9861 7899 9919 7905
rect 10254 7905 10266 7908
rect 10300 7905 10312 7939
rect 10254 7899 10312 7905
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10778 7936 10784 7948
rect 10459 7908 10784 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 16025 7939 16083 7945
rect 13648 7908 15884 7936
rect 13648 7880 13676 7908
rect 9324 7840 9536 7868
rect 9217 7831 9275 7837
rect 3878 7760 3884 7812
rect 3936 7760 3942 7812
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 2556 7704 3249 7732
rect 2556 7692 2562 7704
rect 3237 7701 3249 7704
rect 3283 7701 3295 7735
rect 3237 7695 3295 7701
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 4982 7692 4988 7744
rect 5040 7732 5046 7744
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 5040 7704 5273 7732
rect 5040 7692 5046 7704
rect 5261 7701 5273 7704
rect 5307 7701 5319 7735
rect 9232 7732 9260 7831
rect 10134 7828 10140 7880
rect 10192 7828 10198 7880
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11416 7871 11474 7877
rect 11416 7837 11428 7871
rect 11462 7868 11474 7871
rect 12158 7868 12164 7880
rect 11462 7840 12164 7868
rect 11462 7837 11474 7840
rect 11416 7831 11474 7837
rect 11164 7744 11192 7831
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13630 7868 13636 7880
rect 13495 7840 13636 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13188 7800 13216 7831
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 15028 7877 15056 7908
rect 14921 7871 14979 7877
rect 14921 7837 14933 7871
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15470 7868 15476 7880
rect 15335 7840 15476 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 14936 7800 14964 7831
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15856 7877 15884 7908
rect 16025 7905 16037 7939
rect 16071 7936 16083 7939
rect 16298 7936 16304 7948
rect 16071 7908 16304 7936
rect 16071 7905 16083 7908
rect 16025 7899 16083 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 15102 7800 15108 7812
rect 13188 7772 15108 7800
rect 10042 7732 10048 7744
rect 9232 7704 10048 7732
rect 5261 7695 5319 7701
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 11054 7692 11060 7744
rect 11112 7692 11118 7744
rect 11146 7692 11152 7744
rect 11204 7692 11210 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13188 7732 13216 7772
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 12860 7704 13216 7732
rect 12860 7692 12866 7704
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15672 7732 15700 7831
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 17954 7828 17960 7880
rect 18012 7828 18018 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19889 7871 19947 7877
rect 19889 7868 19901 7871
rect 19116 7840 19901 7868
rect 19116 7828 19122 7840
rect 19889 7837 19901 7840
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20156 7871 20214 7877
rect 20156 7837 20168 7871
rect 20202 7868 20214 7871
rect 20898 7868 20904 7880
rect 20202 7840 20904 7868
rect 20202 7837 20214 7840
rect 20156 7831 20214 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21284 7840 21373 7868
rect 18322 7760 18328 7812
rect 18380 7800 18386 7812
rect 21284 7800 21312 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 18380 7772 21312 7800
rect 18380 7760 18386 7772
rect 14976 7704 15700 7732
rect 14976 7692 14982 7704
rect 17678 7692 17684 7744
rect 17736 7692 17742 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 21284 7741 21312 7772
rect 18509 7735 18567 7741
rect 18509 7732 18521 7735
rect 18104 7704 18521 7732
rect 18104 7692 18110 7704
rect 18509 7701 18521 7704
rect 18555 7701 18567 7735
rect 18509 7695 18567 7701
rect 21269 7735 21327 7741
rect 21269 7701 21281 7735
rect 21315 7701 21327 7735
rect 21269 7695 21327 7701
rect 22002 7692 22008 7744
rect 22060 7692 22066 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3243 7531 3301 7537
rect 3243 7528 3255 7531
rect 2740 7500 3255 7528
rect 2740 7488 2746 7500
rect 3243 7497 3255 7500
rect 3289 7497 3301 7531
rect 3243 7491 3301 7497
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3418 7528 3424 7540
rect 3375 7500 3424 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 3418 7488 3424 7500
rect 3476 7528 3482 7540
rect 3970 7528 3976 7540
rect 3476 7500 3976 7528
rect 3476 7488 3482 7500
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 4672 7500 4997 7528
rect 4672 7488 4678 7500
rect 4985 7497 4997 7500
rect 5031 7497 5043 7531
rect 4985 7491 5043 7497
rect 8294 7488 8300 7540
rect 8352 7488 8358 7540
rect 8757 7531 8815 7537
rect 8757 7497 8769 7531
rect 8803 7528 8815 7531
rect 9398 7528 9404 7540
rect 8803 7500 9404 7528
rect 8803 7497 8815 7500
rect 8757 7491 8815 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9766 7488 9772 7540
rect 9824 7488 9830 7540
rect 10134 7488 10140 7540
rect 10192 7488 10198 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11054 7528 11060 7540
rect 10735 7500 11060 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 11606 7528 11612 7540
rect 11563 7500 11612 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12894 7528 12900 7540
rect 12023 7500 12900 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 18012 7500 18061 7528
rect 18012 7488 18018 7500
rect 18049 7497 18061 7500
rect 18095 7528 18107 7531
rect 19150 7528 19156 7540
rect 18095 7500 19156 7528
rect 18095 7497 18107 7500
rect 18049 7491 18107 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 20254 7488 20260 7540
rect 20312 7488 20318 7540
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 22002 7528 22008 7540
rect 20763 7500 22008 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 6454 7460 6460 7472
rect 1688 7432 6460 7460
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 1688 7333 1716 7432
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 6546 7420 6552 7472
rect 6604 7460 6610 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 6604 7432 8217 7460
rect 6604 7420 6610 7432
rect 8205 7429 8217 7432
rect 8251 7460 8263 7463
rect 9784 7460 9812 7488
rect 8251 7432 9812 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 1940 7395 1998 7401
rect 1940 7361 1952 7395
rect 1986 7392 1998 7395
rect 2498 7392 2504 7404
rect 1986 7364 2504 7392
rect 1986 7361 1998 7364
rect 1940 7355 1998 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3467 7364 3556 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3528 7336 3556 7364
rect 3878 7352 3884 7404
rect 3936 7352 3942 7404
rect 4614 7352 4620 7404
rect 4672 7352 4678 7404
rect 4771 7395 4829 7401
rect 4771 7361 4783 7395
rect 4817 7392 4829 7395
rect 4982 7392 4988 7404
rect 4817 7364 4988 7392
rect 4817 7361 4829 7364
rect 4771 7355 4829 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6365 7395 6423 7401
rect 6043 7364 6316 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1452 7296 1685 7324
rect 1452 7284 1458 7296
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 3510 7284 3516 7336
rect 3568 7284 3574 7336
rect 3053 7259 3111 7265
rect 3053 7225 3065 7259
rect 3099 7256 3111 7259
rect 3896 7256 3924 7352
rect 3099 7228 3924 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 5500 7160 6193 7188
rect 5500 7148 5506 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 6288 7188 6316 7364
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6472 7392 6500 7420
rect 6411 7364 6500 7392
rect 6632 7395 6690 7401
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6632 7361 6644 7395
rect 6678 7392 6690 7395
rect 6914 7392 6920 7404
rect 6678 7364 6920 7392
rect 6678 7361 6690 7364
rect 6632 7355 6690 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 10152 7392 10180 7488
rect 10597 7463 10655 7469
rect 10597 7429 10609 7463
rect 10643 7460 10655 7463
rect 16936 7463 16994 7469
rect 10643 7432 16252 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 9364 7364 10180 7392
rect 9364 7352 9370 7364
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11296 7364 11897 7392
rect 11296 7352 11302 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7361 12495 7395
rect 12437 7355 12495 7361
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7392 12771 7395
rect 13081 7395 13139 7401
rect 12759 7364 12940 7392
rect 12759 7361 12771 7364
rect 12713 7355 12771 7361
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 8956 7256 8984 7287
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10652 7296 10793 7324
rect 10652 7284 10658 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7293 12219 7327
rect 12452 7324 12480 7355
rect 12802 7324 12808 7336
rect 12452 7296 12808 7324
rect 12161 7287 12219 7293
rect 9214 7256 9220 7268
rect 8956 7228 9220 7256
rect 9214 7216 9220 7228
rect 9272 7256 9278 7268
rect 12176 7256 12204 7287
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 12912 7324 12940 7364
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13630 7392 13636 7404
rect 13127 7364 13636 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 12986 7324 12992 7336
rect 12912 7296 12992 7324
rect 12986 7284 12992 7296
rect 13044 7324 13050 7336
rect 14366 7324 14372 7336
rect 13044 7296 14372 7324
rect 13044 7284 13050 7296
rect 14366 7284 14372 7296
rect 14424 7324 14430 7336
rect 15028 7324 15056 7355
rect 15102 7352 15108 7404
rect 15160 7392 15166 7404
rect 15197 7395 15255 7401
rect 15197 7392 15209 7395
rect 15160 7364 15209 7392
rect 15160 7352 15166 7364
rect 15197 7361 15209 7364
rect 15243 7392 15255 7395
rect 15378 7392 15384 7404
rect 15243 7364 15384 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 15488 7324 15516 7352
rect 14424 7296 15516 7324
rect 14424 7284 14430 7296
rect 13078 7256 13084 7268
rect 9272 7228 11376 7256
rect 12176 7228 13084 7256
rect 9272 7216 9278 7228
rect 6730 7188 6736 7200
rect 6288 7160 6736 7188
rect 6181 7151 6239 7157
rect 6730 7148 6736 7160
rect 6788 7188 6794 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 6788 7160 7757 7188
rect 6788 7148 6794 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 7745 7151 7803 7157
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 10226 7148 10232 7200
rect 10284 7148 10290 7200
rect 11238 7148 11244 7200
rect 11296 7148 11302 7200
rect 11348 7188 11376 7228
rect 13078 7216 13084 7228
rect 13136 7216 13142 7268
rect 12529 7191 12587 7197
rect 12529 7188 12541 7191
rect 11348 7160 12541 7188
rect 12529 7157 12541 7160
rect 12575 7157 12587 7191
rect 12529 7151 12587 7157
rect 14918 7148 14924 7200
rect 14976 7188 14982 7200
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14976 7160 15025 7188
rect 14976 7148 14982 7160
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 16224 7188 16252 7432
rect 16936 7429 16948 7463
rect 16982 7460 16994 7463
rect 17696 7460 17724 7488
rect 16982 7432 17724 7460
rect 16982 7429 16994 7432
rect 16936 7423 16994 7429
rect 18322 7352 18328 7404
rect 18380 7352 18386 7404
rect 19150 7352 19156 7404
rect 19208 7401 19214 7404
rect 19208 7395 19236 7401
rect 19224 7361 19236 7395
rect 19208 7355 19236 7361
rect 19208 7352 19214 7355
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 19978 7352 19984 7404
rect 20036 7392 20042 7404
rect 20625 7395 20683 7401
rect 20625 7392 20637 7395
rect 20036 7364 20637 7392
rect 20036 7352 20042 7364
rect 20625 7361 20637 7364
rect 20671 7392 20683 7395
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 20671 7364 21281 7392
rect 20671 7361 20683 7364
rect 20625 7355 20683 7361
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 18138 7284 18144 7336
rect 18196 7284 18202 7336
rect 18506 7284 18512 7336
rect 18564 7324 18570 7336
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18564 7296 19073 7324
rect 18564 7284 18570 7296
rect 19061 7293 19073 7296
rect 19107 7293 19119 7327
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 19061 7287 19119 7293
rect 20640 7296 20821 7324
rect 20640 7268 20668 7296
rect 20809 7293 20821 7296
rect 20855 7293 20867 7327
rect 20809 7287 20867 7293
rect 18782 7216 18788 7268
rect 18840 7216 18846 7268
rect 20622 7216 20628 7268
rect 20680 7216 20686 7268
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 16224 7160 19993 7188
rect 15013 7151 15071 7157
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 2869 6987 2927 6993
rect 2869 6953 2881 6987
rect 2915 6984 2927 6987
rect 3142 6984 3148 6996
rect 2915 6956 3148 6984
rect 2915 6953 2927 6956
rect 2869 6947 2927 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 6972 6956 7297 6984
rect 6972 6944 6978 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 15344 6956 16804 6984
rect 15344 6944 15350 6956
rect 2590 6876 2596 6928
rect 2648 6916 2654 6928
rect 4614 6916 4620 6928
rect 2648 6888 4620 6916
rect 2648 6876 2654 6888
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 9640 6888 9812 6916
rect 9640 6876 9646 6888
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5399 6820 5641 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 9490 6848 9496 6860
rect 8720 6820 9496 6848
rect 8720 6808 8726 6820
rect 9490 6808 9496 6820
rect 9548 6848 9554 6860
rect 9784 6857 9812 6888
rect 14918 6876 14924 6928
rect 14976 6916 14982 6928
rect 14976 6888 16712 6916
rect 14976 6876 14982 6888
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9548 6820 9689 6848
rect 9548 6808 9554 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6848 9827 6851
rect 9815 6820 9996 6848
rect 9815 6817 9827 6820
rect 9769 6811 9827 6817
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3418 6780 3424 6792
rect 3099 6752 3424 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 2884 6712 2912 6743
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 3510 6740 3516 6792
rect 3568 6740 3574 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 3528 6712 3556 6740
rect 2884 6684 3556 6712
rect 5276 6712 5304 6743
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 9585 6783 9643 6789
rect 8251 6752 9260 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 5552 6712 5580 6740
rect 5276 6684 5580 6712
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 8754 6604 8760 6656
rect 8812 6604 8818 6656
rect 9232 6653 9260 6752
rect 9585 6749 9597 6783
rect 9631 6780 9643 6783
rect 9858 6780 9864 6792
rect 9631 6752 9864 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 9968 6712 9996 6820
rect 10042 6808 10048 6860
rect 10100 6808 10106 6860
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 13998 6848 14004 6860
rect 11204 6820 14004 6848
rect 11204 6808 11210 6820
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14292 6820 15884 6848
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10376 6752 10793 6780
rect 10376 6740 10382 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 14292 6780 14320 6820
rect 14660 6792 14688 6820
rect 12768 6752 14320 6780
rect 12768 6740 12774 6752
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14642 6740 14648 6792
rect 14700 6740 14706 6792
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 15654 6740 15660 6792
rect 15712 6740 15718 6792
rect 15856 6789 15884 6820
rect 16684 6789 16712 6888
rect 16776 6848 16804 6956
rect 17126 6944 17132 6996
rect 17184 6944 17190 6996
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 20438 6984 20444 6996
rect 18196 6956 20444 6984
rect 18196 6944 18202 6956
rect 20438 6944 20444 6956
rect 20496 6944 20502 6996
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 16776 6820 17693 6848
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 17954 6808 17960 6860
rect 18012 6808 18018 6860
rect 18230 6808 18236 6860
rect 18288 6808 18294 6860
rect 18506 6808 18512 6860
rect 18564 6808 18570 6860
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17972 6780 18000 6808
rect 17635 6752 18000 6780
rect 18049 6783 18107 6789
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18138 6780 18144 6792
rect 18095 6752 18144 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 9968 6684 10824 6712
rect 10796 6656 10824 6684
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 10928 6684 14228 6712
rect 10928 6672 10934 6684
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6613 9275 6647
rect 9217 6607 9275 6613
rect 10686 6604 10692 6656
rect 10744 6604 10750 6656
rect 10778 6604 10784 6656
rect 10836 6604 10842 6656
rect 11422 6604 11428 6656
rect 11480 6604 11486 6656
rect 12434 6604 12440 6656
rect 12492 6604 12498 6656
rect 14200 6653 14228 6684
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6613 14243 6647
rect 15120 6644 15148 6740
rect 16132 6644 16160 6743
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 16393 6715 16451 6721
rect 16393 6681 16405 6715
rect 16439 6712 16451 6715
rect 20162 6712 20168 6724
rect 16439 6684 20168 6712
rect 16439 6681 16451 6684
rect 16393 6675 16451 6681
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 15120 6616 16160 6644
rect 14185 6607 14243 6613
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 17092 6616 17509 6644
rect 17092 6604 17098 6616
rect 17497 6613 17509 6616
rect 17543 6644 17555 6647
rect 17770 6644 17776 6656
rect 17543 6616 17776 6644
rect 17543 6613 17555 6616
rect 17497 6607 17555 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19061 6647 19119 6653
rect 19061 6644 19073 6647
rect 18564 6616 19073 6644
rect 18564 6604 18570 6616
rect 19061 6613 19073 6616
rect 19107 6613 19119 6647
rect 19061 6607 19119 6613
rect 20070 6604 20076 6656
rect 20128 6604 20134 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 6270 6400 6276 6452
rect 6328 6400 6334 6452
rect 6638 6400 6644 6452
rect 6696 6400 6702 6452
rect 8754 6400 8760 6452
rect 8812 6400 8818 6452
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9306 6440 9312 6452
rect 9171 6412 9312 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 10045 6443 10103 6449
rect 9548 6412 9674 6440
rect 9548 6400 9554 6412
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 5552 6344 5733 6372
rect 5552 6316 5580 6344
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 5626 6264 5632 6316
rect 5684 6264 5690 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6288 6304 6316 6400
rect 5951 6276 6316 6304
rect 6365 6307 6423 6313
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6454 6304 6460 6316
rect 6411 6276 6460 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 4672 6208 6009 6236
rect 4672 6196 4678 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6656 6236 6684 6400
rect 8012 6375 8070 6381
rect 8012 6341 8024 6375
rect 8058 6372 8070 6375
rect 8772 6372 8800 6400
rect 8058 6344 8800 6372
rect 9646 6372 9674 6412
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10318 6440 10324 6452
rect 10091 6412 10324 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10686 6440 10692 6452
rect 10459 6412 10692 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 10836 6412 12081 6440
rect 10836 6400 10842 6412
rect 12069 6409 12081 6412
rect 12115 6409 12127 6443
rect 12069 6403 12127 6409
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 17034 6440 17040 6452
rect 12492 6412 17040 6440
rect 12492 6400 12498 6412
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6409 17739 6443
rect 17681 6403 17739 6409
rect 18049 6443 18107 6449
rect 18049 6409 18061 6443
rect 18095 6440 18107 6443
rect 18506 6440 18512 6452
rect 18095 6412 18512 6440
rect 18095 6409 18107 6412
rect 18049 6403 18107 6409
rect 9769 6375 9827 6381
rect 9769 6372 9781 6375
rect 9646 6344 9781 6372
rect 8058 6341 8070 6344
rect 8012 6335 8070 6341
rect 9769 6341 9781 6344
rect 9815 6372 9827 6375
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 9815 6344 10517 6372
rect 9815 6341 9827 6344
rect 9769 6335 9827 6341
rect 10505 6341 10517 6344
rect 10551 6372 10563 6375
rect 11149 6375 11207 6381
rect 11149 6372 11161 6375
rect 10551 6344 11161 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 11149 6341 11161 6344
rect 11195 6372 11207 6375
rect 11238 6372 11244 6384
rect 11195 6344 11244 6372
rect 11195 6341 11207 6344
rect 11149 6335 11207 6341
rect 11238 6332 11244 6344
rect 11296 6372 11302 6384
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11296 6344 11805 6372
rect 11296 6332 11302 6344
rect 11793 6341 11805 6344
rect 11839 6372 11851 6375
rect 12452 6372 12480 6400
rect 12986 6372 12992 6384
rect 11839 6344 12480 6372
rect 12728 6344 12992 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7432 6276 7757 6304
rect 7432 6264 7438 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 7745 6267 7803 6273
rect 7852 6276 11989 6304
rect 7098 6236 7104 6248
rect 6135 6208 6684 6236
rect 6748 6208 7104 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6012 6168 6040 6199
rect 6748 6168 6776 6208
rect 7098 6196 7104 6208
rect 7156 6236 7162 6248
rect 7852 6236 7880 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 7156 6208 7880 6236
rect 10689 6239 10747 6245
rect 7156 6196 7162 6208
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 10870 6236 10876 6248
rect 10735 6208 10876 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 6012 6140 6776 6168
rect 11992 6168 12020 6267
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 12728 6313 12756 6344
rect 12986 6332 12992 6344
rect 13044 6372 13050 6384
rect 13262 6372 13268 6384
rect 13044 6344 13268 6372
rect 13044 6332 13050 6344
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 12124 6276 12265 6304
rect 12124 6264 12130 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12719 6307 12777 6313
rect 12719 6273 12731 6307
rect 12765 6273 12777 6307
rect 12719 6267 12777 6273
rect 12894 6264 12900 6316
rect 12952 6264 12958 6316
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 17037 6307 17095 6313
rect 14967 6276 16988 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12483 6208 12848 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12710 6168 12716 6180
rect 11992 6140 12716 6168
rect 12710 6128 12716 6140
rect 12768 6128 12774 6180
rect 6362 6060 6368 6112
rect 6420 6060 6426 6112
rect 12820 6109 12848 6208
rect 14660 6168 14688 6264
rect 15102 6196 15108 6248
rect 15160 6196 15166 6248
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6205 15255 6239
rect 15197 6199 15255 6205
rect 15212 6168 15240 6199
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 15470 6236 15476 6248
rect 15427 6208 15476 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 16960 6236 16988 6276
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17696 6304 17724 6403
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 20438 6400 20444 6452
rect 20496 6400 20502 6452
rect 17770 6332 17776 6384
rect 17828 6372 17834 6384
rect 18141 6375 18199 6381
rect 18141 6372 18153 6375
rect 17828 6344 18153 6372
rect 17828 6332 17834 6344
rect 18141 6341 18153 6344
rect 18187 6372 18199 6375
rect 19328 6375 19386 6381
rect 18187 6344 18828 6372
rect 18187 6341 18199 6344
rect 18141 6335 18199 6341
rect 18800 6313 18828 6344
rect 19328 6341 19340 6375
rect 19374 6372 19386 6375
rect 20088 6372 20116 6400
rect 19374 6344 20116 6372
rect 19374 6341 19386 6344
rect 19328 6335 19386 6341
rect 17083 6276 17724 6304
rect 18785 6307 18843 6313
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 18785 6273 18797 6307
rect 18831 6304 18843 6307
rect 19886 6304 19892 6316
rect 18831 6276 19892 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 20456 6304 20484 6400
rect 20533 6307 20591 6313
rect 20533 6304 20545 6307
rect 20456 6276 20545 6304
rect 20533 6273 20545 6276
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 18138 6236 18144 6248
rect 16960 6208 18144 6236
rect 18138 6196 18144 6208
rect 18196 6236 18202 6248
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 18196 6208 18245 6236
rect 18196 6196 18202 6208
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 19058 6196 19064 6248
rect 19116 6196 19122 6248
rect 14660 6140 15240 6168
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 12894 6100 12900 6112
rect 12851 6072 12900 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 15212 6100 15240 6140
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 19076 6168 19104 6196
rect 16724 6140 19104 6168
rect 16724 6128 16730 6140
rect 15286 6100 15292 6112
rect 15212 6072 15292 6100
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 17586 6060 17592 6112
rect 17644 6060 17650 6112
rect 21174 6060 21180 6112
rect 21232 6060 21238 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5350 5896 5356 5908
rect 5215 5868 5356 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7374 5896 7380 5908
rect 6779 5868 7380 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10192 5868 10885 5896
rect 10192 5856 10198 5868
rect 10873 5865 10885 5868
rect 10919 5865 10931 5899
rect 10873 5859 10931 5865
rect 11422 5856 11428 5908
rect 11480 5856 11486 5908
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15654 5896 15660 5908
rect 15611 5868 15660 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 18877 5899 18935 5905
rect 18877 5896 18889 5899
rect 18656 5868 18889 5896
rect 18656 5856 18662 5868
rect 18877 5865 18889 5868
rect 18923 5865 18935 5899
rect 18877 5859 18935 5865
rect 19426 5856 19432 5908
rect 19484 5856 19490 5908
rect 21174 5896 21180 5908
rect 19812 5868 21180 5896
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 5534 5828 5540 5840
rect 3568 5800 5540 5828
rect 3568 5788 3574 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 3418 5760 3424 5772
rect 2593 5723 2651 5729
rect 2700 5732 3424 5760
rect 2608 5624 2636 5723
rect 2700 5701 2728 5732
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 6546 5760 6552 5772
rect 4264 5732 6552 5760
rect 4264 5704 4292 5732
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 6604 5732 7113 5760
rect 6604 5720 6610 5732
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 7101 5723 7159 5729
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 2832 5664 3801 5692
rect 2832 5652 2838 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 4246 5652 4252 5704
rect 4304 5652 4310 5704
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 5166 5692 5172 5704
rect 4663 5664 5172 5692
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 5166 5652 5172 5664
rect 5224 5652 5230 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 11146 5692 11152 5704
rect 9539 5664 11152 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 3970 5624 3976 5636
rect 2608 5596 3976 5624
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 6472 5624 6500 5652
rect 7300 5624 7328 5655
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 6472 5596 7328 5624
rect 9760 5627 9818 5633
rect 9760 5593 9772 5627
rect 9806 5624 9818 5627
rect 11440 5624 11468 5856
rect 12986 5828 12992 5840
rect 11716 5800 12992 5828
rect 11716 5701 11744 5800
rect 12986 5788 12992 5800
rect 13044 5828 13050 5840
rect 13044 5800 13492 5828
rect 13044 5788 13050 5800
rect 11992 5732 13124 5760
rect 11992 5704 12020 5732
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 11974 5692 11980 5704
rect 11931 5664 11980 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12452 5624 12480 5655
rect 12710 5652 12716 5704
rect 12768 5652 12774 5704
rect 13096 5701 13124 5732
rect 13464 5701 13492 5800
rect 13630 5788 13636 5840
rect 13688 5788 13694 5840
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13449 5695 13507 5701
rect 13449 5661 13461 5695
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14185 5695 14243 5701
rect 14185 5692 14197 5695
rect 14056 5664 14197 5692
rect 14056 5652 14062 5664
rect 14185 5661 14197 5664
rect 14231 5692 14243 5695
rect 14231 5664 15148 5692
rect 14231 5661 14243 5664
rect 14185 5655 14243 5661
rect 9806 5596 11468 5624
rect 11716 5596 12480 5624
rect 14452 5627 14510 5633
rect 9806 5593 9818 5596
rect 9760 5587 9818 5593
rect 11716 5568 11744 5596
rect 14452 5593 14464 5627
rect 14498 5624 14510 5627
rect 15120 5624 15148 5664
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15657 5695 15715 5701
rect 15657 5692 15669 5695
rect 15252 5664 15669 5692
rect 15252 5652 15258 5664
rect 15657 5661 15669 5664
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 16666 5624 16672 5636
rect 14498 5596 15056 5624
rect 15120 5596 16672 5624
rect 14498 5593 14510 5596
rect 14452 5587 14510 5593
rect 3050 5516 3056 5568
rect 3108 5516 3114 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 4433 5559 4491 5565
rect 4433 5556 4445 5559
rect 4212 5528 4445 5556
rect 4212 5516 4218 5528
rect 4433 5525 4445 5528
rect 4479 5525 4491 5559
rect 4433 5519 4491 5525
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7469 5559 7527 5565
rect 7469 5556 7481 5559
rect 6972 5528 7481 5556
rect 6972 5516 6978 5528
rect 7469 5525 7481 5528
rect 7515 5525 7527 5559
rect 7469 5519 7527 5525
rect 11698 5516 11704 5568
rect 11756 5516 11762 5568
rect 11790 5516 11796 5568
rect 11848 5516 11854 5568
rect 15028 5556 15056 5596
rect 16666 5584 16672 5596
rect 16724 5624 16730 5636
rect 17512 5624 17540 5655
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 19812 5701 19840 5868
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 20441 5831 20499 5837
rect 20441 5828 20453 5831
rect 19904 5800 20453 5828
rect 19904 5772 19932 5800
rect 20441 5797 20453 5800
rect 20487 5797 20499 5831
rect 20441 5791 20499 5797
rect 19886 5720 19892 5772
rect 19944 5720 19950 5772
rect 20073 5763 20131 5769
rect 20073 5729 20085 5763
rect 20119 5760 20131 5763
rect 20162 5760 20168 5772
rect 20119 5732 20168 5760
rect 20119 5729 20131 5732
rect 20073 5723 20131 5729
rect 20162 5720 20168 5732
rect 20220 5720 20226 5772
rect 17753 5695 17811 5701
rect 17753 5692 17765 5695
rect 17644 5664 17765 5692
rect 17644 5652 17650 5664
rect 17753 5661 17765 5664
rect 17799 5661 17811 5695
rect 17753 5655 17811 5661
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 16724 5596 17540 5624
rect 20456 5624 20484 5791
rect 38197 5695 38255 5701
rect 38197 5661 38209 5695
rect 38243 5692 38255 5695
rect 38243 5664 38792 5692
rect 38243 5661 38255 5664
rect 38197 5655 38255 5661
rect 20456 5596 22094 5624
rect 16724 5584 16730 5596
rect 15378 5556 15384 5568
rect 15028 5528 15384 5556
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 16960 5565 16988 5596
rect 16945 5559 17003 5565
rect 16945 5525 16957 5559
rect 16991 5525 17003 5559
rect 22066 5556 22094 5596
rect 38764 5568 38792 5664
rect 38381 5559 38439 5565
rect 38381 5556 38393 5559
rect 22066 5528 38393 5556
rect 16945 5519 17003 5525
rect 38381 5525 38393 5528
rect 38427 5525 38439 5559
rect 38381 5519 38439 5525
rect 38746 5516 38752 5568
rect 38804 5516 38810 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3329 5355 3387 5361
rect 3329 5352 3341 5355
rect 3108 5324 3341 5352
rect 3108 5312 3114 5324
rect 3329 5321 3341 5324
rect 3375 5321 3387 5355
rect 3329 5315 3387 5321
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 3476 5324 4261 5352
rect 3476 5312 3482 5324
rect 4249 5321 4261 5324
rect 4295 5352 4307 5355
rect 4295 5324 4476 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 3237 5287 3295 5293
rect 3237 5253 3249 5287
rect 3283 5284 3295 5287
rect 4154 5284 4160 5296
rect 3283 5256 4160 5284
rect 3283 5253 3295 5256
rect 3237 5247 3295 5253
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 1664 5219 1722 5225
rect 1664 5185 1676 5219
rect 1710 5216 1722 5219
rect 2130 5216 2136 5228
rect 1710 5188 2136 5216
rect 1710 5185 1722 5188
rect 1664 5179 1722 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 4448 5225 4476 5324
rect 5442 5312 5448 5364
rect 5500 5312 5506 5364
rect 6362 5312 6368 5364
rect 6420 5312 6426 5364
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 14553 5355 14611 5361
rect 14553 5352 14565 5355
rect 12860 5324 14565 5352
rect 12860 5312 12866 5324
rect 14553 5321 14565 5324
rect 14599 5321 14611 5355
rect 14553 5315 14611 5321
rect 15378 5312 15384 5364
rect 15436 5312 15442 5364
rect 15654 5352 15660 5364
rect 15488 5324 15660 5352
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3804 5188 4077 5216
rect 3510 5108 3516 5160
rect 3568 5108 3574 5160
rect 3804 5024 3832 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 4663 5188 5365 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 5353 5185 5365 5188
rect 5399 5216 5411 5219
rect 5460 5216 5488 5312
rect 6380 5284 6408 5312
rect 6549 5287 6607 5293
rect 6549 5284 6561 5287
rect 6380 5256 6561 5284
rect 6549 5253 6561 5256
rect 6595 5253 6607 5287
rect 6549 5247 6607 5253
rect 6822 5244 6828 5296
rect 6880 5244 6886 5296
rect 5399 5188 5488 5216
rect 6365 5219 6423 5225
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6365 5185 6377 5219
rect 6411 5216 6423 5219
rect 6840 5216 6868 5244
rect 6411 5188 6868 5216
rect 11517 5219 11575 5225
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4246 5148 4252 5160
rect 3927 5120 4252 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 4356 5080 4384 5179
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 5132 5120 5273 5148
rect 5132 5108 5138 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 6733 5151 6791 5157
rect 6733 5148 6745 5151
rect 5684 5120 6745 5148
rect 5684 5108 5690 5120
rect 6733 5117 6745 5120
rect 6779 5117 6791 5151
rect 11532 5148 11560 5179
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11848 5188 11989 5216
rect 11848 5176 11854 5188
rect 11977 5185 11989 5188
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 15488 5216 15516 5324
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16485 5287 16543 5293
rect 16485 5284 16497 5287
rect 15580 5256 16497 5284
rect 15580 5225 15608 5256
rect 16485 5253 16497 5256
rect 16531 5253 16543 5287
rect 16485 5247 16543 5253
rect 14415 5188 15516 5216
rect 15565 5219 15623 5225
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 11532 5120 12434 5148
rect 6733 5111 6791 5117
rect 4890 5080 4896 5092
rect 4120 5052 4384 5080
rect 4448 5052 4896 5080
rect 4120 5040 4126 5052
rect 2866 4972 2872 5024
rect 2924 4972 2930 5024
rect 3786 4972 3792 5024
rect 3844 4972 3850 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4448 5021 4476 5052
rect 4890 5040 4896 5052
rect 4948 5040 4954 5092
rect 5721 5083 5779 5089
rect 5721 5049 5733 5083
rect 5767 5080 5779 5083
rect 6454 5080 6460 5092
rect 5767 5052 6460 5080
rect 5767 5049 5779 5052
rect 5721 5043 5779 5049
rect 6454 5040 6460 5052
rect 6512 5040 6518 5092
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 4212 4984 4445 5012
rect 4212 4972 4218 4984
rect 4433 4981 4445 4984
rect 4479 4981 4491 5015
rect 4433 4975 4491 4981
rect 4798 4972 4804 5024
rect 4856 4972 4862 5024
rect 11882 4972 11888 5024
rect 11940 4972 11946 5024
rect 12406 5012 12434 5120
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12584 5120 13093 5148
rect 12584 5108 12590 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15764 5148 15792 5179
rect 16666 5176 16672 5228
rect 16724 5176 16730 5228
rect 14884 5120 15792 5148
rect 14884 5108 14890 5120
rect 15838 5108 15844 5160
rect 15896 5108 15902 5160
rect 16942 5108 16948 5160
rect 17000 5108 17006 5160
rect 12618 5012 12624 5024
rect 12406 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 13722 4972 13728 5024
rect 13780 4972 13786 5024
rect 15562 4972 15568 5024
rect 15620 4972 15626 5024
rect 18046 4972 18052 5024
rect 18104 4972 18110 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2130 4768 2136 4820
rect 2188 4768 2194 4820
rect 2866 4808 2872 4820
rect 2746 4780 2872 4808
rect 2041 4743 2099 4749
rect 2041 4709 2053 4743
rect 2087 4740 2099 4743
rect 2746 4740 2774 4780
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3970 4768 3976 4820
rect 4028 4768 4034 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4120 4780 4261 4808
rect 4120 4768 4126 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4249 4771 4307 4777
rect 4356 4780 4905 4808
rect 2087 4712 2774 4740
rect 2087 4709 2099 4712
rect 2041 4703 2099 4709
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 2590 4672 2596 4684
rect 1728 4644 2596 4672
rect 1728 4632 1734 4644
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3943 4607 4001 4613
rect 3943 4573 3955 4607
rect 3989 4604 4001 4607
rect 4080 4604 4108 4768
rect 3989 4576 4108 4604
rect 3989 4573 4001 4576
rect 3943 4567 4001 4573
rect 3804 4536 3832 4564
rect 4356 4536 4384 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 11882 4768 11888 4820
rect 11940 4768 11946 4820
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13722 4808 13728 4820
rect 13403 4780 13728 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 14734 4768 14740 4820
rect 14792 4768 14798 4820
rect 15562 4768 15568 4820
rect 15620 4768 15626 4820
rect 15838 4768 15844 4820
rect 15896 4768 15902 4820
rect 16942 4768 16948 4820
rect 17000 4808 17006 4820
rect 17681 4811 17739 4817
rect 17681 4808 17693 4811
rect 17000 4780 17693 4808
rect 17000 4768 17006 4780
rect 17681 4777 17693 4780
rect 17727 4777 17739 4811
rect 17681 4771 17739 4777
rect 9769 4743 9827 4749
rect 4724 4712 5304 4740
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4604 4583 4607
rect 4614 4604 4620 4616
rect 4571 4576 4620 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 3804 4508 4384 4536
rect 4448 4536 4476 4567
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4724 4613 4752 4712
rect 4890 4632 4896 4684
rect 4948 4632 4954 4684
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 4908 4604 4936 4632
rect 5276 4613 5304 4712
rect 9769 4709 9781 4743
rect 9815 4740 9827 4743
rect 10226 4740 10232 4752
rect 9815 4712 10232 4740
rect 9815 4709 9827 4712
rect 9769 4703 9827 4709
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 6730 4632 6736 4684
rect 6788 4632 6794 4684
rect 11900 4672 11928 4768
rect 11974 4700 11980 4752
rect 12032 4740 12038 4752
rect 12710 4740 12716 4752
rect 12032 4712 12716 4740
rect 12032 4700 12038 4712
rect 12710 4700 12716 4712
rect 12768 4700 12774 4752
rect 13541 4743 13599 4749
rect 13541 4709 13553 4743
rect 13587 4740 13599 4743
rect 14752 4740 14780 4768
rect 13587 4712 14780 4740
rect 15580 4740 15608 4768
rect 15580 4712 17080 4740
rect 13587 4709 13599 4712
rect 13541 4703 13599 4709
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 11900 4644 12265 4672
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12253 4635 12311 4641
rect 12406 4644 13001 4672
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 4847 4576 5089 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 6917 4607 6975 4613
rect 5399 4576 5488 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 5276 4536 5304 4567
rect 5460 4548 5488 4576
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7558 4604 7564 4616
rect 6963 4576 7564 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9490 4604 9496 4616
rect 9447 4576 9496 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9490 4564 9496 4576
rect 9548 4604 9554 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 9548 4576 10425 4604
rect 9548 4564 9554 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 11238 4564 11244 4616
rect 11296 4564 11302 4616
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12406 4604 12434 4644
rect 12989 4641 13001 4644
rect 13035 4672 13047 4675
rect 15102 4672 15108 4684
rect 13035 4644 14228 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 14200 4616 14228 4644
rect 14292 4644 15108 4672
rect 11664 4576 12434 4604
rect 11664 4564 11670 4576
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13596 4576 14105 4604
rect 13596 4564 13602 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 14182 4564 14188 4616
rect 14240 4564 14246 4616
rect 4448 4508 4844 4536
rect 5276 4508 5396 4536
rect 4816 4480 4844 4508
rect 5368 4480 5396 4508
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 8113 4539 8171 4545
rect 5500 4508 7972 4536
rect 5500 4496 5506 4508
rect 7944 4480 7972 4508
rect 8113 4505 8125 4539
rect 8159 4536 8171 4539
rect 9214 4536 9220 4548
rect 8159 4508 9220 4536
rect 8159 4505 8171 4508
rect 8113 4499 8171 4505
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 11974 4536 11980 4548
rect 10612 4508 11980 4536
rect 10612 4480 10640 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 12066 4496 12072 4548
rect 12124 4536 12130 4548
rect 14292 4536 14320 4644
rect 15102 4632 15108 4644
rect 15160 4672 15166 4684
rect 17052 4681 17080 4712
rect 15381 4675 15439 4681
rect 15381 4672 15393 4675
rect 15160 4644 15393 4672
rect 15160 4632 15166 4644
rect 15381 4641 15393 4644
rect 15427 4641 15439 4675
rect 15381 4635 15439 4641
rect 17037 4675 17095 4681
rect 17037 4641 17049 4675
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 15470 4564 15476 4616
rect 15528 4604 15534 4616
rect 18046 4604 18052 4616
rect 15528 4576 18052 4604
rect 15528 4564 15534 4576
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 12124 4508 14320 4536
rect 12124 4496 12130 4508
rect 4798 4428 4804 4480
rect 4856 4428 4862 4480
rect 5350 4428 5356 4480
rect 5408 4428 5414 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 7064 4440 7113 4468
rect 7064 4428 7070 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 7101 4431 7159 4437
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 7984 4440 8217 4468
rect 7984 4428 7990 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 9858 4428 9864 4480
rect 9916 4428 9922 4480
rect 10594 4428 10600 4480
rect 10652 4428 10658 4480
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 11020 4440 11805 4468
rect 11020 4428 11026 4440
rect 11793 4437 11805 4440
rect 11839 4437 11851 4471
rect 11793 4431 11851 4437
rect 12526 4428 12532 4480
rect 12584 4468 12590 4480
rect 12897 4471 12955 4477
rect 12897 4468 12909 4471
rect 12584 4440 12909 4468
rect 12584 4428 12590 4440
rect 12897 4437 12909 4440
rect 12943 4437 12955 4471
rect 12897 4431 12955 4437
rect 13354 4428 13360 4480
rect 13412 4428 13418 4480
rect 14292 4477 14320 4508
rect 14277 4471 14335 4477
rect 14277 4437 14289 4471
rect 14323 4437 14335 4471
rect 14277 4431 14335 4437
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 7006 4264 7012 4276
rect 6564 4236 7012 4264
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5350 4128 5356 4140
rect 5215 4100 5356 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 6564 4137 6592 4236
rect 7006 4224 7012 4236
rect 7064 4264 7070 4276
rect 7190 4264 7196 4276
rect 7064 4236 7196 4264
rect 7064 4224 7070 4236
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7653 4267 7711 4273
rect 7653 4264 7665 4267
rect 7340 4236 7665 4264
rect 7340 4224 7346 4236
rect 7653 4233 7665 4236
rect 7699 4233 7711 4267
rect 7653 4227 7711 4233
rect 9214 4224 9220 4276
rect 9272 4224 9278 4276
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11296 4236 12173 4264
rect 11296 4224 11302 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14240 4236 14749 4264
rect 14240 4224 14246 4236
rect 14737 4233 14749 4236
rect 14783 4264 14795 4267
rect 14826 4264 14832 4276
rect 14783 4236 14832 4264
rect 14783 4233 14795 4236
rect 14737 4227 14795 4233
rect 14826 4224 14832 4236
rect 14884 4224 14890 4276
rect 7742 4196 7748 4208
rect 6748 4168 7748 4196
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6748 4137 6776 4168
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 8036 4168 8248 4196
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6696 4100 6745 4128
rect 6696 4088 6702 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7432 4100 7849 4128
rect 7432 4088 7438 4100
rect 7837 4097 7849 4100
rect 7883 4128 7895 4131
rect 8036 4128 8064 4168
rect 8110 4137 8116 4140
rect 7883 4100 8064 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8104 4091 8116 4137
rect 8110 4088 8116 4091
rect 8168 4088 8174 4140
rect 8220 4128 8248 4168
rect 10962 4156 10968 4208
rect 11020 4156 11026 4208
rect 11977 4199 12035 4205
rect 11977 4165 11989 4199
rect 12023 4196 12035 4199
rect 12066 4196 12072 4208
rect 12023 4168 12072 4196
rect 12023 4165 12035 4168
rect 11977 4159 12035 4165
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 12618 4196 12624 4208
rect 12452 4168 12624 4196
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 8220 4100 9873 4128
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 10128 4131 10186 4137
rect 10128 4097 10140 4131
rect 10174 4128 10186 4131
rect 10980 4128 11008 4156
rect 10174 4100 11008 4128
rect 10174 4097 10186 4100
rect 10128 4091 10186 4097
rect 11606 4088 11612 4140
rect 11664 4088 11670 4140
rect 12452 4137 12480 4168
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 12894 4156 12900 4208
rect 12952 4156 12958 4208
rect 13541 4199 13599 4205
rect 13541 4196 13553 4199
rect 13188 4168 13553 4196
rect 13188 4140 13216 4168
rect 13541 4165 13553 4168
rect 13587 4196 13599 4199
rect 13587 4168 14872 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12575 4100 13124 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 4614 4020 4620 4072
rect 4672 4060 4678 4072
rect 4982 4060 4988 4072
rect 4672 4032 4988 4060
rect 4672 4020 4678 4032
rect 4982 4020 4988 4032
rect 5040 4060 5046 4072
rect 7101 4063 7159 4069
rect 5040 4032 5488 4060
rect 5040 4020 5046 4032
rect 5460 4004 5488 4032
rect 6748 4032 6960 4060
rect 6748 4004 6776 4032
rect 2590 3952 2596 4004
rect 2648 3992 2654 4004
rect 3050 3992 3056 4004
rect 2648 3964 3056 3992
rect 2648 3952 2654 3964
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 5442 3952 5448 4004
rect 5500 3952 5506 4004
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 6641 3995 6699 4001
rect 5592 3964 6500 3992
rect 5592 3952 5598 3964
rect 5074 3884 5080 3936
rect 5132 3884 5138 3936
rect 6362 3884 6368 3936
rect 6420 3884 6426 3936
rect 6472 3924 6500 3964
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 6730 3992 6736 4004
rect 6687 3964 6736 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 6932 3992 6960 4032
rect 7101 4029 7113 4063
rect 7147 4060 7159 4063
rect 7742 4060 7748 4072
rect 7147 4032 7748 4060
rect 7147 4029 7159 4032
rect 7101 4023 7159 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 12544 4060 12572 4091
rect 11716 4032 12572 4060
rect 12621 4063 12679 4069
rect 11716 4004 11744 4032
rect 12621 4029 12633 4063
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 12802 4060 12808 4072
rect 12759 4032 12808 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 7374 3992 7380 4004
rect 6932 3964 7380 3992
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 7558 3952 7564 4004
rect 7616 3992 7622 4004
rect 11241 3995 11299 4001
rect 7616 3964 7788 3992
rect 7616 3952 7622 3964
rect 6822 3924 6828 3936
rect 6472 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3924 6886 3936
rect 7466 3924 7472 3936
rect 6880 3896 7472 3924
rect 6880 3884 6886 3896
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7760 3924 7788 3964
rect 11241 3961 11253 3995
rect 11287 3992 11299 3995
rect 11698 3992 11704 4004
rect 11287 3964 11704 3992
rect 11287 3961 11299 3964
rect 11241 3955 11299 3961
rect 11698 3952 11704 3964
rect 11756 3952 11762 4004
rect 12526 3992 12532 4004
rect 11992 3964 12532 3992
rect 10134 3924 10140 3936
rect 7760 3896 10140 3924
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 11992 3933 12020 3964
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12636 3992 12664 4023
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12986 4020 12992 4072
rect 13044 4020 13050 4072
rect 13096 4060 13124 4100
rect 13170 4088 13176 4140
rect 13228 4088 13234 4140
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 14369 4131 14427 4137
rect 14369 4097 14381 4131
rect 14415 4128 14427 4131
rect 14550 4128 14556 4140
rect 14415 4100 14556 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 13464 4060 13492 4091
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 14844 4134 14872 4168
rect 15102 4156 15108 4208
rect 15160 4196 15166 4208
rect 15160 4168 15424 4196
rect 15160 4156 15166 4168
rect 15013 4134 15071 4137
rect 14844 4131 15071 4134
rect 14691 4100 14780 4128
rect 14844 4106 15025 4131
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 13096 4032 13492 4060
rect 14752 4060 14780 4100
rect 15013 4097 15025 4106
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4126 15255 4131
rect 15286 4126 15292 4140
rect 15243 4098 15292 4126
rect 15243 4097 15255 4098
rect 15197 4091 15255 4097
rect 15286 4088 15292 4098
rect 15344 4088 15350 4140
rect 15396 4137 15424 4168
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4128 15439 4131
rect 16758 4128 16764 4140
rect 15427 4100 16764 4128
rect 15427 4097 15439 4100
rect 15381 4091 15439 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 14752 4032 14872 4060
rect 13262 3992 13268 4004
rect 12636 3964 13268 3992
rect 13262 3952 13268 3964
rect 13320 3952 13326 4004
rect 13354 3952 13360 4004
rect 13412 3992 13418 4004
rect 14844 3992 14872 4032
rect 14918 4020 14924 4072
rect 14976 4020 14982 4072
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 13412 3964 14320 3992
rect 14844 3964 15516 3992
rect 13412 3952 13418 3964
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3893 12035 3927
rect 11977 3887 12035 3893
rect 12253 3927 12311 3933
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 12342 3924 12348 3936
rect 12299 3896 12348 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12768 3896 12909 3924
rect 12768 3884 12774 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 14182 3884 14188 3936
rect 14240 3884 14246 3936
rect 14292 3924 14320 3964
rect 15488 3936 15516 3964
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 14292 3896 14565 3924
rect 14553 3893 14565 3896
rect 14599 3924 14611 3927
rect 15286 3924 15292 3936
rect 14599 3896 15292 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15470 3884 15476 3936
rect 15528 3884 15534 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 6362 3680 6368 3732
rect 6420 3680 6426 3732
rect 7208 3692 7512 3720
rect 4433 3655 4491 3661
rect 4433 3621 4445 3655
rect 4479 3652 4491 3655
rect 5166 3652 5172 3664
rect 4479 3624 5172 3652
rect 4479 3621 4491 3624
rect 4433 3615 4491 3621
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5534 3612 5540 3664
rect 5592 3612 5598 3664
rect 1670 3544 1676 3596
rect 1728 3544 1734 3596
rect 4706 3584 4712 3596
rect 2700 3556 4712 3584
rect 1026 3476 1032 3528
rect 1084 3516 1090 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1084 3488 1409 3516
rect 1084 3476 1090 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1762 3476 1768 3528
rect 1820 3516 1826 3528
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 1820 3488 2145 3516
rect 1820 3476 1826 3488
rect 2133 3485 2145 3488
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2406 3476 2412 3528
rect 2464 3476 2470 3528
rect 2700 3525 2728 3556
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 5092 3556 6101 3584
rect 5092 3528 5120 3556
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 6089 3547 6147 3553
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 2778 3519 2836 3525
rect 2778 3485 2790 3519
rect 2824 3485 2836 3519
rect 2778 3479 2836 3485
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 2792 3448 2820 3479
rect 3602 3476 3608 3528
rect 3660 3476 3666 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 2096 3420 2820 3448
rect 3053 3451 3111 3457
rect 2096 3408 2102 3420
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 2130 3380 2136 3392
rect 1995 3352 2136 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 2240 3389 2268 3420
rect 3053 3417 3065 3451
rect 3099 3448 3111 3451
rect 4062 3448 4068 3460
rect 3099 3420 4068 3448
rect 3099 3417 3111 3420
rect 3053 3411 3111 3417
rect 4062 3408 4068 3420
rect 4120 3408 4126 3460
rect 4632 3448 4660 3479
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5442 3476 5448 3528
rect 5500 3476 5506 3528
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 6380 3516 6408 3680
rect 7208 3652 7236 3692
rect 7484 3661 7512 3692
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 7800 3692 7972 3720
rect 7800 3680 7806 3692
rect 6840 3624 7236 3652
rect 7469 3655 7527 3661
rect 6840 3525 6868 3624
rect 7469 3621 7481 3655
rect 7515 3621 7527 3655
rect 7834 3652 7840 3664
rect 7469 3615 7527 3621
rect 7576 3624 7840 3652
rect 7098 3544 7104 3596
rect 7156 3544 7162 3596
rect 7190 3544 7196 3596
rect 7248 3544 7254 3596
rect 7576 3593 7604 3624
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3584 7803 3587
rect 7944 3584 7972 3692
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8168 3692 8769 3720
rect 8168 3680 8174 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 12529 3723 12587 3729
rect 12529 3720 12541 3723
rect 8757 3683 8815 3689
rect 10060 3692 12541 3720
rect 7791 3556 7972 3584
rect 7791 3553 7803 3556
rect 7745 3547 7803 3553
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6380 3488 6745 3516
rect 5997 3479 6055 3485
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3485 6883 3519
rect 6825 3479 6883 3485
rect 5368 3448 5396 3476
rect 4632 3420 5396 3448
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 3418 3340 3424 3392
rect 3476 3340 3482 3392
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 6012 3380 6040 3479
rect 7006 3476 7012 3528
rect 7064 3476 7070 3528
rect 7208 3516 7236 3544
rect 7286 3519 7344 3525
rect 7286 3516 7298 3519
rect 7208 3488 7298 3516
rect 7286 3485 7298 3488
rect 7332 3485 7344 3519
rect 7286 3479 7344 3485
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 7524 3488 7665 3516
rect 7524 3476 7530 3488
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 7926 3516 7932 3528
rect 7883 3488 7932 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 10060 3516 10088 3692
rect 12529 3689 12541 3692
rect 12575 3689 12587 3723
rect 12529 3683 12587 3689
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13538 3720 13544 3732
rect 13035 3692 13544 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14240 3692 14320 3720
rect 14240 3680 14246 3692
rect 10134 3612 10140 3664
rect 10192 3652 10198 3664
rect 12894 3652 12900 3664
rect 10192 3624 12900 3652
rect 10192 3612 10198 3624
rect 12636 3593 12664 3624
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 14292 3593 14320 3692
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14608 3692 15025 3720
rect 14608 3680 14614 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15013 3683 15071 3689
rect 16025 3723 16083 3729
rect 16025 3689 16037 3723
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 16040 3652 16068 3683
rect 16758 3680 16764 3732
rect 16816 3680 16822 3732
rect 14568 3624 16068 3652
rect 16316 3624 22094 3652
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 13081 3587 13139 3593
rect 12667 3556 12701 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 14277 3587 14335 3593
rect 13127 3556 14228 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 8113 3479 8171 3485
rect 9876 3488 10088 3516
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 8128 3448 8156 3479
rect 7239 3420 8156 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 9876 3392 9904 3488
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 12805 3519 12863 3525
rect 10468 3488 12756 3516
rect 10468 3476 10474 3488
rect 11330 3448 11336 3460
rect 10428 3420 11336 3448
rect 6914 3380 6920 3392
rect 5224 3352 6920 3380
rect 5224 3340 5230 3352
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 9858 3380 9864 3392
rect 7156 3352 9864 3380
rect 7156 3340 7162 3352
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 10428 3380 10456 3420
rect 11330 3408 11336 3420
rect 11388 3408 11394 3460
rect 12526 3408 12532 3460
rect 12584 3408 12590 3460
rect 12728 3448 12756 3488
rect 12805 3485 12817 3519
rect 12851 3516 12863 3519
rect 13170 3516 13176 3528
rect 12851 3488 13176 3516
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 14200 3516 14228 3556
rect 14277 3553 14289 3587
rect 14323 3553 14335 3587
rect 14277 3547 14335 3553
rect 14568 3516 14596 3624
rect 16114 3544 16120 3596
rect 16172 3544 16178 3596
rect 14200 3488 14596 3516
rect 14936 3488 15240 3516
rect 13357 3479 13415 3485
rect 13372 3448 13400 3479
rect 14936 3448 14964 3488
rect 12728 3420 14964 3448
rect 15010 3408 15016 3460
rect 15068 3408 15074 3460
rect 15212 3448 15240 3488
rect 15286 3476 15292 3528
rect 15344 3476 15350 3528
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 15473 3519 15531 3525
rect 15473 3516 15485 3519
rect 15436 3488 15485 3516
rect 15436 3476 15442 3488
rect 15473 3485 15485 3488
rect 15519 3516 15531 3519
rect 16206 3516 16212 3528
rect 15519 3488 16212 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 16316 3448 16344 3624
rect 20162 3584 20168 3596
rect 15212 3420 16344 3448
rect 17052 3556 20168 3584
rect 10376 3352 10456 3380
rect 10376 3340 10382 3352
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 14826 3380 14832 3392
rect 10560 3352 14832 3380
rect 10560 3340 10566 3352
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 14918 3340 14924 3392
rect 14976 3340 14982 3392
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 15470 3380 15476 3392
rect 15243 3352 15476 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 17052 3389 17080 3556
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 19334 3476 19340 3528
rect 19392 3476 19398 3528
rect 17037 3383 17095 3389
rect 17037 3380 17049 3383
rect 15712 3352 17049 3380
rect 15712 3340 15718 3352
rect 17037 3349 17049 3352
rect 17083 3349 17095 3383
rect 17037 3343 17095 3349
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 17644 3352 19901 3380
rect 17644 3340 17650 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 22066 3380 22094 3624
rect 32122 3584 32128 3596
rect 28460 3556 32128 3584
rect 28074 3476 28080 3528
rect 28132 3476 28138 3528
rect 28460 3460 28488 3556
rect 32122 3544 32128 3556
rect 32180 3544 32186 3596
rect 28442 3408 28448 3460
rect 28500 3408 28506 3460
rect 28534 3408 28540 3460
rect 28592 3448 28598 3460
rect 28592 3420 35894 3448
rect 28592 3408 28598 3420
rect 26510 3380 26516 3392
rect 22066 3352 26516 3380
rect 19889 3343 19947 3349
rect 26510 3340 26516 3352
rect 26568 3340 26574 3392
rect 27522 3340 27528 3392
rect 27580 3380 27586 3392
rect 28629 3383 28687 3389
rect 28629 3380 28641 3383
rect 27580 3352 28641 3380
rect 27580 3340 27586 3352
rect 28629 3349 28641 3352
rect 28675 3349 28687 3383
rect 35866 3380 35894 3420
rect 36998 3380 37004 3392
rect 35866 3352 37004 3380
rect 28629 3343 28687 3349
rect 36998 3340 37004 3352
rect 37056 3340 37062 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3878 3136 3884 3188
rect 3936 3136 3942 3188
rect 4062 3136 4068 3188
rect 4120 3136 4126 3188
rect 5074 3136 5080 3188
rect 5132 3136 5138 3188
rect 5258 3136 5264 3188
rect 5316 3136 5322 3188
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5408 3148 5733 3176
rect 5408 3136 5414 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 6638 3136 6644 3188
rect 6696 3136 6702 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6972 3148 7113 3176
rect 6972 3136 6978 3148
rect 7101 3145 7113 3148
rect 7147 3176 7159 3179
rect 7374 3176 7380 3188
rect 7147 3148 7380 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7484 3148 8064 3176
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 3896 3040 3924 3136
rect 3835 3012 3924 3040
rect 4080 3040 4108 3136
rect 5092 3108 5120 3136
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 5092 3080 5181 3108
rect 5169 3077 5181 3080
rect 5215 3077 5227 3111
rect 5169 3071 5227 3077
rect 5534 3068 5540 3120
rect 5592 3068 5598 3120
rect 7484 3117 7512 3148
rect 7469 3111 7527 3117
rect 7469 3077 7481 3111
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 7558 3068 7564 3120
rect 7616 3108 7622 3120
rect 8036 3108 8064 3148
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 8168 3148 9413 3176
rect 8168 3136 8174 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9401 3139 9459 3145
rect 9784 3148 10793 3176
rect 9674 3108 9680 3120
rect 7616 3080 7788 3108
rect 8036 3080 9680 3108
rect 7616 3068 7622 3080
rect 4080 3012 5212 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1673 2975 1731 2981
rect 1673 2972 1685 2975
rect 1443 2944 1685 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1673 2941 1685 2944
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2774 2972 2780 2984
rect 1903 2944 2780 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2941 2927 2975
rect 2869 2935 2927 2941
rect 1578 2864 1584 2916
rect 1636 2904 1642 2916
rect 2884 2904 2912 2935
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 3936 2944 4169 2972
rect 3936 2932 3942 2944
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 5184 2972 5212 3012
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5316 3012 5641 3040
rect 5316 3000 5322 3012
rect 5629 3009 5641 3012
rect 5675 3040 5687 3043
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 5675 3012 7021 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7650 3040 7656 3052
rect 7009 3003 7067 3009
rect 7484 3012 7656 3040
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 5184 2944 5365 2972
rect 4157 2935 4215 2941
rect 5353 2941 5365 2944
rect 5399 2972 5411 2975
rect 7098 2972 7104 2984
rect 5399 2944 7104 2972
rect 5399 2941 5411 2944
rect 5353 2935 5411 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7484 2972 7512 3012
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7760 3049 7788 3080
rect 9674 3068 9680 3080
rect 9732 3068 9738 3120
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8435 3012 8953 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8941 3009 8953 3012
rect 8987 3040 8999 3043
rect 9490 3040 9496 3052
rect 8987 3012 9496 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 7331 2944 7512 2972
rect 7561 2975 7619 2981
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 8220 2972 8248 3003
rect 9490 3000 9496 3012
rect 9548 3040 9554 3052
rect 9784 3040 9812 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 12253 3179 12311 3185
rect 10781 3139 10839 3145
rect 11716 3148 12204 3176
rect 9858 3068 9864 3120
rect 9916 3068 9922 3120
rect 9548 3012 9812 3040
rect 9876 3040 9904 3068
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 9876 3012 10425 3040
rect 9548 3000 9554 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10502 3000 10508 3052
rect 10560 3000 10566 3052
rect 11716 3040 11744 3148
rect 11790 3068 11796 3120
rect 11848 3068 11854 3120
rect 10612 3012 11744 3040
rect 10612 2972 10640 3012
rect 12066 3000 12072 3052
rect 12124 3000 12130 3052
rect 12176 3040 12204 3148
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12299 3148 12434 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12406 3108 12434 3148
rect 14918 3136 14924 3188
rect 14976 3136 14982 3188
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 16114 3176 16120 3188
rect 15427 3148 16120 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 16206 3136 16212 3188
rect 16264 3176 16270 3188
rect 17865 3179 17923 3185
rect 17865 3176 17877 3179
rect 16264 3148 17877 3176
rect 16264 3136 16270 3148
rect 17865 3145 17877 3148
rect 17911 3145 17923 3179
rect 17865 3139 17923 3145
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 19392 3148 20085 3176
rect 19392 3136 19398 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 20220 3148 26556 3176
rect 20220 3136 20226 3148
rect 14268 3111 14326 3117
rect 12406 3080 14228 3108
rect 12176 3012 13952 3040
rect 7561 2935 7619 2941
rect 7659 2944 8248 2972
rect 8680 2944 10640 2972
rect 1636 2876 2912 2904
rect 1636 2864 1642 2876
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 7576 2904 7604 2935
rect 7064 2876 7604 2904
rect 7064 2864 7070 2876
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 5258 2836 5264 2848
rect 2556 2808 5264 2836
rect 2556 2796 2562 2808
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5442 2796 5448 2848
rect 5500 2796 5506 2848
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 7659 2836 7687 2944
rect 8021 2907 8079 2913
rect 8021 2904 8033 2907
rect 7760 2876 8033 2904
rect 7760 2845 7788 2876
rect 8021 2873 8033 2876
rect 8067 2873 8079 2907
rect 8021 2867 8079 2873
rect 7340 2808 7687 2836
rect 7745 2839 7803 2845
rect 7340 2796 7346 2808
rect 7745 2805 7757 2839
rect 7791 2805 7803 2839
rect 7745 2799 7803 2805
rect 7929 2839 7987 2845
rect 7929 2805 7941 2839
rect 7975 2836 7987 2839
rect 8680 2836 8708 2944
rect 11882 2932 11888 2984
rect 11940 2932 11946 2984
rect 8754 2864 8760 2916
rect 8812 2864 8818 2916
rect 9309 2907 9367 2913
rect 9309 2873 9321 2907
rect 9355 2904 9367 2907
rect 9766 2904 9772 2916
rect 9355 2876 9772 2904
rect 9355 2873 9367 2876
rect 9309 2867 9367 2873
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 9861 2907 9919 2913
rect 9861 2873 9873 2907
rect 9907 2904 9919 2907
rect 10318 2904 10324 2916
rect 9907 2876 10324 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 7975 2808 8708 2836
rect 7975 2805 7987 2808
rect 7929 2799 7987 2805
rect 8846 2796 8852 2848
rect 8904 2796 8910 2848
rect 9950 2796 9956 2848
rect 10008 2796 10014 2848
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12158 2836 12164 2848
rect 12115 2808 12164 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 13924 2836 13952 3012
rect 13998 3000 14004 3052
rect 14056 3000 14062 3052
rect 14200 3040 14228 3080
rect 14268 3077 14280 3111
rect 14314 3108 14326 3111
rect 14936 3108 14964 3136
rect 21450 3108 21456 3120
rect 14314 3080 14964 3108
rect 15028 3080 17724 3108
rect 14314 3077 14326 3080
rect 14268 3071 14326 3077
rect 15028 3040 15056 3080
rect 16301 3043 16359 3049
rect 16301 3040 16313 3043
rect 14200 3012 15056 3040
rect 15120 3012 16313 3040
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15120 2972 15148 3012
rect 16301 3009 16313 3012
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3040 17463 3043
rect 17586 3040 17592 3052
rect 17451 3012 17592 3040
rect 17451 3009 17463 3012
rect 17405 3003 17463 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 17696 3049 17724 3080
rect 19628 3080 21456 3108
rect 19628 3049 19656 3080
rect 21450 3068 21456 3080
rect 21508 3068 21514 3120
rect 26418 3108 26424 3120
rect 25056 3080 26424 3108
rect 25056 3049 25084 3080
rect 26418 3068 26424 3080
rect 26476 3068 26482 3120
rect 26528 3108 26556 3148
rect 26786 3136 26792 3188
rect 26844 3136 26850 3188
rect 27433 3179 27491 3185
rect 27433 3176 27445 3179
rect 26896 3148 27445 3176
rect 26896 3108 26924 3148
rect 27433 3145 27445 3148
rect 27479 3145 27491 3179
rect 27433 3139 27491 3145
rect 28074 3136 28080 3188
rect 28132 3176 28138 3188
rect 28905 3179 28963 3185
rect 28905 3176 28917 3179
rect 28132 3148 28917 3176
rect 28132 3136 28138 3148
rect 28905 3145 28917 3148
rect 28951 3145 28963 3179
rect 28905 3139 28963 3145
rect 28994 3136 29000 3188
rect 29052 3176 29058 3188
rect 29641 3179 29699 3185
rect 29641 3176 29653 3179
rect 29052 3148 29653 3176
rect 29052 3136 29058 3148
rect 29641 3145 29653 3148
rect 29687 3145 29699 3179
rect 33873 3179 33931 3185
rect 33873 3176 33885 3179
rect 29641 3139 29699 3145
rect 32232 3148 33885 3176
rect 26528 3080 26924 3108
rect 26973 3111 27031 3117
rect 26973 3077 26985 3111
rect 27019 3108 27031 3111
rect 32232 3108 32260 3148
rect 33873 3145 33885 3148
rect 33919 3176 33931 3179
rect 33919 3148 35480 3176
rect 33919 3145 33931 3148
rect 33873 3139 33931 3145
rect 27019 3080 32260 3108
rect 33229 3111 33287 3117
rect 27019 3077 27031 3080
rect 26973 3071 27031 3077
rect 33229 3077 33241 3111
rect 33275 3108 33287 3111
rect 35342 3108 35348 3120
rect 33275 3080 35348 3108
rect 33275 3077 33287 3080
rect 33229 3071 33287 3077
rect 35342 3068 35348 3080
rect 35400 3068 35406 3120
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3009 19671 3043
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19613 3003 19671 3009
rect 19720 3012 19901 3040
rect 15068 2944 15148 2972
rect 15068 2932 15074 2944
rect 15654 2932 15660 2984
rect 15712 2932 15718 2984
rect 16758 2932 16764 2984
rect 16816 2932 16822 2984
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 17359 2944 17509 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19720 2972 19748 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 25041 3043 25099 3049
rect 25041 3009 25053 3043
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 25317 3043 25375 3049
rect 25317 3009 25329 3043
rect 25363 3009 25375 3043
rect 25317 3003 25375 3009
rect 26329 3043 26387 3049
rect 26329 3009 26341 3043
rect 26375 3009 26387 3043
rect 26329 3003 26387 3009
rect 18840 2944 19748 2972
rect 19797 2975 19855 2981
rect 18840 2932 18846 2944
rect 19797 2941 19809 2975
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 19812 2904 19840 2935
rect 20162 2932 20168 2984
rect 20220 2932 20226 2984
rect 25130 2932 25136 2984
rect 25188 2932 25194 2984
rect 20809 2907 20867 2913
rect 20809 2904 20821 2907
rect 14936 2876 17448 2904
rect 19812 2876 20821 2904
rect 14936 2836 14964 2876
rect 17420 2845 17448 2876
rect 20809 2873 20821 2876
rect 20855 2873 20867 2907
rect 20809 2867 20867 2873
rect 23658 2864 23664 2916
rect 23716 2904 23722 2916
rect 25332 2904 25360 3003
rect 26344 2972 26372 3003
rect 26510 3000 26516 3052
rect 26568 3000 26574 3052
rect 26605 3043 26663 3049
rect 26605 3009 26617 3043
rect 26651 3040 26663 3043
rect 27249 3043 27307 3049
rect 27249 3040 27261 3043
rect 26651 3012 27261 3040
rect 26651 3009 26663 3012
rect 26605 3003 26663 3009
rect 27249 3009 27261 3012
rect 27295 3040 27307 3043
rect 27522 3040 27528 3052
rect 27295 3012 27528 3040
rect 27295 3009 27307 3012
rect 27249 3003 27307 3009
rect 27522 3000 27528 3012
rect 27580 3000 27586 3052
rect 28442 3000 28448 3052
rect 28500 3000 28506 3052
rect 28534 3000 28540 3052
rect 28592 3000 28598 3052
rect 28718 3000 28724 3052
rect 28776 3000 28782 3052
rect 28902 3000 28908 3052
rect 28960 3000 28966 3052
rect 32306 3000 32312 3052
rect 32364 3040 32370 3052
rect 33689 3043 33747 3049
rect 33689 3040 33701 3043
rect 32364 3012 33701 3040
rect 32364 3000 32370 3012
rect 33689 3009 33701 3012
rect 33735 3009 33747 3043
rect 35452 3040 35480 3148
rect 36998 3136 37004 3188
rect 37056 3136 37062 3188
rect 35713 3111 35771 3117
rect 35713 3077 35725 3111
rect 35759 3108 35771 3111
rect 35759 3080 36492 3108
rect 35759 3077 35771 3080
rect 35713 3071 35771 3077
rect 36464 3052 36492 3080
rect 35989 3043 36047 3049
rect 35989 3040 36001 3043
rect 35452 3012 36001 3040
rect 33689 3003 33747 3009
rect 35989 3009 36001 3012
rect 36035 3009 36047 3043
rect 35989 3003 36047 3009
rect 36173 3043 36231 3049
rect 36173 3009 36185 3043
rect 36219 3009 36231 3043
rect 36173 3003 36231 3009
rect 27157 2975 27215 2981
rect 26344 2944 27108 2972
rect 27080 2904 27108 2944
rect 27157 2941 27169 2975
rect 27203 2972 27215 2975
rect 28552 2972 28580 3000
rect 27203 2944 28580 2972
rect 28629 2975 28687 2981
rect 27203 2941 27215 2944
rect 27157 2935 27215 2941
rect 28629 2941 28641 2975
rect 28675 2972 28687 2975
rect 28920 2972 28948 3000
rect 28675 2944 28948 2972
rect 28675 2941 28687 2944
rect 28629 2935 28687 2941
rect 29086 2932 29092 2984
rect 29144 2932 29150 2984
rect 33502 2932 33508 2984
rect 33560 2932 33566 2984
rect 36188 2972 36216 3003
rect 36446 3000 36452 3052
rect 36504 3000 36510 3052
rect 36725 2975 36783 2981
rect 36725 2972 36737 2975
rect 36188 2944 36737 2972
rect 36725 2941 36737 2944
rect 36771 2972 36783 2975
rect 38010 2972 38016 2984
rect 36771 2944 38016 2972
rect 36771 2941 36783 2944
rect 36725 2935 36783 2941
rect 38010 2932 38016 2944
rect 38068 2932 38074 2984
rect 36357 2907 36415 2913
rect 36357 2904 36369 2907
rect 23716 2876 25360 2904
rect 26344 2876 27016 2904
rect 27080 2876 36369 2904
rect 23716 2864 23722 2876
rect 13924 2808 14964 2836
rect 17405 2839 17463 2845
rect 17405 2805 17417 2839
rect 17451 2805 17463 2839
rect 17405 2799 17463 2805
rect 19889 2839 19947 2845
rect 19889 2805 19901 2839
rect 19935 2836 19947 2839
rect 20990 2836 20996 2848
rect 19935 2808 20996 2836
rect 19935 2805 19947 2808
rect 19889 2799 19947 2805
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 25317 2839 25375 2845
rect 25317 2805 25329 2839
rect 25363 2836 25375 2839
rect 25406 2836 25412 2848
rect 25363 2808 25412 2836
rect 25363 2805 25375 2808
rect 25317 2799 25375 2805
rect 25406 2796 25412 2808
rect 25464 2796 25470 2848
rect 26344 2845 26372 2876
rect 26988 2845 27016 2876
rect 36357 2873 36369 2876
rect 36403 2873 36415 2907
rect 36357 2867 36415 2873
rect 36832 2876 37596 2904
rect 25501 2839 25559 2845
rect 25501 2805 25513 2839
rect 25547 2836 25559 2839
rect 26329 2839 26387 2845
rect 26329 2836 26341 2839
rect 25547 2808 26341 2836
rect 25547 2805 25559 2808
rect 25501 2799 25559 2805
rect 26329 2805 26341 2808
rect 26375 2805 26387 2839
rect 26329 2799 26387 2805
rect 26973 2839 27031 2845
rect 26973 2805 26985 2839
rect 27019 2805 27031 2839
rect 26973 2799 27031 2805
rect 28721 2839 28779 2845
rect 28721 2805 28733 2839
rect 28767 2836 28779 2839
rect 30098 2836 30104 2848
rect 28767 2808 30104 2836
rect 28767 2805 28779 2808
rect 28721 2799 28779 2805
rect 30098 2796 30104 2808
rect 30156 2796 30162 2848
rect 33686 2796 33692 2848
rect 33744 2796 33750 2848
rect 36832 2845 36860 2876
rect 37568 2848 37596 2876
rect 36173 2839 36231 2845
rect 36173 2805 36185 2839
rect 36219 2836 36231 2839
rect 36817 2839 36875 2845
rect 36817 2836 36829 2839
rect 36219 2808 36829 2836
rect 36219 2805 36231 2808
rect 36173 2799 36231 2805
rect 36817 2805 36829 2808
rect 36863 2805 36875 2839
rect 36817 2799 36875 2805
rect 37550 2796 37556 2848
rect 37608 2796 37614 2848
rect 38473 2839 38531 2845
rect 38473 2805 38485 2839
rect 38519 2836 38531 2839
rect 39298 2836 39304 2848
rect 38519 2808 39304 2836
rect 38519 2805 38531 2808
rect 38473 2799 38531 2805
rect 39298 2796 39304 2808
rect 39356 2796 39362 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 2498 2632 2504 2644
rect 1811 2604 2504 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 2498 2592 2504 2604
rect 2556 2592 2562 2644
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 2639 2604 3004 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 2774 2524 2780 2576
rect 2832 2524 2838 2576
rect 2976 2496 3004 2604
rect 3602 2592 3608 2644
rect 3660 2592 3666 2644
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4706 2632 4712 2644
rect 4479 2604 4712 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 7006 2632 7012 2644
rect 6411 2604 7012 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 8297 2635 8355 2641
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 8343 2604 9628 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 7392 2564 7420 2592
rect 4571 2536 7420 2564
rect 8757 2567 8815 2573
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 8757 2533 8769 2567
rect 8803 2564 8815 2567
rect 9490 2564 9496 2576
rect 8803 2536 9496 2564
rect 8803 2533 8815 2536
rect 8757 2527 8815 2533
rect 9490 2524 9496 2536
rect 9548 2524 9554 2576
rect 9600 2564 9628 2604
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 9732 2604 10425 2632
rect 9732 2592 9738 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11882 2632 11888 2644
rect 11103 2604 11888 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12158 2592 12164 2644
rect 12216 2592 12222 2644
rect 16669 2635 16727 2641
rect 16669 2601 16681 2635
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 12066 2564 12072 2576
rect 9600 2536 12072 2564
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 14369 2567 14427 2573
rect 14369 2533 14381 2567
rect 14415 2533 14427 2567
rect 14369 2527 14427 2533
rect 15197 2567 15255 2573
rect 15197 2533 15209 2567
rect 15243 2564 15255 2567
rect 16684 2564 16712 2595
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 16816 2604 17141 2632
rect 16816 2592 16822 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 17129 2595 17187 2601
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 18782 2632 18788 2644
rect 17727 2604 18788 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 19613 2635 19671 2641
rect 19613 2601 19625 2635
rect 19659 2632 19671 2635
rect 20162 2632 20168 2644
rect 19659 2604 20168 2632
rect 19659 2601 19671 2604
rect 19613 2595 19671 2601
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20990 2592 20996 2644
rect 21048 2592 21054 2644
rect 21450 2592 21456 2644
rect 21508 2592 21514 2644
rect 22097 2635 22155 2641
rect 22097 2601 22109 2635
rect 22143 2632 22155 2635
rect 23658 2632 23664 2644
rect 22143 2604 23664 2632
rect 22143 2601 22155 2604
rect 22097 2595 22155 2601
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 24397 2635 24455 2641
rect 24397 2601 24409 2635
rect 24443 2632 24455 2635
rect 25130 2632 25136 2644
rect 24443 2604 25136 2632
rect 24443 2601 24455 2604
rect 24397 2595 24455 2601
rect 25130 2592 25136 2604
rect 25188 2592 25194 2644
rect 25406 2592 25412 2644
rect 25464 2592 25470 2644
rect 26418 2592 26424 2644
rect 26476 2632 26482 2644
rect 27617 2635 27675 2641
rect 27617 2632 27629 2635
rect 26476 2604 27629 2632
rect 26476 2592 26482 2604
rect 27617 2601 27629 2604
rect 27663 2601 27675 2635
rect 27617 2595 27675 2601
rect 28718 2592 28724 2644
rect 28776 2592 28782 2644
rect 29086 2592 29092 2644
rect 29144 2632 29150 2644
rect 29549 2635 29607 2641
rect 29549 2632 29561 2635
rect 29144 2604 29561 2632
rect 29144 2592 29150 2604
rect 29549 2601 29561 2604
rect 29595 2601 29607 2635
rect 29549 2595 29607 2601
rect 30098 2592 30104 2644
rect 30156 2592 30162 2644
rect 30929 2635 30987 2641
rect 30929 2601 30941 2635
rect 30975 2632 30987 2635
rect 32306 2632 32312 2644
rect 30975 2604 32312 2632
rect 30975 2601 30987 2604
rect 30929 2595 30987 2601
rect 32306 2592 32312 2604
rect 32364 2592 32370 2644
rect 33137 2635 33195 2641
rect 33137 2601 33149 2635
rect 33183 2632 33195 2635
rect 33502 2632 33508 2644
rect 33183 2604 33508 2632
rect 33183 2601 33195 2604
rect 33137 2595 33195 2601
rect 33502 2592 33508 2604
rect 33560 2592 33566 2644
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 34241 2635 34299 2641
rect 34241 2632 34253 2635
rect 33744 2604 34253 2632
rect 33744 2592 33750 2604
rect 34241 2601 34253 2604
rect 34287 2601 34299 2635
rect 34241 2595 34299 2601
rect 35342 2592 35348 2644
rect 35400 2592 35406 2644
rect 36446 2592 36452 2644
rect 36504 2592 36510 2644
rect 37550 2592 37556 2644
rect 37608 2592 37614 2644
rect 38010 2592 38016 2644
rect 38068 2592 38074 2644
rect 17957 2567 18015 2573
rect 17957 2564 17969 2567
rect 15243 2536 16574 2564
rect 16684 2536 17969 2564
rect 15243 2533 15255 2536
rect 15197 2527 15255 2533
rect 2976 2468 3096 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1596 2360 1624 2391
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 1728 2400 1961 2428
rect 1728 2388 1734 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 2130 2388 2136 2440
rect 2188 2388 2194 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2363 2400 2421 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 3068 2428 3096 2468
rect 3418 2456 3424 2508
rect 3476 2496 3482 2508
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 3476 2468 3801 2496
rect 3476 2456 3482 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 5258 2456 5264 2508
rect 5316 2456 5322 2508
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6880 2468 7113 2496
rect 6880 2456 6886 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 8260 2468 9413 2496
rect 8260 2456 8266 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 14384 2496 14412 2527
rect 16117 2499 16175 2505
rect 16117 2496 16129 2499
rect 11848 2468 14412 2496
rect 15396 2468 16129 2496
rect 11848 2456 11854 2468
rect 4246 2428 4252 2440
rect 3068 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4396 2400 4721 2428
rect 4396 2388 4402 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5000 2360 5028 2391
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5868 2400 6561 2428
rect 5868 2388 5874 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 8110 2428 8116 2440
rect 6779 2400 8116 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 8938 2388 8944 2440
rect 8996 2388 9002 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 10042 2388 10048 2440
rect 10100 2428 10106 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10100 2400 10609 2428
rect 10100 2388 10106 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10870 2388 10876 2440
rect 10928 2388 10934 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11020 2400 11253 2428
rect 11020 2388 11026 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11756 2400 11989 2428
rect 11756 2388 11762 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12124 2400 12357 2428
rect 12124 2388 12130 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12860 2400 13093 2428
rect 12860 2388 12866 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 13228 2400 13461 2428
rect 13228 2388 13234 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13964 2400 14289 2428
rect 13964 2388 13970 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 15396 2437 15424 2468
rect 16117 2465 16129 2468
rect 16163 2465 16175 2499
rect 16546 2496 16574 2536
rect 17957 2533 17969 2536
rect 18003 2533 18015 2567
rect 21468 2564 21496 2592
rect 23201 2567 23259 2573
rect 23201 2564 23213 2567
rect 21468 2536 23213 2564
rect 17957 2527 18015 2533
rect 23201 2533 23213 2536
rect 23247 2533 23259 2567
rect 23201 2527 23259 2533
rect 26513 2567 26571 2573
rect 26513 2533 26525 2567
rect 26559 2564 26571 2567
rect 28736 2564 28764 2592
rect 26559 2536 28764 2564
rect 26559 2533 26571 2536
rect 26513 2527 26571 2533
rect 29362 2524 29368 2576
rect 29420 2564 29426 2576
rect 30009 2567 30067 2573
rect 30009 2564 30021 2567
rect 29420 2536 30021 2564
rect 29420 2524 29426 2536
rect 30009 2533 30021 2536
rect 30055 2533 30067 2567
rect 30009 2527 30067 2533
rect 32122 2524 32128 2576
rect 32180 2524 32186 2576
rect 16761 2499 16819 2505
rect 16761 2496 16773 2499
rect 16546 2468 16773 2496
rect 16117 2459 16175 2465
rect 16761 2465 16773 2468
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14424 2400 14565 2428
rect 14424 2388 14430 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16264 2400 16497 2428
rect 16264 2388 16270 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16485 2391 16543 2397
rect 16592 2400 16957 2428
rect 9784 2360 9812 2388
rect 16592 2360 16620 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17276 2400 17509 2428
rect 17276 2388 17282 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 17586 2388 17592 2440
rect 17644 2428 17650 2440
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17644 2400 17877 2428
rect 17644 2388 17650 2400
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 18138 2388 18144 2440
rect 18196 2388 18202 2440
rect 18322 2388 18328 2440
rect 18380 2428 18386 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18380 2400 18613 2428
rect 18380 2388 18386 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 18748 2400 18981 2428
rect 18748 2388 18754 2400
rect 18969 2397 18981 2400
rect 19015 2397 19027 2431
rect 18969 2391 19027 2397
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 1596 2332 2544 2360
rect 5000 2332 9812 2360
rect 13280 2332 16620 2360
rect 16669 2363 16727 2369
rect 2516 2304 2544 2332
rect 2498 2252 2504 2304
rect 2556 2252 2562 2304
rect 13280 2301 13308 2332
rect 16669 2329 16681 2363
rect 16715 2360 16727 2363
rect 19812 2360 19840 2391
rect 19886 2388 19892 2440
rect 19944 2388 19950 2440
rect 20806 2388 20812 2440
rect 20864 2388 20870 2440
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 21177 2431 21235 2437
rect 21177 2428 21189 2431
rect 20956 2400 21189 2428
rect 20956 2388 20962 2400
rect 21177 2397 21189 2400
rect 21223 2397 21235 2431
rect 21177 2391 21235 2397
rect 21634 2388 21640 2440
rect 21692 2428 21698 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21692 2400 22017 2428
rect 21692 2388 21698 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22278 2388 22284 2440
rect 22336 2388 22342 2440
rect 22738 2388 22744 2440
rect 22796 2428 22802 2440
rect 23017 2431 23075 2437
rect 23017 2428 23029 2431
rect 22796 2400 23029 2428
rect 22796 2388 22802 2400
rect 23017 2397 23029 2400
rect 23063 2397 23075 2431
rect 23017 2391 23075 2397
rect 23106 2388 23112 2440
rect 23164 2428 23170 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23164 2400 23397 2428
rect 23164 2388 23170 2400
rect 23385 2397 23397 2400
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24121 2431 24179 2437
rect 24121 2428 24133 2431
rect 23900 2400 24133 2428
rect 23900 2388 23906 2400
rect 24121 2397 24133 2400
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 24210 2388 24216 2440
rect 24268 2428 24274 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24268 2400 24593 2428
rect 24268 2388 24274 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 24946 2388 24952 2440
rect 25004 2428 25010 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 25004 2400 25237 2428
rect 25004 2388 25010 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 25314 2388 25320 2440
rect 25372 2428 25378 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25372 2400 25605 2428
rect 25372 2388 25378 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26142 2388 26148 2440
rect 26200 2428 26206 2440
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 26200 2400 26341 2428
rect 26200 2388 26206 2400
rect 26329 2397 26341 2400
rect 26375 2397 26387 2431
rect 26329 2391 26387 2397
rect 26418 2388 26424 2440
rect 26476 2428 26482 2440
rect 26697 2431 26755 2437
rect 26697 2428 26709 2431
rect 26476 2400 26709 2428
rect 26476 2388 26482 2400
rect 26697 2397 26709 2400
rect 26743 2397 26755 2431
rect 26697 2391 26755 2397
rect 27154 2388 27160 2440
rect 27212 2428 27218 2440
rect 27433 2431 27491 2437
rect 27433 2428 27445 2431
rect 27212 2400 27445 2428
rect 27212 2388 27218 2400
rect 27433 2397 27445 2400
rect 27479 2397 27491 2431
rect 27433 2391 27491 2397
rect 27522 2388 27528 2440
rect 27580 2428 27586 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27580 2400 27813 2428
rect 27580 2388 27586 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28258 2388 28264 2440
rect 28316 2428 28322 2440
rect 28537 2431 28595 2437
rect 28537 2428 28549 2431
rect 28316 2400 28549 2428
rect 28316 2388 28322 2400
rect 28537 2397 28549 2400
rect 28583 2397 28595 2431
rect 28537 2391 28595 2397
rect 28718 2388 28724 2440
rect 28776 2388 28782 2440
rect 29365 2431 29423 2437
rect 29365 2397 29377 2431
rect 29411 2428 29423 2431
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29411 2400 29745 2428
rect 29411 2397 29423 2400
rect 29365 2391 29423 2397
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 16715 2332 18828 2360
rect 19812 2332 20545 2360
rect 16715 2329 16727 2332
rect 16669 2323 16727 2329
rect 13265 2295 13323 2301
rect 13265 2261 13277 2295
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 14918 2252 14924 2304
rect 14976 2252 14982 2304
rect 18800 2301 18828 2332
rect 20533 2329 20545 2332
rect 20579 2329 20591 2363
rect 20533 2323 20591 2329
rect 29914 2320 29920 2372
rect 29972 2360 29978 2372
rect 30300 2360 30328 2391
rect 30466 2388 30472 2440
rect 30524 2428 30530 2440
rect 30745 2431 30803 2437
rect 30745 2428 30757 2431
rect 30524 2400 30757 2428
rect 30524 2388 30530 2400
rect 30745 2397 30757 2400
rect 30791 2397 30803 2431
rect 30745 2391 30803 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30892 2400 31125 2428
rect 30892 2388 30898 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 31849 2431 31907 2437
rect 31849 2428 31861 2431
rect 31628 2400 31861 2428
rect 31628 2388 31634 2400
rect 31849 2397 31861 2400
rect 31895 2397 31907 2431
rect 31849 2391 31907 2397
rect 31938 2388 31944 2440
rect 31996 2428 32002 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31996 2400 32321 2428
rect 31996 2388 32002 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32674 2388 32680 2440
rect 32732 2428 32738 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32732 2400 32965 2428
rect 32732 2388 32738 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 33042 2388 33048 2440
rect 33100 2428 33106 2440
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 33100 2400 33333 2428
rect 33100 2388 33106 2400
rect 33321 2397 33333 2400
rect 33367 2397 33379 2431
rect 33321 2391 33379 2397
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34057 2431 34115 2437
rect 34057 2428 34069 2431
rect 33836 2400 34069 2428
rect 33836 2388 33842 2400
rect 34057 2397 34069 2400
rect 34103 2397 34115 2431
rect 34057 2391 34115 2397
rect 34146 2388 34152 2440
rect 34204 2428 34210 2440
rect 34425 2431 34483 2437
rect 34425 2428 34437 2431
rect 34204 2400 34437 2428
rect 34204 2388 34210 2400
rect 34425 2397 34437 2400
rect 34471 2397 34483 2431
rect 34425 2391 34483 2397
rect 34882 2388 34888 2440
rect 34940 2428 34946 2440
rect 35161 2431 35219 2437
rect 35161 2428 35173 2431
rect 34940 2400 35173 2428
rect 34940 2388 34946 2400
rect 35161 2397 35173 2400
rect 35207 2397 35219 2431
rect 35161 2391 35219 2397
rect 35250 2388 35256 2440
rect 35308 2428 35314 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35308 2400 35541 2428
rect 35308 2388 35314 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 35986 2388 35992 2440
rect 36044 2428 36050 2440
rect 36265 2431 36323 2437
rect 36265 2428 36277 2431
rect 36044 2400 36277 2428
rect 36044 2388 36050 2400
rect 36265 2397 36277 2400
rect 36311 2397 36323 2431
rect 36265 2391 36323 2397
rect 36354 2388 36360 2440
rect 36412 2428 36418 2440
rect 36633 2431 36691 2437
rect 36633 2428 36645 2431
rect 36412 2400 36645 2428
rect 36412 2388 36418 2400
rect 36633 2397 36645 2400
rect 36679 2397 36691 2431
rect 36633 2391 36691 2397
rect 37090 2388 37096 2440
rect 37148 2428 37154 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 37148 2400 37473 2428
rect 37148 2388 37154 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 37550 2388 37556 2440
rect 37608 2428 37614 2440
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 37608 2400 37749 2428
rect 37608 2388 37614 2400
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38197 2431 38255 2437
rect 38197 2397 38209 2431
rect 38243 2397 38255 2431
rect 38197 2391 38255 2397
rect 29972 2332 30328 2360
rect 38212 2360 38240 2391
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 38473 2431 38531 2437
rect 38473 2428 38485 2431
rect 38344 2400 38485 2428
rect 38344 2388 38350 2400
rect 38473 2397 38485 2400
rect 38519 2397 38531 2431
rect 38473 2391 38531 2397
rect 38562 2360 38568 2372
rect 38212 2332 38568 2360
rect 29972 2320 29978 2332
rect 38562 2320 38568 2332
rect 38620 2320 38626 2372
rect 18785 2295 18843 2301
rect 18785 2261 18797 2295
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 4246 2048 4252 2100
rect 4304 2088 4310 2100
rect 15378 2088 15384 2100
rect 4304 2060 15384 2088
rect 4304 2048 4310 2060
rect 15378 2048 15384 2060
rect 15436 2048 15442 2100
rect 16482 1368 16488 1420
rect 16540 1408 16546 1420
rect 18138 1408 18144 1420
rect 16540 1380 18144 1408
rect 16540 1368 16546 1380
rect 18138 1368 18144 1380
rect 18196 1368 18202 1420
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 38108 35003 38160 35012
rect 38108 34969 38117 35003
rect 38117 34969 38151 35003
rect 38151 34969 38160 35003
rect 38108 34960 38160 34969
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 38016 25100 38068 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 39028 25032 39080 25084
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 14464 15988 14516 16040
rect 14740 15895 14792 15904
rect 14740 15861 14749 15895
rect 14749 15861 14783 15895
rect 14783 15861 14792 15895
rect 14740 15852 14792 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 14556 15487 14608 15496
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 12532 15308 12584 15360
rect 15108 15351 15160 15360
rect 15108 15317 15117 15351
rect 15117 15317 15151 15351
rect 15151 15317 15160 15351
rect 15108 15308 15160 15317
rect 38384 15351 38436 15360
rect 38384 15317 38393 15351
rect 38393 15317 38427 15351
rect 38427 15317 38436 15351
rect 38384 15308 38436 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 38936 15172 38988 15224
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 14740 15104 14792 15156
rect 12532 14968 12584 15020
rect 14096 15036 14148 15088
rect 15108 15036 15160 15088
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 10600 14900 10652 14952
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8852 14764 8904 14816
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 11336 14764 11388 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 16120 14900 16172 14952
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 17316 14807 17368 14816
rect 17316 14773 17325 14807
rect 17325 14773 17359 14807
rect 17359 14773 17368 14807
rect 17316 14764 17368 14773
rect 17592 14807 17644 14816
rect 17592 14773 17601 14807
rect 17601 14773 17635 14807
rect 17635 14773 17644 14807
rect 17592 14764 17644 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 8852 14560 8904 14612
rect 9956 14560 10008 14612
rect 10876 14560 10928 14612
rect 11796 14603 11848 14612
rect 11796 14569 11805 14603
rect 11805 14569 11839 14603
rect 11839 14569 11848 14603
rect 11796 14560 11848 14569
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 16764 14535 16816 14544
rect 16764 14501 16773 14535
rect 16773 14501 16807 14535
rect 16807 14501 16816 14535
rect 16764 14492 16816 14501
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 12348 14467 12400 14476
rect 12348 14433 12357 14467
rect 12357 14433 12391 14467
rect 12391 14433 12400 14467
rect 12348 14424 12400 14433
rect 12900 14424 12952 14476
rect 14096 14424 14148 14476
rect 17316 14560 17368 14612
rect 19432 14424 19484 14476
rect 20536 14424 20588 14476
rect 38016 14424 38068 14476
rect 8668 14288 8720 14340
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 19340 14399 19392 14408
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 11244 14288 11296 14340
rect 17316 14288 17368 14340
rect 9312 14220 9364 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 10692 14263 10744 14272
rect 10692 14229 10701 14263
rect 10701 14229 10735 14263
rect 10735 14229 10744 14263
rect 10692 14220 10744 14229
rect 11428 14220 11480 14272
rect 13084 14220 13136 14272
rect 15200 14220 15252 14272
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 16580 14220 16632 14272
rect 17592 14220 17644 14272
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 19064 14263 19116 14272
rect 19064 14229 19073 14263
rect 19073 14229 19107 14263
rect 19107 14229 19116 14263
rect 19064 14220 19116 14229
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 38200 14220 38252 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 8116 14016 8168 14068
rect 9404 14016 9456 14068
rect 10692 14016 10744 14068
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 9496 13812 9548 13864
rect 11428 13812 11480 13864
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 16580 14016 16632 14068
rect 16764 14016 16816 14068
rect 17316 14059 17368 14068
rect 17316 14025 17325 14059
rect 17325 14025 17359 14059
rect 17359 14025 17368 14059
rect 17316 14016 17368 14025
rect 17684 14059 17736 14068
rect 17684 14025 17693 14059
rect 17693 14025 17727 14059
rect 17727 14025 17736 14059
rect 17684 14016 17736 14025
rect 19064 14016 19116 14068
rect 19984 14016 20036 14068
rect 17776 13948 17828 14000
rect 20536 13948 20588 14000
rect 12348 13744 12400 13796
rect 9588 13676 9640 13728
rect 12716 13719 12768 13728
rect 12716 13685 12725 13719
rect 12725 13685 12759 13719
rect 12759 13685 12768 13719
rect 12716 13676 12768 13685
rect 13084 13719 13136 13728
rect 13084 13685 13093 13719
rect 13093 13685 13127 13719
rect 13127 13685 13136 13719
rect 13084 13676 13136 13685
rect 18144 13676 18196 13728
rect 20444 13719 20496 13728
rect 20444 13685 20453 13719
rect 20453 13685 20487 13719
rect 20487 13685 20496 13719
rect 20444 13676 20496 13685
rect 21180 13719 21232 13728
rect 21180 13685 21189 13719
rect 21189 13685 21223 13719
rect 21223 13685 21232 13719
rect 21180 13676 21232 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 9404 13472 9456 13524
rect 9312 13336 9364 13388
rect 14464 13472 14516 13524
rect 16580 13472 16632 13524
rect 18512 13472 18564 13524
rect 19340 13515 19392 13524
rect 19340 13481 19349 13515
rect 19349 13481 19383 13515
rect 19383 13481 19392 13515
rect 19340 13472 19392 13481
rect 20536 13472 20588 13524
rect 12164 13404 12216 13456
rect 12624 13336 12676 13388
rect 15936 13404 15988 13456
rect 14096 13336 14148 13388
rect 11888 13200 11940 13252
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 10048 13132 10100 13184
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 15844 13200 15896 13252
rect 19432 13336 19484 13388
rect 20168 13336 20220 13388
rect 17776 13268 17828 13320
rect 18236 13268 18288 13320
rect 21180 13268 21232 13320
rect 13820 13132 13872 13184
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 16580 13132 16632 13184
rect 20536 13200 20588 13252
rect 18144 13132 18196 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 10048 12928 10100 12980
rect 10232 12928 10284 12980
rect 12716 12928 12768 12980
rect 13912 12928 13964 12980
rect 15752 12928 15804 12980
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 16120 12928 16172 12980
rect 13268 12860 13320 12912
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 8760 12792 8812 12844
rect 9956 12835 10008 12844
rect 9956 12801 9965 12835
rect 9965 12801 9999 12835
rect 9999 12801 10008 12835
rect 9956 12792 10008 12801
rect 10048 12835 10100 12844
rect 10048 12801 10082 12835
rect 10082 12801 10100 12835
rect 10048 12792 10100 12801
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 11152 12724 11204 12776
rect 11244 12724 11296 12776
rect 12624 12724 12676 12776
rect 9404 12656 9456 12708
rect 20444 12928 20496 12980
rect 12808 12656 12860 12708
rect 18512 12792 18564 12844
rect 13728 12724 13780 12776
rect 15936 12724 15988 12776
rect 10600 12588 10652 12640
rect 10692 12588 10744 12640
rect 11612 12631 11664 12640
rect 11612 12597 11621 12631
rect 11621 12597 11655 12631
rect 11655 12597 11664 12631
rect 11612 12588 11664 12597
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 13084 12631 13136 12640
rect 12716 12588 12768 12597
rect 13084 12597 13093 12631
rect 13093 12597 13127 12631
rect 13127 12597 13136 12631
rect 13084 12588 13136 12597
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 17040 12656 17092 12708
rect 15844 12588 15896 12640
rect 18236 12631 18288 12640
rect 18236 12597 18245 12631
rect 18245 12597 18279 12631
rect 18279 12597 18288 12631
rect 18236 12588 18288 12597
rect 18512 12588 18564 12640
rect 19432 12767 19484 12776
rect 19432 12733 19466 12767
rect 19466 12733 19484 12767
rect 19432 12724 19484 12733
rect 19616 12767 19668 12776
rect 19616 12733 19625 12767
rect 19625 12733 19659 12767
rect 19659 12733 19668 12767
rect 19616 12724 19668 12733
rect 18696 12656 18748 12708
rect 20076 12588 20128 12640
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 11428 12384 11480 12436
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 9220 12248 9272 12300
rect 9772 12248 9824 12300
rect 9496 12112 9548 12164
rect 12716 12359 12768 12368
rect 12716 12325 12725 12359
rect 12725 12325 12759 12359
rect 12759 12325 12768 12359
rect 12716 12316 12768 12325
rect 13452 12359 13504 12368
rect 13452 12325 13461 12359
rect 13461 12325 13495 12359
rect 13495 12325 13504 12359
rect 13452 12316 13504 12325
rect 15844 12359 15896 12368
rect 15844 12325 15853 12359
rect 15853 12325 15887 12359
rect 15887 12325 15896 12359
rect 15844 12316 15896 12325
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 20260 12316 20312 12368
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 10692 12248 10744 12300
rect 11612 12248 11664 12300
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 16120 12291 16172 12300
rect 16120 12257 16129 12291
rect 16129 12257 16163 12291
rect 16163 12257 16172 12291
rect 16120 12248 16172 12257
rect 19616 12248 19668 12300
rect 20076 12248 20128 12300
rect 20536 12248 20588 12300
rect 11244 12112 11296 12164
rect 9864 12044 9916 12096
rect 10600 12044 10652 12096
rect 13728 12112 13780 12164
rect 16212 12223 16264 12232
rect 16212 12189 16246 12223
rect 16246 12189 16264 12223
rect 16212 12180 16264 12189
rect 18788 12180 18840 12232
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 16672 12044 16724 12096
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4620 11500 4672 11552
rect 20628 11840 20680 11892
rect 6920 11772 6972 11824
rect 10232 11772 10284 11824
rect 9772 11636 9824 11688
rect 10140 11679 10192 11688
rect 10140 11645 10149 11679
rect 10149 11645 10183 11679
rect 10183 11645 10192 11679
rect 10140 11636 10192 11645
rect 11888 11679 11940 11688
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 12900 11636 12952 11645
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 16212 11636 16264 11688
rect 17500 11679 17552 11688
rect 17500 11645 17509 11679
rect 17509 11645 17543 11679
rect 17543 11645 17552 11679
rect 17500 11636 17552 11645
rect 17776 11636 17828 11688
rect 5264 11500 5316 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 11796 11500 11848 11552
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 15660 11500 15712 11552
rect 17868 11500 17920 11552
rect 20536 11500 20588 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3884 11296 3936 11348
rect 4620 11296 4672 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 4712 11160 4764 11212
rect 5264 11092 5316 11144
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 7288 11135 7340 11144
rect 5540 11092 5592 11101
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 9680 11296 9732 11348
rect 10232 11296 10284 11348
rect 10784 11296 10836 11348
rect 11152 11296 11204 11348
rect 11612 11296 11664 11348
rect 13452 11296 13504 11348
rect 13820 11296 13872 11348
rect 14832 11296 14884 11348
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 18604 11339 18656 11348
rect 18604 11305 18613 11339
rect 18613 11305 18647 11339
rect 18647 11305 18656 11339
rect 18604 11296 18656 11305
rect 19248 11296 19300 11348
rect 19984 11339 20036 11348
rect 19984 11305 19993 11339
rect 19993 11305 20027 11339
rect 20027 11305 20036 11339
rect 19984 11296 20036 11305
rect 10968 11228 11020 11280
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 14096 11160 14148 11212
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 5448 11024 5500 11076
rect 6184 11024 6236 11076
rect 8300 11024 8352 11076
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 5172 10956 5224 11008
rect 5632 10956 5684 11008
rect 9772 11024 9824 11076
rect 10324 11024 10376 11076
rect 11796 11024 11848 11076
rect 13544 11024 13596 11076
rect 15200 11160 15252 11212
rect 21364 11296 21416 11348
rect 20628 11203 20680 11212
rect 20628 11169 20637 11203
rect 20637 11169 20671 11203
rect 20671 11169 20680 11203
rect 20628 11160 20680 11169
rect 14924 11092 14976 11144
rect 17776 11092 17828 11144
rect 17868 11092 17920 11144
rect 20352 11135 20404 11144
rect 20352 11101 20361 11135
rect 20361 11101 20395 11135
rect 20395 11101 20404 11135
rect 20352 11092 20404 11101
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 10876 10999 10928 11008
rect 10876 10965 10885 10999
rect 10885 10965 10919 10999
rect 10919 10965 10928 10999
rect 10876 10956 10928 10965
rect 15568 11067 15620 11076
rect 15568 11033 15602 11067
rect 15602 11033 15620 11067
rect 15568 11024 15620 11033
rect 15660 11024 15712 11076
rect 16580 11024 16632 11076
rect 16120 10956 16172 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 8300 10752 8352 10804
rect 10140 10752 10192 10804
rect 10876 10752 10928 10804
rect 11428 10752 11480 10804
rect 11888 10752 11940 10804
rect 5540 10684 5592 10736
rect 10692 10684 10744 10736
rect 5172 10659 5224 10668
rect 5172 10625 5181 10659
rect 5181 10625 5215 10659
rect 5215 10625 5224 10659
rect 5172 10616 5224 10625
rect 5264 10616 5316 10668
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 4804 10548 4856 10600
rect 6000 10616 6052 10668
rect 6920 10616 6972 10668
rect 8944 10616 8996 10668
rect 15476 10684 15528 10736
rect 16212 10795 16264 10804
rect 16212 10761 16221 10795
rect 16221 10761 16255 10795
rect 16255 10761 16264 10795
rect 16212 10752 16264 10761
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 17868 10727 17920 10736
rect 17868 10693 17877 10727
rect 17877 10693 17911 10727
rect 17911 10693 17920 10727
rect 17868 10684 17920 10693
rect 13176 10616 13228 10668
rect 14096 10616 14148 10668
rect 14924 10616 14976 10668
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 18604 10616 18656 10668
rect 4712 10480 4764 10532
rect 5264 10480 5316 10532
rect 5356 10480 5408 10532
rect 10968 10548 11020 10600
rect 10876 10480 10928 10532
rect 11336 10548 11388 10600
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 13544 10548 13596 10600
rect 6368 10412 6420 10464
rect 9772 10412 9824 10464
rect 10232 10412 10284 10464
rect 15200 10412 15252 10464
rect 20536 10591 20588 10600
rect 20536 10557 20545 10591
rect 20545 10557 20579 10591
rect 20579 10557 20588 10591
rect 20536 10548 20588 10557
rect 17316 10455 17368 10464
rect 17316 10421 17325 10455
rect 17325 10421 17359 10455
rect 17359 10421 17368 10455
rect 17316 10412 17368 10421
rect 21180 10455 21232 10464
rect 21180 10421 21189 10455
rect 21189 10421 21223 10455
rect 21223 10421 21232 10455
rect 21180 10412 21232 10421
rect 21548 10455 21600 10464
rect 21548 10421 21557 10455
rect 21557 10421 21591 10455
rect 21591 10421 21600 10455
rect 21548 10412 21600 10421
rect 38384 10412 38436 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4712 10208 4764 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 5540 10208 5592 10260
rect 6368 10208 6420 10260
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 9956 10208 10008 10260
rect 11980 10208 12032 10260
rect 12900 10251 12952 10260
rect 12900 10217 12909 10251
rect 12909 10217 12943 10251
rect 12943 10217 12952 10251
rect 12900 10208 12952 10217
rect 13452 10208 13504 10260
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 4620 10004 4672 10056
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 13820 10072 13872 10124
rect 17316 10208 17368 10260
rect 17868 10208 17920 10260
rect 20352 10208 20404 10260
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 20628 10140 20680 10192
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 20168 10072 20220 10124
rect 13912 10004 13964 10056
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 19984 10004 20036 10056
rect 21548 10208 21600 10260
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 5172 9936 5224 9988
rect 5264 9979 5316 9988
rect 5264 9945 5273 9979
rect 5273 9945 5307 9979
rect 5307 9945 5316 9979
rect 5264 9936 5316 9945
rect 13176 9936 13228 9988
rect 20168 9936 20220 9988
rect 5540 9868 5592 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 10968 9868 11020 9920
rect 14832 9868 14884 9920
rect 15752 9911 15804 9920
rect 15752 9877 15761 9911
rect 15761 9877 15795 9911
rect 15795 9877 15804 9911
rect 15752 9868 15804 9877
rect 17040 9868 17092 9920
rect 17960 9868 18012 9920
rect 19432 9868 19484 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4896 9664 4948 9716
rect 7196 9664 7248 9716
rect 10600 9664 10652 9716
rect 16764 9707 16816 9716
rect 16764 9673 16773 9707
rect 16773 9673 16807 9707
rect 16807 9673 16816 9707
rect 16764 9664 16816 9673
rect 5356 9596 5408 9648
rect 5908 9596 5960 9648
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 13176 9596 13228 9648
rect 15568 9596 15620 9648
rect 17776 9596 17828 9648
rect 20168 9707 20220 9716
rect 20168 9673 20177 9707
rect 20177 9673 20211 9707
rect 20211 9673 20220 9707
rect 20168 9664 20220 9673
rect 21364 9664 21416 9716
rect 21180 9596 21232 9648
rect 3976 9460 4028 9512
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 8760 9528 8812 9580
rect 9772 9528 9824 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 13452 9528 13504 9580
rect 14832 9528 14884 9580
rect 15200 9528 15252 9580
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 17960 9528 18012 9580
rect 19800 9528 19852 9580
rect 9588 9503 9640 9512
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 9496 9392 9548 9444
rect 10784 9460 10836 9512
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 9772 9392 9824 9444
rect 9956 9392 10008 9444
rect 17500 9460 17552 9512
rect 3608 9324 3660 9376
rect 4712 9324 4764 9376
rect 5448 9324 5500 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 14740 9367 14792 9376
rect 14740 9333 14749 9367
rect 14749 9333 14783 9367
rect 14783 9333 14792 9367
rect 14740 9324 14792 9333
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 17224 9324 17276 9376
rect 17684 9460 17736 9512
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 18604 9503 18656 9512
rect 18604 9469 18638 9503
rect 18638 9469 18656 9503
rect 18604 9460 18656 9469
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 19524 9503 19576 9512
rect 18328 9392 18380 9444
rect 19524 9469 19533 9503
rect 19533 9469 19567 9503
rect 19567 9469 19576 9503
rect 19524 9460 19576 9469
rect 19340 9324 19392 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4896 9120 4948 9172
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 11244 9120 11296 9172
rect 13912 9120 13964 9172
rect 16764 9120 16816 9172
rect 4620 9052 4672 9104
rect 4988 9052 5040 9104
rect 6000 9052 6052 9104
rect 5356 8984 5408 9036
rect 5448 8984 5500 9036
rect 7748 8984 7800 9036
rect 9220 8984 9272 9036
rect 10048 8984 10100 9036
rect 10600 8984 10652 9036
rect 17684 9120 17736 9172
rect 18604 9120 18656 9172
rect 19524 9120 19576 9172
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 5172 8916 5224 8968
rect 5632 8916 5684 8968
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 13084 8984 13136 9036
rect 13544 8984 13596 9036
rect 13452 8916 13504 8968
rect 16580 8916 16632 8968
rect 17040 8916 17092 8968
rect 19064 8916 19116 8968
rect 19800 8916 19852 8968
rect 5356 8848 5408 8900
rect 10968 8848 11020 8900
rect 3884 8823 3936 8832
rect 3884 8789 3899 8823
rect 3899 8789 3933 8823
rect 3933 8789 3936 8823
rect 3884 8780 3936 8789
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 5080 8780 5132 8832
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 11336 8780 11388 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 15568 8848 15620 8900
rect 20076 8848 20128 8900
rect 17224 8780 17276 8832
rect 19984 8780 20036 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3608 8576 3660 8628
rect 3884 8576 3936 8628
rect 3976 8576 4028 8628
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 4712 8576 4764 8628
rect 4804 8576 4856 8628
rect 4988 8619 5040 8628
rect 4988 8585 4997 8619
rect 4997 8585 5031 8619
rect 5031 8585 5040 8619
rect 4988 8576 5040 8585
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5356 8576 5408 8628
rect 9588 8576 9640 8628
rect 11888 8576 11940 8628
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5080 8440 5132 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 5540 8440 5592 8492
rect 13268 8576 13320 8628
rect 15016 8576 15068 8628
rect 17224 8576 17276 8628
rect 18328 8576 18380 8628
rect 19340 8576 19392 8628
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 14740 8440 14792 8492
rect 19432 8483 19484 8492
rect 19432 8449 19441 8483
rect 19441 8449 19475 8483
rect 19475 8449 19484 8483
rect 19432 8440 19484 8449
rect 1400 8236 1452 8288
rect 5080 8304 5132 8356
rect 8300 8372 8352 8424
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 11612 8415 11664 8424
rect 11612 8381 11621 8415
rect 11621 8381 11655 8415
rect 11655 8381 11664 8415
rect 11612 8372 11664 8381
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 15292 8372 15344 8424
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 20260 8415 20312 8424
rect 20260 8381 20269 8415
rect 20269 8381 20303 8415
rect 20303 8381 20312 8415
rect 20260 8372 20312 8381
rect 5632 8304 5684 8356
rect 10784 8304 10836 8356
rect 18788 8304 18840 8356
rect 19340 8304 19392 8356
rect 5172 8236 5224 8288
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 12164 8236 12216 8245
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 20904 8279 20956 8288
rect 20904 8245 20913 8279
rect 20913 8245 20947 8279
rect 20947 8245 20956 8279
rect 20904 8236 20956 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5172 8032 5224 8084
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 4896 7964 4948 8016
rect 6552 8032 6604 8084
rect 8852 7964 8904 8016
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 5448 7828 5500 7880
rect 6460 7828 6512 7880
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 8668 7828 8720 7880
rect 12256 8032 12308 8084
rect 15292 8032 15344 8084
rect 18328 8032 18380 8084
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 9772 7896 9824 7948
rect 13084 8007 13136 8016
rect 13084 7973 13093 8007
rect 13093 7973 13127 8007
rect 13127 7973 13136 8007
rect 13084 7964 13136 7973
rect 10784 7896 10836 7948
rect 3884 7803 3936 7812
rect 3884 7769 3893 7803
rect 3893 7769 3927 7803
rect 3927 7769 3936 7803
rect 3884 7760 3936 7769
rect 2504 7692 2556 7744
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 4988 7692 5040 7744
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 12164 7828 12216 7880
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13636 7828 13688 7880
rect 15476 7828 15528 7880
rect 16304 7896 16356 7948
rect 10048 7692 10100 7744
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 11152 7692 11204 7744
rect 12808 7692 12860 7744
rect 15108 7760 15160 7812
rect 14924 7692 14976 7744
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 19064 7828 19116 7880
rect 20904 7828 20956 7880
rect 18328 7760 18380 7812
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 18052 7692 18104 7744
rect 22008 7735 22060 7744
rect 22008 7701 22017 7735
rect 22017 7701 22051 7735
rect 22051 7701 22060 7735
rect 22008 7692 22060 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2688 7488 2740 7540
rect 3424 7488 3476 7540
rect 3976 7488 4028 7540
rect 4620 7488 4672 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 9404 7488 9456 7540
rect 9772 7488 9824 7540
rect 10140 7488 10192 7540
rect 11060 7488 11112 7540
rect 11612 7488 11664 7540
rect 12900 7488 12952 7540
rect 17684 7488 17736 7540
rect 17960 7488 18012 7540
rect 19156 7488 19208 7540
rect 20260 7531 20312 7540
rect 20260 7497 20269 7531
rect 20269 7497 20303 7531
rect 20303 7497 20312 7531
rect 20260 7488 20312 7497
rect 22008 7488 22060 7540
rect 1400 7284 1452 7336
rect 6460 7420 6512 7472
rect 6552 7420 6604 7472
rect 2504 7352 2556 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3884 7352 3936 7404
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 4988 7352 5040 7404
rect 3516 7284 3568 7336
rect 5448 7148 5500 7200
rect 6920 7352 6972 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 11244 7352 11296 7404
rect 10600 7284 10652 7336
rect 9220 7216 9272 7268
rect 12808 7284 12860 7336
rect 13636 7352 13688 7404
rect 12992 7284 13044 7336
rect 14372 7284 14424 7336
rect 15108 7352 15160 7404
rect 15384 7352 15436 7404
rect 15476 7352 15528 7404
rect 6736 7148 6788 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10232 7191 10284 7200
rect 10232 7157 10241 7191
rect 10241 7157 10275 7191
rect 10275 7157 10284 7191
rect 10232 7148 10284 7157
rect 11244 7191 11296 7200
rect 11244 7157 11253 7191
rect 11253 7157 11287 7191
rect 11287 7157 11296 7191
rect 11244 7148 11296 7157
rect 13084 7216 13136 7268
rect 14924 7148 14976 7200
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 19156 7395 19208 7404
rect 19156 7361 19190 7395
rect 19190 7361 19208 7395
rect 19156 7352 19208 7361
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 19984 7352 20036 7404
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18512 7284 18564 7336
rect 18788 7259 18840 7268
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 20628 7216 20680 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3148 6944 3200 6996
rect 6920 6944 6972 6996
rect 15292 6944 15344 6996
rect 2596 6919 2648 6928
rect 2596 6885 2605 6919
rect 2605 6885 2639 6919
rect 2639 6885 2648 6919
rect 2596 6876 2648 6885
rect 4620 6876 4672 6928
rect 9588 6876 9640 6928
rect 8668 6808 8720 6860
rect 9496 6808 9548 6860
rect 14924 6876 14976 6928
rect 3424 6740 3476 6792
rect 3516 6740 3568 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 5540 6740 5592 6792
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 9864 6740 9916 6792
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 11152 6808 11204 6860
rect 14004 6808 14056 6860
rect 10324 6740 10376 6792
rect 12716 6740 12768 6792
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 14648 6783 14700 6792
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 17132 6987 17184 6996
rect 17132 6953 17141 6987
rect 17141 6953 17175 6987
rect 17175 6953 17184 6987
rect 17132 6944 17184 6953
rect 18144 6944 18196 6996
rect 20444 6944 20496 6996
rect 17960 6808 18012 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 10876 6672 10928 6724
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 10784 6604 10836 6656
rect 11428 6647 11480 6656
rect 11428 6613 11437 6647
rect 11437 6613 11471 6647
rect 11471 6613 11480 6647
rect 11428 6604 11480 6613
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 18144 6740 18196 6792
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 20168 6672 20220 6724
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 17776 6604 17828 6656
rect 18512 6604 18564 6656
rect 20076 6647 20128 6656
rect 20076 6613 20085 6647
rect 20085 6613 20119 6647
rect 20119 6613 20128 6647
rect 20076 6604 20128 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 6276 6400 6328 6452
rect 6644 6400 6696 6452
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 9496 6400 9548 6452
rect 5540 6264 5592 6316
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 6460 6264 6512 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 4620 6196 4672 6248
rect 10324 6400 10376 6452
rect 10692 6400 10744 6452
rect 10784 6400 10836 6452
rect 12440 6400 12492 6452
rect 17040 6400 17092 6452
rect 11244 6332 11296 6384
rect 7380 6264 7432 6316
rect 7104 6196 7156 6248
rect 10876 6196 10928 6248
rect 12072 6264 12124 6316
rect 12992 6332 13044 6384
rect 13268 6332 13320 6384
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 14648 6264 14700 6316
rect 12716 6128 12768 6180
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 15292 6239 15344 6248
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 15476 6196 15528 6248
rect 18512 6400 18564 6452
rect 20076 6400 20128 6452
rect 20444 6443 20496 6452
rect 20444 6409 20453 6443
rect 20453 6409 20487 6443
rect 20487 6409 20496 6443
rect 20444 6400 20496 6409
rect 17776 6332 17828 6384
rect 19892 6264 19944 6316
rect 18144 6196 18196 6248
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 12900 6060 12952 6112
rect 16672 6128 16724 6180
rect 15292 6060 15344 6112
rect 17592 6103 17644 6112
rect 17592 6069 17601 6103
rect 17601 6069 17635 6103
rect 17635 6069 17644 6103
rect 17592 6060 17644 6069
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5356 5856 5408 5908
rect 7380 5856 7432 5908
rect 10140 5856 10192 5908
rect 11428 5856 11480 5908
rect 15660 5856 15712 5908
rect 18604 5856 18656 5908
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 3516 5788 3568 5840
rect 5540 5788 5592 5840
rect 3424 5720 3476 5772
rect 6552 5720 6604 5772
rect 2780 5652 2832 5704
rect 4252 5652 4304 5704
rect 5172 5652 5224 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 6460 5652 6512 5704
rect 3976 5584 4028 5636
rect 11152 5652 11204 5704
rect 12992 5788 13044 5840
rect 11980 5652 12032 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 13636 5831 13688 5840
rect 13636 5797 13645 5831
rect 13645 5797 13679 5831
rect 13679 5797 13688 5831
rect 13636 5788 13688 5797
rect 14004 5652 14056 5704
rect 15200 5652 15252 5704
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 4160 5516 4212 5568
rect 6920 5516 6972 5568
rect 11704 5516 11756 5568
rect 11796 5559 11848 5568
rect 11796 5525 11805 5559
rect 11805 5525 11839 5559
rect 11839 5525 11848 5559
rect 11796 5516 11848 5525
rect 16672 5584 16724 5636
rect 17592 5652 17644 5704
rect 21180 5856 21232 5908
rect 19892 5763 19944 5772
rect 19892 5729 19901 5763
rect 19901 5729 19935 5763
rect 19935 5729 19944 5763
rect 19892 5720 19944 5729
rect 20168 5720 20220 5772
rect 15384 5516 15436 5568
rect 38752 5516 38804 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 3056 5312 3108 5364
rect 3424 5312 3476 5364
rect 4160 5244 4212 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2136 5176 2188 5228
rect 5448 5312 5500 5364
rect 6368 5312 6420 5364
rect 12808 5312 12860 5364
rect 15384 5355 15436 5364
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 6828 5244 6880 5296
rect 4252 5108 4304 5160
rect 4068 5040 4120 5092
rect 5080 5108 5132 5160
rect 5632 5108 5684 5160
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11796 5176 11848 5228
rect 15660 5312 15712 5364
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 3792 4972 3844 5024
rect 4160 4972 4212 5024
rect 4896 5040 4948 5092
rect 6460 5040 6512 5092
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 12532 5108 12584 5160
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 14832 5108 14884 5160
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 2872 4768 2924 4820
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 4068 4768 4120 4820
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 2596 4632 2648 4684
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 11888 4768 11940 4820
rect 13728 4768 13780 4820
rect 14740 4768 14792 4820
rect 15568 4768 15620 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 16948 4768 17000 4820
rect 4620 4564 4672 4616
rect 4896 4632 4948 4684
rect 10232 4700 10284 4752
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 11980 4700 12032 4752
rect 12716 4700 12768 4752
rect 7564 4564 7616 4616
rect 9496 4564 9548 4616
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 11612 4564 11664 4616
rect 13544 4564 13596 4616
rect 14188 4564 14240 4616
rect 5448 4496 5500 4548
rect 9220 4496 9272 4548
rect 11980 4496 12032 4548
rect 12072 4496 12124 4548
rect 15108 4632 15160 4684
rect 15476 4607 15528 4616
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 18052 4564 18104 4616
rect 4804 4428 4856 4480
rect 5356 4428 5408 4480
rect 7012 4428 7064 4480
rect 7932 4428 7984 4480
rect 9864 4471 9916 4480
rect 9864 4437 9873 4471
rect 9873 4437 9907 4471
rect 9907 4437 9916 4471
rect 9864 4428 9916 4437
rect 10600 4471 10652 4480
rect 10600 4437 10609 4471
rect 10609 4437 10643 4471
rect 10643 4437 10652 4471
rect 10600 4428 10652 4437
rect 10968 4428 11020 4480
rect 12532 4428 12584 4480
rect 13360 4471 13412 4480
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 5356 4088 5408 4140
rect 7012 4224 7064 4276
rect 7196 4224 7248 4276
rect 7288 4224 7340 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 11244 4224 11296 4276
rect 14188 4224 14240 4276
rect 14832 4224 14884 4276
rect 6644 4088 6696 4140
rect 7748 4156 7800 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7380 4088 7432 4140
rect 8116 4131 8168 4140
rect 8116 4097 8150 4131
rect 8150 4097 8168 4131
rect 8116 4088 8168 4097
rect 10968 4156 11020 4208
rect 12072 4156 12124 4208
rect 11612 4131 11664 4140
rect 11612 4097 11621 4131
rect 11621 4097 11655 4131
rect 11655 4097 11664 4131
rect 11612 4088 11664 4097
rect 12624 4156 12676 4208
rect 12900 4199 12952 4208
rect 12900 4165 12909 4199
rect 12909 4165 12943 4199
rect 12943 4165 12952 4199
rect 12900 4156 12952 4165
rect 4620 4020 4672 4072
rect 4988 4063 5040 4072
rect 4988 4029 4997 4063
rect 4997 4029 5031 4063
rect 5031 4029 5040 4063
rect 4988 4020 5040 4029
rect 2596 3952 2648 4004
rect 3056 3995 3108 4004
rect 3056 3961 3065 3995
rect 3065 3961 3099 3995
rect 3099 3961 3108 3995
rect 3056 3952 3108 3961
rect 5448 3952 5500 4004
rect 5540 3952 5592 4004
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6736 3952 6788 4004
rect 7748 4020 7800 4072
rect 7380 3952 7432 4004
rect 7564 3952 7616 4004
rect 6828 3884 6880 3936
rect 7472 3884 7524 3936
rect 11704 3952 11756 4004
rect 10140 3884 10192 3936
rect 12532 3952 12584 4004
rect 12808 4020 12860 4072
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 14556 4088 14608 4140
rect 15108 4156 15160 4208
rect 15292 4088 15344 4140
rect 16764 4088 16816 4140
rect 13268 3952 13320 4004
rect 13360 3995 13412 4004
rect 13360 3961 13369 3995
rect 13369 3961 13403 3995
rect 13403 3961 13412 3995
rect 14924 4063 14976 4072
rect 14924 4029 14934 4063
rect 14934 4029 14968 4063
rect 14968 4029 14976 4063
rect 14924 4020 14976 4029
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 13360 3952 13412 3961
rect 12348 3884 12400 3936
rect 12716 3884 12768 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 15292 3884 15344 3936
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 6368 3680 6420 3732
rect 5172 3612 5224 3664
rect 5540 3655 5592 3664
rect 5540 3621 5549 3655
rect 5549 3621 5583 3655
rect 5583 3621 5592 3655
rect 5540 3612 5592 3621
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 1032 3476 1084 3528
rect 1768 3476 1820 3528
rect 2412 3519 2464 3528
rect 2412 3485 2421 3519
rect 2421 3485 2455 3519
rect 2455 3485 2464 3519
rect 2412 3476 2464 3485
rect 4712 3544 4764 3596
rect 2044 3408 2096 3460
rect 3608 3519 3660 3528
rect 3608 3485 3617 3519
rect 3617 3485 3651 3519
rect 3651 3485 3660 3519
rect 3608 3476 3660 3485
rect 2136 3340 2188 3392
rect 4068 3408 4120 3460
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5080 3476 5132 3528
rect 5356 3476 5408 3528
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 7748 3680 7800 3732
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 7196 3544 7248 3596
rect 7840 3612 7892 3664
rect 8116 3680 8168 3732
rect 3424 3383 3476 3392
rect 3424 3349 3433 3383
rect 3433 3349 3467 3383
rect 3467 3349 3476 3383
rect 3424 3340 3476 3349
rect 5172 3340 5224 3392
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7472 3476 7524 3528
rect 7932 3476 7984 3528
rect 13544 3680 13596 3732
rect 14188 3680 14240 3732
rect 10140 3612 10192 3664
rect 12900 3612 12952 3664
rect 14556 3680 14608 3732
rect 16764 3723 16816 3732
rect 16764 3689 16773 3723
rect 16773 3689 16807 3723
rect 16807 3689 16816 3723
rect 16764 3680 16816 3689
rect 10416 3476 10468 3528
rect 6920 3340 6972 3392
rect 7104 3340 7156 3392
rect 9864 3340 9916 3392
rect 10324 3340 10376 3392
rect 11336 3408 11388 3460
rect 12532 3451 12584 3460
rect 12532 3417 12541 3451
rect 12541 3417 12575 3451
rect 12575 3417 12584 3451
rect 12532 3408 12584 3417
rect 13176 3476 13228 3528
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 15016 3451 15068 3460
rect 15016 3417 15025 3451
rect 15025 3417 15059 3451
rect 15059 3417 15068 3451
rect 15016 3408 15068 3417
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15384 3476 15436 3528
rect 16212 3476 16264 3528
rect 10508 3340 10560 3392
rect 14832 3340 14884 3392
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 15476 3340 15528 3392
rect 15660 3340 15712 3392
rect 20168 3544 20220 3596
rect 19340 3519 19392 3528
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 17592 3340 17644 3392
rect 28080 3519 28132 3528
rect 28080 3485 28089 3519
rect 28089 3485 28123 3519
rect 28123 3485 28132 3519
rect 28080 3476 28132 3485
rect 32128 3544 32180 3596
rect 28448 3408 28500 3460
rect 28540 3408 28592 3460
rect 26516 3340 26568 3392
rect 27528 3340 27580 3392
rect 37004 3340 37056 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3884 3136 3936 3188
rect 4068 3136 4120 3188
rect 5080 3136 5132 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 5356 3136 5408 3188
rect 6644 3179 6696 3188
rect 6644 3145 6653 3179
rect 6653 3145 6687 3179
rect 6687 3145 6696 3179
rect 6644 3136 6696 3145
rect 6920 3136 6972 3188
rect 7380 3136 7432 3188
rect 5540 3111 5592 3120
rect 5540 3077 5549 3111
rect 5549 3077 5583 3111
rect 5583 3077 5592 3111
rect 5540 3068 5592 3077
rect 7564 3068 7616 3120
rect 8116 3136 8168 3188
rect 2780 2932 2832 2984
rect 1584 2864 1636 2916
rect 3884 2932 3936 2984
rect 5264 3000 5316 3052
rect 7104 2932 7156 2984
rect 7656 3000 7708 3052
rect 9680 3068 9732 3120
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9864 3068 9916 3120
rect 9496 3000 9548 3009
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 11796 3111 11848 3120
rect 11796 3077 11805 3111
rect 11805 3077 11839 3111
rect 11839 3077 11848 3111
rect 11796 3068 11848 3077
rect 12072 3043 12124 3052
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 14924 3136 14976 3188
rect 16120 3136 16172 3188
rect 16212 3136 16264 3188
rect 19340 3136 19392 3188
rect 20168 3136 20220 3188
rect 7012 2864 7064 2916
rect 2504 2796 2556 2848
rect 5264 2796 5316 2848
rect 5448 2839 5500 2848
rect 5448 2805 5457 2839
rect 5457 2805 5491 2839
rect 5491 2805 5500 2839
rect 5448 2796 5500 2805
rect 7288 2796 7340 2848
rect 11888 2975 11940 2984
rect 11888 2941 11897 2975
rect 11897 2941 11931 2975
rect 11931 2941 11940 2975
rect 11888 2932 11940 2941
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 9772 2864 9824 2916
rect 10324 2864 10376 2916
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 12164 2796 12216 2848
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 15016 2932 15068 2984
rect 17592 3000 17644 3052
rect 21456 3068 21508 3120
rect 26424 3068 26476 3120
rect 26792 3179 26844 3188
rect 26792 3145 26801 3179
rect 26801 3145 26835 3179
rect 26835 3145 26844 3179
rect 26792 3136 26844 3145
rect 28080 3136 28132 3188
rect 29000 3136 29052 3188
rect 35348 3068 35400 3120
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 18788 2932 18840 2984
rect 20168 2975 20220 2984
rect 20168 2941 20177 2975
rect 20177 2941 20211 2975
rect 20211 2941 20220 2975
rect 20168 2932 20220 2941
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 23664 2864 23716 2916
rect 26516 3043 26568 3052
rect 26516 3009 26525 3043
rect 26525 3009 26559 3043
rect 26559 3009 26568 3043
rect 26516 3000 26568 3009
rect 27528 3000 27580 3052
rect 28448 3043 28500 3052
rect 28448 3009 28457 3043
rect 28457 3009 28491 3043
rect 28491 3009 28500 3043
rect 28448 3000 28500 3009
rect 28540 3000 28592 3052
rect 28724 3043 28776 3052
rect 28724 3009 28733 3043
rect 28733 3009 28767 3043
rect 28767 3009 28776 3043
rect 28724 3000 28776 3009
rect 28908 3000 28960 3052
rect 32312 3000 32364 3052
rect 37004 3179 37056 3188
rect 37004 3145 37013 3179
rect 37013 3145 37047 3179
rect 37047 3145 37056 3179
rect 37004 3136 37056 3145
rect 29092 2975 29144 2984
rect 29092 2941 29101 2975
rect 29101 2941 29135 2975
rect 29135 2941 29144 2975
rect 29092 2932 29144 2941
rect 33508 2975 33560 2984
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 38016 2932 38068 2984
rect 20996 2796 21048 2848
rect 25412 2796 25464 2848
rect 30104 2796 30156 2848
rect 33692 2839 33744 2848
rect 33692 2805 33701 2839
rect 33701 2805 33735 2839
rect 33735 2805 33744 2839
rect 33692 2796 33744 2805
rect 37556 2796 37608 2848
rect 39304 2796 39356 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2504 2592 2556 2644
rect 2780 2567 2832 2576
rect 2780 2533 2789 2567
rect 2789 2533 2823 2567
rect 2823 2533 2832 2567
rect 2780 2524 2832 2533
rect 3608 2635 3660 2644
rect 3608 2601 3617 2635
rect 3617 2601 3651 2635
rect 3651 2601 3660 2635
rect 3608 2592 3660 2601
rect 4712 2592 4764 2644
rect 7012 2592 7064 2644
rect 7380 2592 7432 2644
rect 9496 2524 9548 2576
rect 9680 2592 9732 2644
rect 11888 2592 11940 2644
rect 12164 2635 12216 2644
rect 12164 2601 12173 2635
rect 12173 2601 12207 2635
rect 12207 2601 12216 2635
rect 12164 2592 12216 2601
rect 12072 2524 12124 2576
rect 16764 2592 16816 2644
rect 18788 2592 18840 2644
rect 20168 2592 20220 2644
rect 20996 2635 21048 2644
rect 20996 2601 21005 2635
rect 21005 2601 21039 2635
rect 21039 2601 21048 2635
rect 20996 2592 21048 2601
rect 21456 2592 21508 2644
rect 23664 2592 23716 2644
rect 25136 2592 25188 2644
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 26424 2592 26476 2644
rect 28724 2592 28776 2644
rect 29092 2592 29144 2644
rect 30104 2635 30156 2644
rect 30104 2601 30113 2635
rect 30113 2601 30147 2635
rect 30147 2601 30156 2635
rect 30104 2592 30156 2601
rect 32312 2592 32364 2644
rect 33508 2592 33560 2644
rect 33692 2592 33744 2644
rect 35348 2635 35400 2644
rect 35348 2601 35357 2635
rect 35357 2601 35391 2635
rect 35391 2601 35400 2635
rect 35348 2592 35400 2601
rect 36452 2635 36504 2644
rect 36452 2601 36461 2635
rect 36461 2601 36495 2635
rect 36495 2601 36504 2635
rect 36452 2592 36504 2601
rect 37556 2635 37608 2644
rect 37556 2601 37565 2635
rect 37565 2601 37599 2635
rect 37599 2601 37608 2635
rect 37556 2592 37608 2601
rect 38016 2635 38068 2644
rect 38016 2601 38025 2635
rect 38025 2601 38059 2635
rect 38059 2601 38068 2635
rect 38016 2592 38068 2601
rect 1676 2388 1728 2440
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 3424 2456 3476 2508
rect 5264 2499 5316 2508
rect 5264 2465 5273 2499
rect 5273 2465 5307 2499
rect 5307 2465 5316 2499
rect 5264 2456 5316 2465
rect 6828 2456 6880 2508
rect 8208 2456 8260 2508
rect 11796 2456 11848 2508
rect 4252 2388 4304 2440
rect 4344 2388 4396 2440
rect 5816 2388 5868 2440
rect 8116 2388 8168 2440
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 8944 2431 8996 2440
rect 8944 2397 8953 2431
rect 8953 2397 8987 2431
rect 8987 2397 8996 2431
rect 8944 2388 8996 2397
rect 9772 2388 9824 2440
rect 10048 2388 10100 2440
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 10968 2388 11020 2440
rect 11704 2388 11756 2440
rect 12072 2388 12124 2440
rect 12808 2388 12860 2440
rect 13176 2388 13228 2440
rect 13912 2388 13964 2440
rect 14372 2388 14424 2440
rect 29368 2524 29420 2576
rect 32128 2567 32180 2576
rect 32128 2533 32137 2567
rect 32137 2533 32171 2567
rect 32171 2533 32180 2567
rect 32128 2524 32180 2533
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16212 2388 16264 2440
rect 17224 2388 17276 2440
rect 17592 2388 17644 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 18328 2388 18380 2440
rect 18696 2388 18748 2440
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 2504 2252 2556 2304
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 20812 2431 20864 2440
rect 20812 2397 20821 2431
rect 20821 2397 20855 2431
rect 20855 2397 20864 2431
rect 20812 2388 20864 2397
rect 20904 2388 20956 2440
rect 21640 2388 21692 2440
rect 22284 2431 22336 2440
rect 22284 2397 22293 2431
rect 22293 2397 22327 2431
rect 22327 2397 22336 2431
rect 22284 2388 22336 2397
rect 22744 2388 22796 2440
rect 23112 2388 23164 2440
rect 23848 2388 23900 2440
rect 24216 2388 24268 2440
rect 24952 2388 25004 2440
rect 25320 2388 25372 2440
rect 26148 2388 26200 2440
rect 26424 2388 26476 2440
rect 27160 2388 27212 2440
rect 27528 2388 27580 2440
rect 28264 2388 28316 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 29920 2320 29972 2372
rect 30472 2388 30524 2440
rect 30840 2388 30892 2440
rect 31576 2388 31628 2440
rect 31944 2388 31996 2440
rect 32680 2388 32732 2440
rect 33048 2388 33100 2440
rect 33784 2388 33836 2440
rect 34152 2388 34204 2440
rect 34888 2388 34940 2440
rect 35256 2388 35308 2440
rect 35992 2388 36044 2440
rect 36360 2388 36412 2440
rect 37096 2388 37148 2440
rect 37556 2388 37608 2440
rect 38292 2388 38344 2440
rect 38568 2320 38620 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 4252 2048 4304 2100
rect 15384 2048 15436 2100
rect 16488 1368 16540 1420
rect 18144 1368 18196 1420
<< metal2 >>
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 38108 35012 38160 35018
rect 38108 34954 38160 34960
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 38120 34649 38148 34954
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38106 34640 38162 34649
rect 38106 34575 38162 34584
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 38016 25152 38068 25158
rect 38016 25094 38068 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 7392 12850 7420 14350
rect 8128 14074 8156 14894
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 8680 14346 8708 14758
rect 8864 14618 8892 14758
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 9324 13394 9352 14214
rect 9416 14074 9444 14758
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 7392 12434 7420 12786
rect 8772 12442 8800 12786
rect 9416 12714 9444 13466
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9416 12458 9444 12650
rect 7300 12406 7420 12434
rect 8760 12436 8812 12442
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 3896 11354 3924 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 11494
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10062 4660 11290
rect 4724 11218 4752 11698
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 5276 11150 5304 11494
rect 6932 11354 6960 11766
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4816 10606 4844 10950
rect 5184 10674 5212 10950
rect 5276 10674 5304 11086
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 5276 10538 5304 10610
rect 5368 10538 5396 11086
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 10674 5488 11018
rect 5552 10742 5580 11086
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 4724 10266 4752 10474
rect 5276 10418 5304 10474
rect 5276 10390 5396 10418
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 8634 3648 9318
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8634 3924 8774
rect 3988 8634 4016 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9110 4660 9998
rect 4908 9722 4936 10202
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 8634 4200 8910
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7342 1440 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7410 2544 7686
rect 2700 7546 2728 7822
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 5234 1440 7278
rect 3160 7002 3188 7346
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 2596 6928 2648 6934
rect 2596 6870 2648 6876
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 2148 4826 2176 5170
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2608 4690 2636 6870
rect 3436 6798 3464 7482
rect 3896 7410 3924 7754
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7546 4016 7686
rect 4632 7546 4660 9046
rect 4724 8634 4752 9318
rect 4908 9178 4936 9454
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8634 4844 8774
rect 5000 8634 5028 9046
rect 5184 8974 5212 9930
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4908 8022 4936 8434
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 5000 7954 5028 8570
rect 5092 8498 5120 8774
rect 5184 8634 5212 8910
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5184 8378 5212 8570
rect 5092 8362 5212 8378
rect 5080 8356 5212 8362
rect 5132 8350 5212 8356
rect 5080 8298 5132 8304
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 8090 5212 8230
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 5000 7410 5028 7686
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3528 6798 3556 7278
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6934 4660 7346
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3436 5778 3464 6734
rect 3528 5846 3556 6734
rect 4632 6254 4660 6870
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5370 2820 5646
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5370 3096 5510
rect 3436 5370 3464 5714
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3528 5166 3556 5782
rect 5276 5710 5304 9930
rect 5368 9654 5396 10390
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5460 9382 5488 10610
rect 5552 10266 5580 10678
rect 5644 10674 5672 10950
rect 6196 10810 6224 11018
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6932 10674 6960 11290
rect 7300 11150 7328 12406
rect 8760 12378 8812 12384
rect 9324 12430 9444 12458
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8312 10810 8340 11018
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8956 10674 8984 10950
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9586 5580 9862
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 9194 5488 9318
rect 5368 9166 5488 9194
rect 5368 9042 5396 9166
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8650 5396 8842
rect 5460 8786 5488 8978
rect 5920 8974 5948 9590
rect 6012 9110 6040 10610
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10266 6408 10406
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6380 9586 6408 10202
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9722 7236 9998
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 6012 8974 6040 9046
rect 7760 9042 7788 9862
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 9178 8800 9522
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 9232 9042 9260 12242
rect 9324 10266 9352 12430
rect 9508 12170 9536 13806
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9600 11234 9628 13670
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12306 9812 13126
rect 9968 12850 9996 14554
rect 10612 14278 10640 14894
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10888 14618 10916 14758
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 11348 14482 11376 14758
rect 11808 14618 11836 15438
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15026 12572 15302
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 12912 14482 12940 14758
rect 14108 14482 14136 15030
rect 14476 14822 14504 15982
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15162 14596 15438
rect 14752 15162 14780 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15120 15094 15148 15302
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12986 10088 13126
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10060 12850 10088 12922
rect 10244 12850 10272 12922
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11354 9720 11494
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9508 11218 9628 11234
rect 9496 11212 9628 11218
rect 9548 11206 9628 11212
rect 9496 11154 9548 11160
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9508 10146 9536 11154
rect 9784 11082 9812 11630
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9416 10118 9536 10146
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5460 8758 5580 8786
rect 5368 8634 5488 8650
rect 5356 8628 5488 8634
rect 5408 8622 5488 8628
rect 5356 8570 5408 8576
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5368 5914 5396 8434
rect 5460 7886 5488 8622
rect 5552 8498 5580 8758
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5644 8362 5672 8910
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 6564 8090 6592 8774
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6472 7478 6500 7822
rect 6564 7478 6592 8026
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 5460 6798 5488 7142
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 2884 4826 2912 4966
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 1688 3602 1716 4626
rect 3804 4622 3832 4966
rect 3988 4826 4016 5578
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5302 4200 5510
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4080 4826 4108 5034
rect 4172 5030 4200 5238
rect 4264 5166 4292 5646
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4632 4078 4660 4558
rect 4816 4486 4844 4966
rect 4908 4690 4936 5034
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4146 4844 4422
rect 5092 4196 5120 5102
rect 5184 4298 5212 5646
rect 5460 5370 5488 6734
rect 5552 6322 5580 6734
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6458 6316 6598
rect 6656 6458 6684 6734
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 5552 5846 5580 6258
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5184 4270 5304 4298
rect 5092 4168 5212 4196
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4620 4072 4672 4078
rect 3054 4040 3110 4049
rect 2596 4004 2648 4010
rect 4620 4014 4672 4020
rect 3054 3975 3056 3984
rect 2596 3946 2648 3952
rect 3108 3975 3110 3984
rect 3056 3946 3108 3952
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1032 3528 1084 3534
rect 1032 3470 1084 3476
rect 662 3360 718 3369
rect 662 3295 718 3304
rect 676 800 704 3295
rect 1044 800 1072 3470
rect 1584 2916 1636 2922
rect 1584 2858 1636 2864
rect 1596 1578 1624 2858
rect 1688 2446 1716 3538
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1412 1550 1624 1578
rect 1412 800 1440 1550
rect 1780 800 1808 3470
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2056 2446 2084 3402
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2148 2446 2176 3334
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2148 870 2268 898
rect 2148 800 2176 870
rect 662 0 718 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2240 762 2268 870
rect 2424 762 2452 3470
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 2650 2544 2790
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 2608 2446 2636 3946
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3882 3632 3938 3641
rect 3882 3567 3938 3576
rect 4712 3596 4764 3602
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2792 2582 2820 2926
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 3436 2514 3464 3334
rect 3620 2650 3648 3470
rect 3896 3194 3924 3567
rect 4712 3538 4764 3544
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 3194 4108 3402
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3896 2774 3924 2926
rect 3712 2746 3924 2774
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 2596 2440 2648 2446
rect 2964 2440 3016 2446
rect 2596 2382 2648 2388
rect 2884 2400 2964 2428
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 800 2544 2246
rect 2884 800 2912 2400
rect 2964 2382 3016 2388
rect 3712 1442 3740 2746
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2650 4752 3538
rect 4816 3534 4844 4082
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5000 3534 5028 4014
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5092 3534 5120 3878
rect 5184 3670 5212 4168
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5092 3194 5120 3470
rect 5184 3398 5212 3606
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5276 3194 5304 4270
rect 5368 4146 5396 4422
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5368 3534 5396 4082
rect 5460 4010 5488 4490
rect 5552 4010 5580 5782
rect 5644 5166 5672 6258
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5370 6408 6054
rect 6472 5710 6500 6258
rect 6564 5778 6592 6258
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 6472 5098 6500 5646
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6748 4690 6776 7142
rect 6932 7002 6960 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7392 6322 7420 7822
rect 8312 7546 8340 8366
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7886 8708 8230
rect 8864 8022 8892 8366
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 6866 8708 7346
rect 9232 7274 9260 8978
rect 9416 8514 9444 10118
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9450 9536 9998
rect 9784 9586 9812 10406
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9600 8634 9628 9454
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9416 8486 9628 8514
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7546 9444 8230
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6458 8800 6598
rect 9324 6458 9352 7346
rect 9600 6934 9628 8486
rect 9784 7954 9812 9386
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7546 9812 7890
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9876 7324 9904 12038
rect 10244 11830 10272 12786
rect 10612 12646 10640 14214
rect 10704 14074 10732 14214
rect 11256 14074 11284 14282
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 12306 10732 12582
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10612 12102 10640 12242
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10152 10810 10180 11630
rect 10244 11354 10272 11766
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10244 10470 10272 11086
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9968 9450 9996 10202
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10060 9042 10088 9862
rect 10336 9586 10364 11018
rect 10612 9722 10640 12038
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 10742 10732 11494
rect 11164 11354 11192 12718
rect 11256 12170 11284 12718
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10612 9042 10640 9658
rect 10796 9518 10824 11290
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10810 10916 10950
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10980 10606 11008 11222
rect 11348 10606 11376 14418
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11440 13870 11468 14214
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11440 12442 11468 13806
rect 12176 13462 12204 13806
rect 12360 13802 12388 14418
rect 12912 14226 12940 14418
rect 13084 14272 13136 14278
rect 12912 14198 13032 14226
rect 13084 14214 13136 14220
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11440 10810 11468 12378
rect 11624 12306 11652 12582
rect 11900 12442 11928 13194
rect 12636 12782 12664 13330
rect 12728 12986 12756 13670
rect 13004 13326 13032 14198
rect 13096 13734 13124 14214
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12624 12776 12676 12782
rect 12676 12724 12848 12730
rect 12624 12718 12848 12724
rect 12636 12714 12848 12718
rect 12636 12708 12860 12714
rect 12636 12702 12808 12708
rect 12808 12650 12860 12656
rect 13096 12646 13124 13670
rect 14108 13394 14136 14418
rect 14476 13530 14504 14758
rect 16132 14278 16160 14894
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17328 14618 17356 14758
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13280 12918 13308 13262
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 12728 12374 12756 12582
rect 12716 12368 12768 12374
rect 12716 12310 12768 12316
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9784 7296 9904 7324
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6458 9536 6802
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5386 6960 5510
rect 6840 5358 6960 5386
rect 6840 5302 6868 5358
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6840 4298 6868 5238
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6748 4270 6868 4298
rect 7024 4282 7052 4422
rect 7012 4276 7064 4282
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5446 3768 5502 3777
rect 5446 3703 5502 3712
rect 5460 3534 5488 3703
rect 5552 3670 5580 3946
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3738 6408 3878
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5368 3194 5396 3470
rect 6656 3194 6684 4082
rect 6748 4010 6776 4270
rect 7012 4218 7064 4224
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6840 3942 6868 4082
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 7116 3602 7144 6190
rect 7392 5914 7420 6258
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7208 3602 7236 4218
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7012 3528 7064 3534
rect 7300 3482 7328 4218
rect 7392 4146 7420 5850
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7576 4010 7604 4558
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7748 4208 7800 4214
rect 7800 4168 7880 4196
rect 7748 4150 7800 4156
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7392 3534 7420 3946
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3534 7512 3878
rect 7064 3476 7328 3482
rect 7012 3470 7328 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7024 3454 7328 3470
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6932 3194 6960 3334
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 5540 3120 5592 3126
rect 5538 3088 5540 3097
rect 5592 3088 5594 3097
rect 5264 3052 5316 3058
rect 5538 3023 5594 3032
rect 5264 2994 5316 3000
rect 5276 2854 5304 2994
rect 7116 2990 7144 3334
rect 7576 3210 7604 3946
rect 7760 3738 7788 4014
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7852 3670 7880 4168
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7944 3534 7972 4422
rect 9232 4282 9260 4490
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8128 3738 8156 4082
rect 8758 3904 8814 3913
rect 8758 3839 8814 3848
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 7932 3528 7984 3534
rect 7392 3194 7604 3210
rect 7380 3188 7604 3194
rect 7432 3182 7604 3188
rect 7668 3488 7932 3516
rect 7380 3130 7432 3136
rect 7564 3120 7616 3126
rect 7392 3068 7564 3074
rect 7392 3062 7616 3068
rect 7392 3046 7604 3062
rect 7668 3058 7696 3488
rect 7932 3470 7984 3476
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7656 3052 7708 3058
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 5264 2848 5316 2854
rect 5448 2848 5500 2854
rect 5264 2790 5316 2796
rect 5446 2816 5448 2825
rect 5500 2816 5502 2825
rect 5446 2751 5502 2760
rect 7024 2650 7052 2858
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4264 2106 4292 2382
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 3620 1414 3740 1442
rect 3620 800 3648 1414
rect 4356 800 4384 2382
rect 5276 1170 5304 2450
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5092 1142 5304 1170
rect 5092 800 5120 1142
rect 5828 800 5856 2382
rect 6564 870 6684 898
rect 6564 800 6592 870
rect 2240 734 2452 762
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6656 762 6684 870
rect 6840 762 6868 2450
rect 7300 800 7328 2790
rect 7392 2650 7420 3046
rect 7656 2994 7708 3000
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 8128 2446 8156 3130
rect 8772 2922 8800 3839
rect 9508 3058 9536 4558
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8220 1170 8248 2450
rect 8484 2440 8536 2446
rect 8864 2428 8892 2790
rect 9692 2650 9720 3062
rect 9784 2922 9812 7296
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6798 9904 7142
rect 10060 6866 10088 7686
rect 10152 7546 10180 7822
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10612 7342 10640 8978
rect 10796 8362 10824 9454
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10796 7954 10824 8298
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 10060 5930 10088 6802
rect 10060 5914 10180 5930
rect 10060 5908 10192 5914
rect 10060 5902 10140 5908
rect 10140 5850 10192 5856
rect 10244 4758 10272 7142
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6458 10364 6734
rect 10888 6730 10916 10474
rect 10980 9926 11008 10542
rect 11624 10130 11652 11290
rect 11808 11082 11836 11494
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11900 10810 11928 11630
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10266 12020 10542
rect 12912 10266 12940 11630
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 13188 9994 13216 10610
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 8906 11008 9862
rect 13188 9654 13216 9930
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9178 11284 9318
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11072 7546 11100 7686
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 6866 11192 7686
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11256 7206 11284 7346
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10704 6458 10732 6598
rect 10796 6458 10824 6598
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10888 6254 10916 6666
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 11164 5710 11192 6802
rect 11256 6390 11284 7142
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 9876 3641 9904 4422
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3670 10180 3878
rect 10612 3777 10640 4422
rect 10980 4214 11008 4422
rect 11256 4282 11284 4558
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 10598 3768 10654 3777
rect 10598 3703 10654 3712
rect 10140 3664 10192 3670
rect 9862 3632 9918 3641
rect 10140 3606 10192 3612
rect 9862 3567 9918 3576
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 9876 3126 9904 3334
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 10336 2922 10364 3334
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10428 2854 10456 3470
rect 11348 3466 11376 8774
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11440 5914 11468 6598
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 10508 3392 10560 3398
rect 11532 3369 11560 9522
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8634 11928 8774
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 11624 7546 11652 8366
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7886 12204 8230
rect 12268 8090 12296 8366
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 12820 7342 12848 7686
rect 12912 7546 12940 8230
rect 13096 8022 13124 8978
rect 13280 8922 13308 12582
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13464 11354 13492 12310
rect 13740 12170 13768 12718
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13464 10266 13492 11290
rect 13556 11082 13584 11494
rect 13832 11354 13860 13126
rect 13924 12986 13952 13126
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13556 10130 13584 10542
rect 13832 10130 13860 11290
rect 14108 11218 14136 13330
rect 15212 12306 15240 14214
rect 16592 14074 16620 14214
rect 16776 14074 16804 14486
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17328 14074 17356 14282
rect 17604 14278 17632 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 38028 14482 38056 25094
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 38016 14476 38068 14482
rect 38016 14418 38068 14424
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17696 14074 17724 14350
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 16592 13530 16620 14010
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12986 15792 13126
rect 15856 12986 15884 13194
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15948 12782 15976 13398
rect 16592 13190 16620 13466
rect 17788 13326 17816 13942
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 18156 13190 18184 13670
rect 18248 13326 18276 14214
rect 18524 13530 18552 14350
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19076 14074 19104 14214
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19352 13530 19380 14350
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 16132 12986 16160 13126
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 12374 15884 12582
rect 15948 12434 15976 12718
rect 15948 12406 16160 12434
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 16132 12306 16160 12406
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16224 11694 16252 12174
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 14844 11354 14872 11630
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 14108 10674 14136 11154
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14936 10674 14964 11086
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 15212 10470 15240 11154
rect 15488 10742 15516 11494
rect 15672 11082 15700 11494
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13464 8974 13492 9522
rect 13556 9042 13584 10066
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9178 13952 9998
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14844 9586 14872 9862
rect 15212 9738 15240 10406
rect 15212 9710 15332 9738
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13188 8894 13308 8922
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13004 7342 13032 7822
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 6458 12480 6598
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11716 5234 11744 5510
rect 11808 5234 11836 5510
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4146 11652 4558
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11716 4010 11744 5170
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4826 11928 4966
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11992 4758 12020 5646
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11992 4554 12020 4694
rect 12084 4554 12112 6258
rect 12728 6186 12756 6734
rect 12820 6304 12848 7278
rect 13004 6390 13032 7278
rect 13096 7274 13124 7958
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12900 6316 12952 6322
rect 12820 6276 12900 6304
rect 12716 6180 12768 6186
rect 12716 6122 12768 6128
rect 12728 5710 12756 6122
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12820 5370 12848 6276
rect 12900 6258 12952 6264
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 4570 12572 5102
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 12360 4542 12572 4570
rect 12084 4214 12112 4490
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 12360 3942 12388 4542
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4010 12572 4422
rect 12636 4214 12664 4966
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12728 3942 12756 4694
rect 12820 4078 12848 5306
rect 12912 4214 12940 6054
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 13004 4078 13032 5782
rect 13188 4298 13216 8894
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8634 13308 8774
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 14752 8498 14780 9318
rect 15028 8634 15056 9454
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7410 13676 7822
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13096 4270 13216 4298
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 13004 3754 13032 4014
rect 13096 3913 13124 4270
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13082 3904 13138 3913
rect 13082 3839 13138 3848
rect 12912 3726 13032 3754
rect 12912 3670 12940 3726
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 13188 3534 13216 4082
rect 13280 4010 13308 6326
rect 13648 5846 13676 7346
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 14016 5710 14044 6802
rect 14384 6798 14412 7278
rect 14936 7206 14964 7686
rect 15120 7410 15148 7754
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14936 6934 14964 7142
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14660 6322 14688 6734
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13740 4826 13768 4966
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13372 4010 13400 4422
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13556 3738 13584 4558
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13176 3528 13228 3534
rect 12530 3496 12586 3505
rect 13176 3470 13228 3476
rect 12530 3431 12532 3440
rect 12584 3431 12586 3440
rect 12532 3402 12584 3408
rect 10508 3334 10560 3340
rect 11518 3360 11574 3369
rect 10520 3097 10548 3334
rect 11518 3295 11574 3304
rect 11796 3120 11848 3126
rect 10506 3088 10562 3097
rect 11796 3062 11848 3068
rect 10506 3023 10508 3032
rect 10560 3023 10562 3032
rect 10508 2994 10560 3000
rect 9956 2848 10008 2854
rect 10416 2848 10468 2854
rect 9956 2790 10008 2796
rect 10414 2816 10416 2825
rect 10468 2816 10470 2825
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9496 2576 9548 2582
rect 9968 2530 9996 2790
rect 10414 2751 10470 2760
rect 9496 2518 9548 2524
rect 8944 2440 8996 2446
rect 8864 2400 8944 2428
rect 8484 2382 8536 2388
rect 8944 2382 8996 2388
rect 8036 1142 8248 1170
rect 8036 800 8064 1142
rect 6656 734 6868 762
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8496 762 8524 2382
rect 8680 870 8800 898
rect 8680 762 8708 870
rect 8772 800 8800 870
rect 9508 800 9536 2518
rect 9784 2502 9996 2530
rect 11808 2514 11836 3062
rect 14016 3058 14044 5646
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14752 4826 14780 5102
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 4282 14228 4558
rect 14844 4282 14872 5102
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3738 14228 3878
rect 14568 3738 14596 4082
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14844 3482 14872 4218
rect 14936 4078 14964 6870
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 6254 15148 6734
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 4690 15148 6190
rect 15212 5710 15240 9522
rect 15304 8430 15332 9710
rect 15580 9654 15608 11018
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16132 10062 16160 10950
rect 16224 10810 16252 11630
rect 16592 11082 16620 13126
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 17052 12442 17080 12650
rect 17040 12436 17092 12442
rect 18156 12434 18184 13126
rect 18524 12850 18552 13466
rect 19444 13394 19472 14418
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 14074 20024 14214
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20548 14006 20576 14418
rect 38212 14278 38240 34886
rect 39028 25084 39080 25090
rect 39028 25026 39080 25032
rect 39040 24857 39068 25026
rect 39026 24848 39082 24857
rect 39026 24783 39082 24792
rect 38384 15360 38436 15366
rect 38384 15302 38436 15308
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 19432 12776 19484 12782
rect 18524 12714 18736 12730
rect 19260 12724 19432 12730
rect 19260 12718 19484 12724
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 18524 12708 18748 12714
rect 18524 12702 18696 12708
rect 18524 12646 18552 12702
rect 18696 12650 18748 12656
rect 19260 12702 19472 12718
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 17040 12378 17092 12384
rect 17972 12406 18184 12434
rect 18248 12434 18276 12582
rect 18248 12406 18368 12434
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11354 16712 12038
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16684 10674 16712 11290
rect 17512 10810 17540 11630
rect 17788 11150 17816 11630
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 11150 17908 11494
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17328 10266 17356 10406
rect 17880 10266 17908 10678
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17972 10146 18000 12406
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 17604 10118 18276 10146
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15764 9586 15792 9862
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 8906 15608 9318
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15304 8090 15332 8366
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15304 7002 15332 8026
rect 16316 7954 16344 10066
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16776 9722 16804 9998
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16580 8968 16632 8974
rect 16632 8916 16712 8922
rect 16580 8910 16712 8916
rect 16592 8894 16712 8910
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7410 15516 7822
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15292 6248 15344 6254
rect 15396 6236 15424 7346
rect 15488 6254 15516 7346
rect 16684 7342 16712 8894
rect 16776 8430 16804 9114
rect 17052 8974 17080 9862
rect 17604 9602 17632 10118
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17512 9574 17632 9602
rect 17512 9518 17540 9574
rect 17696 9518 17724 9998
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17788 9518 17816 9590
rect 17972 9586 18000 9862
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17236 8838 17264 9318
rect 17696 9178 17724 9454
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8634 17264 8774
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15344 6208 15424 6236
rect 15476 6248 15528 6254
rect 15292 6190 15344 6196
rect 15476 6190 15528 6196
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 15120 4078 15148 4150
rect 15304 4146 15332 6054
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5370 15424 5510
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15488 4622 15516 6190
rect 15672 5914 15700 6734
rect 16684 6186 16712 7278
rect 17144 7002 17172 7822
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17696 7546 17724 7686
rect 17972 7546 18000 7822
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 18064 6882 18092 7686
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 7002 18184 7278
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17972 6866 18092 6882
rect 18248 6866 18276 10118
rect 18340 9450 18368 12406
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18616 10674 18644 11290
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18800 9518 18828 12174
rect 19260 11354 19288 12702
rect 19628 12306 19656 12718
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12306 20116 12582
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11354 20024 12174
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20180 10146 20208 13330
rect 20456 12986 20484 13670
rect 20548 13530 20576 13942
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20548 13258 20576 13466
rect 21192 13326 21220 13670
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20272 12374 20300 12582
rect 20548 12458 20576 13194
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 20456 12434 20576 12458
rect 20364 12430 20576 12434
rect 20364 12406 20484 12430
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20364 11150 20392 12406
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20548 11558 20576 12242
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 20640 11898 20668 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 21376 11354 21404 12038
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20364 10266 20392 11086
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 10266 20576 10542
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20640 10198 20668 11154
rect 38396 10470 38424 15302
rect 38936 15224 38988 15230
rect 38936 15166 38988 15172
rect 38948 15065 38976 15166
rect 38934 15056 38990 15065
rect 38934 14991 38990 15000
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 38384 10464 38436 10470
rect 38384 10406 38436 10412
rect 20628 10192 20680 10198
rect 20180 10130 20300 10146
rect 20628 10134 20680 10140
rect 20168 10124 20300 10130
rect 20220 10118 20300 10124
rect 20168 10066 20220 10072
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 8634 18368 9386
rect 18616 9178 18644 9454
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18340 8090 18368 8570
rect 18800 8362 18828 9454
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18340 7410 18368 7754
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18524 6866 18552 7278
rect 18800 7274 18828 8026
rect 19076 7886 19104 8910
rect 19352 8634 19380 9318
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19444 8498 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19536 9178 19564 9454
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19812 8974 19840 9522
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19996 8838 20024 9998
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20180 9722 20208 9930
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20088 8634 20116 8842
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20272 8514 20300 10118
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 20180 8486 20300 8514
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 17960 6860 18092 6866
rect 18012 6854 18092 6860
rect 18236 6860 18288 6866
rect 17960 6802 18012 6808
rect 18236 6802 18288 6808
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18524 6746 18552 6802
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17052 6458 17080 6598
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17788 6390 17816 6598
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 18156 6254 18184 6734
rect 18524 6718 18644 6746
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 6458 18552 6598
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15672 5370 15700 5850
rect 16684 5642 16712 6122
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 5710 17632 6054
rect 18616 5914 18644 6718
rect 19076 6254 19104 7822
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19168 7410 19196 7482
rect 19352 7410 19380 8298
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19444 5914 19472 6734
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19892 6316 19944 6322
rect 19996 6304 20024 7346
rect 20180 6730 20208 8486
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20272 7546 20300 8366
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20640 7274 20668 10134
rect 21192 9654 21220 10406
rect 21560 10266 21588 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21376 9722 21404 9998
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7886 20944 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 22020 7546 22048 7686
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20088 6458 20116 6598
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19944 6276 20024 6304
rect 19892 6258 19944 6264
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19904 5778 19932 6258
rect 20180 5778 20208 6666
rect 20456 6458 20484 6938
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21192 5914 21220 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 16684 5234 16712 5578
rect 38752 5568 38804 5574
rect 38752 5510 38804 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 38764 5273 38792 5510
rect 38750 5264 38806 5273
rect 16672 5228 16724 5234
rect 38750 5199 38806 5208
rect 16672 5170 16724 5176
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4826 15608 4966
rect 15856 4826 15884 5102
rect 16960 4826 16988 5102
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 18064 4622 18092 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15658 4040 15714 4049
rect 15658 3975 15714 3984
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15304 3534 15332 3878
rect 15292 3528 15344 3534
rect 14844 3466 15056 3482
rect 15292 3470 15344 3476
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 14844 3460 15068 3466
rect 14844 3454 15016 3460
rect 15016 3402 15068 3408
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14844 3074 14872 3334
rect 14936 3194 14964 3334
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 14004 3052 14056 3058
rect 14844 3046 15056 3074
rect 14004 2994 14056 3000
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11900 2650 11928 2926
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12084 2582 12112 2994
rect 15028 2990 15056 3046
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 12176 2650 12204 2790
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 11796 2508 11848 2514
rect 9784 2446 9812 2502
rect 11796 2450 11848 2456
rect 14292 2502 14412 2530
rect 9772 2440 9824 2446
rect 10048 2440 10100 2446
rect 9772 2382 9824 2388
rect 9876 2400 10048 2428
rect 9876 800 9904 2400
rect 10048 2382 10100 2388
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 10612 870 10732 898
rect 10612 800 10640 870
rect 8496 734 8708 762
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10704 762 10732 870
rect 10888 762 10916 2382
rect 10980 800 11008 2382
rect 11716 800 11744 2382
rect 12084 800 12112 2382
rect 12820 800 12848 2382
rect 13188 800 13216 2382
rect 13924 800 13952 2382
rect 14292 800 14320 2502
rect 14384 2446 14412 2502
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14936 1170 14964 2246
rect 15396 2106 15424 3470
rect 15488 3398 15516 3878
rect 15672 3398 15700 3975
rect 16776 3738 16804 4082
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 32128 3596 32180 3602
rect 32128 3538 32180 3544
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15672 2990 15700 3334
rect 16132 3194 16160 3538
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 16224 3194 16252 3470
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 17604 3058 17632 3334
rect 19352 3194 19380 3470
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20180 3194 20208 3538
rect 28080 3528 28132 3534
rect 26790 3496 26846 3505
rect 28080 3470 28132 3476
rect 26790 3431 26846 3440
rect 26516 3392 26568 3398
rect 26516 3334 26568 3340
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 26424 3120 26476 3126
rect 26424 3062 26476 3068
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 16776 2650 16804 2926
rect 18800 2650 18828 2926
rect 20180 2650 20208 2926
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21008 2650 21036 2790
rect 21468 2650 21496 3062
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 23664 2916 23716 2922
rect 23664 2858 23716 2864
rect 23676 2650 23704 2858
rect 25148 2650 25176 2926
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 25424 2650 25452 2790
rect 26436 2650 26464 3062
rect 26528 3058 26556 3334
rect 26804 3194 26832 3431
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 27540 3058 27568 3334
rect 28092 3194 28120 3470
rect 28448 3460 28500 3466
rect 28448 3402 28500 3408
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 28460 3058 28488 3402
rect 28552 3058 28580 3402
rect 28920 3194 29040 3210
rect 28920 3188 29052 3194
rect 28920 3182 29000 3188
rect 28920 3058 28948 3182
rect 29000 3130 29052 3136
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28724 3052 28776 3058
rect 28724 2994 28776 3000
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 28736 2650 28764 2994
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29104 2650 29132 2926
rect 30104 2848 30156 2854
rect 30104 2790 30156 2796
rect 30116 2650 30144 2790
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 26424 2644 26476 2650
rect 26424 2586 26476 2592
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 30104 2644 30156 2650
rect 30104 2586 30156 2592
rect 32140 2582 32168 3538
rect 37004 3392 37056 3398
rect 37004 3334 37056 3340
rect 37016 3194 37044 3334
rect 37004 3188 37056 3194
rect 37004 3130 37056 3136
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 32312 3052 32364 3058
rect 32312 2994 32364 3000
rect 32324 2650 32352 2994
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 33520 2650 33548 2926
rect 33692 2848 33744 2854
rect 33692 2790 33744 2796
rect 33704 2650 33732 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2650 35388 3062
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36464 2650 36492 2994
rect 38016 2984 38068 2990
rect 38016 2926 38068 2932
rect 37556 2848 37608 2854
rect 37556 2790 37608 2796
rect 37568 2650 37596 2790
rect 38028 2650 38056 2926
rect 39304 2848 39356 2854
rect 39304 2790 39356 2796
rect 32312 2644 32364 2650
rect 32312 2586 32364 2592
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 35348 2644 35400 2650
rect 35348 2586 35400 2592
rect 36452 2644 36504 2650
rect 36452 2586 36504 2592
rect 37556 2644 37608 2650
rect 37556 2586 37608 2592
rect 38016 2644 38068 2650
rect 38016 2586 38068 2592
rect 29368 2576 29420 2582
rect 29368 2518 29420 2524
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18696 2440 18748 2446
rect 19524 2440 19576 2446
rect 18696 2382 18748 2388
rect 19444 2400 19524 2428
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15488 1306 15516 2382
rect 16224 1306 16252 2382
rect 16488 1420 16540 1426
rect 16488 1362 16540 1368
rect 15396 1278 15516 1306
rect 16132 1278 16252 1306
rect 14936 1142 15056 1170
rect 15028 800 15056 1142
rect 15396 800 15424 1278
rect 16132 800 16160 1278
rect 16500 800 16528 1362
rect 17236 800 17264 2382
rect 17604 800 17632 2382
rect 18156 1426 18184 2382
rect 18144 1420 18196 1426
rect 18144 1362 18196 1368
rect 18340 800 18368 2382
rect 18708 800 18736 2382
rect 19444 800 19472 2400
rect 19524 2382 19576 2388
rect 19892 2440 19944 2446
rect 20812 2440 20864 2446
rect 19944 2400 20024 2428
rect 19892 2382 19944 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 1306 20024 2400
rect 19812 1278 20024 1306
rect 20548 2400 20812 2428
rect 19812 800 19840 1278
rect 20548 800 20576 2400
rect 20812 2382 20864 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 21640 2440 21692 2446
rect 22284 2440 22336 2446
rect 21640 2382 21692 2388
rect 22020 2400 22284 2428
rect 20916 800 20944 2382
rect 21652 800 21680 2382
rect 22020 800 22048 2400
rect 22284 2382 22336 2388
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 25320 2440 25372 2446
rect 26148 2440 26200 2446
rect 25320 2382 25372 2388
rect 26068 2400 26148 2428
rect 22756 800 22784 2382
rect 23124 800 23152 2382
rect 23860 800 23888 2382
rect 24228 800 24256 2382
rect 24964 800 24992 2382
rect 25332 800 25360 2382
rect 26068 800 26096 2400
rect 26148 2382 26200 2388
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 28264 2440 28316 2446
rect 28724 2440 28776 2446
rect 28264 2382 28316 2388
rect 28644 2400 28724 2428
rect 26436 800 26464 2382
rect 27172 800 27200 2382
rect 27540 800 27568 2382
rect 28276 800 28304 2382
rect 28644 800 28672 2400
rect 28724 2382 28776 2388
rect 29380 800 29408 2518
rect 37476 2502 37596 2530
rect 30472 2440 30524 2446
rect 30472 2382 30524 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 33048 2440 33100 2446
rect 33048 2382 33100 2388
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 37096 2440 37148 2446
rect 37096 2382 37148 2388
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 1306 29960 2314
rect 29748 1278 29960 1306
rect 29748 800 29776 1278
rect 30484 800 30512 2382
rect 30852 800 30880 2382
rect 31588 800 31616 2382
rect 31956 800 31984 2382
rect 32692 800 32720 2382
rect 33060 800 33088 2382
rect 33796 800 33824 2382
rect 34164 800 34192 2382
rect 34900 800 34928 2382
rect 35268 800 35296 2382
rect 36004 800 36032 2382
rect 36372 800 36400 2382
rect 37108 800 37136 2382
rect 37476 800 37504 2502
rect 37568 2446 37596 2502
rect 38212 2502 38332 2530
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 38212 800 38240 2502
rect 38304 2446 38332 2502
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 38568 2372 38620 2378
rect 38568 2314 38620 2320
rect 38580 800 38608 2314
rect 39316 800 39344 2790
rect 10704 734 10916 762
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 38106 34584 38162 34640
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3054 4004 3110 4040
rect 3054 3984 3056 4004
rect 3056 3984 3108 4004
rect 3108 3984 3110 4004
rect 662 3304 718 3360
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3882 3576 3938 3632
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5446 3712 5502 3768
rect 5538 3068 5540 3088
rect 5540 3068 5592 3088
rect 5592 3068 5594 3088
rect 5538 3032 5594 3068
rect 8758 3848 8814 3904
rect 5446 2796 5448 2816
rect 5448 2796 5500 2816
rect 5500 2796 5502 2816
rect 5446 2760 5502 2796
rect 10598 3712 10654 3768
rect 9862 3576 9918 3632
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 13082 3848 13138 3904
rect 12530 3460 12586 3496
rect 12530 3440 12532 3460
rect 12532 3440 12584 3460
rect 12584 3440 12586 3460
rect 11518 3304 11574 3360
rect 10506 3052 10562 3088
rect 10506 3032 10508 3052
rect 10508 3032 10560 3052
rect 10560 3032 10562 3052
rect 10414 2796 10416 2816
rect 10416 2796 10468 2816
rect 10468 2796 10470 2816
rect 10414 2760 10470 2796
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 39026 24792 39082 24848
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38934 15000 38990 15056
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 38750 5208 38806 5264
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 15658 3984 15714 4040
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 26790 3440 26846 3496
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38101 34642 38167 34645
rect 39200 34642 40000 34672
rect 38101 34640 40000 34642
rect 38101 34584 38106 34640
rect 38162 34584 40000 34640
rect 38101 34582 40000 34584
rect 38101 34579 38167 34582
rect 39200 34552 40000 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 39021 24850 39087 24853
rect 39200 24850 40000 24880
rect 39021 24848 40000 24850
rect 39021 24792 39026 24848
rect 39082 24792 40000 24848
rect 39021 24790 40000 24792
rect 39021 24787 39087 24790
rect 39200 24760 40000 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 38929 15058 38995 15061
rect 39200 15058 40000 15088
rect 38929 15056 40000 15058
rect 38929 15000 38934 15056
rect 38990 15000 40000 15056
rect 38929 14998 40000 15000
rect 38929 14995 38995 14998
rect 39200 14968 40000 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 38745 5266 38811 5269
rect 39200 5266 40000 5296
rect 38745 5264 40000 5266
rect 38745 5208 38750 5264
rect 38806 5208 40000 5264
rect 38745 5206 40000 5208
rect 38745 5203 38811 5206
rect 39200 5176 40000 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 3049 4042 3115 4045
rect 15653 4042 15719 4045
rect 3049 4040 15719 4042
rect 3049 3984 3054 4040
rect 3110 3984 15658 4040
rect 15714 3984 15719 4040
rect 3049 3982 15719 3984
rect 3049 3979 3115 3982
rect 15653 3979 15719 3982
rect 8753 3906 8819 3909
rect 13077 3906 13143 3909
rect 8753 3904 13143 3906
rect 8753 3848 8758 3904
rect 8814 3848 13082 3904
rect 13138 3848 13143 3904
rect 8753 3846 13143 3848
rect 8753 3843 8819 3846
rect 13077 3843 13143 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 5441 3770 5507 3773
rect 10593 3770 10659 3773
rect 5441 3768 10659 3770
rect 5441 3712 5446 3768
rect 5502 3712 10598 3768
rect 10654 3712 10659 3768
rect 5441 3710 10659 3712
rect 5441 3707 5507 3710
rect 10593 3707 10659 3710
rect 3877 3634 3943 3637
rect 9857 3634 9923 3637
rect 3877 3632 9923 3634
rect 3877 3576 3882 3632
rect 3938 3576 9862 3632
rect 9918 3576 9923 3632
rect 3877 3574 9923 3576
rect 3877 3571 3943 3574
rect 9857 3571 9923 3574
rect 12525 3498 12591 3501
rect 26785 3498 26851 3501
rect 12525 3496 26851 3498
rect 12525 3440 12530 3496
rect 12586 3440 26790 3496
rect 26846 3440 26851 3496
rect 12525 3438 26851 3440
rect 12525 3435 12591 3438
rect 26785 3435 26851 3438
rect 657 3362 723 3365
rect 11513 3362 11579 3365
rect 657 3360 11579 3362
rect 657 3304 662 3360
rect 718 3304 11518 3360
rect 11574 3304 11579 3360
rect 657 3302 11579 3304
rect 657 3299 723 3302
rect 11513 3299 11579 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 5533 3090 5599 3093
rect 10501 3090 10567 3093
rect 5533 3088 10567 3090
rect 5533 3032 5538 3088
rect 5594 3032 10506 3088
rect 10562 3032 10567 3088
rect 5533 3030 10567 3032
rect 5533 3027 5599 3030
rect 10501 3027 10567 3030
rect 5441 2818 5507 2821
rect 10409 2818 10475 2821
rect 5441 2816 10475 2818
rect 5441 2760 5446 2816
rect 5502 2760 10414 2816
rect 10470 2760 10475 2816
rect 5441 2758 10475 2760
rect 5441 2755 5507 2758
rect 10409 2755 10475 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _125_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 1688980957
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _128_
timestamp 1688980957
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _129_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _130_
timestamp 1688980957
transform 1 0 25024 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _131_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36432 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _132_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _133_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _134_
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _135_
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _136_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _137_
timestamp 1688980957
transform 1 0 19596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _138_
timestamp 1688980957
transform 1 0 17388 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _139_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _140_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _141_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _142_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _143_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _144_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _145_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _146_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _147_
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _148_
timestamp 1688980957
transform 1 0 17572 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _149_
timestamp 1688980957
transform 1 0 11500 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _150_
timestamp 1688980957
transform 1 0 9476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _151_
timestamp 1688980957
transform 1 0 9016 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _152_
timestamp 1688980957
transform 1 0 18400 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _153_
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _154_
timestamp 1688980957
transform 1 0 8924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _155_
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _156_
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1688980957
transform 1 0 13248 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _158_
timestamp 1688980957
transform 1 0 8372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _159_
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_4  _160_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _161_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _162_
timestamp 1688980957
transform 1 0 35696 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _163_
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _164_
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _165_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1688980957
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp 1688980957
transform 1 0 16744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _168_
timestamp 1688980957
transform 1 0 17664 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 1688980957
transform 1 0 15732 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _170_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__nand3b_2  _171_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _172_
timestamp 1688980957
transform 1 0 17112 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1688980957
transform 1 0 15088 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1688980957
transform 1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _175_
timestamp 1688980957
transform 1 0 14444 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _176_
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _177_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 1688980957
transform 1 0 19412 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _179_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _180_
timestamp 1688980957
transform 1 0 19320 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _181_
timestamp 1688980957
transform 1 0 16744 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _182_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _183_
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1688980957
transform 1 0 20516 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _185_
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1688980957
transform 1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _187_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _188_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _189_
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _190_
timestamp 1688980957
transform 1 0 4600 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _191_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _192_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _193_
timestamp 1688980957
transform 1 0 5152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _194_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _195_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _196_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _197_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _198_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _199_
timestamp 1688980957
transform 1 0 4232 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _200_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _201_
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _202_
timestamp 1688980957
transform 1 0 11592 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _203_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _204_
timestamp 1688980957
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _205_
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _206_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _207_
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _208_
timestamp 1688980957
transform 1 0 12972 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_
timestamp 1688980957
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _210_
timestamp 1688980957
transform 1 0 14168 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _211_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_1  _212_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _213_
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _214_
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _215_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _216_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _217_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _219_
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _220_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _221_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _222_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _223_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _225_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _226_
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _227_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1688980957
transform 1 0 6624 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _229_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _230_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _231_
timestamp 1688980957
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _232_
timestamp 1688980957
transform 1 0 6716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _233_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _238_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1688980957
transform 1 0 11592 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor4b_4  _243_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _246_
timestamp 1688980957
transform 1 0 10672 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _247_
timestamp 1688980957
transform 1 0 14536 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _248_
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _250_
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _252_
timestamp 1688980957
transform 1 0 12880 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _253_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _254_
timestamp 1688980957
transform 1 0 16468 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _255_
timestamp 1688980957
transform 1 0 17204 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _256_
timestamp 1688980957
transform 1 0 14260 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _257_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _258_
timestamp 1688980957
transform 1 0 14720 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _259_
timestamp 1688980957
transform 1 0 17204 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _260_
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _261_
timestamp 1688980957
transform 1 0 19044 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _262_
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _263_
timestamp 1688980957
transform 1 0 19044 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _264_
timestamp 1688980957
transform 1 0 14720 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _265_
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _266_
timestamp 1688980957
transform 1 0 20240 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _267_
timestamp 1688980957
transform 1 0 19596 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _268_
timestamp 1688980957
transform 1 0 15272 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _269_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _270_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _271_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _272_
timestamp 1688980957
transform 1 0 2760 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _273_
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _274_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _275_
timestamp 1688980957
transform 1 0 14168 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _276_
timestamp 1688980957
transform 1 0 13984 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _277_
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _278_
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _279_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _280_
timestamp 1688980957
transform 1 0 7820 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _281_
timestamp 1688980957
transform 1 0 7728 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _282_
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _283_
timestamp 1688980957
transform 1 0 7360 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _284_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _285_
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _286_
timestamp 1688980957
transform 1 0 7912 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _287_
timestamp 1688980957
transform 1 0 7360 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _288_
timestamp 1688980957
transform 1 0 10580 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _289_
timestamp 1688980957
transform 1 0 9476 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _290_
timestamp 1688980957
transform 1 0 9108 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _291_
timestamp 1688980957
transform 1 0 9200 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _292_
timestamp 1688980957
transform 1 0 13064 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _293_
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _294_
timestamp 1688980957
transform 1 0 13340 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _295_
timestamp 1688980957
transform 1 0 10948 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _296_
timestamp 1688980957
transform 1 0 12512 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _326__74 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _326_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 13064 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 14168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1688980957
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__S0
timestamp 1688980957
transform 1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__S0
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__S0
timestamp 1688980957
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__S0
timestamp 1688980957
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__S0
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__S0
timestamp 1688980957
transform 1 0 18216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__S0
timestamp 1688980957
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__S0
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A1
timestamp 1688980957
transform 1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A1
timestamp 1688980957
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A1
timestamp 1688980957
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A1
timestamp 1688980957
transform 1 0 16744 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A0
timestamp 1688980957
transform 1 0 16928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A0
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A0
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A0
timestamp 1688980957
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A1
timestamp 1688980957
transform 1 0 20424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A1
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A1
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A1
timestamp 1688980957
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A0
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A0
timestamp 1688980957
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A0
timestamp 1688980957
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A0
timestamp 1688980957
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__D
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A1
timestamp 1688980957
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A1
timestamp 1688980957
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A1
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 1688980957
transform 1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A2
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__C
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1688980957
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A1
timestamp 1688980957
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A1
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A0
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A0
timestamp 1688980957
transform 1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A0
timestamp 1688980957
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A0
timestamp 1688980957
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A1
timestamp 1688980957
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A1
timestamp 1688980957
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A1
timestamp 1688980957
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 1688980957
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A0
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A0
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A0
timestamp 1688980957
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A0
timestamp 1688980957
transform 1 0 12696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold17_A
timestamp 1688980957
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1688980957
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_107 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_123 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_131
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_147
timestamp 1688980957
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_164
timestamp 1688980957
transform 1 0 16192 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_175
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_179
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_186
timestamp 1688980957
transform 1 0 18216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_191
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_219
timestamp 1688980957
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_231
timestamp 1688980957
transform 1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_235
timestamp 1688980957
transform 1 0 22724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_239
timestamp 1688980957
transform 1 0 23092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_243
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_247
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_256
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_263
timestamp 1688980957
transform 1 0 25300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_267
timestamp 1688980957
transform 1 0 25668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_271
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_275
timestamp 1688980957
transform 1 0 26404 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_287
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_291
timestamp 1688980957
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_295
timestamp 1688980957
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_318
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_323
timestamp 1688980957
transform 1 0 30820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_327
timestamp 1688980957
transform 1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_331
timestamp 1688980957
transform 1 0 31556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_340
timestamp 1688980957
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_347
timestamp 1688980957
transform 1 0 33028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_351
timestamp 1688980957
transform 1 0 33396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_355
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_359
timestamp 1688980957
transform 1 0 34132 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_371
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_375
timestamp 1688980957
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_379
timestamp 1688980957
transform 1 0 35972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_383
timestamp 1688980957
transform 1 0 36340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_387
timestamp 1688980957
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 1688980957
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_78
timestamp 1688980957
transform 1 0 8280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_97
timestamp 1688980957
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_106 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_122 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_134
timestamp 1688980957
transform 1 0 13432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_184
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_196
timestamp 1688980957
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_200
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_215 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_257
timestamp 1688980957
transform 1 0 24748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_266
timestamp 1688980957
transform 1 0 25576 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_288
timestamp 1688980957
transform 1 0 27600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_296
timestamp 1688980957
transform 1 0 28336 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_311
timestamp 1688980957
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_323
timestamp 1688980957
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_357
timestamp 1688980957
transform 1 0 33948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_369
timestamp 1688980957
transform 1 0 35052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_375
timestamp 1688980957
transform 1 0 35604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_401
timestamp 1688980957
transform 1 0 37996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_22
timestamp 1688980957
transform 1 0 3128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_58
timestamp 1688980957
transform 1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_74
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_171
timestamp 1688980957
transform 1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_175
timestamp 1688980957
transform 1 0 17204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_187
timestamp 1688980957
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_217
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_229
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_241
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_300
timestamp 1688980957
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_19
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_22
timestamp 1688980957
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_34
timestamp 1688980957
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_45
timestamp 1688980957
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_72
timestamp 1688980957
transform 1 0 7728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_89
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_158
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_12
timestamp 1688980957
transform 1 0 2208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_24
timestamp 1688980957
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_47
timestamp 1688980957
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_59
timestamp 1688980957
transform 1 0 6532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_66
timestamp 1688980957
transform 1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_74
timestamp 1688980957
transform 1 0 7912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1688980957
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_89
timestamp 1688980957
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_96
timestamp 1688980957
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_105
timestamp 1688980957
transform 1 0 10764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_117
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1688980957
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_145
timestamp 1688980957
transform 1 0 14444 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_161
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_28
timestamp 1688980957
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_42
timestamp 1688980957
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_62
timestamp 1688980957
transform 1 0 6808 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_74
timestamp 1688980957
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_98
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1688980957
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_126
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_138
timestamp 1688980957
transform 1 0 13800 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_156
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_188
timestamp 1688980957
transform 1 0 18400 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_200
timestamp 1688980957
transform 1 0 19504 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_212
timestamp 1688980957
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 1688980957
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_70
timestamp 1688980957
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_107
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_118
timestamp 1688980957
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1688980957
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_208
timestamp 1688980957
transform 1 0 20240 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_212
timestamp 1688980957
transform 1 0 20608 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_224
timestamp 1688980957
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_236
timestamp 1688980957
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_248
timestamp 1688980957
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_60
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_88
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_92
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_95
timestamp 1688980957
transform 1 0 9844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1688980957
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_129
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_141
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_157
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_189
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_219
timestamp 1688980957
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_22
timestamp 1688980957
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_48
timestamp 1688980957
transform 1 0 5520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_57
timestamp 1688980957
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_68
timestamp 1688980957
transform 1 0 7360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_113
timestamp 1688980957
transform 1 0 11500 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_124
timestamp 1688980957
transform 1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 1688980957
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_170
timestamp 1688980957
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_187
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_207
timestamp 1688980957
transform 1 0 20148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_219
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_231
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_243
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_26
timestamp 1688980957
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_43
timestamp 1688980957
transform 1 0 5060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_87
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_96
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_108
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_122
timestamp 1688980957
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_131
timestamp 1688980957
transform 1 0 13156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_143
timestamp 1688980957
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_154
timestamp 1688980957
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_206
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_24
timestamp 1688980957
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_33
timestamp 1688980957
transform 1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_46
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_50
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_62
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_125
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_163
timestamp 1688980957
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_171
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_181
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_203
timestamp 1688980957
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_228
timestamp 1688980957
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_240
timestamp 1688980957
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_91
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_103
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_129
timestamp 1688980957
transform 1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_207
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_56
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_60
timestamp 1688980957
transform 1 0 6624 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_72
timestamp 1688980957
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_94
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_98
timestamp 1688980957
transform 1 0 10120 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_110
timestamp 1688980957
transform 1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_122
timestamp 1688980957
transform 1 0 12328 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_126
timestamp 1688980957
transform 1 0 12696 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_136
timestamp 1688980957
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_147
timestamp 1688980957
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_164
timestamp 1688980957
transform 1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_183
timestamp 1688980957
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_187
timestamp 1688980957
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_213
timestamp 1688980957
transform 1 0 20700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_225
timestamp 1688980957
transform 1 0 21804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_237
timestamp 1688980957
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1688980957
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_35
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1688980957
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_44
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1688980957
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_98
timestamp 1688980957
transform 1 0 10120 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_110
timestamp 1688980957
transform 1 0 11224 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_125
timestamp 1688980957
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_178
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_187
timestamp 1688980957
transform 1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_191
timestamp 1688980957
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_206
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_210
timestamp 1688980957
transform 1 0 20424 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_228
timestamp 1688980957
transform 1 0 22080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_240
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_401
timestamp 1688980957
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_42
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_67
timestamp 1688980957
transform 1 0 7268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_75
timestamp 1688980957
transform 1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_86
timestamp 1688980957
transform 1 0 9016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_122
timestamp 1688980957
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_126
timestamp 1688980957
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1688980957
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_177
timestamp 1688980957
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_195
timestamp 1688980957
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_207
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_219
timestamp 1688980957
transform 1 0 21252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1688980957
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1688980957
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_405
timestamp 1688980957
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_94
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 1688980957
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_123
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_174
timestamp 1688980957
transform 1 0 17112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_214
timestamp 1688980957
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_218
timestamp 1688980957
transform 1 0 21160 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_230
timestamp 1688980957
transform 1 0 22264 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_242
timestamp 1688980957
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_401
timestamp 1688980957
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_40
timestamp 1688980957
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_44
timestamp 1688980957
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_85
timestamp 1688980957
transform 1 0 8924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_94
timestamp 1688980957
transform 1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_136
timestamp 1688980957
transform 1 0 13616 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_148
timestamp 1688980957
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_186
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_198
timestamp 1688980957
transform 1 0 19320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1688980957
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_73
timestamp 1688980957
transform 1 0 7820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_94
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_106
timestamp 1688980957
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_118
timestamp 1688980957
transform 1 0 11960 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_128
timestamp 1688980957
transform 1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_132
timestamp 1688980957
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_136
timestamp 1688980957
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_174
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 1688980957
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_401
timestamp 1688980957
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_65
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_84
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_107
timestamp 1688980957
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_123
timestamp 1688980957
transform 1 0 12420 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_141
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_177
timestamp 1688980957
transform 1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_185
timestamp 1688980957
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_209
timestamp 1688980957
transform 1 0 20332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_221
timestamp 1688980957
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1688980957
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_81
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_95
timestamp 1688980957
transform 1 0 9844 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_168
timestamp 1688980957
transform 1 0 16560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_172
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_191
timestamp 1688980957
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_207
timestamp 1688980957
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_211
timestamp 1688980957
transform 1 0 20516 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_223
timestamp 1688980957
transform 1 0 21620 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_235
timestamp 1688980957
transform 1 0 22724 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 1688980957
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_401
timestamp 1688980957
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_77
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_87
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_91
timestamp 1688980957
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_117
timestamp 1688980957
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_127
timestamp 1688980957
transform 1 0 12788 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_132
timestamp 1688980957
transform 1 0 13248 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_136
timestamp 1688980957
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_140
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_144
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_148
timestamp 1688980957
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_152
timestamp 1688980957
transform 1 0 15088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_156
timestamp 1688980957
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_160
timestamp 1688980957
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_177
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_189
timestamp 1688980957
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_219
timestamp 1688980957
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1688980957
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1688980957
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_405
timestamp 1688980957
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_113
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_147
timestamp 1688980957
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_164
timestamp 1688980957
transform 1 0 16192 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_168
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_187
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_206
timestamp 1688980957
transform 1 0 20056 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_218
timestamp 1688980957
transform 1 0 21160 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_230
timestamp 1688980957
transform 1 0 22264 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_242
timestamp 1688980957
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_401
timestamp 1688980957
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_91
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 1688980957
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_155
timestamp 1688980957
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_159
timestamp 1688980957
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_177
timestamp 1688980957
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 1688980957
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 1688980957
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_115
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_124
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1688980957
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 1688980957
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_405
timestamp 1688980957
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1688980957
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_401
timestamp 1688980957
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 1688980957
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 1688980957
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_401
timestamp 1688980957
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1688980957
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_405
timestamp 1688980957
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1688980957
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1688980957
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_401
timestamp 1688980957
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1688980957
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_401
timestamp 1688980957
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_405
timestamp 1688980957
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1688980957
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_401
timestamp 1688980957
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1688980957
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_405
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1688980957
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_401
timestamp 1688980957
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1688980957
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1688980957
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1688980957
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1688980957
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_401
timestamp 1688980957
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 1688980957
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 1688980957
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_405
timestamp 1688980957
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_401
timestamp 1688980957
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_405
timestamp 1688980957
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1688980957
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_401
timestamp 1688980957
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1688980957
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1688980957
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_405
timestamp 1688980957
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1688980957
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1688980957
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_401
timestamp 1688980957
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1688980957
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1688980957
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_405
timestamp 1688980957
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1688980957
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_401
timestamp 1688980957
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1688980957
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1688980957
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_405
timestamp 1688980957
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_401
timestamp 1688980957
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1688980957
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1688980957
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1688980957
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1688980957
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_401
timestamp 1688980957
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1688980957
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1688980957
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1688980957
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_405
timestamp 1688980957
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1688980957
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_401
timestamp 1688980957
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1688980957
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1688980957
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1688980957
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_405
timestamp 1688980957
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1688980957
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1688980957
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_401
timestamp 1688980957
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_401
timestamp 1688980957
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1688980957
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1688980957
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1688980957
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1688980957
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1688980957
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1688980957
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1688980957
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 1688980957
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 1688980957
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1688980957
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_225
timestamp 1688980957
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_237
timestamp 1688980957
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_249
timestamp 1688980957
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 1688980957
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_293
timestamp 1688980957
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 1688980957
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 1688980957
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 1688980957
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 1688980957
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 1688980957
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_405
timestamp 1688980957
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 19872 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 20148 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold9 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  hold10
timestamp 1688980957
transform 1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 28980 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 27968 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 4140 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold20 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold22
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold24
timestamp 1688980957
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 6992 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold27 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform 1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 16100 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 14260 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 10764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 14076 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 10212 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 10028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 20516 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 19412 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 19412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 20516 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 19320 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 8004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 9016 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 8280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold64
timestamp 1688980957
transform 1 0 14352 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 13064 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 21344 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 20516 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 21344 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 20700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 12052 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 11224 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 9384 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 9108 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 18308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 17480 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 17572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 16744 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform 1 0 15364 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1688980957
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1688980957
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input6 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 19596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 20976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 26496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 33120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 34224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 37996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap45
timestamp 1688980957
transform 1 0 17940 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output41 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 1688980957
transform 1 0 4784 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  wire46
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_47
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_48
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_49
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_50
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_51
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_52
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_53
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_54
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_55
timestamp 1688980957
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_56
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_57
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_58
timestamp 1688980957
transform 1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_59
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_60
timestamp 1688980957
transform 1 0 25024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_61
timestamp 1688980957
transform 1 0 26128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_62
timestamp 1688980957
transform 1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_63
timestamp 1688980957
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_64
timestamp 1688980957
transform 1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_65
timestamp 1688980957
transform 1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_66
timestamp 1688980957
transform 1 0 31648 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_67
timestamp 1688980957
transform 1 0 32752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_68
timestamp 1688980957
transform 1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_69
timestamp 1688980957
transform 1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_70
timestamp 1688980957
transform 1 0 36064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_71
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_72
timestamp 1688980957
transform 1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_73
timestamp 1688980957
transform 1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_nn_75
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal3 s 39200 5176 40000 5296 0 FreeSans 480 0 0 0 nn_ids[0]
port 0 nsew signal input
flabel metal3 s 39200 14968 40000 15088 0 FreeSans 480 0 0 0 nn_ids[1]
port 1 nsew signal input
flabel metal3 s 39200 24760 40000 24880 0 FreeSans 480 0 0 0 nn_ids[2]
port 2 nsew signal input
flabel metal3 s 39200 34552 40000 34672 0 FreeSans 480 0 0 0 nn_ids[3]
port 3 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 4 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 5 nsew ground bidirectional
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 wb_clk_i
port 6 nsew signal input
flabel metal2 s 1030 0 1086 800 0 FreeSans 224 90 0 0 wb_rst_i
port 7 nsew signal input
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 8 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 9 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 10 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 11 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 12 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 13 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 14 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 15 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 16 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 17 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 18 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 19 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 20 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 21 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 22 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 23 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 24 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 25 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 26 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 27 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 28 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 29 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 30 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 31 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 32 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 33 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 34 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 35 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 36 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 37 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 38 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 39 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 40 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 41 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 42 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 43 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 44 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 45 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 46 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 47 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 48 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 49 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 50 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 51 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 52 nsew signal input
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 53 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 54 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 55 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 56 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 57 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 58 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 59 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 60 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 61 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 62 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 63 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 64 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 65 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 66 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 67 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 68 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 69 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 70 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 71 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 72 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 73 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 74 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 75 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 76 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 77 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 78 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 79 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 80 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 81 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 82 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 83 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 84 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 85 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 86 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 87 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 88 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 89 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 90 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 91 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 92 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 93 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 94 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 95 nsew signal tristate
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 96 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 97 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 98 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 99 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 100 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 101 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 102 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 103 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 104 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 105 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 106 nsew signal input
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 107 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 108 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 109 nsew signal input
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 110 nsew signal input
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 wbs_we_i
port 111 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
