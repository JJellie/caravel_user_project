// This is the unpowered netlist.
module wishbone_nn (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \fifo_in.FIFO[0][0] ;
 wire \fifo_in.FIFO[0][10] ;
 wire \fifo_in.FIFO[0][11] ;
 wire \fifo_in.FIFO[0][12] ;
 wire \fifo_in.FIFO[0][13] ;
 wire \fifo_in.FIFO[0][14] ;
 wire \fifo_in.FIFO[0][15] ;
 wire \fifo_in.FIFO[0][16] ;
 wire \fifo_in.FIFO[0][17] ;
 wire \fifo_in.FIFO[0][18] ;
 wire \fifo_in.FIFO[0][19] ;
 wire \fifo_in.FIFO[0][1] ;
 wire \fifo_in.FIFO[0][20] ;
 wire \fifo_in.FIFO[0][21] ;
 wire \fifo_in.FIFO[0][22] ;
 wire \fifo_in.FIFO[0][23] ;
 wire \fifo_in.FIFO[0][24] ;
 wire \fifo_in.FIFO[0][25] ;
 wire \fifo_in.FIFO[0][26] ;
 wire \fifo_in.FIFO[0][27] ;
 wire \fifo_in.FIFO[0][28] ;
 wire \fifo_in.FIFO[0][29] ;
 wire \fifo_in.FIFO[0][2] ;
 wire \fifo_in.FIFO[0][30] ;
 wire \fifo_in.FIFO[0][31] ;
 wire \fifo_in.FIFO[0][3] ;
 wire \fifo_in.FIFO[0][4] ;
 wire \fifo_in.FIFO[0][5] ;
 wire \fifo_in.FIFO[0][6] ;
 wire \fifo_in.FIFO[0][7] ;
 wire \fifo_in.FIFO[0][8] ;
 wire \fifo_in.FIFO[0][9] ;
 wire \fifo_in.FIFO[1][0] ;
 wire \fifo_in.FIFO[1][10] ;
 wire \fifo_in.FIFO[1][11] ;
 wire \fifo_in.FIFO[1][12] ;
 wire \fifo_in.FIFO[1][13] ;
 wire \fifo_in.FIFO[1][14] ;
 wire \fifo_in.FIFO[1][15] ;
 wire \fifo_in.FIFO[1][16] ;
 wire \fifo_in.FIFO[1][17] ;
 wire \fifo_in.FIFO[1][18] ;
 wire \fifo_in.FIFO[1][19] ;
 wire \fifo_in.FIFO[1][1] ;
 wire \fifo_in.FIFO[1][20] ;
 wire \fifo_in.FIFO[1][21] ;
 wire \fifo_in.FIFO[1][22] ;
 wire \fifo_in.FIFO[1][23] ;
 wire \fifo_in.FIFO[1][24] ;
 wire \fifo_in.FIFO[1][25] ;
 wire \fifo_in.FIFO[1][26] ;
 wire \fifo_in.FIFO[1][27] ;
 wire \fifo_in.FIFO[1][28] ;
 wire \fifo_in.FIFO[1][29] ;
 wire \fifo_in.FIFO[1][2] ;
 wire \fifo_in.FIFO[1][30] ;
 wire \fifo_in.FIFO[1][31] ;
 wire \fifo_in.FIFO[1][3] ;
 wire \fifo_in.FIFO[1][4] ;
 wire \fifo_in.FIFO[1][5] ;
 wire \fifo_in.FIFO[1][6] ;
 wire \fifo_in.FIFO[1][7] ;
 wire \fifo_in.FIFO[1][8] ;
 wire \fifo_in.FIFO[1][9] ;
 wire \fifo_in.FIFO[2][0] ;
 wire \fifo_in.FIFO[2][10] ;
 wire \fifo_in.FIFO[2][11] ;
 wire \fifo_in.FIFO[2][12] ;
 wire \fifo_in.FIFO[2][13] ;
 wire \fifo_in.FIFO[2][14] ;
 wire \fifo_in.FIFO[2][15] ;
 wire \fifo_in.FIFO[2][16] ;
 wire \fifo_in.FIFO[2][17] ;
 wire \fifo_in.FIFO[2][18] ;
 wire \fifo_in.FIFO[2][19] ;
 wire \fifo_in.FIFO[2][1] ;
 wire \fifo_in.FIFO[2][20] ;
 wire \fifo_in.FIFO[2][21] ;
 wire \fifo_in.FIFO[2][22] ;
 wire \fifo_in.FIFO[2][23] ;
 wire \fifo_in.FIFO[2][24] ;
 wire \fifo_in.FIFO[2][25] ;
 wire \fifo_in.FIFO[2][26] ;
 wire \fifo_in.FIFO[2][27] ;
 wire \fifo_in.FIFO[2][28] ;
 wire \fifo_in.FIFO[2][29] ;
 wire \fifo_in.FIFO[2][2] ;
 wire \fifo_in.FIFO[2][30] ;
 wire \fifo_in.FIFO[2][31] ;
 wire \fifo_in.FIFO[2][3] ;
 wire \fifo_in.FIFO[2][4] ;
 wire \fifo_in.FIFO[2][5] ;
 wire \fifo_in.FIFO[2][6] ;
 wire \fifo_in.FIFO[2][7] ;
 wire \fifo_in.FIFO[2][8] ;
 wire \fifo_in.FIFO[2][9] ;
 wire \fifo_in.FIFO[3][0] ;
 wire \fifo_in.FIFO[3][10] ;
 wire \fifo_in.FIFO[3][11] ;
 wire \fifo_in.FIFO[3][12] ;
 wire \fifo_in.FIFO[3][13] ;
 wire \fifo_in.FIFO[3][14] ;
 wire \fifo_in.FIFO[3][15] ;
 wire \fifo_in.FIFO[3][16] ;
 wire \fifo_in.FIFO[3][17] ;
 wire \fifo_in.FIFO[3][18] ;
 wire \fifo_in.FIFO[3][19] ;
 wire \fifo_in.FIFO[3][1] ;
 wire \fifo_in.FIFO[3][20] ;
 wire \fifo_in.FIFO[3][21] ;
 wire \fifo_in.FIFO[3][22] ;
 wire \fifo_in.FIFO[3][23] ;
 wire \fifo_in.FIFO[3][24] ;
 wire \fifo_in.FIFO[3][25] ;
 wire \fifo_in.FIFO[3][26] ;
 wire \fifo_in.FIFO[3][27] ;
 wire \fifo_in.FIFO[3][28] ;
 wire \fifo_in.FIFO[3][29] ;
 wire \fifo_in.FIFO[3][2] ;
 wire \fifo_in.FIFO[3][30] ;
 wire \fifo_in.FIFO[3][31] ;
 wire \fifo_in.FIFO[3][3] ;
 wire \fifo_in.FIFO[3][4] ;
 wire \fifo_in.FIFO[3][5] ;
 wire \fifo_in.FIFO[3][6] ;
 wire \fifo_in.FIFO[3][7] ;
 wire \fifo_in.FIFO[3][8] ;
 wire \fifo_in.FIFO[3][9] ;
 wire \fifo_in.FIFO[4][0] ;
 wire \fifo_in.FIFO[4][10] ;
 wire \fifo_in.FIFO[4][11] ;
 wire \fifo_in.FIFO[4][12] ;
 wire \fifo_in.FIFO[4][13] ;
 wire \fifo_in.FIFO[4][14] ;
 wire \fifo_in.FIFO[4][15] ;
 wire \fifo_in.FIFO[4][16] ;
 wire \fifo_in.FIFO[4][17] ;
 wire \fifo_in.FIFO[4][18] ;
 wire \fifo_in.FIFO[4][19] ;
 wire \fifo_in.FIFO[4][1] ;
 wire \fifo_in.FIFO[4][20] ;
 wire \fifo_in.FIFO[4][21] ;
 wire \fifo_in.FIFO[4][22] ;
 wire \fifo_in.FIFO[4][23] ;
 wire \fifo_in.FIFO[4][24] ;
 wire \fifo_in.FIFO[4][25] ;
 wire \fifo_in.FIFO[4][26] ;
 wire \fifo_in.FIFO[4][27] ;
 wire \fifo_in.FIFO[4][28] ;
 wire \fifo_in.FIFO[4][29] ;
 wire \fifo_in.FIFO[4][2] ;
 wire \fifo_in.FIFO[4][30] ;
 wire \fifo_in.FIFO[4][31] ;
 wire \fifo_in.FIFO[4][3] ;
 wire \fifo_in.FIFO[4][4] ;
 wire \fifo_in.FIFO[4][5] ;
 wire \fifo_in.FIFO[4][6] ;
 wire \fifo_in.FIFO[4][7] ;
 wire \fifo_in.FIFO[4][8] ;
 wire \fifo_in.FIFO[4][9] ;
 wire \fifo_in.FIFO[5][0] ;
 wire \fifo_in.FIFO[5][10] ;
 wire \fifo_in.FIFO[5][11] ;
 wire \fifo_in.FIFO[5][12] ;
 wire \fifo_in.FIFO[5][13] ;
 wire \fifo_in.FIFO[5][14] ;
 wire \fifo_in.FIFO[5][15] ;
 wire \fifo_in.FIFO[5][16] ;
 wire \fifo_in.FIFO[5][17] ;
 wire \fifo_in.FIFO[5][18] ;
 wire \fifo_in.FIFO[5][19] ;
 wire \fifo_in.FIFO[5][1] ;
 wire \fifo_in.FIFO[5][20] ;
 wire \fifo_in.FIFO[5][21] ;
 wire \fifo_in.FIFO[5][22] ;
 wire \fifo_in.FIFO[5][23] ;
 wire \fifo_in.FIFO[5][24] ;
 wire \fifo_in.FIFO[5][25] ;
 wire \fifo_in.FIFO[5][26] ;
 wire \fifo_in.FIFO[5][27] ;
 wire \fifo_in.FIFO[5][28] ;
 wire \fifo_in.FIFO[5][29] ;
 wire \fifo_in.FIFO[5][2] ;
 wire \fifo_in.FIFO[5][30] ;
 wire \fifo_in.FIFO[5][31] ;
 wire \fifo_in.FIFO[5][3] ;
 wire \fifo_in.FIFO[5][4] ;
 wire \fifo_in.FIFO[5][5] ;
 wire \fifo_in.FIFO[5][6] ;
 wire \fifo_in.FIFO[5][7] ;
 wire \fifo_in.FIFO[5][8] ;
 wire \fifo_in.FIFO[5][9] ;
 wire \fifo_in.FIFO[6][0] ;
 wire \fifo_in.FIFO[6][10] ;
 wire \fifo_in.FIFO[6][11] ;
 wire \fifo_in.FIFO[6][12] ;
 wire \fifo_in.FIFO[6][13] ;
 wire \fifo_in.FIFO[6][14] ;
 wire \fifo_in.FIFO[6][15] ;
 wire \fifo_in.FIFO[6][16] ;
 wire \fifo_in.FIFO[6][17] ;
 wire \fifo_in.FIFO[6][18] ;
 wire \fifo_in.FIFO[6][19] ;
 wire \fifo_in.FIFO[6][1] ;
 wire \fifo_in.FIFO[6][20] ;
 wire \fifo_in.FIFO[6][21] ;
 wire \fifo_in.FIFO[6][22] ;
 wire \fifo_in.FIFO[6][23] ;
 wire \fifo_in.FIFO[6][24] ;
 wire \fifo_in.FIFO[6][25] ;
 wire \fifo_in.FIFO[6][26] ;
 wire \fifo_in.FIFO[6][27] ;
 wire \fifo_in.FIFO[6][28] ;
 wire \fifo_in.FIFO[6][29] ;
 wire \fifo_in.FIFO[6][2] ;
 wire \fifo_in.FIFO[6][30] ;
 wire \fifo_in.FIFO[6][31] ;
 wire \fifo_in.FIFO[6][3] ;
 wire \fifo_in.FIFO[6][4] ;
 wire \fifo_in.FIFO[6][5] ;
 wire \fifo_in.FIFO[6][6] ;
 wire \fifo_in.FIFO[6][7] ;
 wire \fifo_in.FIFO[6][8] ;
 wire \fifo_in.FIFO[6][9] ;
 wire \fifo_in.FIFO[7][0] ;
 wire \fifo_in.FIFO[7][10] ;
 wire \fifo_in.FIFO[7][11] ;
 wire \fifo_in.FIFO[7][12] ;
 wire \fifo_in.FIFO[7][13] ;
 wire \fifo_in.FIFO[7][14] ;
 wire \fifo_in.FIFO[7][15] ;
 wire \fifo_in.FIFO[7][16] ;
 wire \fifo_in.FIFO[7][17] ;
 wire \fifo_in.FIFO[7][18] ;
 wire \fifo_in.FIFO[7][19] ;
 wire \fifo_in.FIFO[7][1] ;
 wire \fifo_in.FIFO[7][20] ;
 wire \fifo_in.FIFO[7][21] ;
 wire \fifo_in.FIFO[7][22] ;
 wire \fifo_in.FIFO[7][23] ;
 wire \fifo_in.FIFO[7][24] ;
 wire \fifo_in.FIFO[7][25] ;
 wire \fifo_in.FIFO[7][26] ;
 wire \fifo_in.FIFO[7][27] ;
 wire \fifo_in.FIFO[7][28] ;
 wire \fifo_in.FIFO[7][29] ;
 wire \fifo_in.FIFO[7][2] ;
 wire \fifo_in.FIFO[7][30] ;
 wire \fifo_in.FIFO[7][31] ;
 wire \fifo_in.FIFO[7][3] ;
 wire \fifo_in.FIFO[7][4] ;
 wire \fifo_in.FIFO[7][5] ;
 wire \fifo_in.FIFO[7][6] ;
 wire \fifo_in.FIFO[7][7] ;
 wire \fifo_in.FIFO[7][8] ;
 wire \fifo_in.FIFO[7][9] ;
 wire \fifo_in.count[0] ;
 wire \fifo_in.count[1] ;
 wire \fifo_in.count[2] ;
 wire \fifo_in.read_addr[0] ;
 wire \fifo_in.read_addr[1] ;
 wire \fifo_in.read_addr[2] ;
 wire \fifo_in.write_addr[0] ;
 wire \fifo_in.write_addr[1] ;
 wire \fifo_in.write_addr[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__0422__B (.DIODE(_0281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0424__A (.DIODE(_0281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0425__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0425__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0426__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0426__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0427__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0428__B (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0429__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0429__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0430__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0430__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0431__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0433__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0433__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0434__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0434__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0435__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0437__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0437__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0438__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0438__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0439__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0441__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0441__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0442__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0442__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0443__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0444__B (.DIODE(_0305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0445__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0445__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0446__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0446__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0447__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0449__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0449__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0450__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0450__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0451__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0453__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0453__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0454__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0454__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0455__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0457__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0457__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0458__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0459__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0461__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0461__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0462__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0462__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0463__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0464__B (.DIODE(_0320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0465__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0465__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0466__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0467__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0469__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0470__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0470__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0471__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0473__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0473__S1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0474__S0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0474__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0475__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0477__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0477__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0478__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0478__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0479__S (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0481__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0481__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0482__S0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0482__S1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0483__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0484__B (.DIODE(_0335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0486__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0486__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0487__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0489__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0489__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0490__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0490__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0491__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0493__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0495__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0498__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0498__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0499__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0503__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0507__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0509__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0509__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0510__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0510__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0511__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0514__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0514__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0515__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0517__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0517__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0518__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0518__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0519__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0521__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0521__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__B (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0531__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0533__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0533__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0535__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0537__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0537__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0539__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__B (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__S0 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0543__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__S0 (.DIODE(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__S0 (.DIODE(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0547__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0549__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0549__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__S0 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0551__S (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0555__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0558__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0559__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0561__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0563__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0565__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0566__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0568__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0570__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__S (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0578__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0589__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0601__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0602__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__S (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0620__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0624__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0644__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__S (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0666__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__S (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__S (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0734__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__S (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0764__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0777__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__S (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__D (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__B (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__S (.DIODE(_0275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0846__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_0393_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(_0275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold561_A (.DIODE(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold563_A (.DIODE(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__inv_2 _0409_ (.A(net1),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _0410_ (.A(net34),
    .Y(_0277_));
 sky130_fd_sc_hd__or4bb_1 _0411_ (.A(net26),
    .B(net25),
    .C_N(net23),
    .D_N(net22),
    .X(_0278_));
 sky130_fd_sc_hd__or4_1 _0412_ (.A(net19),
    .B(net18),
    .C(net21),
    .D(net20),
    .X(_0279_));
 sky130_fd_sc_hd__or4_1 _0413_ (.A(net15),
    .B(net14),
    .C(net17),
    .D(net16),
    .X(_0280_));
 sky130_fd_sc_hd__or3_2 _0414_ (.A(_0278_),
    .B(_0279_),
    .C(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__or4_1 _0415_ (.A(net33),
    .B(net32),
    .C(net4),
    .D(net3),
    .X(_0282_));
 sky130_fd_sc_hd__or4_1 _0416_ (.A(net29),
    .B(net28),
    .C(net31),
    .D(net30),
    .X(_0283_));
 sky130_fd_sc_hd__or4_1 _0417_ (.A(net6),
    .B(net5),
    .C(net8),
    .D(net7),
    .X(_0284_));
 sky130_fd_sc_hd__or4_1 _0418_ (.A(net10),
    .B(net9),
    .C(net12),
    .D(net11),
    .X(_0285_));
 sky130_fd_sc_hd__or4_2 _0419_ (.A(_0282_),
    .B(_0283_),
    .C(_0284_),
    .D(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__or3_1 _0420_ (.A(net13),
    .B(net27),
    .C(net24),
    .X(_0287_));
 sky130_fd_sc_hd__or3b_1 _0421_ (.A(net1),
    .B(_0287_),
    .C_N(net67),
    .X(_0288_));
 sky130_fd_sc_hd__nor4_1 _0422_ (.A(_0277_),
    .B(_0281_),
    .C(_0286_),
    .D(_0288_),
    .Y(net69));
 sky130_fd_sc_hd__or2_1 _0423_ (.A(net68),
    .B(net2),
    .X(_0289_));
 sky130_fd_sc_hd__nor4_2 _0424_ (.A(_0281_),
    .B(_0286_),
    .C(_0288_),
    .D(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__mux4_1 _0425_ (.A0(\fifo_in.FIFO[4][0] ),
    .A1(\fifo_in.FIFO[5][0] ),
    .A2(\fifo_in.FIFO[6][0] ),
    .A3(\fifo_in.FIFO[7][0] ),
    .S0(net129),
    .S1(net124),
    .X(_0291_));
 sky130_fd_sc_hd__mux4_1 _0426_ (.A0(\fifo_in.FIFO[0][0] ),
    .A1(\fifo_in.FIFO[1][0] ),
    .A2(\fifo_in.FIFO[2][0] ),
    .A3(\fifo_in.FIFO[3][0] ),
    .S0(net129),
    .S1(net124),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _0427_ (.A0(_0292_),
    .A1(_0291_),
    .S(net121),
    .X(_0293_));
 sky130_fd_sc_hd__and2_1 _0428_ (.A(_0290_),
    .B(_0293_),
    .X(net70));
 sky130_fd_sc_hd__mux4_1 _0429_ (.A0(\fifo_in.FIFO[4][1] ),
    .A1(\fifo_in.FIFO[5][1] ),
    .A2(\fifo_in.FIFO[6][1] ),
    .A3(\fifo_in.FIFO[7][1] ),
    .S0(net129),
    .S1(net124),
    .X(_0294_));
 sky130_fd_sc_hd__mux4_1 _0430_ (.A0(\fifo_in.FIFO[0][1] ),
    .A1(\fifo_in.FIFO[1][1] ),
    .A2(\fifo_in.FIFO[2][1] ),
    .A3(\fifo_in.FIFO[3][1] ),
    .S0(net129),
    .S1(net124),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _0431_ (.A0(_0295_),
    .A1(_0294_),
    .S(net121),
    .X(_0296_));
 sky130_fd_sc_hd__and2_1 _0432_ (.A(_0290_),
    .B(_0296_),
    .X(net81));
 sky130_fd_sc_hd__mux4_1 _0433_ (.A0(\fifo_in.FIFO[4][2] ),
    .A1(\fifo_in.FIFO[5][2] ),
    .A2(\fifo_in.FIFO[6][2] ),
    .A3(\fifo_in.FIFO[7][2] ),
    .S0(net128),
    .S1(net123),
    .X(_0297_));
 sky130_fd_sc_hd__mux4_1 _0434_ (.A0(\fifo_in.FIFO[0][2] ),
    .A1(\fifo_in.FIFO[1][2] ),
    .A2(\fifo_in.FIFO[2][2] ),
    .A3(\fifo_in.FIFO[3][2] ),
    .S0(net128),
    .S1(net123),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _0435_ (.A0(_0298_),
    .A1(_0297_),
    .S(net121),
    .X(_0299_));
 sky130_fd_sc_hd__and2_1 _0436_ (.A(_0290_),
    .B(_0299_),
    .X(net92));
 sky130_fd_sc_hd__mux4_1 _0437_ (.A0(\fifo_in.FIFO[4][3] ),
    .A1(\fifo_in.FIFO[5][3] ),
    .A2(\fifo_in.FIFO[6][3] ),
    .A3(\fifo_in.FIFO[7][3] ),
    .S0(net129),
    .S1(net124),
    .X(_0300_));
 sky130_fd_sc_hd__mux4_1 _0438_ (.A0(\fifo_in.FIFO[0][3] ),
    .A1(\fifo_in.FIFO[1][3] ),
    .A2(\fifo_in.FIFO[2][3] ),
    .A3(\fifo_in.FIFO[3][3] ),
    .S0(net129),
    .S1(net127),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _0439_ (.A0(_0301_),
    .A1(_0300_),
    .S(net121),
    .X(_0302_));
 sky130_fd_sc_hd__and2_1 _0440_ (.A(_0290_),
    .B(_0302_),
    .X(net95));
 sky130_fd_sc_hd__mux4_1 _0441_ (.A0(\fifo_in.FIFO[4][4] ),
    .A1(\fifo_in.FIFO[5][4] ),
    .A2(\fifo_in.FIFO[6][4] ),
    .A3(\fifo_in.FIFO[7][4] ),
    .S0(net129),
    .S1(net127),
    .X(_0303_));
 sky130_fd_sc_hd__mux4_1 _0442_ (.A0(\fifo_in.FIFO[0][4] ),
    .A1(\fifo_in.FIFO[1][4] ),
    .A2(\fifo_in.FIFO[2][4] ),
    .A3(\fifo_in.FIFO[3][4] ),
    .S0(net129),
    .S1(net127),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _0443_ (.A0(_0304_),
    .A1(_0303_),
    .S(net121),
    .X(_0305_));
 sky130_fd_sc_hd__and2_1 _0444_ (.A(_0290_),
    .B(_0305_),
    .X(net96));
 sky130_fd_sc_hd__mux4_1 _0445_ (.A0(\fifo_in.FIFO[4][5] ),
    .A1(\fifo_in.FIFO[5][5] ),
    .A2(\fifo_in.FIFO[6][5] ),
    .A3(\fifo_in.FIFO[7][5] ),
    .S0(net128),
    .S1(net123),
    .X(_0306_));
 sky130_fd_sc_hd__mux4_1 _0446_ (.A0(\fifo_in.FIFO[0][5] ),
    .A1(\fifo_in.FIFO[1][5] ),
    .A2(\fifo_in.FIFO[2][5] ),
    .A3(\fifo_in.FIFO[3][5] ),
    .S0(net128),
    .S1(net123),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _0447_ (.A0(_0307_),
    .A1(_0306_),
    .S(net121),
    .X(_0308_));
 sky130_fd_sc_hd__and2_1 _0448_ (.A(net119),
    .B(_0308_),
    .X(net97));
 sky130_fd_sc_hd__mux4_1 _0449_ (.A0(\fifo_in.FIFO[4][6] ),
    .A1(\fifo_in.FIFO[5][6] ),
    .A2(\fifo_in.FIFO[6][6] ),
    .A3(\fifo_in.FIFO[7][6] ),
    .S0(net128),
    .S1(net123),
    .X(_0309_));
 sky130_fd_sc_hd__mux4_1 _0450_ (.A0(\fifo_in.FIFO[0][6] ),
    .A1(\fifo_in.FIFO[1][6] ),
    .A2(\fifo_in.FIFO[2][6] ),
    .A3(\fifo_in.FIFO[3][6] ),
    .S0(net128),
    .S1(net123),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _0451_ (.A0(_0310_),
    .A1(_0309_),
    .S(net121),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _0452_ (.A(net119),
    .B(_0311_),
    .X(net98));
 sky130_fd_sc_hd__mux4_1 _0453_ (.A0(\fifo_in.FIFO[4][7] ),
    .A1(\fifo_in.FIFO[5][7] ),
    .A2(\fifo_in.FIFO[6][7] ),
    .A3(\fifo_in.FIFO[7][7] ),
    .S0(net129),
    .S1(net124),
    .X(_0312_));
 sky130_fd_sc_hd__mux4_1 _0454_ (.A0(\fifo_in.FIFO[0][7] ),
    .A1(\fifo_in.FIFO[1][7] ),
    .A2(\fifo_in.FIFO[2][7] ),
    .A3(\fifo_in.FIFO[3][7] ),
    .S0(net129),
    .S1(net124),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _0455_ (.A0(_0313_),
    .A1(_0312_),
    .S(net121),
    .X(_0314_));
 sky130_fd_sc_hd__and2_1 _0456_ (.A(net119),
    .B(_0314_),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 _0457_ (.A0(\fifo_in.FIFO[4][8] ),
    .A1(\fifo_in.FIFO[5][8] ),
    .A2(\fifo_in.FIFO[6][8] ),
    .A3(\fifo_in.FIFO[7][8] ),
    .S0(net128),
    .S1(net123),
    .X(_0315_));
 sky130_fd_sc_hd__mux4_1 _0458_ (.A0(\fifo_in.FIFO[0][8] ),
    .A1(\fifo_in.FIFO[1][8] ),
    .A2(\fifo_in.FIFO[2][8] ),
    .A3(\fifo_in.FIFO[3][8] ),
    .S0(net128),
    .S1(net123),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _0459_ (.A0(_0316_),
    .A1(_0315_),
    .S(net121),
    .X(_0317_));
 sky130_fd_sc_hd__and2_1 _0460_ (.A(net119),
    .B(_0317_),
    .X(net100));
 sky130_fd_sc_hd__mux4_1 _0461_ (.A0(\fifo_in.FIFO[4][9] ),
    .A1(\fifo_in.FIFO[5][9] ),
    .A2(\fifo_in.FIFO[6][9] ),
    .A3(\fifo_in.FIFO[7][9] ),
    .S0(net129),
    .S1(net124),
    .X(_0318_));
 sky130_fd_sc_hd__mux4_1 _0462_ (.A0(\fifo_in.FIFO[0][9] ),
    .A1(\fifo_in.FIFO[1][9] ),
    .A2(\fifo_in.FIFO[2][9] ),
    .A3(\fifo_in.FIFO[3][9] ),
    .S0(net129),
    .S1(net124),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _0463_ (.A0(_0319_),
    .A1(_0318_),
    .S(net121),
    .X(_0320_));
 sky130_fd_sc_hd__and2_1 _0464_ (.A(net119),
    .B(_0320_),
    .X(net101));
 sky130_fd_sc_hd__mux4_1 _0465_ (.A0(\fifo_in.FIFO[4][10] ),
    .A1(\fifo_in.FIFO[5][10] ),
    .A2(\fifo_in.FIFO[6][10] ),
    .A3(\fifo_in.FIFO[7][10] ),
    .S0(net128),
    .S1(net123),
    .X(_0321_));
 sky130_fd_sc_hd__mux4_1 _0466_ (.A0(\fifo_in.FIFO[0][10] ),
    .A1(\fifo_in.FIFO[1][10] ),
    .A2(\fifo_in.FIFO[2][10] ),
    .A3(\fifo_in.FIFO[3][10] ),
    .S0(net128),
    .S1(net124),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _0467_ (.A0(_0322_),
    .A1(_0321_),
    .S(net121),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _0468_ (.A(net119),
    .B(_0323_),
    .X(net71));
 sky130_fd_sc_hd__mux4_1 _0469_ (.A0(\fifo_in.FIFO[4][11] ),
    .A1(\fifo_in.FIFO[5][11] ),
    .A2(\fifo_in.FIFO[6][11] ),
    .A3(\fifo_in.FIFO[7][11] ),
    .S0(net128),
    .S1(net123),
    .X(_0324_));
 sky130_fd_sc_hd__mux4_1 _0470_ (.A0(\fifo_in.FIFO[0][11] ),
    .A1(\fifo_in.FIFO[1][11] ),
    .A2(\fifo_in.FIFO[2][11] ),
    .A3(\fifo_in.FIFO[3][11] ),
    .S0(net128),
    .S1(net123),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _0471_ (.A0(_0325_),
    .A1(_0324_),
    .S(net121),
    .X(_0326_));
 sky130_fd_sc_hd__and2_1 _0472_ (.A(net119),
    .B(_0326_),
    .X(net72));
 sky130_fd_sc_hd__mux4_1 _0473_ (.A0(\fifo_in.FIFO[4][12] ),
    .A1(\fifo_in.FIFO[5][12] ),
    .A2(\fifo_in.FIFO[6][12] ),
    .A3(\fifo_in.FIFO[7][12] ),
    .S0(net128),
    .S1(net123),
    .X(_0327_));
 sky130_fd_sc_hd__mux4_1 _0474_ (.A0(\fifo_in.FIFO[0][12] ),
    .A1(\fifo_in.FIFO[1][12] ),
    .A2(\fifo_in.FIFO[2][12] ),
    .A3(\fifo_in.FIFO[3][12] ),
    .S0(net128),
    .S1(net124),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _0475_ (.A0(_0328_),
    .A1(_0327_),
    .S(net121),
    .X(_0329_));
 sky130_fd_sc_hd__and2_1 _0476_ (.A(net119),
    .B(_0329_),
    .X(net73));
 sky130_fd_sc_hd__mux4_1 _0477_ (.A0(\fifo_in.FIFO[4][13] ),
    .A1(\fifo_in.FIFO[5][13] ),
    .A2(\fifo_in.FIFO[6][13] ),
    .A3(\fifo_in.FIFO[7][13] ),
    .S0(net129),
    .S1(net124),
    .X(_0330_));
 sky130_fd_sc_hd__mux4_1 _0478_ (.A0(\fifo_in.FIFO[0][13] ),
    .A1(\fifo_in.FIFO[1][13] ),
    .A2(\fifo_in.FIFO[2][13] ),
    .A3(\fifo_in.FIFO[3][13] ),
    .S0(net129),
    .S1(net124),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _0479_ (.A0(_0331_),
    .A1(_0330_),
    .S(\fifo_in.read_addr[2] ),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _0480_ (.A(net119),
    .B(_0332_),
    .X(net74));
 sky130_fd_sc_hd__mux4_1 _0481_ (.A0(\fifo_in.FIFO[4][14] ),
    .A1(\fifo_in.FIFO[5][14] ),
    .A2(\fifo_in.FIFO[6][14] ),
    .A3(\fifo_in.FIFO[7][14] ),
    .S0(net129),
    .S1(net124),
    .X(_0333_));
 sky130_fd_sc_hd__mux4_1 _0482_ (.A0(\fifo_in.FIFO[0][14] ),
    .A1(\fifo_in.FIFO[1][14] ),
    .A2(\fifo_in.FIFO[2][14] ),
    .A3(\fifo_in.FIFO[3][14] ),
    .S0(net129),
    .S1(net124),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _0483_ (.A0(_0334_),
    .A1(_0333_),
    .S(net121),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _0484_ (.A(net119),
    .B(_0335_),
    .X(net75));
 sky130_fd_sc_hd__mux4_1 _0485_ (.A0(\fifo_in.FIFO[4][15] ),
    .A1(\fifo_in.FIFO[5][15] ),
    .A2(\fifo_in.FIFO[6][15] ),
    .A3(\fifo_in.FIFO[7][15] ),
    .S0(net131),
    .S1(net126),
    .X(_0336_));
 sky130_fd_sc_hd__mux4_1 _0486_ (.A0(\fifo_in.FIFO[0][15] ),
    .A1(\fifo_in.FIFO[1][15] ),
    .A2(\fifo_in.FIFO[2][15] ),
    .A3(\fifo_in.FIFO[3][15] ),
    .S0(net131),
    .S1(net126),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _0487_ (.A0(_0337_),
    .A1(_0336_),
    .S(net122),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _0488_ (.A(net119),
    .B(_0338_),
    .X(net76));
 sky130_fd_sc_hd__mux4_1 _0489_ (.A0(\fifo_in.FIFO[4][16] ),
    .A1(\fifo_in.FIFO[5][16] ),
    .A2(\fifo_in.FIFO[6][16] ),
    .A3(\fifo_in.FIFO[7][16] ),
    .S0(net130),
    .S1(net125),
    .X(_0339_));
 sky130_fd_sc_hd__mux4_1 _0490_ (.A0(\fifo_in.FIFO[0][16] ),
    .A1(\fifo_in.FIFO[1][16] ),
    .A2(\fifo_in.FIFO[2][16] ),
    .A3(\fifo_in.FIFO[3][16] ),
    .S0(net130),
    .S1(net125),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _0491_ (.A0(_0340_),
    .A1(_0339_),
    .S(net122),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _0492_ (.A(net119),
    .B(_0341_),
    .X(net77));
 sky130_fd_sc_hd__mux4_1 _0493_ (.A0(\fifo_in.FIFO[4][17] ),
    .A1(\fifo_in.FIFO[5][17] ),
    .A2(\fifo_in.FIFO[6][17] ),
    .A3(\fifo_in.FIFO[7][17] ),
    .S0(net130),
    .S1(net125),
    .X(_0342_));
 sky130_fd_sc_hd__mux4_1 _0494_ (.A0(\fifo_in.FIFO[0][17] ),
    .A1(\fifo_in.FIFO[1][17] ),
    .A2(\fifo_in.FIFO[2][17] ),
    .A3(\fifo_in.FIFO[3][17] ),
    .S0(net130),
    .S1(net125),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _0495_ (.A0(_0343_),
    .A1(_0342_),
    .S(net122),
    .X(_0344_));
 sky130_fd_sc_hd__and2_1 _0496_ (.A(net119),
    .B(_0344_),
    .X(net78));
 sky130_fd_sc_hd__mux4_1 _0497_ (.A0(\fifo_in.FIFO[4][18] ),
    .A1(\fifo_in.FIFO[5][18] ),
    .A2(\fifo_in.FIFO[6][18] ),
    .A3(\fifo_in.FIFO[7][18] ),
    .S0(net130),
    .S1(net125),
    .X(_0345_));
 sky130_fd_sc_hd__mux4_1 _0498_ (.A0(\fifo_in.FIFO[0][18] ),
    .A1(\fifo_in.FIFO[1][18] ),
    .A2(\fifo_in.FIFO[2][18] ),
    .A3(\fifo_in.FIFO[3][18] ),
    .S0(net130),
    .S1(net125),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _0499_ (.A0(_0346_),
    .A1(_0345_),
    .S(net122),
    .X(_0347_));
 sky130_fd_sc_hd__and2_1 _0500_ (.A(net118),
    .B(_0347_),
    .X(net79));
 sky130_fd_sc_hd__mux4_1 _0501_ (.A0(\fifo_in.FIFO[4][19] ),
    .A1(\fifo_in.FIFO[5][19] ),
    .A2(\fifo_in.FIFO[6][19] ),
    .A3(\fifo_in.FIFO[7][19] ),
    .S0(net131),
    .S1(net126),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _0502_ (.A0(\fifo_in.FIFO[0][19] ),
    .A1(\fifo_in.FIFO[1][19] ),
    .A2(\fifo_in.FIFO[2][19] ),
    .A3(\fifo_in.FIFO[3][19] ),
    .S0(net131),
    .S1(net126),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _0503_ (.A0(_0349_),
    .A1(_0348_),
    .S(net122),
    .X(_0350_));
 sky130_fd_sc_hd__and2_1 _0504_ (.A(net118),
    .B(_0350_),
    .X(net80));
 sky130_fd_sc_hd__mux4_1 _0505_ (.A0(\fifo_in.FIFO[4][20] ),
    .A1(\fifo_in.FIFO[5][20] ),
    .A2(\fifo_in.FIFO[6][20] ),
    .A3(\fifo_in.FIFO[7][20] ),
    .S0(net130),
    .S1(net125),
    .X(_0351_));
 sky130_fd_sc_hd__mux4_1 _0506_ (.A0(\fifo_in.FIFO[0][20] ),
    .A1(\fifo_in.FIFO[1][20] ),
    .A2(\fifo_in.FIFO[2][20] ),
    .A3(\fifo_in.FIFO[3][20] ),
    .S0(net130),
    .S1(net125),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _0507_ (.A0(_0352_),
    .A1(_0351_),
    .S(net122),
    .X(_0353_));
 sky130_fd_sc_hd__and2_1 _0508_ (.A(net118),
    .B(_0353_),
    .X(net82));
 sky130_fd_sc_hd__mux4_1 _0509_ (.A0(\fifo_in.FIFO[4][21] ),
    .A1(\fifo_in.FIFO[5][21] ),
    .A2(\fifo_in.FIFO[6][21] ),
    .A3(\fifo_in.FIFO[7][21] ),
    .S0(net131),
    .S1(net126),
    .X(_0354_));
 sky130_fd_sc_hd__mux4_1 _0510_ (.A0(\fifo_in.FIFO[0][21] ),
    .A1(\fifo_in.FIFO[1][21] ),
    .A2(\fifo_in.FIFO[2][21] ),
    .A3(\fifo_in.FIFO[3][21] ),
    .S0(net131),
    .S1(net126),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _0511_ (.A0(_0355_),
    .A1(_0354_),
    .S(net122),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _0512_ (.A(net118),
    .B(_0356_),
    .X(net83));
 sky130_fd_sc_hd__mux4_1 _0513_ (.A0(\fifo_in.FIFO[4][22] ),
    .A1(\fifo_in.FIFO[5][22] ),
    .A2(\fifo_in.FIFO[6][22] ),
    .A3(\fifo_in.FIFO[7][22] ),
    .S0(net131),
    .S1(net126),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_1 _0514_ (.A0(\fifo_in.FIFO[0][22] ),
    .A1(\fifo_in.FIFO[1][22] ),
    .A2(\fifo_in.FIFO[2][22] ),
    .A3(\fifo_in.FIFO[3][22] ),
    .S0(net131),
    .S1(net126),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _0515_ (.A0(_0358_),
    .A1(_0357_),
    .S(net122),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _0516_ (.A(net118),
    .B(_0359_),
    .X(net84));
 sky130_fd_sc_hd__mux4_1 _0517_ (.A0(\fifo_in.FIFO[4][23] ),
    .A1(\fifo_in.FIFO[5][23] ),
    .A2(\fifo_in.FIFO[6][23] ),
    .A3(\fifo_in.FIFO[7][23] ),
    .S0(net131),
    .S1(net126),
    .X(_0360_));
 sky130_fd_sc_hd__mux4_1 _0518_ (.A0(\fifo_in.FIFO[0][23] ),
    .A1(\fifo_in.FIFO[1][23] ),
    .A2(\fifo_in.FIFO[2][23] ),
    .A3(\fifo_in.FIFO[3][23] ),
    .S0(net131),
    .S1(net126),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _0519_ (.A0(_0361_),
    .A1(_0360_),
    .S(net122),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _0520_ (.A(net118),
    .B(_0362_),
    .X(net85));
 sky130_fd_sc_hd__mux4_1 _0521_ (.A0(\fifo_in.FIFO[4][24] ),
    .A1(\fifo_in.FIFO[5][24] ),
    .A2(\fifo_in.FIFO[6][24] ),
    .A3(\fifo_in.FIFO[7][24] ),
    .S0(net130),
    .S1(net125),
    .X(_0363_));
 sky130_fd_sc_hd__mux4_1 _0522_ (.A0(\fifo_in.FIFO[0][24] ),
    .A1(\fifo_in.FIFO[1][24] ),
    .A2(\fifo_in.FIFO[2][24] ),
    .A3(\fifo_in.FIFO[3][24] ),
    .S0(net130),
    .S1(net125),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _0523_ (.A0(_0364_),
    .A1(_0363_),
    .S(net122),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _0524_ (.A(net118),
    .B(_0365_),
    .X(net86));
 sky130_fd_sc_hd__mux4_1 _0525_ (.A0(\fifo_in.FIFO[4][25] ),
    .A1(\fifo_in.FIFO[5][25] ),
    .A2(\fifo_in.FIFO[6][25] ),
    .A3(\fifo_in.FIFO[7][25] ),
    .S0(net131),
    .S1(net126),
    .X(_0366_));
 sky130_fd_sc_hd__mux4_1 _0526_ (.A0(\fifo_in.FIFO[0][25] ),
    .A1(\fifo_in.FIFO[1][25] ),
    .A2(\fifo_in.FIFO[2][25] ),
    .A3(\fifo_in.FIFO[3][25] ),
    .S0(net131),
    .S1(net126),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _0527_ (.A0(_0367_),
    .A1(_0366_),
    .S(net122),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _0528_ (.A(net118),
    .B(_0368_),
    .X(net87));
 sky130_fd_sc_hd__mux4_1 _0529_ (.A0(\fifo_in.FIFO[4][26] ),
    .A1(\fifo_in.FIFO[5][26] ),
    .A2(\fifo_in.FIFO[6][26] ),
    .A3(\fifo_in.FIFO[7][26] ),
    .S0(net130),
    .S1(net125),
    .X(_0369_));
 sky130_fd_sc_hd__mux4_1 _0530_ (.A0(\fifo_in.FIFO[0][26] ),
    .A1(\fifo_in.FIFO[1][26] ),
    .A2(\fifo_in.FIFO[2][26] ),
    .A3(\fifo_in.FIFO[3][26] ),
    .S0(net130),
    .S1(net125),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _0531_ (.A0(_0370_),
    .A1(_0369_),
    .S(net122),
    .X(_0371_));
 sky130_fd_sc_hd__and2_1 _0532_ (.A(net118),
    .B(_0371_),
    .X(net88));
 sky130_fd_sc_hd__mux4_1 _0533_ (.A0(\fifo_in.FIFO[4][27] ),
    .A1(\fifo_in.FIFO[5][27] ),
    .A2(\fifo_in.FIFO[6][27] ),
    .A3(\fifo_in.FIFO[7][27] ),
    .S0(net130),
    .S1(net125),
    .X(_0372_));
 sky130_fd_sc_hd__mux4_1 _0534_ (.A0(\fifo_in.FIFO[0][27] ),
    .A1(\fifo_in.FIFO[1][27] ),
    .A2(\fifo_in.FIFO[2][27] ),
    .A3(\fifo_in.FIFO[3][27] ),
    .S0(net130),
    .S1(net125),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _0535_ (.A0(_0373_),
    .A1(_0372_),
    .S(net122),
    .X(_0374_));
 sky130_fd_sc_hd__and2_1 _0536_ (.A(net118),
    .B(_0374_),
    .X(net89));
 sky130_fd_sc_hd__mux4_1 _0537_ (.A0(\fifo_in.FIFO[4][28] ),
    .A1(\fifo_in.FIFO[5][28] ),
    .A2(\fifo_in.FIFO[6][28] ),
    .A3(\fifo_in.FIFO[7][28] ),
    .S0(net131),
    .S1(net126),
    .X(_0375_));
 sky130_fd_sc_hd__mux4_1 _0538_ (.A0(\fifo_in.FIFO[0][28] ),
    .A1(\fifo_in.FIFO[1][28] ),
    .A2(\fifo_in.FIFO[2][28] ),
    .A3(\fifo_in.FIFO[3][28] ),
    .S0(net131),
    .S1(net126),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _0539_ (.A0(_0376_),
    .A1(_0375_),
    .S(net122),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _0540_ (.A(net118),
    .B(_0377_),
    .X(net90));
 sky130_fd_sc_hd__mux4_1 _0541_ (.A0(\fifo_in.FIFO[4][29] ),
    .A1(\fifo_in.FIFO[5][29] ),
    .A2(\fifo_in.FIFO[6][29] ),
    .A3(\fifo_in.FIFO[7][29] ),
    .S0(net130),
    .S1(net125),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_1 _0542_ (.A0(\fifo_in.FIFO[0][29] ),
    .A1(\fifo_in.FIFO[1][29] ),
    .A2(\fifo_in.FIFO[2][29] ),
    .A3(\fifo_in.FIFO[3][29] ),
    .S0(net130),
    .S1(net125),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _0543_ (.A0(_0379_),
    .A1(_0378_),
    .S(net122),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _0544_ (.A(net118),
    .B(_0380_),
    .X(net91));
 sky130_fd_sc_hd__mux4_1 _0545_ (.A0(\fifo_in.FIFO[4][30] ),
    .A1(\fifo_in.FIFO[5][30] ),
    .A2(\fifo_in.FIFO[6][30] ),
    .A3(\fifo_in.FIFO[7][30] ),
    .S0(\fifo_in.read_addr[0] ),
    .S1(net127),
    .X(_0381_));
 sky130_fd_sc_hd__mux4_1 _0546_ (.A0(\fifo_in.FIFO[0][30] ),
    .A1(\fifo_in.FIFO[1][30] ),
    .A2(\fifo_in.FIFO[2][30] ),
    .A3(\fifo_in.FIFO[3][30] ),
    .S0(\fifo_in.read_addr[0] ),
    .S1(net127),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _0547_ (.A0(_0382_),
    .A1(_0381_),
    .S(net122),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _0548_ (.A(net118),
    .B(_0383_),
    .X(net93));
 sky130_fd_sc_hd__mux4_1 _0549_ (.A0(\fifo_in.FIFO[4][31] ),
    .A1(\fifo_in.FIFO[5][31] ),
    .A2(\fifo_in.FIFO[6][31] ),
    .A3(\fifo_in.FIFO[7][31] ),
    .S0(net131),
    .S1(net126),
    .X(_0384_));
 sky130_fd_sc_hd__mux4_1 _0550_ (.A0(\fifo_in.FIFO[0][31] ),
    .A1(\fifo_in.FIFO[1][31] ),
    .A2(\fifo_in.FIFO[2][31] ),
    .A3(\fifo_in.FIFO[3][31] ),
    .S0(net131),
    .S1(net126),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(_0385_),
    .A1(_0384_),
    .S(\fifo_in.read_addr[2] ),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _0552_ (.A(net118),
    .B(_0386_),
    .X(net94));
 sky130_fd_sc_hd__nand3_2 _0553_ (.A(net686),
    .B(net68),
    .C(net67),
    .Y(_0387_));
 sky130_fd_sc_hd__or4b_4 _0554_ (.A(\fifo_in.write_addr[1] ),
    .B(net1),
    .C(_0387_),
    .D_N(\fifo_in.write_addr[2] ),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _0555_ (.A0(net643),
    .A1(net654),
    .S(net117),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _0556_ (.A0(net538),
    .A1(net724),
    .S(net117),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _0557_ (.A0(net422),
    .A1(net520),
    .S(net117),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _0558_ (.A0(net525),
    .A1(net540),
    .S(net117),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _0559_ (.A0(net224),
    .A1(net514),
    .S(net117),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _0560_ (.A0(net368),
    .A1(net389),
    .S(net117),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0561_ (.A0(net652),
    .A1(net666),
    .S(net117),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _0562_ (.A0(net535),
    .A1(net583),
    .S(net117),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0563_ (.A0(net329),
    .A1(net606),
    .S(net117),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0564_ (.A0(net326),
    .A1(net391),
    .S(net116),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0565_ (.A0(net154),
    .A1(net162),
    .S(net116),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _0566_ (.A0(net227),
    .A1(net243),
    .S(net116),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _0567_ (.A0(net136),
    .A1(net178),
    .S(net116),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _0568_ (.A0(net398),
    .A1(net416),
    .S(net116),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0569_ (.A0(net217),
    .A1(net237),
    .S(net116),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(net381),
    .A1(net406),
    .S(net116),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0571_ (.A0(net353),
    .A1(net355),
    .S(net116),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0572_ (.A0(net307),
    .A1(net309),
    .S(_0388_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0573_ (.A0(net212),
    .A1(net259),
    .S(net116),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0574_ (.A0(net340),
    .A1(net361),
    .S(net116),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0575_ (.A0(net133),
    .A1(net140),
    .S(net116),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0576_ (.A0(net151),
    .A1(net193),
    .S(net116),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0577_ (.A0(net419),
    .A1(net434),
    .S(net116),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0578_ (.A0(net191),
    .A1(net201),
    .S(net116),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0579_ (.A0(net232),
    .A1(net290),
    .S(net116),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0580_ (.A0(net278),
    .A1(net292),
    .S(net116),
    .X(_0025_));
 sky130_fd_sc_hd__and4b_1 _0581_ (.A_N(\fifo_in.write_addr[0] ),
    .B(net68),
    .C(net67),
    .D(_0276_),
    .X(_0389_));
 sky130_fd_sc_hd__and3b_2 _0582_ (.A_N(\fifo_in.write_addr[1] ),
    .B(_0389_),
    .C(\fifo_in.write_addr[2] ),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _0583_ (.A0(net630),
    .A1(net563),
    .S(net115),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0584_ (.A0(net546),
    .A1(net506),
    .S(net115),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0585_ (.A0(net499),
    .A1(net439),
    .S(net115),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _0586_ (.A0(net622),
    .A1(net588),
    .S(net115),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(net577),
    .A1(net528),
    .S(net115),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0588_ (.A0(net280),
    .A1(net235),
    .S(net115),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0589_ (.A0(net664),
    .A1(net643),
    .S(net115),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0590_ (.A0(net571),
    .A1(net538),
    .S(net115),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0591_ (.A0(net473),
    .A1(net422),
    .S(net115),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0592_ (.A0(net544),
    .A1(net525),
    .S(net115),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0593_ (.A0(net522),
    .A1(net224),
    .S(net115),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net475),
    .A1(net368),
    .S(net115),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0595_ (.A0(net668),
    .A1(net652),
    .S(net115),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net558),
    .A1(net535),
    .S(net115),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0597_ (.A0(net703),
    .A1(net329),
    .S(net115),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(net376),
    .A1(net326),
    .S(net114),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0599_ (.A0(net168),
    .A1(net154),
    .S(net114),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0600_ (.A0(net298),
    .A1(net227),
    .S(net114),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0601_ (.A0(net142),
    .A1(net136),
    .S(net114),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net445),
    .A1(net398),
    .S(net114),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0603_ (.A0(net219),
    .A1(net217),
    .S(net114),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0604_ (.A0(net395),
    .A1(net381),
    .S(net114),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0605_ (.A0(net465),
    .A1(net353),
    .S(net114),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0606_ (.A0(net363),
    .A1(net307),
    .S(_0390_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0607_ (.A0(net344),
    .A1(net212),
    .S(net114),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0608_ (.A0(net408),
    .A1(net340),
    .S(net114),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0609_ (.A0(net184),
    .A1(net133),
    .S(net114),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(net170),
    .A1(net151),
    .S(net114),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0611_ (.A0(net447),
    .A1(net419),
    .S(net114),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0612_ (.A0(net203),
    .A1(net191),
    .S(net114),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0613_ (.A0(net315),
    .A1(net232),
    .S(net114),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(net302),
    .A1(net278),
    .S(net114),
    .X(_0057_));
 sky130_fd_sc_hd__nand4_1 _0615_ (.A(net689),
    .B(net686),
    .C(net68),
    .D(net67),
    .Y(_0391_));
 sky130_fd_sc_hd__or2_1 _0616_ (.A(net676),
    .B(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__or2_4 _0617_ (.A(net1),
    .B(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _0618_ (.A0(net563),
    .A1(net579),
    .S(net103),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0619_ (.A0(net506),
    .A1(net712),
    .S(net103),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0620_ (.A0(net439),
    .A1(net449),
    .S(net103),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0621_ (.A0(net588),
    .A1(net614),
    .S(net103),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0622_ (.A0(net528),
    .A1(net581),
    .S(net103),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0623_ (.A0(net235),
    .A1(net288),
    .S(net103),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0624_ (.A0(net643),
    .A1(net645),
    .S(net103),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0625_ (.A0(net538),
    .A1(net598),
    .S(net103),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0626_ (.A0(net422),
    .A1(net495),
    .S(net103),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0627_ (.A0(net525),
    .A1(net717),
    .S(net103),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0628_ (.A0(net224),
    .A1(net483),
    .S(net103),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0629_ (.A0(net368),
    .A1(net719),
    .S(net103),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(net652),
    .A1(net662),
    .S(net103),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0631_ (.A0(net535),
    .A1(net590),
    .S(net103),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0632_ (.A0(net329),
    .A1(net565),
    .S(net103),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0633_ (.A0(net326),
    .A1(net333),
    .S(net102),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0634_ (.A0(net154),
    .A1(net311),
    .S(net102),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0635_ (.A0(net227),
    .A1(net275),
    .S(net102),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(net136),
    .A1(net188),
    .S(net102),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0637_ (.A0(net398),
    .A1(net469),
    .S(net102),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0638_ (.A0(net217),
    .A1(net273),
    .S(net102),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(net381),
    .A1(net424),
    .S(net102),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0640_ (.A0(net353),
    .A1(net359),
    .S(net102),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0641_ (.A0(net307),
    .A1(net331),
    .S(net102),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0642_ (.A0(net212),
    .A1(net271),
    .S(net102),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(net340),
    .A1(net387),
    .S(net102),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0644_ (.A0(net133),
    .A1(net146),
    .S(net102),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0645_ (.A0(net151),
    .A1(net166),
    .S(net102),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0646_ (.A0(net419),
    .A1(net451),
    .S(net102),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0647_ (.A0(net191),
    .A1(net214),
    .S(net102),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0648_ (.A0(net232),
    .A1(net251),
    .S(_0393_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(net278),
    .A1(net294),
    .S(net102),
    .X(_0089_));
 sky130_fd_sc_hd__and3b_2 _0650_ (.A_N(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(_0389_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _0651_ (.A0(net600),
    .A1(net563),
    .S(net113),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(net510),
    .A1(net506),
    .S(net113),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0653_ (.A0(net481),
    .A1(net439),
    .S(net113),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0654_ (.A0(net624),
    .A1(net588),
    .S(net113),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(net634),
    .A1(net528),
    .S(net113),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0656_ (.A0(net296),
    .A1(net235),
    .S(net113),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0657_ (.A0(net647),
    .A1(net643),
    .S(net113),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(net573),
    .A1(net538),
    .S(net113),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0659_ (.A0(net463),
    .A1(net422),
    .S(net113),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0660_ (.A0(net618),
    .A1(net525),
    .S(net113),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0661_ (.A0(net497),
    .A1(net224),
    .S(net113),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(net443),
    .A1(net368),
    .S(net113),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0663_ (.A0(net674),
    .A1(net652),
    .S(net113),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(net638),
    .A1(net535),
    .S(net113),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0665_ (.A0(net575),
    .A1(net329),
    .S(net113),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0666_ (.A0(net335),
    .A1(net326),
    .S(net112),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(net174),
    .A1(net154),
    .S(net112),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0668_ (.A0(net241),
    .A1(net227),
    .S(net112),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0669_ (.A0(net182),
    .A1(net136),
    .S(net112),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0670_ (.A0(net461),
    .A1(net398),
    .S(net112),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0671_ (.A0(net269),
    .A1(net217),
    .S(net112),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0672_ (.A0(net428),
    .A1(net381),
    .S(net112),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0673_ (.A0(net365),
    .A1(net353),
    .S(net112),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0674_ (.A0(net342),
    .A1(net307),
    .S(net112),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0675_ (.A0(net257),
    .A1(net212),
    .S(net112),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0676_ (.A0(net410),
    .A1(net340),
    .S(net112),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0677_ (.A0(net699),
    .A1(net133),
    .S(net112),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(net160),
    .A1(net151),
    .S(net112),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(net436),
    .A1(net419),
    .S(net112),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0680_ (.A0(net195),
    .A1(net191),
    .S(net112),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0681_ (.A0(net249),
    .A1(net232),
    .S(_0394_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0682_ (.A0(net304),
    .A1(net278),
    .S(net112),
    .X(_0121_));
 sky130_fd_sc_hd__or4_4 _0683_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(net1),
    .D(_0387_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _0684_ (.A0(net563),
    .A1(net594),
    .S(net111),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0685_ (.A0(net506),
    .A1(net512),
    .S(net111),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0686_ (.A0(net439),
    .A1(net709),
    .S(net111),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(net588),
    .A1(net707),
    .S(net111),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0688_ (.A0(net528),
    .A1(net713),
    .S(net111),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0689_ (.A0(net235),
    .A1(net722),
    .S(net111),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(net643),
    .A1(net658),
    .S(net111),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0691_ (.A0(net538),
    .A1(net602),
    .S(net111),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(net422),
    .A1(net432),
    .S(net111),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0693_ (.A0(net525),
    .A1(net612),
    .S(net111),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(net224),
    .A1(net720),
    .S(net111),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0695_ (.A0(net368),
    .A1(net378),
    .S(net111),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(net652),
    .A1(net670),
    .S(net111),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(net535),
    .A1(net550),
    .S(net111),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(net329),
    .A1(net383),
    .S(net111),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(net326),
    .A1(net385),
    .S(net110),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(net154),
    .A1(net176),
    .S(net110),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0701_ (.A0(net227),
    .A1(net282),
    .S(net110),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(net136),
    .A1(net197),
    .S(net110),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0703_ (.A0(net398),
    .A1(net471),
    .S(net110),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(net217),
    .A1(net245),
    .S(net110),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(net381),
    .A1(net704),
    .S(net110),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0706_ (.A0(net353),
    .A1(net402),
    .S(net110),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(net307),
    .A1(net706),
    .S(net110),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(net212),
    .A1(net701),
    .S(net110),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0709_ (.A0(net340),
    .A1(net708),
    .S(net110),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0710_ (.A0(net133),
    .A1(net138),
    .S(net110),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(net151),
    .A1(net164),
    .S(net110),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0712_ (.A0(net419),
    .A1(net453),
    .S(net110),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(net191),
    .A1(net207),
    .S(net110),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0714_ (.A0(net232),
    .A1(net239),
    .S(_0395_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(net278),
    .A1(net357),
    .S(net110),
    .X(_0153_));
 sky130_fd_sc_hd__nor3b_4 _0716_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C_N(_0389_),
    .Y(_0396_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(net596),
    .A1(net563),
    .S(net109),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(net530),
    .A1(net506),
    .S(net109),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(net501),
    .A1(net439),
    .S(net109),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _0720_ (.A0(net626),
    .A1(net588),
    .S(net109),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(net554),
    .A1(net528),
    .S(net109),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0722_ (.A0(net267),
    .A1(net235),
    .S(net109),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(net660),
    .A1(net643),
    .S(net109),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0724_ (.A0(net610),
    .A1(net538),
    .S(net109),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0725_ (.A0(net491),
    .A1(net422),
    .S(net109),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(net632),
    .A1(net525),
    .S(net109),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(net263),
    .A1(net224),
    .S(net109),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(net459),
    .A1(net368),
    .S(net109),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _0729_ (.A0(net672),
    .A1(net652),
    .S(net109),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(net556),
    .A1(net535),
    .S(net109),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _0731_ (.A0(net393),
    .A1(net329),
    .S(net109),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net695),
    .A1(net326),
    .S(net108),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _0733_ (.A0(net158),
    .A1(net154),
    .S(net108),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(net350),
    .A1(net227),
    .S(net108),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(net697),
    .A1(net136),
    .S(net108),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(net489),
    .A1(net398),
    .S(net108),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _0737_ (.A0(net323),
    .A1(net217),
    .S(net108),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(net487),
    .A1(net381),
    .S(net108),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _0739_ (.A0(net485),
    .A1(net353),
    .S(net108),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(net313),
    .A1(net307),
    .S(net108),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(net221),
    .A1(net212),
    .S(net108),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(net346),
    .A1(net340),
    .S(net108),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _0743_ (.A0(net148),
    .A1(net133),
    .S(net108),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(net702),
    .A1(net151),
    .S(net108),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _0745_ (.A0(net467),
    .A1(net419),
    .S(net108),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(net255),
    .A1(net191),
    .S(net108),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _0747_ (.A0(net715),
    .A1(net232),
    .S(_0396_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(net300),
    .A1(net278),
    .S(net108),
    .X(_0185_));
 sky130_fd_sc_hd__o41a_2 _0749_ (.A1(net684),
    .A2(net679),
    .A3(net681),
    .A4(net68),
    .B1(net67),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _0750_ (.A(net681),
    .B(net67),
    .Y(_0398_));
 sky130_fd_sc_hd__o211a_1 _0751_ (.A1(net681),
    .A2(_0397_),
    .B1(net682),
    .C1(_0276_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2b_1 _0752_ (.A_N(net68),
    .B(net679),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2b_1 _0753_ (.A_N(net679),
    .B(net68),
    .Y(_0400_));
 sky130_fd_sc_hd__a21oi_1 _0754_ (.A1(_0399_),
    .A2(_0400_),
    .B1(\fifo_in.count[0] ),
    .Y(_0401_));
 sky130_fd_sc_hd__and3_1 _0755_ (.A(\fifo_in.count[0] ),
    .B(_0399_),
    .C(_0400_),
    .X(_0402_));
 sky130_fd_sc_hd__o21ai_1 _0756_ (.A1(_0401_),
    .A2(_0402_),
    .B1(_0397_),
    .Y(_0403_));
 sky130_fd_sc_hd__o211a_1 _0757_ (.A1(net679),
    .A2(_0397_),
    .B1(_0403_),
    .C1(_0276_),
    .X(_0187_));
 sky130_fd_sc_hd__a21bo_1 _0758_ (.A1(net681),
    .A2(_0400_),
    .B1_N(_0399_),
    .X(_0404_));
 sky130_fd_sc_hd__xnor2_1 _0759_ (.A(net684),
    .B(net68),
    .Y(_0405_));
 sky130_fd_sc_hd__xnor2_1 _0760_ (.A(_0404_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__nor2_1 _0761_ (.A(net684),
    .B(_0397_),
    .Y(_0407_));
 sky130_fd_sc_hd__a211oi_1 _0762_ (.A1(_0397_),
    .A2(_0406_),
    .B1(_0407_),
    .C1(net1),
    .Y(_0188_));
 sky130_fd_sc_hd__or4bb_4 _0763_ (.A(net1),
    .B(_0387_),
    .C_N(\fifo_in.write_addr[2] ),
    .D_N(\fifo_in.write_addr[1] ),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(net563),
    .A1(net567),
    .S(net107),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(net506),
    .A1(net508),
    .S(net107),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _0766_ (.A0(net439),
    .A1(net493),
    .S(net107),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(net588),
    .A1(net636),
    .S(net107),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(net528),
    .A1(net620),
    .S(net107),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(net235),
    .A1(net284),
    .S(net107),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(net643),
    .A1(net721),
    .S(net107),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(net538),
    .A1(net585),
    .S(net107),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(net422),
    .A1(net718),
    .S(net107),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(net525),
    .A1(net548),
    .S(net107),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _0774_ (.A0(net224),
    .A1(net441),
    .S(net107),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0775_ (.A0(net368),
    .A1(net430),
    .S(net107),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(net652),
    .A1(net705),
    .S(net107),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(net535),
    .A1(net710),
    .S(net107),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(net329),
    .A1(net569),
    .S(net107),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(net326),
    .A1(net532),
    .S(net106),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(net154),
    .A1(net180),
    .S(net106),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _0781_ (.A0(net227),
    .A1(net261),
    .S(net106),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(net136),
    .A1(net172),
    .S(net106),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(net398),
    .A1(net725),
    .S(net106),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(net217),
    .A1(net726),
    .S(net106),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(net381),
    .A1(net412),
    .S(net106),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _0786_ (.A0(net353),
    .A1(net714),
    .S(net106),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(net307),
    .A1(net321),
    .S(_0408_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(net212),
    .A1(net265),
    .S(net106),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(net340),
    .A1(net374),
    .S(net106),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(net133),
    .A1(net186),
    .S(net106),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(net151),
    .A1(net209),
    .S(net106),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(net419),
    .A1(net477),
    .S(net106),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(net191),
    .A1(net711),
    .S(net106),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _0794_ (.A0(net232),
    .A1(net319),
    .S(net106),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(net278),
    .A1(net723),
    .S(net106),
    .X(_0220_));
 sky130_fd_sc_hd__a21o_1 _0796_ (.A1(net68),
    .A2(net67),
    .B1(net686),
    .X(_0265_));
 sky130_fd_sc_hd__and3_1 _0797_ (.A(_0276_),
    .B(_0387_),
    .C(net687),
    .X(_0221_));
 sky130_fd_sc_hd__a31o_1 _0798_ (.A1(net686),
    .A2(net68),
    .A3(net67),
    .B1(net689),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _0799_ (.A(_0276_),
    .B(_0391_),
    .C(net690),
    .X(_0222_));
 sky130_fd_sc_hd__nand2_1 _0800_ (.A(net676),
    .B(_0391_),
    .Y(_0267_));
 sky130_fd_sc_hd__a21oi_1 _0801_ (.A1(_0392_),
    .A2(net677),
    .B1(net1),
    .Y(_0223_));
 sky130_fd_sc_hd__or3_1 _0802_ (.A(net684),
    .B(net679),
    .C(net681),
    .X(_0268_));
 sky130_fd_sc_hd__and3b_1 _0803_ (.A_N(net68),
    .B(net67),
    .C(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__and4b_2 _0804_ (.A_N(net68),
    .B(net67),
    .C(_0268_),
    .D(net128),
    .X(_0270_));
 sky130_fd_sc_hd__nor2_1 _0805_ (.A(net1),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o21a_1 _0806_ (.A1(net128),
    .A2(_0269_),
    .B1(_0271_),
    .X(_0224_));
 sky130_fd_sc_hd__a21oi_1 _0807_ (.A1(net123),
    .A2(_0270_),
    .B1(net1),
    .Y(_0272_));
 sky130_fd_sc_hd__o21a_1 _0808_ (.A1(net123),
    .A2(_0270_),
    .B1(_0272_),
    .X(_0225_));
 sky130_fd_sc_hd__nand3_1 _0809_ (.A(net121),
    .B(net123),
    .C(_0270_),
    .Y(_0273_));
 sky130_fd_sc_hd__a21o_1 _0810_ (.A1(net123),
    .A2(_0270_),
    .B1(net121),
    .X(_0274_));
 sky130_fd_sc_hd__and3_1 _0811_ (.A(_0276_),
    .B(_0273_),
    .C(_0274_),
    .X(_0226_));
 sky130_fd_sc_hd__and3_2 _0812_ (.A(\fifo_in.write_addr[2] ),
    .B(\fifo_in.write_addr[1] ),
    .C(_0389_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(net640),
    .A1(net563),
    .S(net105),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(net516),
    .A1(net506),
    .S(net105),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _0815_ (.A0(net479),
    .A1(net439),
    .S(net105),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(net628),
    .A1(net588),
    .S(net105),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0817_ (.A0(net592),
    .A1(net528),
    .S(net105),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0818_ (.A0(net247),
    .A1(net235),
    .S(net105),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0819_ (.A0(net649),
    .A1(net643),
    .S(net105),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(net604),
    .A1(net538),
    .S(net105),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0821_ (.A0(net503),
    .A1(net422),
    .S(net105),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0822_ (.A0(net542),
    .A1(net525),
    .S(net105),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(net455),
    .A1(net224),
    .S(net105),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0824_ (.A0(net426),
    .A1(net368),
    .S(net105),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(net656),
    .A1(net652),
    .S(net105),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0826_ (.A0(net552),
    .A1(net535),
    .S(net105),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _0827_ (.A0(net616),
    .A1(net329),
    .S(net105),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(net337),
    .A1(net326),
    .S(net104),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(net700),
    .A1(net154),
    .S(net104),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0830_ (.A0(net698),
    .A1(net227),
    .S(net104),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(net156),
    .A1(net136),
    .S(net104),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(net400),
    .A1(net398),
    .S(net104),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0833_ (.A0(net229),
    .A1(net217),
    .S(net104),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _0834_ (.A0(net414),
    .A1(net381),
    .S(net104),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _0835_ (.A0(net404),
    .A1(net353),
    .S(net104),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _0836_ (.A0(net372),
    .A1(net307),
    .S(_0275_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(net253),
    .A1(net212),
    .S(net104),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(net370),
    .A1(net340),
    .S(net104),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _0839_ (.A0(net144),
    .A1(net133),
    .S(net104),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(net199),
    .A1(net151),
    .S(net104),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _0841_ (.A0(net696),
    .A1(net419),
    .S(net104),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _0842_ (.A0(net205),
    .A1(net191),
    .S(net104),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _0843_ (.A0(net348),
    .A1(net232),
    .S(net104),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(net286),
    .A1(net278),
    .S(net104),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(net563),
    .A1(net716),
    .S(net117),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(net506),
    .A1(net518),
    .S(net117),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _0847_ (.A0(net439),
    .A1(net457),
    .S(net117),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(net588),
    .A1(net608),
    .S(net117),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(net528),
    .A1(net560),
    .S(net117),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _0850_ (.A0(net235),
    .A1(net317),
    .S(net117),
    .X(_0264_));
 sky130_fd_sc_hd__dfxtp_1 _0851_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net655),
    .Q(\fifo_in.FIFO[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0852_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net539),
    .Q(\fifo_in.FIFO[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0853_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net521),
    .Q(\fifo_in.FIFO[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0854_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net541),
    .Q(\fifo_in.FIFO[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0855_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net515),
    .Q(\fifo_in.FIFO[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0856_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net390),
    .Q(\fifo_in.FIFO[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0857_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net667),
    .Q(\fifo_in.FIFO[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0858_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net584),
    .Q(\fifo_in.FIFO[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0859_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net607),
    .Q(\fifo_in.FIFO[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0860_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net392),
    .Q(\fifo_in.FIFO[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0861_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net163),
    .Q(\fifo_in.FIFO[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0862_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net244),
    .Q(\fifo_in.FIFO[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0863_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net179),
    .Q(\fifo_in.FIFO[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0864_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net417),
    .Q(\fifo_in.FIFO[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0865_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net238),
    .Q(\fifo_in.FIFO[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0866_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net407),
    .Q(\fifo_in.FIFO[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0867_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net356),
    .Q(\fifo_in.FIFO[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0868_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net310),
    .Q(\fifo_in.FIFO[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0869_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net260),
    .Q(\fifo_in.FIFO[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0870_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net362),
    .Q(\fifo_in.FIFO[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0871_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net141),
    .Q(\fifo_in.FIFO[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0872_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net194),
    .Q(\fifo_in.FIFO[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0873_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net435),
    .Q(\fifo_in.FIFO[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0874_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net202),
    .Q(\fifo_in.FIFO[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0875_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net291),
    .Q(\fifo_in.FIFO[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0876_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net293),
    .Q(\fifo_in.FIFO[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0877_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net631),
    .Q(\fifo_in.FIFO[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0878_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net547),
    .Q(\fifo_in.FIFO[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0879_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net500),
    .Q(\fifo_in.FIFO[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0880_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net623),
    .Q(\fifo_in.FIFO[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0881_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net578),
    .Q(\fifo_in.FIFO[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0882_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net281),
    .Q(\fifo_in.FIFO[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0883_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net665),
    .Q(\fifo_in.FIFO[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0884_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net572),
    .Q(\fifo_in.FIFO[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0885_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net474),
    .Q(\fifo_in.FIFO[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0886_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net545),
    .Q(\fifo_in.FIFO[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0887_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net523),
    .Q(\fifo_in.FIFO[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0888_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net476),
    .Q(\fifo_in.FIFO[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0889_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net669),
    .Q(\fifo_in.FIFO[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0890_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net559),
    .Q(\fifo_in.FIFO[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0891_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net330),
    .Q(\fifo_in.FIFO[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0892_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net377),
    .Q(\fifo_in.FIFO[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0893_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net169),
    .Q(\fifo_in.FIFO[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0894_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net299),
    .Q(\fifo_in.FIFO[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0895_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net143),
    .Q(\fifo_in.FIFO[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0896_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net446),
    .Q(\fifo_in.FIFO[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0897_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net220),
    .Q(\fifo_in.FIFO[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0898_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net396),
    .Q(\fifo_in.FIFO[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0899_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net466),
    .Q(\fifo_in.FIFO[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0900_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net364),
    .Q(\fifo_in.FIFO[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0901_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net345),
    .Q(\fifo_in.FIFO[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0902_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net409),
    .Q(\fifo_in.FIFO[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0903_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net185),
    .Q(\fifo_in.FIFO[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0904_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net171),
    .Q(\fifo_in.FIFO[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0905_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net448),
    .Q(\fifo_in.FIFO[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0906_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net204),
    .Q(\fifo_in.FIFO[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0907_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net316),
    .Q(\fifo_in.FIFO[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0908_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net303),
    .Q(\fifo_in.FIFO[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0909_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net580),
    .Q(\fifo_in.FIFO[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0910_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net507),
    .Q(\fifo_in.FIFO[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0911_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net450),
    .Q(\fifo_in.FIFO[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0912_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net615),
    .Q(\fifo_in.FIFO[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0913_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net582),
    .Q(\fifo_in.FIFO[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0914_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net289),
    .Q(\fifo_in.FIFO[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0915_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net646),
    .Q(\fifo_in.FIFO[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0916_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net599),
    .Q(\fifo_in.FIFO[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0917_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net496),
    .Q(\fifo_in.FIFO[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0918_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net526),
    .Q(\fifo_in.FIFO[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0919_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net484),
    .Q(\fifo_in.FIFO[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0920_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net369),
    .Q(\fifo_in.FIFO[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0921_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net663),
    .Q(\fifo_in.FIFO[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0922_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net591),
    .Q(\fifo_in.FIFO[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0923_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net566),
    .Q(\fifo_in.FIFO[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0924_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net334),
    .Q(\fifo_in.FIFO[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0925_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net312),
    .Q(\fifo_in.FIFO[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0926_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net276),
    .Q(\fifo_in.FIFO[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0927_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net189),
    .Q(\fifo_in.FIFO[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0928_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net470),
    .Q(\fifo_in.FIFO[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0929_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net274),
    .Q(\fifo_in.FIFO[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0930_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net425),
    .Q(\fifo_in.FIFO[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0931_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net360),
    .Q(\fifo_in.FIFO[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0932_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net332),
    .Q(\fifo_in.FIFO[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0933_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net272),
    .Q(\fifo_in.FIFO[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0934_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net388),
    .Q(\fifo_in.FIFO[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0935_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net147),
    .Q(\fifo_in.FIFO[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0936_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net167),
    .Q(\fifo_in.FIFO[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0937_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net452),
    .Q(\fifo_in.FIFO[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0938_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net215),
    .Q(\fifo_in.FIFO[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0939_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net252),
    .Q(\fifo_in.FIFO[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0940_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net295),
    .Q(\fifo_in.FIFO[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0941_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net601),
    .Q(\fifo_in.FIFO[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0942_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net511),
    .Q(\fifo_in.FIFO[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0943_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net482),
    .Q(\fifo_in.FIFO[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0944_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net625),
    .Q(\fifo_in.FIFO[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0945_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net635),
    .Q(\fifo_in.FIFO[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0946_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net297),
    .Q(\fifo_in.FIFO[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0947_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net648),
    .Q(\fifo_in.FIFO[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0948_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net574),
    .Q(\fifo_in.FIFO[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0949_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net464),
    .Q(\fifo_in.FIFO[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0950_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net619),
    .Q(\fifo_in.FIFO[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0951_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net498),
    .Q(\fifo_in.FIFO[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0952_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net444),
    .Q(\fifo_in.FIFO[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0953_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net675),
    .Q(\fifo_in.FIFO[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0954_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net639),
    .Q(\fifo_in.FIFO[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0955_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net576),
    .Q(\fifo_in.FIFO[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0956_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net336),
    .Q(\fifo_in.FIFO[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0957_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net175),
    .Q(\fifo_in.FIFO[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0958_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net242),
    .Q(\fifo_in.FIFO[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0959_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net183),
    .Q(\fifo_in.FIFO[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0960_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net462),
    .Q(\fifo_in.FIFO[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0961_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net270),
    .Q(\fifo_in.FIFO[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net429),
    .Q(\fifo_in.FIFO[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net366),
    .Q(\fifo_in.FIFO[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net343),
    .Q(\fifo_in.FIFO[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net258),
    .Q(\fifo_in.FIFO[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net411),
    .Q(\fifo_in.FIFO[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net134),
    .Q(\fifo_in.FIFO[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net161),
    .Q(\fifo_in.FIFO[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net437),
    .Q(\fifo_in.FIFO[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _0970_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net196),
    .Q(\fifo_in.FIFO[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _0971_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net250),
    .Q(\fifo_in.FIFO[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _0972_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net305),
    .Q(\fifo_in.FIFO[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _0973_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net595),
    .Q(\fifo_in.FIFO[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0974_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net513),
    .Q(\fifo_in.FIFO[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0975_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net440),
    .Q(\fifo_in.FIFO[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0976_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net589),
    .Q(\fifo_in.FIFO[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0977_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net529),
    .Q(\fifo_in.FIFO[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0978_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net236),
    .Q(\fifo_in.FIFO[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0979_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net659),
    .Q(\fifo_in.FIFO[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0980_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net603),
    .Q(\fifo_in.FIFO[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0981_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net433),
    .Q(\fifo_in.FIFO[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _0982_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net613),
    .Q(\fifo_in.FIFO[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _0983_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net225),
    .Q(\fifo_in.FIFO[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net379),
    .Q(\fifo_in.FIFO[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net671),
    .Q(\fifo_in.FIFO[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net551),
    .Q(\fifo_in.FIFO[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net384),
    .Q(\fifo_in.FIFO[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net386),
    .Q(\fifo_in.FIFO[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net177),
    .Q(\fifo_in.FIFO[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net283),
    .Q(\fifo_in.FIFO[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net198),
    .Q(\fifo_in.FIFO[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net472),
    .Q(\fifo_in.FIFO[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net246),
    .Q(\fifo_in.FIFO[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net382),
    .Q(\fifo_in.FIFO[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net403),
    .Q(\fifo_in.FIFO[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net308),
    .Q(\fifo_in.FIFO[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net213),
    .Q(\fifo_in.FIFO[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net341),
    .Q(\fifo_in.FIFO[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net139),
    .Q(\fifo_in.FIFO[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net165),
    .Q(\fifo_in.FIFO[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net454),
    .Q(\fifo_in.FIFO[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net208),
    .Q(\fifo_in.FIFO[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net240),
    .Q(\fifo_in.FIFO[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net358),
    .Q(\fifo_in.FIFO[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net597),
    .Q(\fifo_in.FIFO[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net531),
    .Q(\fifo_in.FIFO[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net502),
    .Q(\fifo_in.FIFO[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net627),
    .Q(\fifo_in.FIFO[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net555),
    .Q(\fifo_in.FIFO[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net268),
    .Q(\fifo_in.FIFO[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net661),
    .Q(\fifo_in.FIFO[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net611),
    .Q(\fifo_in.FIFO[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net492),
    .Q(\fifo_in.FIFO[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net633),
    .Q(\fifo_in.FIFO[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net264),
    .Q(\fifo_in.FIFO[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net460),
    .Q(\fifo_in.FIFO[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net673),
    .Q(\fifo_in.FIFO[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net557),
    .Q(\fifo_in.FIFO[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net394),
    .Q(\fifo_in.FIFO[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net327),
    .Q(\fifo_in.FIFO[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net159),
    .Q(\fifo_in.FIFO[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net351),
    .Q(\fifo_in.FIFO[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net137),
    .Q(\fifo_in.FIFO[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net490),
    .Q(\fifo_in.FIFO[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net324),
    .Q(\fifo_in.FIFO[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net488),
    .Q(\fifo_in.FIFO[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net486),
    .Q(\fifo_in.FIFO[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net314),
    .Q(\fifo_in.FIFO[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net222),
    .Q(\fifo_in.FIFO[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net347),
    .Q(\fifo_in.FIFO[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net149),
    .Q(\fifo_in.FIFO[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net152),
    .Q(\fifo_in.FIFO[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net468),
    .Q(\fifo_in.FIFO[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net256),
    .Q(\fifo_in.FIFO[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net233),
    .Q(\fifo_in.FIFO[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net301),
    .Q(\fifo_in.FIFO[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net683),
    .Q(\fifo_in.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net680),
    .Q(\fifo_in.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net685),
    .Q(\fifo_in.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net568),
    .Q(\fifo_in.FIFO[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net509),
    .Q(\fifo_in.FIFO[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net494),
    .Q(\fifo_in.FIFO[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net637),
    .Q(\fifo_in.FIFO[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net621),
    .Q(\fifo_in.FIFO[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net285),
    .Q(\fifo_in.FIFO[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net644),
    .Q(\fifo_in.FIFO[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net586),
    .Q(\fifo_in.FIFO[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net423),
    .Q(\fifo_in.FIFO[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net549),
    .Q(\fifo_in.FIFO[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net442),
    .Q(\fifo_in.FIFO[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net431),
    .Q(\fifo_in.FIFO[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net653),
    .Q(\fifo_in.FIFO[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net536),
    .Q(\fifo_in.FIFO[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net570),
    .Q(\fifo_in.FIFO[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net533),
    .Q(\fifo_in.FIFO[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net181),
    .Q(\fifo_in.FIFO[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net262),
    .Q(\fifo_in.FIFO[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net173),
    .Q(\fifo_in.FIFO[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net399),
    .Q(\fifo_in.FIFO[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net218),
    .Q(\fifo_in.FIFO[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net413),
    .Q(\fifo_in.FIFO[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net354),
    .Q(\fifo_in.FIFO[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net322),
    .Q(\fifo_in.FIFO[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net266),
    .Q(\fifo_in.FIFO[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net375),
    .Q(\fifo_in.FIFO[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net187),
    .Q(\fifo_in.FIFO[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net210),
    .Q(\fifo_in.FIFO[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net478),
    .Q(\fifo_in.FIFO[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net192),
    .Q(\fifo_in.FIFO[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net320),
    .Q(\fifo_in.FIFO[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net279),
    .Q(\fifo_in.FIFO[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net688),
    .Q(\fifo_in.write_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1073_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net691),
    .Q(\fifo_in.write_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1074_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net678),
    .Q(\fifo_in.write_addr[2] ));
 sky130_fd_sc_hd__dfxtp_4 _1075_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net693),
    .Q(\fifo_in.read_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0225_),
    .Q(\fifo_in.read_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1077_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0226_),
    .Q(\fifo_in.read_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net641),
    .Q(\fifo_in.FIFO[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net517),
    .Q(\fifo_in.FIFO[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net480),
    .Q(\fifo_in.FIFO[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net629),
    .Q(\fifo_in.FIFO[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net593),
    .Q(\fifo_in.FIFO[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net248),
    .Q(\fifo_in.FIFO[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net650),
    .Q(\fifo_in.FIFO[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net605),
    .Q(\fifo_in.FIFO[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net504),
    .Q(\fifo_in.FIFO[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net543),
    .Q(\fifo_in.FIFO[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net456),
    .Q(\fifo_in.FIFO[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net427),
    .Q(\fifo_in.FIFO[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net657),
    .Q(\fifo_in.FIFO[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net553),
    .Q(\fifo_in.FIFO[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net617),
    .Q(\fifo_in.FIFO[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net338),
    .Q(\fifo_in.FIFO[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net155),
    .Q(\fifo_in.FIFO[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net228),
    .Q(\fifo_in.FIFO[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net157),
    .Q(\fifo_in.FIFO[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net401),
    .Q(\fifo_in.FIFO[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net230),
    .Q(\fifo_in.FIFO[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net415),
    .Q(\fifo_in.FIFO[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net405),
    .Q(\fifo_in.FIFO[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net373),
    .Q(\fifo_in.FIFO[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net254),
    .Q(\fifo_in.FIFO[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net371),
    .Q(\fifo_in.FIFO[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net145),
    .Q(\fifo_in.FIFO[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net200),
    .Q(\fifo_in.FIFO[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net420),
    .Q(\fifo_in.FIFO[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net206),
    .Q(\fifo_in.FIFO[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net349),
    .Q(\fifo_in.FIFO[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net287),
    .Q(\fifo_in.FIFO[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net564),
    .Q(\fifo_in.FIFO[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net519),
    .Q(\fifo_in.FIFO[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net458),
    .Q(\fifo_in.FIFO[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net609),
    .Q(\fifo_in.FIFO[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net561),
    .Q(\fifo_in.FIFO[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net318),
    .Q(\fifo_in.FIFO[5][5] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_8 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_0393_),
    .X(net103));
 sky130_fd_sc_hd__buf_8 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(_0275_),
    .X(net105));
 sky130_fd_sc_hd__buf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_0408_),
    .X(net107));
 sky130_fd_sc_hd__buf_8 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_8 fanout109 (.A(_0396_),
    .X(net109));
 sky130_fd_sc_hd__buf_6 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_8 fanout111 (.A(_0395_),
    .X(net111));
 sky130_fd_sc_hd__buf_8 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_8 fanout113 (.A(_0394_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(_0390_),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(_0388_),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout121 (.A(net694),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(\fifo_in.read_addr[2] ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_6 fanout124 (.A(net127),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net127),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(\fifo_in.read_addr[1] ),
    .X(net127));
 sky130_fd_sc_hd__buf_6 fanout128 (.A(net692),
    .X(net128));
 sky130_fd_sc_hd__buf_8 fanout129 (.A(\fifo_in.read_addr[0] ),
    .X(net129));
 sky130_fd_sc_hd__buf_8 fanout130 (.A(\fifo_in.read_addr[0] ),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(\fifo_in.read_addr[0] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wbs_dat_i[26]),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0020_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(wbs_dat_i[30]),
    .X(net231));
 sky130_fd_sc_hd__buf_2 hold101 (.A(net58),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0184_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(wbs_dat_i[5]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 hold104 (.A(net62),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0127_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\fifo_in.FIFO[5][20] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0014_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\fifo_in.FIFO[1][30] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0152_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\fifo_in.FIFO[4][18] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\fifo_in.FIFO[2][17] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0107_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\fifo_in.FIFO[5][17] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0011_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\fifo_in.FIFO[1][20] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0142_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\fifo_in.FIFO[6][5] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0232_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\fifo_in.FIFO[2][30] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0120_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0044_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\fifo_in.FIFO[3][30] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0088_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\fifo_in.FIFO[6][24] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0251_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\fifo_in.FIFO[0][29] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0183_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\fifo_in.FIFO[2][24] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0114_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\fifo_in.FIFO[5][24] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0018_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\fifo_in.FIFO[6][26] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\fifo_in.FIFO[7][17] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0206_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\fifo_in.FIFO[0][10] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0164_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\fifo_in.FIFO[7][24] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0213_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\fifo_in.FIFO[0][5] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0159_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\fifo_in.FIFO[2][20] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0110_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0253_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\fifo_in.FIFO[3][24] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0082_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\fifo_in.FIFO[3][20] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0078_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\fifo_in.FIFO[3][17] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0075_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(wbs_dat_i[31]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 hold147 (.A(net59),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0220_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\fifo_in.FIFO[4][5] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\fifo_in.FIFO[3][26] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0031_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\fifo_in.FIFO[1][17] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0139_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\fifo_in.FIFO[7][5] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0194_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\fifo_in.FIFO[6][31] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0258_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\fifo_in.FIFO[3][5] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0063_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\fifo_in.FIFO[5][30] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0084_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0024_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\fifo_in.FIFO[5][31] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0025_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\fifo_in.FIFO[3][31] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0089_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\fifo_in.FIFO[2][5] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0095_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\fifo_in.FIFO[4][17] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0043_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\fifo_in.FIFO[0][31] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\fifo_in.FIFO[0][26] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0185_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\fifo_in.FIFO[4][31] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0057_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\fifo_in.FIFO[2][31] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0121_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(wbs_dat_i[23]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 hold176 (.A(net50),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0145_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\fifo_in.FIFO[5][23] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0017_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0180_),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\fifo_in.FIFO[3][16] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0074_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\fifo_in.FIFO[0][23] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_0177_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\fifo_in.FIFO[4][30] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0056_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\fifo_in.FIFO[5][5] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0264_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\fifo_in.FIFO[7][30] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0219_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(wbs_dat_i[27]),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\fifo_in.FIFO[7][23] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0212_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\fifo_in.FIFO[0][20] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0174_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(wbs_dat_i[15]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_2 hold195 (.A(net41),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0169_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(wbs_dat_i[14]),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 hold198 (.A(net40),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0040_),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 hold2 (.A(net53),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 hold20 (.A(net54),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\fifo_in.FIFO[3][23] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0081_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\fifo_in.FIFO[3][15] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0073_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\fifo_in.FIFO[2][15] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0105_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\fifo_in.FIFO[6][15] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0242_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(wbs_dat_i[25]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 hold209 (.A(net52),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0181_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0147_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\fifo_in.FIFO[2][23] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0113_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\fifo_in.FIFO[4][24] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0050_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\fifo_in.FIFO[0][25] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0179_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\fifo_in.FIFO[6][30] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0257_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\fifo_in.FIFO[0][17] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(wbs_dat_i[16]),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0171_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(wbs_dat_i[22]),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 hold222 (.A(net49),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0211_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\fifo_in.FIFO[5][22] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0016_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\fifo_in.FIFO[1][31] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0153_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\fifo_in.FIFO[3][22] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0080_),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 hold23 (.A(net42),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\fifo_in.FIFO[5][25] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0019_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\fifo_in.FIFO[4][23] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0049_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\fifo_in.FIFO[2][22] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0112_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(wbs_dat_i[11]),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_2 hold237 (.A(net37),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0069_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\fifo_in.FIFO[6][25] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0243_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0252_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\fifo_in.FIFO[6][23] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0250_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\fifo_in.FIFO[7][25] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0214_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\fifo_in.FIFO[4][15] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0041_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\fifo_in.FIFO[1][11] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0133_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(wbs_dat_i[21]),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\fifo_in.FIFO[6][18] ),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 hold250 (.A(net48),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0143_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\fifo_in.FIFO[1][14] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_0136_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\fifo_in.FIFO[1][15] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0137_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\fifo_in.FIFO[3][25] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0083_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\fifo_in.FIFO[5][11] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_0005_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0245_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\fifo_in.FIFO[5][15] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0009_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\fifo_in.FIFO[0][14] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0168_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\fifo_in.FIFO[4][21] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_0047_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(wbs_dat_i[19]),
    .X(net397));
 sky130_fd_sc_hd__buf_2 hold267 (.A(net45),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0208_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\fifo_in.FIFO[6][19] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\fifo_in.FIFO[0][16] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0246_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\fifo_in.FIFO[1][22] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0144_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\fifo_in.FIFO[6][22] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0249_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\fifo_in.FIFO[5][21] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0015_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\fifo_in.FIFO[4][25] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0051_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\fifo_in.FIFO[2][25] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0170_),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0115_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\fifo_in.FIFO[7][21] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0210_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\fifo_in.FIFO[6][21] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0248_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\fifo_in.FIFO[5][19] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0013_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(wbs_dat_i[28]),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 hold288 (.A(net55),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0255_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\fifo_in.FIFO[2][27] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(wbs_dat_i[8]),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_2 hold291 (.A(net65),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0197_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\fifo_in.FIFO[3][21] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0079_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\fifo_in.FIFO[6][11] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0238_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\fifo_in.FIFO[2][21] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0111_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\fifo_in.FIFO[7][11] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0116_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0117_),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0200_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\fifo_in.FIFO[1][8] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0130_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\fifo_in.FIFO[5][28] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0022_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\fifo_in.FIFO[2][28] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0118_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(wbs_dat_i[2]),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_2 hold308 (.A(net57),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0124_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\fifo_in.FIFO[5][16] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\fifo_in.FIFO[7][10] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0199_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\fifo_in.FIFO[2][11] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0101_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\fifo_in.FIFO[4][19] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_0045_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\fifo_in.FIFO[4][28] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0054_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\fifo_in.FIFO[3][2] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0060_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0010_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\fifo_in.FIFO[3][28] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0086_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\fifo_in.FIFO[1][28] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0150_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\fifo_in.FIFO[6][10] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_0237_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\fifo_in.FIFO[5][2] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0261_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\fifo_in.FIFO[0][11] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0165_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\fifo_in.FIFO[1][27] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\fifo_in.FIFO[2][19] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0109_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\fifo_in.FIFO[2][8] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0098_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\fifo_in.FIFO[4][22] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0048_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\fifo_in.FIFO[0][28] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0182_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\fifo_in.FIFO[3][19] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0077_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0149_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\fifo_in.FIFO[1][19] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0141_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\fifo_in.FIFO[4][8] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_0034_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\fifo_in.FIFO[4][11] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0037_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\fifo_in.FIFO[7][28] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0217_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\fifo_in.FIFO[6][2] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0229_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\fifo_in.FIFO[3][27] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\fifo_in.FIFO[2][2] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_0092_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\fifo_in.FIFO[3][10] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_0068_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\fifo_in.FIFO[0][22] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_0176_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\fifo_in.FIFO[0][21] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_0175_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\fifo_in.FIFO[0][19] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(_0173_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0085_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\fifo_in.FIFO[0][8] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_0162_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\fifo_in.FIFO[7][2] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_0191_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\fifo_in.FIFO[3][8] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(_0066_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\fifo_in.FIFO[2][10] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(_0100_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\fifo_in.FIFO[4][2] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_0028_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\fifo_in.FIFO[4][16] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\fifo_in.FIFO[0][2] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(_0156_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\fifo_in.FIFO[6][8] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(_0235_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(wbs_dat_i[1]),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_2 hold375 (.A(net46),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0059_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\fifo_in.FIFO[7][1] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0190_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\fifo_in.FIFO[2][1] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0042_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0091_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\fifo_in.FIFO[1][1] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0123_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\fifo_in.FIFO[5][10] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0004_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\fifo_in.FIFO[6][1] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0228_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\fifo_in.FIFO[5][1] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0260_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\fifo_in.FIFO[5][8] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\fifo_in.FIFO[4][27] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0002_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\fifo_in.FIFO[4][10] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0036_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(wbs_dat_i[9]),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_2 hold394 (.A(net66),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_0067_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(wbs_dat_i[4]),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_2 hold397 (.A(net61),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0126_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\fifo_in.FIFO[0][1] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(wbs_dat_i[18]),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0053_),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0155_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\fifo_in.FIFO[7][15] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0204_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(wbs_dat_i[13]),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 hold404 (.A(net39),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_0202_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(wbs_dat_i[7]),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_2 hold407 (.A(net64),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0001_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\fifo_in.FIFO[5][9] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\fifo_in.FIFO[7][18] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0003_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\fifo_in.FIFO[6][9] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0236_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\fifo_in.FIFO[4][9] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0035_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\fifo_in.FIFO[4][1] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0027_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\fifo_in.FIFO[7][9] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0198_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\fifo_in.FIFO[1][13] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0207_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0135_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\fifo_in.FIFO[6][13] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0240_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\fifo_in.FIFO[0][4] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0158_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\fifo_in.FIFO[0][13] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0167_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\fifo_in.FIFO[4][13] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0039_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\fifo_in.FIFO[5][4] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\fifo_in.FIFO[2][16] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0263_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(wbs_dat_i[0]),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_2 hold432 (.A(net35),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_0259_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\fifo_in.FIFO[3][14] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(_0072_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\fifo_in.FIFO[7][0] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_0189_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\fifo_in.FIFO[7][14] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_0203_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0106_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\fifo_in.FIFO[4][7] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_0033_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\fifo_in.FIFO[2][7] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(_0097_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\fifo_in.FIFO[2][14] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_0104_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\fifo_in.FIFO[4][4] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_0030_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\fifo_in.FIFO[3][0] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(_0058_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\fifo_in.FIFO[1][16] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\fifo_in.FIFO[3][4] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_0062_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\fifo_in.FIFO[5][13] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_0007_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\fifo_in.FIFO[7][7] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_0196_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(wbs_dat_i[3]),
    .X(net587));
 sky130_fd_sc_hd__buf_2 hold457 (.A(net60),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0125_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\fifo_in.FIFO[3][13] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0138_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0071_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\fifo_in.FIFO[6][4] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0231_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\fifo_in.FIFO[1][0] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0122_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\fifo_in.FIFO[0][0] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0154_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\fifo_in.FIFO[3][7] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0065_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\fifo_in.FIFO[2][0] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\fifo_in.FIFO[5][18] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_0090_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\fifo_in.FIFO[1][7] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_0129_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\fifo_in.FIFO[6][7] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_0234_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\fifo_in.FIFO[5][14] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_0008_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\fifo_in.FIFO[5][3] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_0262_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\fifo_in.FIFO[0][7] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0012_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_0161_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\fifo_in.FIFO[1][9] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0131_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\fifo_in.FIFO[3][3] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_0061_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\fifo_in.FIFO[6][14] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0241_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\fifo_in.FIFO[2][9] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0099_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\fifo_in.FIFO[7][4] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\fifo_in.FIFO[7][16] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_0193_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\fifo_in.FIFO[4][3] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0029_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\fifo_in.FIFO[2][3] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0093_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\fifo_in.FIFO[0][3] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_0157_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\fifo_in.FIFO[6][3] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_0230_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\fifo_in.FIFO[4][0] ),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_2 hold5 (.A(net44),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0205_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0026_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\fifo_in.FIFO[0][9] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0163_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\fifo_in.FIFO[2][4] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0094_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\fifo_in.FIFO[7][3] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0192_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\fifo_in.FIFO[2][13] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0103_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\fifo_in.FIFO[6][0] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\fifo_in.FIFO[2][18] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0227_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(wbs_dat_i[6]),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_2 hold512 (.A(net63),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0195_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\fifo_in.FIFO[3][6] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0064_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\fifo_in.FIFO[2][6] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_0096_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\fifo_in.FIFO[6][6] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_0233_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0108_),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(wbs_dat_i[12]),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_2 hold521 (.A(net38),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0201_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\fifo_in.FIFO[5][6] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0000_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\fifo_in.FIFO[6][12] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0239_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\fifo_in.FIFO[1][6] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0128_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\fifo_in.FIFO[0][6] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\fifo_in.FIFO[4][26] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0160_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\fifo_in.FIFO[3][12] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0070_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\fifo_in.FIFO[4][6] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0032_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\fifo_in.FIFO[5][12] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0006_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\fifo_in.FIFO[4][12] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0038_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\fifo_in.FIFO[1][12] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0052_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0134_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\fifo_in.FIFO[0][12] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0166_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\fifo_in.FIFO[2][12] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0102_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\fifo_in.write_addr[2] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0267_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_0223_),
    .X(net678));
 sky130_fd_sc_hd__buf_1 hold548 (.A(\fifo_in.count[1] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_0187_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\fifo_in.FIFO[7][26] ),
    .X(net186));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold550 (.A(\fifo_in.count[0] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_0398_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0186_),
    .X(net683));
 sky130_fd_sc_hd__buf_1 hold553 (.A(\fifo_in.count[2] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0188_),
    .X(net685));
 sky130_fd_sc_hd__buf_1 hold555 (.A(\fifo_in.write_addr[0] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_0265_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0221_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\fifo_in.write_addr[1] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0266_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0215_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0222_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\fifo_in.read_addr[0] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0224_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\fifo_in.read_addr[2] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\fifo_in.FIFO[0][15] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\fifo_in.FIFO[6][28] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\fifo_in.FIFO[0][18] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\fifo_in.FIFO[6][17] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\fifo_in.FIFO[2][26] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\fifo_in.FIFO[6][16] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\fifo_in.FIFO[3][18] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\fifo_in.FIFO[1][24] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\fifo_in.FIFO[0][27] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\fifo_in.FIFO[4][14] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\fifo_in.FIFO[1][21] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\fifo_in.FIFO[7][12] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\fifo_in.FIFO[1][23] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\fifo_in.FIFO[1][3] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\fifo_in.FIFO[1][25] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\fifo_in.FIFO[1][2] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\fifo_in.FIFO[7][13] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0076_),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\fifo_in.FIFO[7][29] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\fifo_in.FIFO[3][1] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\fifo_in.FIFO[1][4] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\fifo_in.FIFO[7][22] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\fifo_in.FIFO[0][30] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\fifo_in.FIFO[5][0] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\fifo_in.FIFO[3][9] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\fifo_in.FIFO[7][8] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\fifo_in.FIFO[3][11] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\fifo_in.FIFO[1][10] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(wbs_dat_i[29]),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\fifo_in.FIFO[7][6] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\fifo_in.FIFO[1][5] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\fifo_in.FIFO[7][31] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\fifo_in.FIFO[5][7] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\fifo_in.FIFO[7][19] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\fifo_in.FIFO[7][20] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0172_),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 hold60 (.A(net56),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0218_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\fifo_in.FIFO[5][27] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0021_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\fifo_in.FIFO[2][29] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0119_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\fifo_in.FIFO[1][18] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0140_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\fifo_in.FIFO[6][27] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0254_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\fifo_in.FIFO[1][26] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\fifo_in.FIFO[5][29] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0023_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\fifo_in.FIFO[4][29] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0055_),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\fifo_in.FIFO[6][29] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0256_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\fifo_in.FIFO[1][29] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0151_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\fifo_in.FIFO[7][27] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0216_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0148_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(wbs_dat_i[24]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 hold81 (.A(net51),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0146_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\fifo_in.FIFO[3][29] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0087_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(wbs_dat_i[20]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 hold86 (.A(net47),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0209_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\fifo_in.FIFO[4][20] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0046_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\fifo_in.FIFO[5][26] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\fifo_in.FIFO[0][24] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_0178_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(wbs_dat_i[10]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 hold93 (.A(net36),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0132_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(wbs_dat_i[17]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 hold96 (.A(net43),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0244_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\fifo_in.FIFO[6][20] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0247_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(wbs_adr_i[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wbs_adr_i[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(wbs_adr_i[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(wbs_adr_i[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(wbs_adr_i[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(wbs_adr_i[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(wbs_adr_i[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(wbs_adr_i[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(wbs_adr_i[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(wbs_adr_i[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(wbs_adr_i[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(wbs_adr_i[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(wbs_adr_i[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(wbs_adr_i[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(wbs_adr_i[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(wbs_adr_i[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(wbs_adr_i[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(wbs_adr_i[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(wbs_adr_i[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(wbs_adr_i[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(wbs_adr_i[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(wbs_adr_i[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(wbs_adr_i[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(wbs_adr_i[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(wbs_adr_i[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(wbs_adr_i[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(wbs_cyc_i),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(net562),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(net223),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(net367),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(net651),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(net534),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(wbs_adr_i[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(net328),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(net325),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(net153),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(net226),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(net135),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(net397),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(net505),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(net216),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(net380),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(net352),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(wbs_adr_i[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(net306),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(net211),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(net339),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(net132),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(net150),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(net418),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(net190),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(net438),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(net231),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(net277),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(wbs_adr_i[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(net587),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(net527),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(net234),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(net642),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(net537),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(net421),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(net524),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(wbs_stb_i),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(wbs_we_i),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(wbs_adr_i[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(wbs_adr_i[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(wbs_adr_i[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 max_cap118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 max_cap119 (.A(_0290_),
    .X(net119));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net120),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_1 wire120 (.A(net69),
    .X(net120));
endmodule

